-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HLT1Qw/HpdDFjcTFSa2lA1LPig6lNANd7YW+1y3uigsvr22670oGyIe4iHR0I+qbZFoMPGQpOSyJ
rEzn89LTnhJ39hxn3/X1mKkGi1nMkFDRM3/LS7KQ2z3GEAWRSadQxMPJbFEbog2IxX796a4wCJqs
slUzdUoQxJAIpCVmVegB8z5Zd+gbCL+nYjiKl6xQ9BXADSuCX+rzWRevH23OrqiL3KMKd1R8LSaG
SgihbHeMqGtiRNDkN/C0Gr010o6CZ56rgU6hhnYf0yLgmVRVNkXde3G9vvZo/+XEzBHfijGfDxvr
KUsLCzbp/O0mQvLn0EYIzX0UBz/eI5wZV0VQOg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9616)
`protect data_block
98Cr0etAQc7Y3KnahKSgZ3fVCvVsNh5A8fVomIiL1dVF1TcncP+bOuzVDTeHjviPcUv/8TJ4KPQE
DmXeK6LOTnnbOjBvYlptfjNxEw9fg6FOkiSKZurYSunHrAhQuMjklqhpuD0Q6AY8grsNtu21/0Yh
Tz8N/teu7056BdTFjFYSqQ2iKTilRkoAuJMYJSB3FE/IqWO7w2Edbx7vpTYgk1ncyJtrLbnrMNG7
f3RquOj+Xi9Dz78cwxxH87lECmmangpX+FfpRXsCF8756Fpp3l1Ap5063Mb0gnc89S4YX4g/n6Wo
Kw+NDCwnns4phXucrQgnubECzsFAbomYsLl4mNVIQ1f18D0IBuN/UJdzLh4G4736wws6bxiL3L98
iKpJelnME0Ef3/1Wo6k0B0ZgD2lMWfJyVBBkdsh1Dn64nLvst/Udy6T4mJHmMVZbN/bqulLTge1M
iDZJWgXydI2i9SW/r1nr21FcpmRJWMMpX980Vcqu9gykckz+WwnqIeuUMxi432uAWysMl0q55+l0
kIjxoDuCVR3hWunXVd8ywmwooBNUK+q+cr4FnoWggRuxkWwyoI8ndCzUOc3yE+okqd1fWnRaVLp8
U4e5maPSwCOjwhXazTo2aQXdbg+RxB91dq8ZQoJHcz8eanJF+m0pPxLRpQPfIJPQGXFqNE4p5wrs
MJHjJYtIgLOIciJelNLQ/jaHgxOepBkvECfOZIxCnq7C9uFHmpr1o7mYq82V0k0LuIGTS6HBwJy4
5vrzuFhCkeVpt3ewGz+tDE7K/A28hMBpVPuU/0yAmGO4Al4lY3iXyLS5yzJFGHw/cK6rrw0AIN6m
I/3ZSqItdSkFnnFZEv3bPOC4YVCxgZW3nZdOmkov7atqMf2TSS9yKNfvMs8kxKh+0KGpio5QW9+b
G8tjF4Q/+YjYmZ+t9iDCKPEiJdzaJ3RoA4soFoTJup1Bw2nUjzzRoQemOdXR2x8ksPeIqZUrLhbg
wC9GzwaRh7AdrxYIIJPVHO3eAoXAFLz8Au3bqZr0HTvtNqMirBZTaOob9a6Ur2LNrbkrPM0c7/da
umd88cWmxVgyCEkEh0RSjbE235BQnfBUR6A0cr+BCfNsBBkKXdcAGQkSml1qF37k78v92FfJqGz6
RLZoAIhQVjXbw7pWoQxLp52wEVGM7qKs41t8xXMF5FukhX1RtWxCL13we/LyFpGzgF9NZVTHc3e8
KxCn485j++SX7by1JKecWHMJg+uaeADmDSvxXqT0BzYhnPMGkdgoOuvpKUtfTN3Nz7sZG+ir6Pg2
aWVP2LRwv5IcNmieTAH1OWIAW7dSKfTEcV8pw7mk7KoYYBCdXNH6zXKT81ljhxcrN0TrJBycPP8t
z2aG2GqXWMsQ3iWCfrpoo8DmGeILeSsRxgbzKMHPWl94QC3fk9SeYN+Mw6IfeR/OJnEGcOpKeIse
srknhqHGipuHxw54UWKqYWjMQVAtVv5MXhDeP/iMwzgL6xmZe7hK9K5mHiLNVIybMRdr92lGPsvh
jrSvp17KcOWzAb9OX8NaSo+EUHCd1/OZY/MKtonYi5QS+HdP7ndQ5sxM/AVyNAiAOAZPrCSTOp4q
9LD1jcb0cXK73oTbx9fpe+AhuC5vugJXphPVHrVwYWK9It5N1F8yqw0p8RWJ9i8ZUjiqL+i/UF55
VJO4NKDzzmjWN2jyqtf7drnUxRqwlBMnUuZUVpJi5WVo+RqaoRm9eYLhCI2k9A0fXQhEKu2ZEHWT
Aq5IqoJLEcs9qc2LDOGp4my6A14ooXnafHeZ9X6xMf/AYpiUi/IKUNSXwZXd+TYoEvES2OqEOm2F
bXqlVwkwHOS+C0H1pOQl6X2tSNhNIVQqx62nsTR9e7hAfzX1F6gjv0UziCIIRFF4iIfqY+4ALTp+
oc50mlrNNFGPCkhuRlxjQQCxAbsbH5wGxmtG1ecO0G0l7+krs4kiInsSMJwt26PDHX2U055+PwJy
QowoGIohL1ckIutSwsAisJXZchqfjJHSi6+gBzXd8FyV0e9nWoCF6wlQLB6WDTixIsJYG1qxCflH
bkE+IPkbv2byvRwKlFcnKu+U7LSvmLDC1BULfLTz4pElXu5gagmdQwFUr+2QmWEelAfMxVid7zox
03ZJ22CQBI7YHzsc9X+DnlnC6aPMZKborp+IbUbZ4G/AzcEZxdyhyD7ACr/ASTpApHD0NJwKkGB5
RaIKHg3OriV27rNi9fk73ewKIuKIs1rRIH4ldSArTvUCuSOK1Cp8igW559SF6V0xdv7WiDMLXCKZ
fmFmZvJaAZGQdJ/gyjqma7OCEGpJ26KxpKZomyVaF0aG1xTMEV5BuXCJ7jVFs7i2nBJL6AnPiJ25
HMvxoLdU51x0mSwGLDhF4A6sM3DUgxuONNjeckCrb+TTbfy5ZVVuDvWutazt2D5TNze0Wke1JWYk
HfqHgOAe5azQkEWGw0gZxULIuxXtln07pJbTk/MzwKoMR4J03scFTpCp7QP8dXVkjBu5ySJnuakk
M1LZVPKDOzb9tiCpkJgl3R/PwiwriFfEQYIDrAyZQhzt/5kpjpkNGttPJPWU6io+VI8lkFsZwjjT
0c+b7ZNeX+AfZCZM8rEqhvoGWhqxwtKs4tLsDuAoG279aAJXfUgjLBXpAKSwRDGR3TqdqvAMUcni
QiEHZcUSIApDecoj9TiNXYH6U6Ya1FwM0jfVyA/69sUekYpmPo3leSPzFCyoRxBfvB6ZWh+b/BFY
4SUhxBSSmSCaNIYJ+TriK2/zL3d1BH1S27VRH5HgixfFjsiV2v3VfXCpe3jZUIaQcOamQoaPv4ta
nBPqMBvUqrqIno8uv1tr+8uNaRf8v//YJ+EJtGr9ZDboTaqftyoozcSjJjY77QNmOt6cESlMrfYQ
IRp2fI+jPIs03PdFtGjmsS6bnWz3u3mhBQM1Iebgsl3i6S8lu8sfQlexfBVsUGFhwyj4nE6tpB7F
eehGbGQqy8TJOZmF7nFZ/cMQlyMBvHQwlLeRBC1Ot31GpRq7VTS4WSCk03GbF/xB9ymElMg3gVUq
uu9hVjVi0PmG4FlIPXaIdFZy6K5y3MgKzeTZBksOtdfyc9xyUDzwUXDF9DUMhVlp42eFZ79B0WU+
+K/xMo0y7KmBHSPIhhfdotDCk1LHmp1oxhTIHLj2kh9S8nQ/OCwiI11ObPJ1So60ETrj6gYrrZV7
V1v1/Ss2X/MNJ0y18ITlbhyalHA8W0KUzPaUlGbq59DnM2XyWiCcKKcmidOMe5tlAsTZi4H4iEQY
yvepDVoDRjTAVeal8brFQdSS4yWNUXH0mNNnOdWiGao9PkHEIhtUp4KRfLlleOstJo/cN/E7HOUw
zq578Z0rlH6ejA7EDR2wqwN5vku/4RC0TWXi+5w4FtnXdtO4fY3m+kZsRpuU0i8zcQwbQRZHmCko
azLhZHUrn7xy/xDwgAAW4gIAY9P/k2e0faxUTqBV59yfyj+pjLtNgCuHm/VNK4hRrTftq05jaiAZ
cwJsUxKS5bbbl/TFsKdrF0QTcqfvvkq39qrIhU0MwlwL05hJ1xkioolD+B6J/dxXwik/ooIm39O6
qoJf/MSOjjDXWBBSr3+O8OIHztwZf8d2wa1rCyBqYBZkOYVJ0N0Lyuar7D3d/cK47nLo0Y7Ym9rU
6br78f1r3icqLP9+aSRLDHw8TgTL6V48SG2FNZdLBtWfolm4+ra8iCinc1hfrXZpGJN5KBLg31T0
1KMmog6UAhL4xk4lEzs+lLHJozZo2UwAUDK0ec5mlI1xWPgse4mXphVlRaQt/62xfrEq2ZrQdmkf
0l+0rUHqO+P6ZTLMM0GnydhWqpjOw/H2C41Eu8MfakAx5/1cWfo++FCmqXM42+/2zfF3d+YntQP5
NbhWVNO5M0Bbi78qDrveduK/4F6uu5DwJNfnoTWZanfAOWjyAOncv5mAz/L9+u7yTZ/y2nwrjd/A
Y3TFi0kiNbSMDaDo2EgNnmSSS1XqPCFz/os4X8dRojr76NWkCwpPVR40QEnElyasPeh9DJQheteq
KG+SFO0QF1Mf9L4GP2fh9hML3PRfUklYrFnCE3IGzb/ufX6VWqE32cLBHmFFW7lT04O9yYgOPOsa
IMBEKShNU/Wiw36W24uo5PUAwH4m6WXW/Wg2e9F8NBb5dYkiIeELKtZMq2iNNTLPYDGyijleuKNX
7asnrpenIlQhC5KJxA1PGr1wJw95Rc4h/di7qxkJtMsaIL+Pr5rFsdRY6jTVnQ4CgndC/dtefyoL
Bb/Emp7YD9oZ+aXOn1A2LFk8oxqnuyaVVEviOkggEfEQyG7MWhWKeJBcoX17puZRwjxpSOtYMnKu
GULsdmuccBSvD0itPITygH4f+3HJt7UabMqYBNXgz0zpOCLwaz+dgchK0WnV1XMOkza8jCRMHuul
CEPJEtXw0PnrQRkuHTZqGY3ktZCQIWUpXzv7QAHeK8gjxp+VX9ofcNJ7bP7mK0r0GxcwhcsPsB2T
nqNy2AcOMwm1S3B373DGM/5BjX6cHCvMqHAe2m76wUUxpJ/EjVk55KPPePJbNf37nw/2iJQSgemK
drZc/XaqBblVttjici7kdhznb0SEsJViopS5pAxDv10ZX54KSOEiFghmYJWnsjTKuhRMyvNcLy1J
iK5lodenIom7VTRZslhUyrkz57hwi+Epqd8c9SPVBUsHpiNcGZdsGQ1R/rxMpwYhIhGpRxerAsLD
XbgiZ+zLyOtV8bDsSIFAoGpfOJWTOw1mVO5tIVc8JJ1qjA2bcfzoBvLd44BdGCYYC8gHWhidXfGg
0KmpiwAQ/smrRXapjVDtgXft4M2H8mQlOr7T2F5d718tkj9rhOWDr1pDY0dSM+JsKXxeWnK9jicT
mhFunOt4eUEDHTaPy19FsKhRO+yINN36g5j1N/kPlmkpXGqDyLmnH/X2OIQzgDSxDYq37q3zff8w
ChosMF3jZ2mw9WhYPilwSphRHoXABLoqOpAdPQX8tVoPnCvlKCBU/DL4MS+DqkE534cP18UbL2Q6
sPaKMAQmU82tnCCDjJgHrvZReWXvQR00e9UfckSNrnEQ/8mfhedV0Eo/4iNMSfOYl+IBTbbP3xkt
aqo1wZIMF8b+yAhdn9t8znytLMqzUBGuHUfaWQar2QyoGYn5UPAuFU/dM68kyNqpkEqJtR0tGt5q
ZqAhYntsSL2j87npoA1jDQ6QFiygYylerhtDVHSjxq0aFA2kv0CMOHZ2w2pzZIWcY68UQgqn3tKN
HXNkY3PWq4CJrpo024w6gWQ7IsoB8QZp1Gnv78Y1PiwCZgF+1voFoS7sRAHjyRbLAqLUS63u8El8
/0Q8tDa1b+JQrsjE6BY6gVSt9KJkwws5oq+DyJzdF4nWH60VzgntzfyTohwKe4dDtqy+yiv3gVlW
JiTqNlQi8RguGE92jScK+LsV/C1GS3QTfZMYSi3lHDQpHymVrlG+7BDuUFLPrHS0JP2/bXe4rnb4
HNIONRw6bFrrtCBrhAZva18prUfdUKbOsPYn71GjR7sR1qUcMs2edE5jlu/TpLgIbIYSqRBdT3gM
PB4f4KMuFEOXS8SC3w5AE1dWTNPShfdnLBXPcNJztY+iR6mlKGtHQxXOM5oQ+oMXErKN/t5agStA
QTM7XcGzFxEOgqy3H3CNJOuIPkFatudAvvAAvWfoOWEyYq8R1X++91xHTbZQQpNFHeZ1dj4RYbOG
Ryrroc41xjjJJK4pbweGXuNtSmaUt4qkqf+emTsK0HNPeQsB8JN8uyseBp3sL9B4xVPYHX1R8UuR
ee9MFLtagkIF3ow1g5DYuD++AOL8l0+LIRyR33bBJ/YtyF43zndG2a+Q8hp2FXTbYGKQPdd1GLRu
rq94IqKD8wRl47i8Xugv03k34biQVzUNXzlYo0gYEL2xhQZfEb88XcTQHISm6i3jvGS0BDTrt5Uf
gYB3hRvItYPuu+wjoStdq4Hf7loaY9yQtAwQyjxoUxw9e30xsPv3Qtf7ScdPiCMhiL2u7lSB2d3o
HG087pUlSpBFHk/8FJhLdqFQulxbc8FBCLR/No+Mvm5VsZy3ktPXO1vAqbaAnz6gVr0QmHiM6qkL
XZ8rMvbVH5ZdprMelAAFo1RH9K/iqNP8DqwCxuAL5x/ZyhU151Uio5/WP3M7Da1hsRc3plqEZMb3
BQgXn19hk0tzJ7432OdCcMfNHYNTuNMoRKMsoEfUmoD5rn2YM3FJNGznNFeqmzDIdSIRIPvQgizd
2+qPd5wLPm7UdWLswX0FEd1sOYXuSnMFpuLboEOh0SDPKk0cncUCmf24dV7s7cMa0v5F5VbxjMcU
1Ua0BtHOy2/FnP8o0fFRQZz5XYNYjrM0VRmEq75tEnN+lU/tx3QVNOut9NryGtJJpNNfky/T8JX0
zhwoagF3AAL/W8o++XNbbAHrUDd2QUX8hJRDwykyTUz9BdV8smX3zvR3vFAAaHVe7wn7zHs0OyvH
yRlOictBhT70mIJQQOcbWFt5CQtuXzuNVSQSZvjw2hXojG6jG7mDdV4EC9FlsbUUmizlCAxKRgNp
3SbRP7z8O/5WTmTbdnFLSHh4N6pgfimTjGDlcRKB1XfQ24Pon8bjXz+ZeKuTwOXJOsW6oMgMkWJz
tvXwkWdh5oNYoWx357y3whcXMH4kegnnMNqrOQV8/Y7SvFkDvu4h8i145DQbt4BDDgiNS80SE0UG
UFkILJfQ7pR4fyw3xodQFXWFUDNl5+xXYIurPUETqKlAjKG9AgLOU5yHhNZ3qtXInY+dpbYPKqRq
VdI2OFF6LoPEel8v/99+cv1EOEr4j7lMvDc2QbFjpVsEPet9b1znNmLMY+P7vjrFux50+2ltUMN1
rXNn+9BQysLjOChhb04kjRgkPYm7LAIoDixV4QXCUWnyzome+6dG60+yEYCCNgVc4ssam9k+L1Nu
hpjpSkWji7Tn2PPNJbkkKhwqWZqKV1vFDWTOmdc4lef6zSHrWIxi0OyWWJr0dz6IOaePdew0MHGf
oWVUx7dM1OGP8ukN3rTwGHjVMz3sFaq0FNPbOieKhq1w+7n4/qtECKsTaXN3JUBCZiAzBFX9eBR5
9Z/o0JNcCv4n0YdOEblJ8h5rBovgHyBqfulw3MNPUQ5BA0tniPSRTphbcNz2weW77R8beZME5LHi
a8HXy/PfNFGP8JgopJsYDwZ2n6bi179r/WcaPuW4KNwUSNwFSPDEJTYSsGjcvqvxo/RVJAb2EG6h
vr/3XCxmnEehZ/mIrKFxnhqFAoeIkPpUV67HuI5BLA9tPdHfkf3uXs0n0PyVqVyVSpl+bl8Mpmi/
P3rHG7AmkLBOPVbTAWH8ukzA9ZdSzVKpsXTfuAVjI0pFuBw8DLAuIG/VTkOBiiziwxEFsP5J9enh
E5fmoVHSO8SiGPHYWYEWYGQV9mj4rsmbqzTzrtJRK8NBAWXUx6KxUGBqDWYYw6YXbUGytka1E0kM
kkwJh5SoSwCIyRSSmO6Vrpzxn6WPdD5B95v0ztdm8cHFoDLHqEDBCE8RAtoDShM4TBrXgpWDL6o6
HK2E7PpZXAQCQaQDkuWFCdFK8esv9LZd+q1ntgarNSF8uG3/rznpw+AK4P9WMjhjt05ma5b4lzng
TYR6MdxYECkH6+RwK7ZyAm9tGBJ1nLiEW9T7m06QAkS2RLxdWFPEcTHleH9Jpk0vYn+fM1Uw5U6d
5Ktumj7BPcl0Qv/T28ZkdaA1aMJAqMFku9iye4cqOIoPKJAGFatNfyjlvAhcQb3Bz18e5w5Sn0ik
sOc+BPZNQCwG/PMkwZeXFvNfuLeJR/L1LcVpr5c0VEejgIpdnKd0QJ3qqV5W0Ijt5q0H0/otZEIr
dON2L928dbnlI4Gn8i8aWXcurv2ET1IH0prHYVtzeGex4hSWIGI+0u3CzUinnMXoZ5ZoPul42VlD
2CNqA7M1s21/VvDwomn9S711KRbmVJzg8EeI+FUp1chiZj76lrCGPTIzJnQ36k72VyuSqKwaaY32
JlCPWRw/AWuQ+UpCMK7aGNvXqmC7JUuk29hlWlVKSuCy7HyJ89XXVmvwyePbh4m2ek8/yCSX21WB
Ap/h1KOK+NFfinkPQKNc/MRfwj+XRUxYpy3HbjnOLyvYFAR6pqb7iNbQKZnMxl3PSun0LyZTABev
rDOQN0OKm1ACMAmjNDrVO++uaJB+t+tykS+DwIKBZnBdav/QgE/93tEA3niMCPL3qBqBOIkp+g6S
1L2s/dnXdst0dfA0WnhnQeDDrk9lwGRGGEWPqb+9qBsUUBP9VrfnwPY2USiOltF/G7Lv41zn6F3q
r76L9H3+eBRdDFRfFJybO/d0O49aMze4VyTS8AwuwNPtM3OVjMV3bRrp96JWKiy+hHOrd+jeTdrg
4Z0gYUMKAM3Yxcu4CH6uwKc2VfguAUNYUgR/9SasNlh+Ti4ez26kGoj9oVPnIxe+vOXMIds54lfy
TGV4LjhtRMOm7fqalavXih6fA+PT7g8gZDrV0lLvcU+Ar0gjPkuPFMCbV+cWclkWPDb1GfMibhyl
Y2VLSFSpvZB2OwHk3gs3V6Vnef16deQZLKOIMgy9HBouN3gEmmx8g1+5WrNDdwMGPYSZZpd3qTH4
bDRrFCm394jaCgrPDsodN/9FCMUCs62utK6dMc3kI+4xoDx8g5VxoHob0yGbqb5YHH8ldWwHGWnb
IrbfvlQD4CoZb3hap6FvxabLvCsi0sCuIIpSi4qOkYThGXDRPsmHXUHf2Qm2TTAk3eOrDkVQcimn
xB+oMs3D+TlPUdwJeOYdeljZspbMgYgfPMCzjATkCtfi8Smk6tccc+QM7hkCS/ggusUHTm9l28Cv
M35LQPIffq2eloipYCyLr2jxAoKnc0ICFCvGsQsfl4g5OFldpVF4i6k1ayor/b3nFO/wDmHRgMgb
SUsnasCrXUE9YyunlHVk2UsbM05gT25l0p+Xs9KACv2+mJGKUZMdYo13SyQzc1RrhMDxQcJNT6fX
8QqEftSeE/XXGgpm9dAonb4c+h7THsNLRWfGDiuuExYMD0oSgRoLmN14A2RpWo0Ky1a/6r3+0ZDw
3anF8OChsvsaPEl8iQj2aOPBgh3VSZbk6QMG4K2ptLwQXjCD7NWFUqIHEui8ozGJAsl1Qjn+18dQ
lcU19+SAnJv3Cedz6aYFvxDqarPJREsq5mfm16zuRZOE67LQpmESPYEFigpehJyIDgOz+inkoNO2
5z7h8lnWs1CjpvfVzICXDfVy72pQhHLcwzsIEeHgqD08f0Rpm3SHjX/xuttOjdTNKhMpuJJSGXYL
vx4+DyNFwn2joGJjToqHXnSh9KdjogRpksBJmnztKXztsSL2cXtRCA5eWGwNtU61HkV1aPNMD4E6
nFy8/YVvyoMOqJtOcV/sXqEt3umyVblbzpryTDzCtV6BeAsqr+BFMA/16Y3ZAKw416XuESYRm46f
EmAsRakyJgdrTa7kuhoNpex7xnuGqyErGzkoHKX7PSoK6T0bY6AiSd93BD5fbHEHtNz65Slg2B7Z
OkjwB2JylFGmaFDXXl8ebOlYJGaD6gJA1Z2Sg+TbIRL4Xj0C5yQDF9YpnNp2zNs2rvA3nUaot0rs
ucTt/hK9Mz84o41vWEF7NPUDZp3xKla844HAzSzhO5LIRonLOjlQ5fmOlbEWtCZY3R5qFil2bIpm
xEMsky7Puu7/kr4687JYB3nxsGxc9jxQ4Jln/52z4uQ3S0L/PiGEJ0xQbOerz7mNCwjczjo7SsCv
eyw4f1k/pvs0IdNvkUusnJwVeeQWOsAV7It9zjwLu0L/WCxrAGRRlgsG3KCaJXblTVVwIPPK5DK7
dhIem6Kf7rp47Qk5p2rKLJpuHyo0mEPJB9aM2ezXTdj3hwpmB6iXTehAv1/LG4wHC4WmlLE2zdtB
kTIpG16bQHgWXbtXWxN+Azo1QczBn81pT/YSfzgyAQjG/ze+VsHz8mf2gj8dBnJZDYXJQsHGxw1k
cC5RpkYJT/HgMZFSznFTM4/0qa9MOa9axYFlLKAjEhC710CfoV2jyddYscZdl+7HcuMa9K/Nn50B
pN8Da4v2AmJ/SLAQ4bPtsFm61WiUQ8s7Jg8+BQ+5xaWbSD/7Cs+RWASqhPHU0Qvz18eUoby5z3yx
LGo/S+e41VWECZuKr9wrwMw+eQb88f0+VMipItf6vuVRgQ8yiHZddiRebSRaGLel2kcCi8HgAWBd
07KFo1qo6umsjdtExBPyedglGV88yZ6YQfcxErw9ikmt9l8Y3ppexgFAYR1+809PsBNmKd+VCd23
Zo8Lh5Qneqrcgij9bcQKtPnZqZeybWk+hXxUgjorKzWsnvgpSPWAmddJgWvZc7H6eYVd8M+Co5FP
htnF969UYhF3aSGzXyyPUnP3g/E1yXHVbdXiNXnwXGzhBbGQkKsc4VvRGzfKHz33WrZpdYflhAbj
RR0laOA2ngP6CY6j904s3MLX6/JLmo2M8zoFKyKOZucGOKIWTdj53+jf6OVLQN65SwDmG3xpk6PL
ClUiXpXGaH8rKl5PistRprVGB1wNt+rPQq73F1cxbQ2YssMznaw3PP+Qay69/yejme2/7bOezZf1
yagacsVaGEHFTA9iFqrHkt2ioyVOKHtgjVIlurZjee45SiwI2OAaKaCOeToRZSwOXSgEHVspeoGF
LdySDR7hWnVSxRsbnKAfv6NT4A7U1rThtXdKHJTZRfcTsggVhSfeeM9ECkH2CyShaB/7AFzBuyHA
k0jg5yoU48BmTAsHuttdYmykMGulvUYm7DndA8AysnQRAVwYV5UHwL4S6kA0jgXg8/d7HWclaz+v
LzbWZPT8JV5od5tdkr+nIZsqcTsOlP9V4ue5djZJplTOUY6nWxW+Hmmth7kDQLWQ2dF6CnyVQEHF
ViTg7ClyTVcLDDfRmDqUWf3WDPF3BUlNgqRQPC/2t85pBCvAzsYCe0BRuVvqJzE3hKFHz+wy/57Y
qe+1/BubhQyQMnR+NQIEHnxkC/aFs1YVPOFEVj1SvEyi8cADys/O2WaNYT71KsvYOih6m15hnOa6
m8oh0lnpryXANwWzKy1ka0JDuKmYfGBAkRnaNrjCYfh+g8VPbyIdP1R3KTsUmfeFfWDaN4ek2yBM
Q20F3HKucbWu0gXbiESqmOavmrNwtFESumImIi0HTZNs/5xttow2yI6NFyH0AhXVrKyaPONkbE7E
/Ugy16zQ8EhOUSj1J4vDf+bvIyE1wPlxj6SkNXO8UP8B5vNefXkcNqD2VvP7baFDAAXiATCLCTPO
gdRJF70P/4oPli6O0/bpFNrZGBUwSQSewDh9hGnG5jiEiqSmL7HKR7r0nobjnfJW8gx21Ph4016u
L6kSj59MVtUBwhCP1qUBufokyg0X9SQ6npGp10e31zW6KYWyFK1UfWaOAD/HT2Ir+k7tPqcFokJB
emxHSwpDRdKJVhvWM0tVgKKfx2AWJOnuWZ/u+NAopB7okQErJOh2S+VzLD/F3u3Z/n6MsEPphQOi
gvFsvFiMmjqqR4BY4pxBuLSEJSbtLFQY8cljusEt3tx7Bh7X1b7qFxZ++8pDHTQxDjs5KhLGIU1i
vdeivW5o2HzDGSdUsKwrJHv2X2cNYYcVXWB1h3DUFlkykqXLu/YpvYkJBM034opeQJyUwsaYg2ve
lnC/19yNEk3bulU6kaVBOF6LlPXza6JUi7ethWnhqR/X6/Vu+n+hw4Eda52zc2V1G8IqqLtk1lk1
tgPfsMfi3V2z7Adl3DKoIgIhhihJVLnBeKkS/y/uGY8/V4py+B9NhiqrFN6QOMxZmI/jCXjAOorY
1PzpnOEEzuJpb02FBktf4eCYax8m6o2ELadCutHTKzbeKvYDdRFskjvdZRBdu7wvgQVWBrKoJsmz
XEe0G4dIuS0pSRqOrahyaFp4zNZUTE995Lae8HERrGPchDB2FzizjolM+A2i8GBGmWVju5cgv935
y1BlQsZpDWuXn5vyemY0nTC5Sh3CXmIquMZpCOOPIbYUTmg1Qb2NIAtCnx71HEodUuBh9EFLMhEG
/iyJGrA+s7GaSjkL0NusigDAGz6+tSvCl+8x7nmVvM9+qvpQJjYVHlXoJeH0bit20ppvNk43swDo
NkW27GxkNGDSHJzepogsQmFmQGpDfioTUIOZyp5Aolc3GPfE/cbTckf3JSQal8pwPtwBwg7U7DoX
1xfsLFUabqGqKkj12QSEDhVeufR9I6Rv0Yiw2sxUEphIrC9yGc3XD2Y/A6V/D5VRCmqizhn6Voeh
xcnwwU1/BgUaucKy9tthmJZuQBrnRqQ4mpDOaxm5MCJfgyGmlLVgUqsqxFNeZCtN5fGvqCE/S0tg
y8waB6hZoVLewtTQ5p03iP/5m8TgDRy+MajHIy6c/LBJIukLgHGYbnwPzqetEwvV8FFDGm0qzxT1
4Si62E6Z79/nnhUT3whjL4B6MwZAil1ujwWlkinvIvQBdyOVjGv8gZeY25VlHtdIGNJZ7T8dmztZ
Q8mDSYO5NsIprBeaqyj1CwWph7XRz3PkS+cD37+VCHNKaeoM38RQC7+qSZAX35NgrfBljCAWIiYk
I0jhYRxmrbAzry9K0CxtiYU1OHtWlfIDxqqr6xSLdIHBH08vxikFR+qR4wo5ssIhqHZ+BOK3SSRU
JBKYBQp0nUVuLsTLuydxQ8rZKhLL/6dvyfJYCulNc3ERZ1SVEmLn+JE7+V7B+Wri2iKRNm4JtnJ/
p3kplJMHvwQ/AeqSBZ87f4/PHF/mbUiT0B9iHjvPQVOvU1XWW//NhLaYjxrveQf2IR1Q0PTNrw0F
0m4qOStJl0Lh47/0TSF9o0ZSxY7TCzFv7nhGOUoJ6gN+vVbbvnFYCQ==
`protect end_protected
