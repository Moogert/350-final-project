-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NZlSwQ9AKMOzctcj2vHhckQfhZlovJwgyiHskOUkati7Lv8RqNV3J7yn4kyjFf9BtRdacgOwoU04
EKrZM6iSfiGf/yGNhv/KGA7SWikGMD0Z2eJGJ8sCSFVfHY9KAy3RxQi/b20L+5EXGFC889w1+QqG
WRa78zDGpAX7EuPaeTVLPimzHDbuKB96CUeaHzj0dmrBqXrEsfSIk03Fo9gDnwHgeeSZd0o6NVMJ
YAW7YpDpo57ssZYm20gecrDXbRtPif9lOoRgt6O8Y1hg2OwIMAcZ0TkBK8c2fsC/zPIyBMiVvNvq
/4E91QhLyGqqWcG1CYKi3V0EShpCpgduwRVrGg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
hkWLNGLmSupcQ3kOfqT8sokh95jCnmFGoFaA+rlAcbaxnvQnZbq+AZAbLwVH0v8KmrfgaM168aa0
XHkONYfevb5v1zN4nmJy+SMjtc5HvjfEd/Nnmex//6dY+xDNu/VKI+8EFu/c4NmykVyIpU/Cbl0P
i7rZbxCkLSUGHnrT1fqNfZ3iP3ZpJDHCRWGjxfyNB2zqCFF4B+OAtkDTmz+YjZP2wDe/AWXJ7J0n
usOx9ycV80nqfPi2aVeD/OPyMw0Tvql0N08EQ66GF6TDvgHNmYA2cmnm4+CE5fG7sZj13tVQ5Ixn
2igXFcFcUhvBNeIk16dL0wau4VIVu0Hdamucd+aW515HNsSRcjCdNqbwmCzigSYLjFJMrUSIehYr
+SiObzagGNwJ457B7ZEgft3XjD01acLiW2FdSBN+18PQLW6E2T/dCRl3oCyKWAYrMPpowg8DpdwP
48MNiySs7MlOtME89b8qLu1snRdpiTBRS7TsZ4ft4A/2D2mZmIENRMmlvk97ot405Dt7XGd/zegw
TckSLUsvjMsY4rYGO5TXk0bldH0PL2WNO7TdlwtBWbNvQLHpcXR1wRDh5siNzBqzTNieFSUNTCtQ
UT1Yb8dm7Iz7NfzM7CNIHhQwodv198Ma497Y590QHC1LkSRb2soB2I5i25MFA0VZEFvGWrdD2bxb
8K+jmg7ELrxR8/iPQso+9XrGnYlfNV34T/lDxnncMdoCLmCee7pqfqQbHd5bEQijrdXyrLF+pQkx
Klp/vDsRtZkGXCjhG7vDpder5VDQBx/uhhQF3tv2CwBMS6S1bm4ByR//EeuGNSnlAJ1Q10fvxJmf
3zlmeIC1xl5A6iK9h88CGopGtfC+PUWW36xYjzJgD568I+ymF+v+uoZaISMRVLXtZMW1aPxsevxV
ACUlnlVxZNBld9hz5acjwYaqIoH54U9DD/hnY3LhKGKhYMNgQsvHk99fBf2p5XG3iyIdZbjUfuNh
dlCwJYgZ2ghgsJNSbWzHHK8TINaIwIpOr2PELrYtGtMDWO5ev/Y9LonQfz6ZotdlqL0/OPehu8gS
J3ELybE4dDUMyz34/qW5cAh09zvvhFjVDXdH3fPXllP90a2Bdm4aGYoAjmYkeWHC0H2c4X/mOzWU
19K7g7MvK7fXMruaQt4Bni/y8V2jKZNckp3XlvmLxKjVPhkkm6xI6UFi5Xl5eE8p1s90iIg0gWOE
ex+Kd7PQ2RKt6mrNnr3Q/ZkdLWXDBRxhsIjXzw29Kpcp9VwcLhGEyzN5hpSb2+4DCixgEGbaosx7
xO9oYlfOtcj+1WCf+p7stmSEdw4uyCpoadsln0GdrfZw1TIF8+CTCyxuuzzSqQz8Ot4Kp6CgbUTE
ZrOHBqgDXrOTw/CxGBPjERUIcJ2jjQRqHd+XbdYNGCaQE3KzHE+lBDDetkBjUs3ttb/AYtIam2ta
C7ZiHu3U23soHJqVK6ZsL+54m6uC0ipmyZtGvIyogC2TmYjdfRwvHiouoxFmaPqxsdMozQbAF7Wp
+HPyij7WQeLH1l7qCC6H9AvNrp0QUIuvmWBuSCegI1lr77VVnBCtw2t8yXSVVdPq9jInPc5A4A6Q
VqGD/VDMQLdAOpBn5mJP6skNnYllOAHhXut8UAcGat8j1DSggb08Ggr3O/t9KJFOkAS8Ws/2E9NP
QlaGzHm3ofUvxDv4Ct0I/QjvaVphrOYdwt7Ib6VL+hwAbhbl4cRFRMPa4Tr2K1HNaNpSf3hu7fav
kM33NfVxrDIOhHlsubsea9lqMZKqjTVIw3qIhojrstOKjUAfTvEq1LuGhDsePhghIoGFWbjdvNnS
bXlfL7yLb2Jjte590jTSPlmw8KGonN+FgL3e3+PxS15r6LLFj8rEA9yRaZZPACCF6pT/Y9boFJwd
jhebigdBxlBG0hcQMgk1AWpwp3J2b4WXlamUEzCuIOARINwJQzvhQ2xVyHlvK4AAJyNA+TMoWzZo
X3F7bjHGRuJilrD9u2nEvZscJJXWD/EDJ/Y+MMQ3C7NkZ61d/duiuAdwZl9Ok1J43/TwDEU9vRmj
yMYM3B0kI8dk27LzjdC+sS3AT+Pk5yg+K28Mf9AcsDsjP0OIptfr/KJn5+JCjCmgDBGaVyP6raAy
e2pHc3lDaJCNl1v97jM9H2Qt2doF5pT4R1gxusmhYHcZgYrx7WnHa1K0WMT2e6DttBjXSdbyP1jW
MkxHkLJi7/gr1Hm2CbZ5mF9bfaDvnoBt/dEwKQEV5qp5D2we0mGsONQdJ0mp0rIOXDzlfWOwt+z2
mSGV9uFC+MP9KZEm0VaS6F6Y9Y8E0n5bDhsbwEqS65c3lqYEWLubcZRdaLooJGMkZkf0HETDz4e0
LHM/3+fkxbAUBOB2dFgN6F+jh5XTWe3ZmX48EjgtFLakXwb625HWlnCLi4MtYpp0JAZT40hLgTOb
Ls9FRpyOY3nQmcbXceaSc5fZv3QD6e4nzK1CmnW+VJlQBWxN76O+Q+KRFdnUmu8j6zb6v5tdJUx4
GBJnKfUnk5cArC2N8YYbbjTyNh1aU4+brmeQr2BDU/oblIB8oJ2GImJ6WBXy+ZiQMO+IQMUzkCzR
Udy+wLjAKPepAkI4g7rqYx/pWKIQ5KZ1BPXDZWoq8q4OjBgUWOSU4BXisOfB4YPWUuJIqoKCiT+5
XPhrSLHbKkSdvyR9VUbiqE8dqJHHE1Oag79aWJYeJzxiegrYs00++h3o6/id+m+I0/Kg+TcT/gLl
wMaROpOxh+fPOTrt27+mHQ2IfyCKv4mXdMkQ4EzuYLgfw+VJtl8zgNmIv33cfTQ1D42LWkHbYVMb
hreip6QW98LqcE4az4BY0oEDiTilbpUb6SofOQDQqPGUEajxpWfqACQFp3sZfe5KgWtd67T0vxLh
RJM0hI5obqnyDJFLT10ZxuWWfnqCmJnhy0kYifuAwFxe4gfnv4eZ+3B8r+rx3p3v5cSC3UwMFEoZ
k/Ef76ltTwf6/JHSQUKKiy9pUBkqZGWwK3V9xKl9kC1UCqGWdraQP+vFSiP1xMTi8pgwoYl74gbr
wagR8/nD3GfWU00QPYiQAPkYvGtyI+R5q/fGONSbtrJniUtOH7nZQN2mbSULuY60fvE3pt1RaWdT
vK7XuohJ5QVgdu1xZcg4za3xk5sZ8znt4Q03+6QBib1Aj1DWQzSASSigySmiSQUmh5ebApLvnJ/c
bd9LgOVz6S9KR6l6qf8FlBUqdI94la+3Z65NAmvQAtb1Z+Aa+2VxvY75o8jH3ofrUxCKTZ51OXPK
PivrZCPbErDUKC6w4idS1Q1QCJQpc3JV5uVn9L4EPYucSZKffGarDYm5NJj6WZyXZPXarC7zWc7i
afst+azoymkwKc3/OPHDU2kJ7BZyjWICVhrBvZrNXKRoCeuERKunDshgTDz5O0IqAooedFj06p1r
01pT0HjPOkSD4qs1LWGP2ju6y6R1JzsL2GqEKWhOq0lhR2RoiQaG7j1r2OMf9c791V7zNDjAg19U
q49RW/u5DlhTPl6mGk2n2G985CC9L6PQp+N9nPtXtdrVkIAw0zDGeQKKCKuWir/WqwiMr4d1AA+w
aUHfSVn06QB4THsGdsRQHn4KKL2N3ZgxZGZF0mN08DFtCg5kLS7W7RZB7KIDlRSDg58tAqsPsgXx
qVqk+FExnQs/kwH2wl1pMvY5zyhhNrTtmPHEABRcE2X2BiYJCyP6b3YWwbZLA4ht+HMcxBmr74Ke
00SU7KU2BtSovY7dE6VGbGlk5b5P3BgoZqbkLHOM5eX4dFAY902SVdx1us9nQ8Xh8rg2D/1i7V5b
GgfjGDE1GXdyMmVr57CyBz90s6Pwf3SmnQCS1+9poEz9Sad22UaMTHoE7/cPxOZwLOe9UkAb1OqC
nPox10/3UiER/o8o+7w2bLof5VnG6BroISj1XUlOGJ+FYbT0A3meqUP0JvUaqWpeK3+3wVQXMMBE
vPJjDJkIjfzJ0rK1IQhuDqBemR4tS2Jm4mMCmue3e4ZSZ+LGd7eeWu+omC1JJ4o6tMnjgJt6NYyh
BlRheZNBO9YWeb3ELBLSiycryxKHNS3SwusvG699tkCa2ZZCxlAhFJmveN4MB/WnZNuNdQ5RuWrQ
xxP8I98UlTGvxWpP397D434QJAHmpWfU2i3sGpbWSj09moCoutcd4dYBlaTuHEy0dkhQ8sf2KncM
MaUOCbrB/YISkV3ANMAozI+aT9UcyFADHjDt+OMzqRzKmoTN/94MwyIXLk8m/hpLk1NDhBzDhkez
Os0qzK9hs5A6n9yaWeouYCIj0EJToEG4LJeQumuP73Ckh8pIHY20/GaqyBBfXPbKeUtPCgv5Plpg
oMfuUhk+OPrhG7YzcYl50b38/dDrgerbU1iANI0ppDkxq22wY0YJkEBnf6BGmAxGx2QJ//xgqNBG
tDSyiqOmviBQUcJgEHSlKiHRpKR9cwl3KVtc4R5SPp26YNo9ma5zNBIFWA+9kei5M470Mg8/J3E1
WUNE4kL1sx/o3Udphl+RnvYH4sTjKR6zB43q/DxpHV+ZDoQxRuJYnCpX9ZcKLSF3zV7UBzwUBqFm
nf48xr81rp86SWgLrC7GtnnPSvZe/rwUNfT9Iq47+17DBxTNeQ++fiELTRfgTzzYgagn8xghrD4u
aK7wrsNnSk1vlp+MafTA/DQ9V7Yf8JfgRWHINfkuv7Az7XOHgMRPIUi+91CgE5nCQUH4wW6oZtwN
whJj3l6Xz5IttNzNEO5fRY7G0xAseA1cQjbbdYJE8Szs794/s7pGiwJ2kw4zVMIRzxEicQedkr7e
fgrbJ76cshO9/HrsLZvslXA6zbhJ3mxRx2xc5e3+6U7tcrlqbdQcsi/dZkJ2Tozz+dROUmyWUD9Q
1BQJk8Mb2Vv6CXunH9HKFRQZ1p+it9Vwa8FX+jPJ0s/EsfR0Q9vBINIn0atG+A/yo54eNKnVwhuZ
tZ81I9s9ozDLKhTIvS84uipOwm8u2Uaco/gQwJm2Mc6x+DWFvGHx8WsPl9e/y0GAaUstH5zKr3sb
lmfUtKgm+dGzhHYCvyD4qkLwvUSTen+VcVXZmXKkS0952wfaHMolCWbDuN2HO/EfuNmuTBmXfsYw
JSnH7l+Ebqqj+KDxgjNx6aY0CN04ehe+IEqWUmRic5K/2HCU+vE82BjhZKD0s32AiMXbvwdOM+Q1
+GHIP7KlUd1YzurSm8tMMA7oLbIR1ikzU5F7QSi1ubpHt8NXCl+dTO5+NKweazQktAU187YZYq2C
UzWcl7amnNCER2CxzTsDkB8svNJPZ/FykJ/9eNLafGlCPRlgC5gQv+pV3kw/A4IjV36tpmLvSlDO
sl87PG3A8r2+wLwaI0qMoEP7w8gANI72M0Pd2MoedJf6cKjfOTuKdErGyuk0iliAf6UbhX2UfBVB
fJTtUyxgfsEcthieM+HaeJWqvzvK1HRhYh5vNDRxDCoU+Y2fRQpiAiVo9aw3mF9l5Kybh3GReN0i
Gt8PZ+HnXXLkRUQr5hV63+cHHraKHa5TMwdrU8x2T/NSk9/wRN21d151zU+GCcrQ28xSJziTIkO1
SH6oVHTrVaACTiJr9m32yJGGZa7Xj0hhK6nYAUdV87u2xD9/UhIaA+5bv6jNGuWhOyyTyFwchRma
j4TrL0LgXYWlVonPVAGKpBwe6hZpQ5ioaoBOh/SpgsfqfvTRhqbyKewSjT1ol0/fk4sUCD7Furia
55+Le32JycJnPxDTxl+KTrCcdzlcl4C5NQAwC6ll8ntvmbTZIxa4/iAzl77f7/jOvniR8XskYtdY
S3/mFuzdk4AtBIlokqg2tbgM6h3f6EKu7kTqxltBKokTWUrNke2hlCeljyKRG0BkJzx0EnUB64H3
oxXPuNvVaBncqFRdb1JgTu6mBcgCACosJDR/jCK1nAKM48q3LGjom/xK5iT8JZWKUraLlzxMjwnZ
ExTiPTOZmQvlz6Vs7mFJ+11br2kFoTwKI/S0RoxyrRnNaFMVYBG1ZDgpN4NQENstEByEFLNFhVk1
HxmH9VQ5H3laPoLdp2Ng2yRg19XldMBFoLYHWkY/QAWa+7WfBE0mYvjuMPvZRZw5trf8rzcxyYIb
jOUKPvD+IRIzGOA2rPonrFc/wCCD8fL4dfVy3xZy1i1m60vrECocFIglVlfrnC9kKc0Nymj1PeiS
oPRhs/uIhq+/Ol4IkkWPtuQoBUUU+jhRvaye9I/WsGNBhHTw84C0YfS+A8A6TVhwqB4Q4cfTq6lu
tdOfVUKddj6eVIJ+6W/DBpJbq3BHhAbl8L2v5oSQ9q8PYzz/s+jfMSf4BMI9016MExaAsA+lbDLK
loIXY7B85UOQvjm/es3N+9VPzLfBYb9g5cDoNdHnXR6cXDs/x6UC3ejShiA7gIpfer8TlqtCar9h
/FSmZeinizt62gZpb6qv8w+87f1EbSW90lCjOGIgVBk6DO5An6j5ZkV1EyancR5CzHhAiRdZgO6h
It1Mo6IpfC1Kc5jfAoyKYeeh17LSxk1V0M+nAG0jqM94S+7MeVe9qsjMnXJYfD14ZrxpCWdYUkCb
tD1PZGNRJTs+4d9V/hCBdQWJvzhd2Vcju1DkG8ElymMmrIX2Yi43A6fyrWlfLGM4rs2XwjJ/Uu8j
pdHPTd8fr9V7jAEHUmyXTcVxg7Fnt0j2ISThFHxIGxoN4hvenmDYu11NyfpNvH52EB67UZjxU4dm
I75r/MzIKQJn7B5S0hh3AgKEUO+wiW6LLg2DsUbEVV6pkFrTfHt/aksLYWhqQCDbpDqK+Z1l+6FB
utwNWfL5CtHZws2zAxhXcathY5zyEJMRzSyO7qZZprUWHpokhqUVSNpQ1yxnslhP+wL30TuAwRgY
nMnvQzvMzAIDg0ya8LC1VjThjVmsrTlhKhmkK11ceLcUcDXzvaLRgXwTi5J+lvbLp/C+SM3U6CnX
r6i027ZUFq85bkX0DsxvZ3NkR+lNnPfSW30k3ak8ArkEQ5ht9veVPxZspNBrexZjr88aEaPmUFip
hZ2ioRk3Nydy5yfDWOc7rwIPdZgb3lnt2IR99pIKeF5E+dOrPGleHjUJfoRomZhfToYfD1jGmUQG
mGjhOBybzFeu/1Imm/rI/XftJt+gR0BWKRFqns6npwwlkkBNpeu08CEWE5FHbNybunHSXwjY8fME
yQudI8WDgGNlrlDvqv3Plr6GznovkZFcJnwdRzAhnakkUZgO2ozaHuMFirb0H8Kl2ZjwuVmfnaLI
AlJ0QMbflZuVEnp23XVTLpNQKnMtLu+oeTXh6fmhsjXEPjkUbScBEXXb6xZ6j1ajSHByEz+hJo5V
v1uNKEdyBuloBxip2Yncj9AlIAazrxVJYPUUoHOal++c6M4ilCiRg5Tc04lAPa2KvYkuGJnDU89t
hHRPMc8umJcPWA0G3iKybSLSlWkL6zuPsLh09feeNzcYapxf3da2Gf45VBP6eXnDrfQwEvosXIWr
R6nOQFr9PJ09LZXKlXiZZKNrgWipKHiTkDfyGo/szb30/YhEDUpoDz7sC3lYr839S8MV01Xqz7aW
P5CmCkDCKqmxERNwoGqsE/TUc3v45D0C92bJNA/PmTIa/2adeBs2T1NXMYr7tnDL6xovEl95m9Ls
z5Cj9fPRI3h4Vir35QRuUKxjPUOvETW2pxqPza9dysS2LLMTlzFpjo49DJXRgd053z1j3BkTxI93
Obr/SHdnkEK0nFCDMEeBxiZq0QePvshgbAA+Zk5p1gpjYoxCvU+GlR/2mUYGFyG1aCzMEV3DuNcg
aqcjB8Ws075w4HdmsqdreDFW0MuMzhKIROIdtQjp/L5EWnwiXv+OHTTYquvQImCjl5+7zQRmI2AM
i+dkZm2LaRzYYHJADtV8lYdeeLwm66wnnfoe+fitRCdk+qarDsk/yMBeQsAYmWZlyOQ18bylYL/M
StrRhO2mNxbbt7JJJKlPsAih86y/KiBhiyPImtbT6ik2e+UQIrTlz0eHbz5XKAo0ka2404yxGV6t
r9r9MzsishsShi3vun7TDw37gdpHdHe941xH/jSrsv9XYlJPmKRlzSOONui3T11leOMWEbfawhcJ
2UGt2Yy5DgsN9p46PotHajvT1qSW34ZbzQn5/82lhI0W3qDmGHFF4D52/reDcJE62rYh28Gh8yeK
1gkS6bIzQqpUzD33HgKCXQBQzAEkpzdRcwFc4qpNDGTaUCxmz+oRYuFF0Y/HLXP13i4WIXeBAQVj
zJnJ6Tr8bl3RINmgORyxjrfMabyoOW4oKPUKx0E0XBj+rDIlYoZm94XjowcccMGBDGJBK1j5f9Nc
a2ijPG3zv+Dp0FICDi0qNYJ3lrNXbBPQnnpjgXe6d9lEVD7a57GIZCj8/Zzxz21PgQXNjwqOM5u3
ODrp+UKhH0NREY4Ep1yOD/2/gqK1ienzeS7+aj+3zzWHv4y5eHtiXtGjgArcGiKDfadq97qsCRk2
npvtiVHzz1o55oTXvx2SeYOMjAnhy9rJWnZNGuXpXp69WNef3jM5sfbxAewKDVI6GkSVuATvL9af
QI3J6G4TCAMu3VlNtCQ+IWi4Y6aPIEdW0neMIVyKVnzRGm+Mtiz8ctwA/gD2Y4LOc/TCqDOYKg3i
GWz/bUhUwooKr5dmvHwn/hQ4Ihw+hzzYuGDrskM/vqwFPcZ31I51E9ZvdRPO7/DAmVZGFiQu3fql
nF8WRCf95g8f00jydnG2ux37O7WkIJC4Bzl0DaVvSreCQitFBcFctrqPGyN2vNGejkmUu1FEAKfm
M0VTsnG0PEWWvxoguijCVLKM0ITqlnBezKsSk4bvqnHD5gvIEtoNJUMMgNBcUitObIrT9S5kBms1
ulUBD7nXzQDg5+yLihVaIx0eF+Eu12JaPcY/heOcgg+dkiX0G1YirOs2yebxmJFLGyuEHc0HIlR1
BmwKNZxpcD6WmQtbxgzlAqlHaoVct3Sm8Uc+FsUQKhpjKAjk0Y6bQ2ETFEGw8GsQPB62VgtlytXE
5rTHRlEWxhJlq2yCmNqfMU5zjSRiTpB93JgoxHCKfWuXUFd+JjvvR0/NqFR2mAdyiNthmKZPHKEc
n+eKgadPM2PQYU42GV843ULvadwdO2NGEnnT+YgCbqRexyg+BA1+HXSlgcC2RsytQrT8KlLqdV7P
NS9Hr70kbhZMCXLKbNATEKy37oXcthygdy8zEu5rF51Dw/pCOu2Ek/4Dey1wLt3JrJq67H+zRBO8
WMmYaTMkMf4uwwc00XVZnBuZeOeV5Va5j9R5I22ZBfA3VGC5mOxaMFYrYly8Ry9/jkmG1CHyuGuF
FDief7QJCs/swj2NJf1mIVSX7iM3n5PPrmkisPiH5og3hxVyUZ25e0V9ctD2LLJ3zlmUvRXqsUIY
cT1msiSN1B1z/kEqaEeUs4Q4UMB4VVobcf0gDqm5vxYCSEvpAwrwIdRE7N3vvxRhznQvz6RqlCmG
3rkay6PJyza+scycOl9mhPo+sa5/JuZdwuPQXd6Pe3HAQCdF3R5c+XxThVnl4IraFuDEOMxsG+8x
ws+srhmc1RjnlMHjWF7lqbVHN8j/fOqszZBTg0PNsrXDCb1O1cgLBbxWdcdgmEsMZ5jrCYbtgsQy
lE7LBewFZqManl8qvE0/2wciYM7vo/7aEvoZNv9hLxIm8E+GBV+TpO3mlsfl+20g47+UGZF+p7mE
KeAnxiYqlhXtaigUZuB1CreowfP3iFr7WgaNR4S65YgACPPfWBJMWBmIzZWRnO8Y+gj18OBKdRgI
pVsWDYap/I3HwE+VsqIiFfUnJYNO3wDgOQeOXV5toayroieCF2e9t8Kce5yypkkHe0EX/4kznowH
Lh9+9dKFciGY/lt90D78+4YUwg/6ccQvGWCTSghIe+KVmanjvB/zLmYJy+UTVGiEHDVy4Q06X5+9
zcpjmCtwYVpilIjqmPdgSkSdWGNQmie7uDPQYpTEbQqTVYeq2yQyX4wVJ1EriyzR8Gu0EIdiB/Cs
tU+qw3+uEMgtQ3qeP3VP2Jh7wH4CbIWqF+UeXfD8t1eaMxNfrH87z7095TtWNy953HcOHru/UVAQ
HeCsqJYV8NsTdsS6TvYfsSmuGQ2hIHeQjsP69iRjnFFIhu6EuPicuWIitJv4ERKgK5D1ccyjicxK
3l6yL0m7BjupXM4WIAjuchh5AMKlySknfZi2ger/b0nINOabMKFFlaxo09zPSJiVBd5vcmZTieE5
HcEgi8lH3qdpTwmDDbahEH9jlsnPBexDE/gC1zQ3apq52BsDIE0ZI/8+z6ziwrZr9CUlWpW37myG
A6c96QTd761mcKljj11sj7yQf6k5tsj7FzpM8UlonnLy2msco/gF7FTYkRn69hIu0+7kZkNlNoq5
WGr8OZsYQCxLkFVUzLlRKwVo+Ow8eB/5F3FQ/H36OgjQUbw7isYBH3cWWnQLr2hFAiUauyvyWk/p
5CkpAWRBDRNpiNQ/MFWqEZbxK/Eo79oPOkRS6ZuKb/btqIo4qmor4yObJQRyPMAeOOP93hJwdthZ
rTkgMud+j3ooTC+I3y0LUcjCuyHM0tbbtjp6127jOK4gyKxWa4eJiEWo+WkVAzZ5UAA9PbQcCYZV
QOVJC/nldARIwqZhU/o/xqJ/kS48Teamh4eDliaP8O8NOXp5YExTSMN5JWq4jTSGydBfbmRfQo8X
v0FsZCcx/4YPwN9FPg6Zq4WoR6/avabXy657omR1UH4okIUUoPgLinCiSakprXKJTJEx9PxeQkHg
RG4v7/hXJF5X5j4lbZZLDJrhO+6cmLDDUZL2kIb4NJSFFcDlJwBoqno3XTsJ1Vg3D1bcfssL4LKw
RvCglcvSd+M8LLIe46q8V06F1UUh6vhU+NOw6egIOfO2bCiwwzcNim/5jEfeAeoHMfJ3cM2JHzou
DxzIQNSs5I+z9J3uO71FvQI7lzArwhVJwxdOjPAHkoDCll+wlKh/R0Ml5ffQkHDP5Jb4rw8a9UPs
OaObWmi6WdKJbG9HsD316Al7H0Lp4zg1uQQb9578u5CExXPiPjbOilPiGXHczqW8ngTpz4LZWgvg
QC5Cs50YuHLEbSP/GLKkcwb/5P1YYb+jDj5qTHeVVmT1LAj9/owJjhIHCNuEUMkg6sC4BO5M0E8c
0XLhqgtettml6zyfcJq1+Y8QlURe7w/RXWeGvKFERKniWQjZXiEc4i5bTWHl34u9qZzcj56zG9tK
OJUzKAh9W7xCjq6cGWUYBmcJplI05OvphwyiGoJITd3owSZ1+tqLnehygGDJJ5ExGXmkJgmuwOjW
sUbV/+cpJryNH+qY/G4RHGm+THBswAAfLT60ys0Vrq+undy1fkcP6Epl/clk6wAlafm29bvNJANo
On/KMZ0sY6iC8M4j4HmJoNtrllj3sbQDy04kdbEmc+5vv0tG6sdx1AqGBnmGX2otZaKCw3tGZ44n
eWgpXAc9MPJS/BAKq77+G1x+mssQMg3sVOsit1l+8jCGfg3pGLWBBky5UyfiuoCMnlvw/FQK7wsI
Lc9tJ/Ws47Q1pyJWC/faYYsVmjtwE3lKmmO1VNh+4saf0EyOxADJNcDiqNzd3HvgiJB2TmSP68s7
eFn7EB48U/anbchIxmlbwsfIqwWOdIMpGn7jrGKqvol7OLhtplwiGL2ndJTxcwVV+KQWww7M91RP
SsrfOhq+WVuAmpk98eP/7FmicqokH1fBXAUwjoEYfb2XOs09bh8CqNt7tA/7gz24h+IGdtS86IdW
5x2hBgNXcpww2wMUXrlVjus9jEiShgv39boy03Fk51xcsvJvmv2RPx2rv/nI26AL9XwZVyATpENo
eRmDp9n8aLHjPPygg7k4bxuhtu0dQJeVAgqT7qCdAbocpedGpRIWNeR37m8htA7kgiljXf+UjTWq
WOIjz2lc8ZIowoiVQDGnZ8/GqUycIurQd+KPVZ6rQfPdOhUAI2yT6LFgJhlCUX9IwLQ5nZkKWXbd
YTff4yd9H5Jw5L4jLW25ZqGHV+T7tFLiQal9Fu2fyYlc4Y/MVfFLncZBD3Nexd6Y+NXuZ3wsIrHV
04kH689IQpKv3a1vTgzZpqP4VmR1T2gL+UEhrV2tMfmhGXtZyIzrJCCS/uq8LRd9BVp12+mgV8kk
jT6qKMjHqEjN45T2Mau1iwINzysXcMuMvs9w7QuouliIUDvMtetFU01t+3xExpbPEjpP3tUlq3T6
SSj23rVNNF4LtajJfGgSSAju+Ch8RkOkaWYaxPvezzPZmNY9Oy1QaCNVaQS5/lf67j5glddag+yS
Sl/0xSR/+abcj8f44gtfbb1VfpwtwiQGnm7QwtOu4EX9ZnfctULin2RE1obuJHD1U7t2pSMrs9Hk
k+9qKr498TZcrYodTB/0pv+XejIrwKZXmizSzYi3yJK9zSjJKCHbR72VRIMeaNv6xJU9sQrmwUQw
3V8pfNtpntk/xgwmg0Tun2ZntC8d5O8nGi1Uq790kJJUPMFJMIP/2nK8zR1VBXuBH2rtnbxa9hiB
Kh3KAJFpyHqIGopuKlrgpRPetG2rs8rGt4moqtYsHUe+PsWeUsDE4SPmX6bhjXaGP2njMYCndpLP
2ly9ryxZhMhKcge1/1lgH+KZu+sBnOjXieiTMc2RiWM2v8d9b1PT5BTmUHp3JrMlAHi3GXBgvwOq
/LajR0Z3pW/LMa96Gm7bTAdhbMeeG9iPIYtktr16uNzd7egOCrTXco9ALDu97uo9p8D7nlqCEDzg
0rG63vjIeuYAEGKJPXuTaQL0ZHZGzdwyPL2lB6iXbzHbSJrrsa/BMM4/AbopwXbn5VJtVTsY5qo1
1/IDPZ3rx0tSexk353vqV1PUpq6acn5+VmQ9xMcBcWecKemMgpjDCIjTrTWk4O5YwD1aJfnsxdLW
9xeqO1EQvFAXfU6abps1GeLZbXssymZ/dATY5/pVQPFTDOmQFvfPv01QBD7h5Q6Z9+khUF/rRiAE
Jj1cK7e/DjSrpCuxlIF/g6IYOpLe71Ks82td4cy5Jxdd6Ut2WihAeYWW5lzZLqgQKZNDi5t3ETKs
sZ8CasQTiGaeOymq3vU4/toNUueqqIoK/tp+MN27FM711tSemtpH724Dtsan2pl3GVccmaOQi4ju
aGxg+tPK0jMTPWIzsn59T65e/9Nh3XZAqUcG84jaJio71r415JkHdi7hsGavEdrnzfwtXSJw1aMk
gTh5GcQGiASie9krAyT+RJOmWZdNVu5bGqOzorZQ2YH41Obdc4BSEPOVEhGY6pJtNIYRCE5Q7dKS
cWjcEpquFMg430ev85Nk18XdcAy9Pw99Pefu5FTgR261YCYTXVUEs4C75Ns+iwhJXu7KpGYwUSa1
EcM8CGIsStRxZAyMgKhEAWVaIknkumd7yradSgtwFZKatQSewejIf6nxJUOohiVeCxggPzPFEpue
1nlEiPfhCFYdNFEIRr/k/fnhU1QjvJmn7FEcnyO4YdfF2a+q8SLnn3rLzN+ST8DWGYnR9fWE2JRT
eRfYiZHDWbrUHVytgp4UfmgndCzApZMMyl1kKLK70mhqOUhJTt8RaDkk0d8+7MxwoWujRU2nrwat
atW/pWhoqYvUIFTGNyvv6PI+AysHpDLyAVEREK6GjIdEHAncl1jM9WsNnD5rXFWg13iV2sQABgG3
9Gq5NujNDeG2yJk4HWShzyqC9v7f/uKMb5ttZEuJ42Zv0pKQA5Jqy9zS262kZWNi2JJtW2cmX3Qz
961lkDJxyHoRK83sB3NJCsH2m7hGt9lkUHGeWPVVlLwGZfpD0HGmFT05LO2VXcklBYmiVfkyT2BN
CM0Dd8KycjGiuaGkwcZ0VKwR0Y3C52e7USYH0d494y1Sdw7c0rkDX0Re8ynv3Mh/oPRO7Im+76qO
tMQYzOVzt8iH8ti3UkJA44ZfKTNF6woDt5W6uLgYf8dGweimblavBhtRVuXcYWck1A+i54TFXlC0
7Ix3PyUnqzCNkeD+roS989tkHO5Rc1HX4M0fBPyqkiautRBE6yxKXvDMou2XpU/IqmxhRlg60yHm
s49gXBkb3VBdXWqET2g8Oe/2aLd6L4yGkM4dEGZiRT5wCH+EirXWhD0uOWGTtPhNsj46LDUERdDz
buPIoxRCrIumfiNJxjT2OEHQw4d2VlV04HzaS5fdOfku6Urpl6ChbBvkXpLcDAA=
`protect end_protected
