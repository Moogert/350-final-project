��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���D��ܨ::��{:�6�4�'���4u@��E�o<#��|��h%w��П�M�:�������6��W����~�H-_B�s+{�LnR���{��q��ʝO���
	Eݴ�5�]-l z�2�zK�Ԟ��� �U��F�Ig��{���;�5��`JJ5;6�M2���Mn��-�+󯂀C��U�
��R%�����oxTO��نw�dI_�� oF]_#��o�o��Bߋ�֬�a�.���H}>w�?���~��i�m�]�����p��s@�⋓k�T<�M����^�L��-����r�V�ހ`4�	XWS���GjZh5��V(�Ǽ��mm�`���3���ު�P��1����#�ҮCǡ<�>��u�U_�F��Aq�8Jy�T��z���kzϴ�YT+�B�I]�t�Ԯg��c�9|���e��|�� r��!�g�~�yS�ψ@vf���6�n����&+�~G@����;m��q��Z\}��u�u�H2<)?Zٹ�d���bTzdL�r4�v���b}>�N ��j�lG�����4��%����7�;���C}t��Tc:> c^���R�`gP�A�:���ߋJ/��\����r�MFf� ۴0��A�L>�k�P�Α���6藒F�A(�"�ǩ����Q#:Y��R���<�߷�
}N�R�z�Kv�WsI�/J����|Kʀ]���]/9���5P�Www;V�:@���ZE�.YW��5��>����>�Kay�+�lS)��:�S|v�M�!��e���N?g�r1��'�*�����rn�>n�,=�!h��U�ML�	�k��R3��ʱ�D��2��SxBe�J���h����-|���;&'d��h5;vz�b�u΢Ot����A��O@�܊K�!$�L{<����8>:'��Zƙ3�d�����G�Y9�kQ�
E�&6�v�����N��|�vh����"t����N�%'�t���7G5x����덼���Jޢ-h����ǤY� G�:�q{�N� _�ˢ�b��:A(.�u!���@-�p��.�L@4d�G��>�Z�3)�[w3���>�J۸|��a�����;���)n/��&Gav�3Wm�舭M�5�y�Qdl���5`��&��P&�`�|y=�"H����a��_�?Ư(�!� ��+I�>t�6�����r=�8�8����y8�C��$�K��K}V�/ǣ�}iX,4�^�z]YT���~d��FM�E`c�|���Lhe��8���E_;�G�������Bt e�.+Y�z��D��Dk^�_A2��
<EzlCl�	��\{�F��a���/�����SH`�J���*H�9�ʶ^ZG������NZ��N�����j�9.�B�f�r}WG��������eJ}����onA*/X�s�>8�.�1WܓE�b֏�?:=��b@��ޘ#7Y��$�;<�K�����*y�[�_�Q6AeA�iq���W �[�FJYDq����E�X�~xaʠ�� 5J��2�bP���@�O�-��&4�p�L�1��.��<�����zN�ys�}g	�:�]�4C,���6`<=�u$���C��Rg��c�K�5��r�<�/F��x��GT�jW�`pF�?۴o���Dc���H:�`i���-HmS>6�?`��컧�Le�`�C�Cش ���A�#B�,�)��$do�jH�w�]�=�G�|Ō9�r�j΃�,���� g�4�>�	�W%V'+@���� ͍P�C��(J�R><����E��Ý
vf�RZ���؍��BG����1y$��M~�!��?�ۺ� .=Wh�@;��at(ο0��6�}Pn,6�i�L��I��e�C@���D*�cvJ�z�ywC��÷V{�y*7Di�P�H��yV�$e`{ׄnI�;�\�AS�-�}}�ؾ�ҟ���;tFP���)��A�"�y_�O�%�a�mo\p���t��3�� :���CT�ℴ��<�o�"&!�͌d^\��W�w&E�jL���(��<�[ZI�G?zˡS���		������ޢ�:W�GiN%S4{�,A�"Tb@����j�5��X �Zc�~_�H�-�u����/��_���C����_�ץ:F�z9kW�%6�c4�`!�1�a��*���<oJ��y��L2E���vB[���N`�f?����j������2��s�t�K5^M� 4�*��]2�L׊�^�(u��:R���_�ql��p��nU�珇�Ϙoxͫ��I+ȯ�P���1|���?��s�أ�Ly��=�ǎC�t�	�|u���x�ʖ8�Hk��lin1��m+G��Xߪ=:6��%����0�F���%�,���C�8�W~3I6;ʛ��LӠ!M�[��ay�)��L@D�>^ucZ�5e���vѝJǭPDu�J�ZG�������q������ '4� rbs���yY7��7�j/�7���P��6��A�R�f0����T���7�=y��+����ɔ��M�XƚE&.Ά�q����S��6��Lv�u��48g�m��qZ�z�,�N�Ǥ�m�oX��˳��/��\�R��$V��hϢd/�ђ[]A9� d�ΪBv�?q�LY����Gk��c݆-��#{��w�ȻF�<�^��rpC�v�
_ݤG�_�����@�#<�Q���l�6��q�L�U�"#��Y��2�ߞ�q�*5��T$ig%jQ�Wh?9܉9��L=�g�{��P�>9�����!��N��0UW�ܷ�u�RWm=��mm��.��rM���/Cl|���`����K�6�;B���56Q�{si�OF�x��|�v��#��Q���W=�r�懲�X���:�I�ng���G�o��)ʍ�?U)m�ä�*o�p�W�.֪̂��o�Ɉ~�.��m�nx1��;#��T�c��l^9T�G��?5s���Sh| �,��� BKl�'��8s��Ɵ�i���/��i����},�8�B�k�2I����O�m�T����d6�Aq_�.�9��]{�HvF:�E
5�0��\7�򘡎�/4o�}��#TF7���yO@13��i���1Â���B�6�吞�y=M�\k�*#Ȏ�4Okn`Ôp$c��@�c��U:�|�,�|�-0�Q���<W��,�`��_�ꦎ2A�+ko8JqG�;��\A5 ��\�QG����S��P�@������T���述���W�-��_��P��<�`����X2�`>�ݗ�Q�-Q��h�Z�Љ��L� ':P�oQ�gH�3�<�U����$�ݼY�X;�5��C���m����	��!�P\"v�����\^�N���f��q���}FCF����>?�M��v*�=�(�tw���ᨁ�L����/��Ú�,ڼH�*p� *=�z�&�G������Wb�*�-�MϝM���{a��
�*S�i*����8���ڙ*���ȍ�9J션��u�c�G��+R.��:�ߜi	�K�DMw�l;�8��F���1E	q".�����)�fB�`��Z-� Üd��է����@*��B������%Pⴙ�ca�k؍_����gF����K���M���Ǎo��)��ٹ@��n�Q"��
�˼�+V�����u��v�S|�4)��Y��?GG�L��Is��hqػ���N�"���0>�KQ��H�z����+W�r�Moo*�Riޫ��1CV1T�X����H�Gxg�Zܘ�s�Q�8�� LG�޻�����4X2�0H��F;�m�N���"/LY�os�����9��[�,�Ŷso�g�(c�'�w	0�V��OѬ�����N6,��x}I4�ϼ L��"� ��;c�r�]��N!�H�e���1g��
e�o�x��B<�Č�32�!+~4��|�>�K�À=��k.C�������Tc�+��� �6��e�t�����s$�ص�=N&���'֨��qk$4�5;��F�h]��	���)Q�a��J��S[�i�#Q�uI�l[��/
��̄�n.z�+4F@}~W>��= �|�yD)�he���&�5S�l�g���R����|�L��'z~�9�ҌP�9Q>D�1��K\fL��5��1�3� W��44=h.L��H:I?pgl��5�U�c��&���gH~,}����
�,i[�� �4�����"{m�]�*:���UmA����9"��10:�5��Z��U��,����>~2l�1�EJ�٣��~�R4i���l�߰�3����_gQxz,�י�QVϾP�̤0!���!�Y�wT[�@�d|$V��/�aWII	�t!(��U�@�����e2�����^oZ�y�U�U��M���8���,�"���D解7�!�`��X<
+%>]����p��?��곪K�y%�	l�ϲ���5�) �b�R�R"�u5�4K�@Tذ*��9*m����#��]��C�KV`{������Qu�=�$!!�#�Ϥ����\�d��uYä���&'�'[at��tЈ�Ed |Xw�CC�L9�W��$B�P@�>�~N8�e�Rbg�z$�q��,��N��0��+���G��P%c�T�aSl]%|�n����[}���ͣ�(��X��E��h��Ͼ�o�Wб�%TU{���H�C�<�� T˷�C��o��	�Ju�n5�Np�&wTa�vZ�j;�i�^H�}@��;�A����Moo��
D��4߭�F.�}�����;-�|�4�NY�&�:�k���Yd�%�a��K�e�{|Z�}�iύ熛6��x'+�M����z�E�$�i�9k#�X��dFU������&�%���Y=��_-t�?�z�^�ɡZr�bM/�,���cno2�����Pd�L!JV�87��G��� �"w�C�U��]�:�=dJ.I�J&��:�U֮���K��`����40��zrs�K�>Ԑ���k�*Z��Vtu��EU�SY�O��V�{�0�8O��-��?��h�~�}��_zOF���Ճ����_	��bJ`�����(#�0,i~A ����L!l�E��P{�2-�bT��d�
�<�v:�2�����E<��{I�r#\��k�YְHj��.����hT�e!��08es{tfbq!��Э#��|�����D�1
��K�E-e-OX`|��t�±M��|����լ.�W0��������y�����+�����7]!����|s�C���+D��Ss�D�Jt|
�]N̏�66��*`�V�S�-�:{�H)���� ��/��y�̲p�$jE�? �0~6��C����(�#;��a��2d�$SN9tS��%$KZ��E`œ�U��:��R�!B�=,��PJjt@�"7�!`q��wOu�Y���K%��AΓ��zQJ��W�pc�W�AA/���ϲ�����dm�3�â������<h�ZS\�w(Q������N����d�C�7�bx���qi���m��
#���=�kV��4�]փ���(f�a��V�:a>���=��$���c�8�=�O�^@��Kv�}��}�.4��t�迓mGǆ��֩9��o�����G�sv�,�/���qȣ����S@kj']:�#]���#b�ӱ��3�w0|8���ע�F�@�)���B@}���-�)<N����X[\��Ի:.u�\ob�%W��Gf�������S��Nf:�}�t�30w�����J�npN#�����Ӎ���2vAOX*e������Ĕ]L�'ހA�Nӎ�������X��k@�gb�Tt�]�Y�����p���GnFNA+�
�ts�'�ˏ��O�/U�c�=Q=�0PK�|I��ϱ�߆���C&���>�v�|<�������J5�a���I�hH-�ͳ
�x�(�>�h�{��e�t�SgY�B�/ҷ���bq�Ƕ0�܉��1=�]k���`~˘��N��J��n�����mõwÔ\�ӑgW9J(���#ۭBB���ٹ��WWaL\7 �c�wĒ��H�3j L�y���?
�N/:+ ��{�/��m,6Gˁ��
���Z?�tEp�l���)(��g�N ps�\d	�/u���\�ƙ ������$��
�(��J9�����A��ZVM��"�уf��1E;��8��a�k�9k�	�QW���;F�=
o"Y�U{�r2�9d�D���̽nĬ�0H���Ү�Q�0�u���?�Z���n��p��b�s���qN����.� Xd���n�3��D��`�-B�[�a�|՗.����ws<��В�q����S�S���1�s27�e�=�va��܍x�|��L�7�K0��[��̾�xY͎�.K%\|�J�����(��`:`�MC`�́b���ɞ���-����E@����{6I�V��O! ��i(Z�1��gƙ�����ʯE</���{8o�HƲ���^�0r���/���x�NOeݠ����-R�^��ův��d��қ�v�z'��|Z޹�a�]m��� }���tz(��i�+��H�0��H���X���zn ���.�ׯ�}�"�'��s�uAbCN;e�>��z��X#-��)���i�M��ۖq�Qt������#��e?�ܘ#F�0��g�qdwޖ!y~�q�_ro���Oa)�k#��\5�������׬�����s#7
�*K��4�kG$��A\�T�������N�;�(��އc]����xL��2�X���Vv�>d�����z�Il��X6q�y�?�,����gsuXj|9(�#B7O��&�aY��H`|j�l�`q����[���C���E\�G���=Oy㝟�8ht]bzm����{��.��#^-� T|'�@��i�O|Z �d��DU�?�V)a�`��+�� �)z��5η�!�͙�+�5���Y/�0΄k��@7<)��Մ�nJ�Yp��Kۨ�qNo��7a�C}��_x�EUZ%�>3w�+�6�I>� � ���)B|q�B��4-�,��ΐ��|\h�"]D��u���������Pw&�~V�ש�`\�o ��*�f����n��IB��Sr��v�N��u�)����5��=MC �!��	oTd���k/�NoV�M�
�	�8t�n���x!�W�p?5���_�֍�
:#I.H.���o����=o�ZP�j\��>$�h�K��C�+��I�� �V�`�sH#�`�B˭U�V �+=Ub3�~�:̉N���$p�r�0���l{1R�c{1��'��Ql��ت�o��V�c|Q��� ~z"DU�T��6l ~V�r�D�O���Z4�W��~jrPf�ق���@oq(�C&�ڴ�"����~(���W�9L/�z������ٳђj��C�~ZR�Ѕ��	l>�`�s����$�~XMT�xaB��E�!�d��4�ʣX��Ӯ�l3��Gx�Ҧ-S,2>����--�r��a�B�@ᙠ����;�1���"���R�"1�����yfx�[���q��QȎ�T4�D�[R#0ƅ;MG�X�]��{�h�ss��TiOk�7�����gVg8�p��9Pؘ�H��ru�7)�Lܠ���$-M;K���8��%�s\�A�]룔;)�N3�	�����K�W;H��g�#�����/�R��,�y��@.��PQ޴y���1K�⧏�h#�Y��5��Vm��/8�H@ӿ���0��@� P��Q�k,��C��"�.?���X$z�� M�q��{�E\�}PX�G95�Y�dT��
{�b��!^��@�<�z&�'����$�}�8�����|\�x��7�dW�Ī�L���͜��ig�xe\	�O���L<��]�v�4	��B�ZE�]�8���4���V�uh�Jn/"x��?@�hB�n%���tm�<)[��v����A�Z	���j.�	!֘d���P��by��W֪��-Z��$T��u˳"����UM)�ddL%����h�z���=�Jj���\"�6����5�y���[��}��&�U����Dt�=�TIdi(�oYh%� kh~�M��]?�� �=Q�jdӑ�dݥ�C}�1��˾�O������;�5�m�?ۥ�2�<0,�lY��Eș��y<(U�c��/:�>	y-H�b��GT۷��g�Y�v��}�}��g��&.�DY("�j r�]â���s�jΝ=J��ݢ�m/�6�^<1�9���M�W�z����N�N�I�Ք]S=��K(�h��������=��݁��/��y�cph���4 ��g~���k����_�L��B���;�<��M�ٟ°�(�F5�*�soz��/��G�/u{BI�O�uk �J���U	�W���M�T���#R%�:|!�~�b�\�Li��WKl#��m�L�f��e���'(���������K"g��>�Á�xۊ���0nȪ_Oe�".v��I�+ �F'�2/g�9�s��\���P].K�9C^�Me���\
@�7=����jp�5^!�ҠժH;q����Ҡ3-t�-����I��/.x�.�C<��/�����be��6�ַԪ`�B�d=�
��
���4�9�1�q�����bI:
U����;��ֿ�:^�/#y���?AjO�_�b5(�zȪ#5D�Q(����HXQ��R#&eP������w"*��s��KM�9S1�oZO#1�E�q:+b��1=��}l�|�QlW�'��U2v�/�c!o���mjiѡ�]%a~Ɔ�Is��
��R�we�×��c�&)�U!S`(2��+b7��\�@?;�F�k��3�\�˜��Hݳ�U�B8(���s�����M�W籯"��ޙ�Z&?�cC�j�让܃6e�)ϲ���$p�~��L���@���t�Z�Ӝy���د����Ԫ���@���m�hAV�/�>��޳C�:5�8"@Yj��{=�.zs_BY0�5������1�X� �Ϫ�=i߿T?�-�D]��ʚV�m����g'� h~���#�O����?ʐ�SI?��J(��Y�T��}r����^5�\�ȌQ��u�rˬ�pK)
�^���|vh]z��n����+������ȁQ�/:��X�9&V���\V�
2O,�����&�5Hȅ���_����-�##���q�1��������2[SV���(HA��g1?+���EiuK,� ����N�IKT�'�J	�W���'�u>�|t|�k쀜�%1��}�2NbV�t_��L��	A��,����W��-�0V�%�w���y4kH�^M���Z~���+.���Qo;�s�؜��g���S8۹s�C��˨����(|E:� ���{�Bl�Ş��� ���:��fLvi*!UU�0�H��"H��6m�w����m�@�ob��4(f�a�&�P�&��r�H5)���m��\ӄ}T}����v�7=#��+#��8��V���p�R	��H[�W26����c�)r`z:��.���۹~�mν�vo�<�1�l�?���m�OA�������bcĔƫ�0�_�T �.�.���
���d���djp�[�\��su:#;�2�OD�V�WU�;��A�zu�(y݇S|gp�[��ˤ۬_ՒA�ӪJ�����,z�r����zS��^���K]F򩟘����	|��X�#Uc��G�~�7̡��B��XZT&GzɃ8t
�Xg���]�0��Yy��=�J��� ]���^��'��Ry.�<�s�,��a��t[h�0*��<xp�����η.59]cI]�h8���Q��]�T���1�(�JE.�a�=�i���(+���T��+��i+Q���8�����RwR`���(_(+�i?QF�UM#�
�`��'ў�:í��=��T�D1!��H���@��Ǐ�=ssx��R��> �A2��U:��G����΋N�z4(��_hY�2	`��ɽ)d_�L��&�L��L��}�hޟ��U��Z�h�w ك�ѐ�4|�t��57��+�%i���Y�)h�@u�)�Tր�SH)�f��R�St>so���B�tD�v'�j+��1���	:�:܎��C��lc��(�]PpM�R� �f�p���6��DW�^�h;�X��;߾�^Z)�4���,78�a/3�+���ҭ��K�DR�O#Vm����S�"�E]M)a�J����+�*��_5' �Jy[���K?��U8$���FUc9�{������
4�\ґ��~G̯�(�L�r $�tK}�FM�fe�U�;N_���� ?�NC
j���<����E1�h��2\��c=�����\6����ǋ@!]0s�LF�L�_'u��Nbd��Y�5��L����:�gFg��$>w��Gf-�2�X  �����]/,�`Y�&�9f?g,��Ƭ�tO��4�/<6r���5�i����~��+&���i��_� �ܬf��HR����w+�-�=�K0�17�M�@����Y�x��]BG��'5<�s0�)&���9�IR�r��>�T�����{�-��c��}�%)3Y�M7���P��2��d�Rn�˜G)��YW�K��a<�0J�7��K����Xs
�f��Z�����߅�L��ȩVFU��Z����=������t�܊��DLwW��*��N��$�����u=�~� w�>`C D�o��%�ZR�s�T#O��Js6hʀp)���ձW3Zẑ��lҮ�.J�_\�LZSbT}���I8�!�N%����4e�X�5�7��}�J�`�ˏv]�j���J��⢂m9su��vO�F�pF�fZ��9��KM�=-	:(��J�K@6-��pe&�2-O�r�����Z݂��ы3M�����%��L���a�^����[\��5�|�����KL[��Z�-�An8��̻�Ku1# L�*y5��8���o��5Ae����H�W��刕lS�2w7Qq���6X�"�j�Ϯ�Os�`7ʷ��&Zu���bj�*f0��Ԕ���W���ej'e��~��[�M?�|X��,�k=}�yi)a�7�������g$�k=$�D�M����5h���ې��а��5�,���X0�fP��- *j:}��D{5ۑbm��NRE�Jې���`��QO�2DF� lL�ܔ�X����x�����+���G�":+ȬS�f�͵Y-#�~����,	�5�p�D��l�F͝#�Jt3w-F���ur8c��}L;�x+1Rn��l��R�l��6ָ �u!�c���R��!�^k��H��g���4� ýֱY���A�5�B��E��^;�����MZ���O-NM��k�ԒOW^ap��4H7v=.��6õ �6����Z�D�}^��Ӡ��_�fF�L��/�!�$TVB78Y�~����YքL�u��ـV5�o_�:<���wϔ����e��!��<R�0tE�ƀ�r"|�C�GWɏqk�D���ԗ)�h�혜��
9%ޓ�X��#v��U5�c��"����[��vL5`A]HًC)k_:亻�̒��"В�
��#�bP�3?����r��}v>��a�ajq�����`# a���kI����侃����aDbb�}���\g,5}{�@A*qR]t�Oĉ5�{�ǟm�C�f�Ā�t��ruX};}Vˠ��a�����%�.��Qs���������U���y$��.?�%&�T���������ͽ��/����O7��rXpQ+��e��M�GA����!�E�O��m���bx%���?Z.�	:�3�X��$7�V�LЏ`Y`�l0mu�˘�v[��Ay���O3z�4Y�R�����a���c��%���Lo��_�vA�4a���˅Hg�OS��\����a�rʵ��
GB�����	�Mk�܏��~l���qEc"��G��a� 2%����k��w.f��1a����Ê�jR�S��P������z.]�5�񘇴��ؐ�� Y�?����#��7��3` H�W6�}I�a��2}�MF������T���IUݭy�CD#�=�#�ǋ��R'��'�4�����*'¡s(; �pd�OAײ�ya�v��0�!?��2b ����y�Y�V�m���<p��>�|��]�]��UY����<e{t�����Q��\A,b*n�ek� ���O��
 ���J6<���Ŭ��J�t��`QЦ�(��m���t���sr��Pr���	�ӤE�7�Z3V
2����t
�y��2Y��n3ڢB�/��X� �a�+&��e�)�&���3�PnC���T�x������򶟣s�K%�҄^(X/��[��k�Z�qlw����I.���s�����&{�޾k�|Z�s���Xen�>uͮM��N��(E�A�,H_�������/R�}���]�랰�%����/����O��o�K(S�=����~��	
�V������TM��1���)l��AB�@���q��M7���<��hŐ80/���M��!�C�u}no6�z4��ZU��ס�2��A6�Zd@�k�6�fK��o(�4��7�a69ZQcr���}SAV�|A `��;��WT�����{ �^����H�;�>a���C~e悠��M2x=�*r���{)z9>�Օ��j�#���lF��!�{��
��ᶝ���ql�b���Z�i�
��X�ߦ�%�w���<�oM}�ܱ��Au�!����E=�}���҃�N�\9�d���*KU�9�[e��Z��ZjP.Iq5`
=�˛�/�o�q;���F�^�9#��K�h��p�m��U�A���ݧe��B+�b׮"�A�W䢀1�豧��%�P͢V��HuA`˻�T�4��H����������g4_���� ��Ʋ]�&�e�l�ĥS�pCq�S����Kqf����5�Fin޳Y�Q��^i��/{���ȿ	,XB ��{�)��*bh=�����w�(�M��q�6SA]iA��^���n��S9$17����Bu�K�h��ށ'v�5`6�6`�(/���J$��O.^9BT���aUu�����1wiv!�b�SO���i)U��A�E�M�/�A&kNB3�ߑ�!��Z�G&]$#-)���>�ٹ�GW���2��>��p��Α3-�Z�Vgg���ߞN�14���'W�o�Mp�G����%�zK�Sy�K��)�9��dB`��}�P�K��q��DR߶f���Tj;Y���j�MPہ� z	n�����-��g�,[�0YMB�Z�qB*3�N(�˙���u����&�q��D���-��w���)*�uW��0x{h_D_;���&�#d��J� Q�Jf��1ِ��2����5���<y��[�=G'�JD疉e f���Y'4�.�K}ÙG۠O�{rj�p(�6��%5Ʒ�б��9��?�:�����<q�[���O����FQ`�"l���X��li���r�F0(�B(���pz��X��S��������gW���𧧛`���;l�mx�]Ԁ�	C�\�j���.G��\��\���R9�ĵ_�4��s����9��=�����v�BYm �QyHM�o^!��M���}	'��������_��lϤ��<���X(M̐�v矞n<�^�i���0�l3�Z�%ށ8P�{hݢ��(��:0(7��^T
ʘ�Ok�6��1־��{KVb����S8����rw؊K������$��zi�Ǆc��"�4du[ou�����z���=F%���[��_>�"V	���'3�i��t4���_���y�eI����������B�Y�LD�M@4}v�,�����E���Jz���'���P2��O�I
�c��D�H5v���Ё�h�Q0�h��#�h���4�~Q
�m-�\ϱM�VKrK�>���b�^JO�o���������Ž>*o=��'�۹�V���Fs�o:�uzK4i������Cj������2T{l������ʣ�����BA����Vԅ�!�=����T3�.Y�4��A�g��GV�^�<��S�3��Q����Ə��Շ�h���=�qɳ?/�$��$Vh�����{�T_�+8d�+`G��j�_���n�� ��@ð�� !��wuz����(W���o�K�eͫw��
k���*��Wd>�@���ۻ�>Ѷ���x��^���|�H��(��e��R�?py���/9����s�j ��r����Z�N,h���$��9�{��ƿ�Ɂ���q>a�Q�-Bp�������dN�b��eM ��#�w[��t��EJr��}�M`ߜB��g��&B�{:[�Z<���zy����!	�e��@s_����'����6��G��֐t��1 ]����F�,<����pB���^�)��EI�6����-#W	���m!t��%���i��H�w�'��^���Q���s�P66����r�i�����OʙA����yN~"�y*N���G�pz��iY��2 L�_����H<F���=T�ڻ���U���x	�y���?����`�ġ������B��$'ۘ �v�HB���>>��C_��|Y���({S�Q/�H�u�!�g�)���c�`���si-)�L�̈́��ِL|���c��,!�5w-��H��9x���A٦Z�?Mz��~��IH1����LV�u1k
Ӑ��i%Gﳚ����T3R!e� �=Lv����S	�=X4M;��.���C�2�u�������G�:�9��B��.�Fڨ`w\�P���LV�z��L1�_3IaS�̞�(vI%�y��^2=�Ͽ��| ^�Ԁu_�a:�ֈ�r�
R~ց\�� �����G�2��gS"Y�i�PH��W> V���! ���������"Ֆ%/�˷���;D���o~=ƶY��ᖦ��������~�qI�lb����fO�7@���&/����Һ,�P|�CAZVу� ��!XL���c]N��L\ P>�HHqH��yaX�A�vX:-���:��3�3�#c�v$����g"K�@������&�������}Y<N���iмl���lS�X_ x��� �/Gؽ+���J9^Rߖ�������ؐ����:�L�m���U�@�ZZ��Nh1�c��Za�{M�� �J8�.E3�p��kW��KJ&|_�o��C��$����)������T#�4�O�V�^�zĭ?�ьC.�|�84���'�.[[[�:V�B%�x����G�� ��a�,rO����	��}��Ӵ�>���P�9/�x��xf��	���Jv�i�&dqJ�������kC o	����0�Hu6mk�vs�FaB�^���/�F���e� VAy�R����������ۖI*�3v�Pr6-�щ����'oh��ːHe�_��g�/7T�2\�Mg�X8��V�����\*�ꪏ~�{h�-Ȏk��&�.`7�鰸��~N&Z�����]�St�$�R�"��qL?8��Y\(�/��.�P���� ��.�뿃{�aC���t�n2�?])��閚�1M��) qdO���hd�v�|��\ټ���E�B��	7$o�$*�e?F�a$k�w�6��O��M���B����p�x�8G����ts)�V&��(������D�H}
�%�pM:*:�t����8�/?��r�p��qe�Dq �2�%�P�W��WB�
��4(�4��*�ρ��w�h�*˛)I�����m,� #���Ń��j���vh�|�<��X��ș��"������E��|�S��H7%�j�C��B��:kA`�EV�,Q)F�2�/���Ƥ��qz(Z�F	|@n�S�G��}�#���xP.�6����:o��/�	�T�&���98���ʨ��f(Mn2�����rz,I�?��J�f�;-Q�(_���& �m���^��d)��*�b('{$N6��D��5� �;wT]���n/�^ӊ�:[�����Y0U�1���(ЩT�}�����5��!#K^}`e�Y�qNc��m�2�Ib	����BE���VL�Z��x%Nɭ�L>��H�=����T,��o.�:�_�c�ZT�ޅ�&Tغ E?([�%��=8�� I�*�a ����7�v2�ɫ����׏������w�:��50�i/��5���{���&
�@�(%-�N�}���O�l9���(XRp������ZQ3�w4��!����B�-A<&�J�C��l&#V�U@by��P� *Hm�X�
9��J��Ǥk%?����#!B.��F�Vj"���L�y�?e��!��c�:mz�����	!��e�cz>��&�o��'*��t�3G���1F��S%2�G�� Ӷ���Z�[���Ǿ���7�g�g���/B���ѥ���N0<\oz5�����z{�(�N�di�5��w�V ���.7��껑�,��V��oc�����[;'�j+Wl��n:��Zh�/���9�p�+��eN0F��%/�扼%A��7����������/B �r�e#U�`Xu�a*.mto�����V/�;���p�Q��x ��%!����$����c��?�1�.Qh���:};ձ����լ}�0勢g�N����Ã1A8t
Ì����۲�C��$���"��w��u��ogƠ��2���* �[HS�4��R!3İ�0��A�zX�l\�vӞ]AiJ�0�'Y�1��\��m���0�6�½z��M���=+�5\n�*�M8�zL��a���/��e�W���<� ��@%^�J,��Hҗ���[��&�_?��ӌK�X�U�y���yE�卿H0��[uG(��m�AB�Ә���XVP :,���)�.蔺����N .��YL���6#s�	�0��&�Oj49�����&d��U����#�r�횤XW�<׻��7|�J��}7�-���\j��~�x6�NA�2~�c)A���E%})d�Þe�2���m�U�ɞJ�x����A~�v�����[毠U�����Ԋ0�ژ�XP�s�J��ƫ7���[�J!�&�CVa�m�o�� ��z�g��S�9�S��s7mZ��N�"	pT_FUb�kύi%q��@Y�zHK�s�@niǿ8/����2*���W$�0���)0\��fj��������U�b��T$�	�hL{v�쥥�{|q�?UA���Im��EŋM!o�W���f�B-α'%��ᶿܰ��ō�p����Q���$��oȰ�PӖ}��� ^��Ƣ!T����f�����6"Y�*:.�Ƕ�=9.<���"|nO�~��vͷ�^�kM�U��ѣ�2��h��Z�cXIӦk����/�/�x�N/����v��h�A��1Jd2P8��H��l��"ɻ�>2�w$���6J���Q�f/8Rx�($��}��	�.<e}pQ���'�;֙U)9�$�_�C�,��G�txFg�{"��ɠ��#�tg���79}�1��N���e4�r
����)�\6qP� �?�9V����q0L�X�櫜�O��_o���?�����(Èv���s�5Z��@k�m|��)�U�x��$�.�4>-{�����!!_U��k�hl�SAg��#�8bٔ��j��ޘ��!�d���C��Ý�%UN����>��(�jG�rc��֓�;�I����㟫 IgU�U�r���Ѡn����; �S��Cp��ڻz̋||��S���WΨq]��l�����p�8S��T�u.p"��&Ü�0���M���ms<4���1��V�� ��m��'���&F����5.W��{���n�i���dh߅�y���o�����Z�Nr:#v'�Z���𨚘7G7� �y�~�#&�o�H�gU�3�(R#���HiR�T&�@eH��3��K"�<%	py>~w(\�̢Y��h��@Ѭ�����	�7�%�@�c¦�N��Re��̳�}�!�x o-YL��eya�i��	4�R{M�_�f��W�S}���O�|�����f���o�0�JDK��f�'w',�����9 �C���N3/��q8�$<jFԠ˛��*�߆��Zg���e���.4�n��P`:���2��	 �Ȓu*��\pG�E]@�^�� Ѳ#"4ـB��{mH/̨�2��E��w�D���D˜3,�4�,�T�o0�L��wh�������8���e�L���)�_�I�@�t0�	�{�� �Bo�᠎�z��MC8QI��&}��j���)��e�����o�'g۳��z!#�s`u0�5�[��vϙ����x֯nl{ОFY��_�G%pڳ&!��N�fYZ�^����Z��c
�g��2�7{�*ܕ0N�,��
{P5��HGm����[�0uC�~]�N���k��MS���}O�+1ɕ�C?_i�p��0���}ҼK��n���l�Py��_wM��w:��ޛu���J���kw��~&����v��o�l�(�P�oX�\�5�)鶭��>�`���c����V��\����?]�~���Ĕ�)�x��a<_�d0�
60�֬��A����I�ԩ�|���gp�s� Y� b�JW�UT�������
�{����v
�@5���v�蹨u3��1f%�6Nۙ>��C��Km�{�Rq��h��0� ����8`;��HE�g's��_!�N.k�U���9:���
EL�����Q����Cu���1HD�����g@�6�s�K�-�����d��t<��}��z��\n	�ܳ���>C�I�PN�0>�A/���3L��"1:M{.a��T�h��|��es��X~��Ʌ��2�h1��!o	u�(�WC�9X{,��j�N��!�P)[���H��@�ALկh�Ӑ��@�h��Z����&z�ևO7o���%c-��IN�k�&�Jā���%���Y�����{�@��o9W��W�R��Ҽޤk�>�d����$��e��0~�Ve.a/!�<2Oy�3�z��!dBCyoZ@[戉�S]�����lxC�}�%��{dC0m�^��;z7Qћ�y��3�P���Ye�&���W�����-�ɺiB�s����#�����?/��5���"p��ا��Y;\ �y�h����-�k�7׵a��D�ӛ�%5<7l[_�ڝ;�V�ݽ*�"bN�00y��ĸ�0P�����8c�r�qyM*�Hk�;�\E*�V�kDd�(���h}�����<��r��چǪH���-�7�h������-����W��ˑ/��6X��R�ӿ�0dx;[ߜб9�a��_�������������M���o�9��J�}�P�[�:�P��T��gO��I&ЃHq͜0Q�\�ET0�mFlsmwZ�1L�P���{�|�������O��\��E�kZ����d9y�Ώe��*�57
���0��>�¨@�i뤙���Z��ZJ��;�Z#s�Ns=ʢ4��lI�cL�*����sʑ��p�.}:�e��9>l%�e�T/c��)��8|~���q�wq�����f�\���R����®���G������f;iR��]���;	��ƞ�ul�n��o�0E'���sg�xy���w)��`�?���m���7���1�Al��=_��<.6�j�lK��zO����\���w���]TK|��K�?�*#���)�S���\�cM�w�~�<nzO�yXA�Ġ^��y8��1��':aK�ԧ�ܟ�(�W�����G�����Qf`���%��`���P�]�4��P��VZ�?���(p�:�� ����RϽ(���))uc�����o 2bʗ�2hhk���/�����gP�,���(���<��˰�����C����'����rЖ��a��)+9��n�ǃu�����%:@�"��Bъ�r�'_�^�*g\~�"9˞����,�߹�{3v�AH$��*��%Cޠ�9s!��rͯ�/_�eWP�#!���˭��躖�<�=��mP�2�~�{�?���X%Lq.�&��͠1`Nqk�����Rp%�� k��$��̱e`�(9�^�4��zt�j"�R6�Xt����@�|�z��k���N����SvNI�+ӭQ��B�Ȣ��X1��!oNM��\K��JAtd@��vu,�.��<�w��{܇c�B�������vΒ��Y>ޚ9)���R_�k 5ŵ?�K��ߞ���?e���.b�����qJr��Wxd��W]7LQ=ؐ�1��"�*Cj��7��Y����&���
F�8���΄�h��3���#�~b؍�Wo�p"$���Ű�O���W�_|Nъ���8�Ѓ�m/�����А�<s(�{|}�V�M���s4�B����V��C�C�\4-�G¥����*��������	�a}N���ζ	�h��!���y��ߤTp Ԑ bZ&��b$Frg�<��`OگH
?��UR}Ԡ�(eN�����a��$��)V�2��ܧ+���4t�|�k�t��.��L�zV��ގ�[�����~bƔԱ���v<#�4e�1"�ţ�4����2z1�0i�vi)BQ�+��(����HBZh#���#�bmX�^6��;F�]|t�WO8[r�sS�(��n�j�]��d�#��;ڦlXP��w̲~�@ز��Im9@�=CC�&�V�j�����rs͉-<�3�!C������=��g�`Kc!�y�1���d�N"8�%����xwmn��ڣ`�3S|�:~��H��
�VN�8���T&}=��8]�����C���� =��K��c����\e�=���'H�����T�l� ����kEwY	���Ĕ�=���(q�4��me�+��b�:i� }�!�`Je
ii)���)�8/��e��4�t��	���p�i�Z��d�Ψ�7�um+�##��6���5�M-���D�-����M��L�C�����Lݬ����gd��[	�'��T%[��,|:=����8����5A���kk�h��(7���Uo�zu/;��@e}2d�9����x��#\���/���#�v:�Y� �))��Vf�A1���Q���Jf�{�Q�S�E�v*�bm��MSj�i�zH-�Qr	��t��}�f-��=�w�0{5��;������K;A�Ո���W5���U8���v1n�8 ٦�ĭ�{��"e��徇h���o|0țϭzٌ���)E+0�{���Vw|Z�|JT�;��?�;�cl�8-A[QuXT���w�[HB�}�����d<�>��H��������_n�?��[�uɀ�)d�#xSnE���-�!�Ge  ^��`�o�QhȚ��d�Z�{�=Z!?���V�߃��j%�'�v@-.�FJp�3��}�1��:��=5K������]{�����9�T��d���#�GC>
�r.�if��d��/�f��eE��6�;��v˕�U_v��b���mH-n�NHUq~r���L�4Q8�v V5�Ḿ��Uq���5�b�ՙ��o��h;��n��,*����v|ɻY�`�"����n�o�:�_�؈X6�������u'F�[��^q�
����w���F@�It�D�Q�Aբ�U�C6�ɻ���H#�'��xR��}.p���j������Mض~y���_�5dx0,0۬OY`EG�]zhp�樂�+%�lY�K~>����FZ�OЕ�ܠɫ��p)O=��5ZST����i`�'�y�h���,��t��{�;Z
����Ặ����6��,<�Ʀ���$(��4�f��0=����0̮��K��^X��<�������E��ʻ~����8��q����n1B����rt��n���.,J��˒e�N@�[��I�v�8��A1�����_>5���i�Me%WA�����\�K���" jn�r+F�x���[����+��������u�#?�y�~���W�W��ɓ�rI�{�4�|\��K6֨@r�+�"o	x�ۡ��<���8�����> {:��w_O����s0�@�O>���xI�A6��n��O�:�Y��m`�Y^���T̹>�y���)��K��w��x�'�D}ȫ�����{�ы7�$)o�H �%�X��6^m����k��VO����Xł����FFN�%�
+woF8~�$�A~������\pT#����&����F�+���m��i�;��T�?�M��Oς9\X���3@�D8�ɵ��	)��/y�g+��M8�Vi�����aǺ�d7��gx&���9�mz������`���T���Á�62?<�0|	���k~"I?<��עG���'l��K���/h�_M�����&+"^n�*- +Ί�$�����50��"�V㤺�N^���p	Q��,c�S�RG�����Z'�_������q�5o�g��.��FW9^��-�;��i�o��ZR��j��ro����M�mpu�T�fd�5%���EX_	�l����ݍ8!%�*��b�j5�k�M��g�yF!�y��x�w0�'h}��+<	"h�����^<���
.ۿn����}�����647t�`eE��$;�!o<�j)�[K&�j�Ģ�|H�>E���`K�W�ˆ9�ym؂� �:�N�,�%�Oo��zǡ,��rfs��A��m�;f�D���
ٝd�:]�>Be7-���imk�W+ؓ�	IDW:
і�w���:�䄼]~A�	B+�{��4�}q;m����8��7(<�$mQ)j,��B��$_���� <�U���t��I�׀��rX �GE��o�3L��5?@uɺ��������u�$/���ݨ��%9���P���&,5͙FPN��BXW�T/�[3�8�V�q�8��0=�wI�:P5 �|� ���e�k�����*���2�h�ߜ�MC��ё�0ƻ���Ai���O�����oX�6��4sT����m�b�`2�k�J!���f%��T$��d����4^��(���d���K�\e���bPO38��vf�I�=5n�N:�\�ɸ۪憏8ʴZ7O����O��Y3��~[n�i�s�����x/΋#@�N��'��>�sipU�xD\1��b���*g-d�����;�ݖG:��$����.�-����z���6!���T�?��&�Rux��Cb�+�X}Ъ#j%�a��ൾ����c����P~���
>PdD���Z�/*ȩ磪�ܬ��{�p�a���P}�_N��t7�%���<��!|�<(������=}�2�>���H*�Ѵ���������I��H% 6H*��m����lhQІͿ��?Ce�nt����_�߆��)w��o��D~1�IR���3�<ѽ��:
�X����)��Ma���ia�S�AAcI�R�7@Oְ�姢o�QWc�6v-�SJ�/�0	�<}Y��hh��f��mc`$Q�wn�b��#t�C#����]g��A5��=�m�Vv�[��X�g�&×�ezh[�ʆr>h��k��v�HzhC�V��Ј �h.�?I�kb
��t���=�0��|i4�1�E%�����	w����կ���C2�a^S�Q}�y�>��.��u8���/FYms�������V����K��s�NZXY���߹��X�>���r�F.��i"%�a�'tz<ѿt�v��y���5��E9]�0y��Dݴ�0K�|�gm��[��0�Ko�_�>���N,��b�5}��]p���)z�ژֵ@�S���TѤ�e��'��Ǯ`!�'��#PżsM?����u�k%)�	p-}�Jz.�e�����_�c���N1o��`Z* ��K�h�X{�|sV�U!.<Z �Y/�8�Č����ا��j���b�X@�]�J�(��*���ҁ����Yv��E��2�`�f脌:u�/�(�����A��85E�$qR+��"ߣtx�����u���z2�����N$�jC������D�^���
3��7�-u~��Gyq4��R"m��(L��пu���6����pL�JSF٦�Wk���.u=8�_�ȑ����\��]�������>0��K*t�
�:&���n.����'ߚ�=��#��E1ᰯ��s�Mu�Ή�K�x��*1�`���JE(9�jQ5̺P($"פ�h��@� I��CRn���sj�1��_�DA�)���UR�(^�o0�F��5 �@h#�r�MC�^�ƼX�2�^bD�96ݹ�������v��z�AJ%���nP�g��ُ1ǟ��8���D\����q��2a�ǌ�D�[�+���������v���Ol��Fq��0���`�X��[z�`lV��͟�*�� �e����g1�_�`���:sT1L�2�FbϹ���(�۷Y*����1.8�s#������^=*6��!���� ��%}w7?f2\�#`d�/q0�=���R
PV����|/�
?R�]��4e�wW�����IB�`�� ���
=�Ә�jv��L��X��T&�?����)'�v�|{tG�U�Z�H�ʉ�"S4N�A�i��c2��e�J�UwhM7}1���XVx�9��IU$�,~��]��3R]3���V��4	�F8m]u�]?��dC��q~��0mi���Zh+�bz�lؽm}�=��v-k��<�$,F����%�*�����«�u\_�[%�i��k*�I/S'�@��u�(/���K�+��DA�&�3�]ş���O��~�E�=ڌ9Ԍ�aI�����@l��-��S�0��ܸ�]K�<��2-�׹�D�YlF9'27��R�,*jl����͊B�Bl3��4�|.h����o_>^�#p,��_�l훗� ���l,�}WƜ��]�q�om� y?�8����1U�N/�����rQ�����u|U�S;�+'y���#���ϛ�.~�q�'(��{�&��Z�����i*�6�u�=�'��\����/�ȭO�M�H���M?Wq���2_]����`J&%�n=x�`�����ɖ���\g�Ҵ�x�!��U}�+M=�xX����o�TJ7�1�4U�^D���RhD�w��&Y����g0�Ĵڊ��Me=����L���q27?B����$҇۾�M���Oj�^ʓ�/�VQ�J}��,7�J�ޚ	׮Km��)I�
�n~��B�Ѥj�،a3�E/�>"��r���,���`侎�2)l��.�E���D�~��b�����Va���<dU4�;�?�ꗓ+d8}�ɪ0؅p'�#�t1��+�Px��A=��i��q�޽S��fP����W(��~={�gg3�(��2'�?�؆�W�7���߹Z����?��]��C iZ��̓\>x�?>չ;��|x0�g+SH�cL!3� �ܫC��g�3�NA�����%��?D�7 ��~�ktX��HɘO��_\�~H�;%o/�3o�DG,�^�MuCع���k!�����u�������m�Y!o��R�|N��m����:���"ΫE�������7�k�1����~�r���٭���_���o6bs�6�;�k�qex����y��Z6-��RHH���2"8��}����A��t��_�'H��ј�B��|HT�H!L�-� `5p��y'�ލ��U�}�`M�v)����v$5l��X��c���Pc��)dj=H8�[�o�W0r�j�����I�@(d�l�	CА|9��R�Į9��J$��3�l�EH��(ުw�^7h:@r7��w	\��\l�Mp��%fkQ���q�	�˨f������YE��K�c����1p�9ܭebC�n\����7��>ϿB�;4�9RUH>x�`�J�����>l�^[R�ٓ��&���ٹM����?��#�=e�w��&Q��Ќn٪ښ�J�h�O��Td��������yf:��;��z��GpxN��Qս�ց�u&-/x����]*��_�E]�����V��K�g���P�LbF@���V��Y��D�/�)_b�]^�#��&���!�.7
� a��eb���AZ������ ׅ7�A%[�!Њ�o�hm�:뵮ةń�1�#��^	�}���ӏg�_��F�SO��������:����ΦX�f�/� ���i�yu�����.��h� �_��h݄x�n`���=�F�w�E�bN���7��ª��/�R�;+�f�8Y��ʜ1!r_ibb!���7wn�7^�Mt����&w�02�J:�|9'{h�*��迍��P������w
�
!$�[�x�n��ӑ���`����)��6h(�
�&L����46�y�V ���ʣX�:������s������������!���(E�o�#å�� kD�Ds�Ju���7�ө�w��\�P�h���H	)�q��ʂ��>_7w�Q RM7�آb���!���@(1���]bԟ-_F0�}�+���S�C|�=�>�/)d��@k�ںkY2�B�.�١|����"���<�z.�?oeZ�*�4>�V��+��`�N�"�N`=��:�3m�E���Gd)����ϔ^ �m��Vy����dee�S���l�-2��ޜJ��XԌ�W:�Y���g����ay��� �˳��0)݁p {"]i-�|��� �;Luz�M�֚�9��P)��uCJھ�����D�Z�Q�}L��u��D�ڇ�0�[>��A2{v���U`v���t�v�L`��8v�.�GA*q�N����l�`��4�%jj����2>�&���Oen�'k� uo"�r��0� ����?�dϖ��[��y�[K�h�r�9�=�I��!M��|H��h')-Y��L<xN�ˏ���z��Wjx�$�7�Y�K�s�q�4qˁnR9.N��y�ziUDm�*W�)�>��x��S����
��Z��z�}2F����;	Vh�>�} Ɛ�(@�䉔Q�kE�׮�NxA{^?0�I��
%�kk�Y����=�=Ɠq�@hom���9~���`;fW��&y?p�Dp��k��!�A=��r��=nԺIlo�&�I�����C�j|s��I�ވ�5C�k��]�姈� t+
ä�� 1	Q��F��X�p���� D2Ƭ�S��V�C�px���!����͌`�G�?B|���~B�
6Y3g���ʏ��l�B�o{ x3_�}� �T��'o@i�q��ߟ���a����	~`��%XP�{�|�c������\���H�z��G^"�~f���8���A
�[�e�e��Z@����t�;G��La��w��\���"�bK�s�g����ٽ����	�gn���jp"�n�C�4-�4��b���#>�i�}J���BQk�#�1R�=aC3
Ҳ0�;�D�,g�X,���^���X��]�a>�K��ў�z�Hy�ǆ�?�"�$(���KTA&�O�L��XM᱿�JY�
��t	����5�G���`o:kŷ|�P�<���
I�u�� �����.b���g��*f'���Ѵ^4u�m���B�����_!���Bw�If�$�{F���5�yɭ~R8 �N�5�S��A�wO7�'t'�!��LR�$m�Aj��,l��QX��-���a�TQn���љ��1��Z3�c$,!@�X��S`�ʐ�2�|��c�=�̾q��?{q���SO�GE+���Α���a�6�^Y8�ΠֺB���fӴ�4%@�Bl��-[c��8)飁��8]x��*jW�a}���(��P�Kz.g,�E���2�o�H*�#4, ��$�o��9�42�/�%�j)�*�5��]��s�r����+�I��P52��+Y�/��(Kk��W�V�,��5�~g�[U�Ϋ"hٵ���L�Ɨ�m81������w�X����������*�|/�o���]�_Z馣��O�V�+����P\M�rE\g�;=��	*�H?H�q�(5܂��C��6R�b��[�u�������Q��Sb�\VTE��|{���x�,��d�v�mc���\΂�_Ԡ݁�-)��v"���*x��(���c8��#���d�z��Nz;yh[��[����m\B�%�4x��������'ίa�R"췏F����#}n�/�q�`Y"�����rc�N�ڄ6Q$mF=�{ݼ&��{�Z!�O�w�X��+�!�E�sC�`�MMaDF곏GMƾ��Q߾H�?j�񴟡������l#�=1�p�@C&����m�=9�v8�xH��H�Xk0�lBUY����˵T���
�j�AT/��$��c4��c�l.�huJ��S�`x�70��=�,,6P����t|�P�W�e��t3٪��c',xi�?���><fC��߆�O'��H��R���E.�z��6�Ω��XWP �=�K�΢2����l3*�u}h�$��fcX���)woVW��jR�ltw؁����m"�A���Y��]�Fޡ�:"�c�.�&="�!��@x��0z{�M��SiJ����Ӹ�X"z�r�oR�bHg��Q��d�ˊ�ӗ6�R��[��.��h'�̇{_�o7�#:ZSS��i�>s�& H:̧.t�s�i��6�N���t��j[/J_�'^��X'�q�I`����P�z����I.��{�A	���<�H���%�ִ�vυ���`y��K�,'��]��� �A�h?���3�B�J�[��o5�tW0 ���F���BÄqW�w��)AY?�A<0W��7�U��Ý���|D1��Թ�\�a0�
�� rnX@Z�~s�g�Rm����{{�_�O&6�q-��I�O��凚,-t��ǒ �wLR��q���J��j[��Rߜx�pV��٩�Hęt;l8��h�yY���_�(%Eׯ:�C����5 J\�Bs�s�غB���+�7௻#$�w�Kr�X���87�y�\U�xB��(�t���mVA���jj{*u���Wrg�X�����P�߿�����ZP�ջz@��5����Ȟ��xB�TGX��w2�#����f�z����NrU~ �@ޮ_�&~��RΌFfz;�AU;�;D��\�UOu��E�Ո��U������,����b���4��y��G��bI�yz�g����������?I�����.
�����[�3�������Td����VO���t&t[Z���������l)Ly�Nmi�B�]�r���j��Rr�;�iN�E�g�f�1�����&�y`�O���Y�J���#��������ѠqH*��C˻�oY�#�W��ݝi��>�Jodyn������l�����2���=����<�MJ6�>��3!ek�Bˬ��Y�~�y8g[玁���Xq��Lj3�}�^̾D�}c�[ī�nxLh�\��8�@Ws�1/' ީ�j�m�_{��ٞ�a�2s���ߊ�[��M�3yhHS4��$�(<�3�w�]'�^O��Ӕ"��&��W�GJ<�s�+T�I'�!V�+�M�r?dz�(��{B0�p܄C����3�&,(�u��!S���m�ZIx�g[�h����s;&P�ͧu�w���y�K�_n�H�!��Z��$������+���B���r�IC⦚��!�Gq	.�����}b��t�d�h#e}�b �6���ڴ �}{'_Q��F��ܦ� �M4wY�#M.Џ�<��L ��ݒ�)���Zm(�w�j~�Ik��c���k'�Ep�� �!��� (���G���Dz.�E��S��/�s^
w�\���\�%(NV���� }�x<P�C�?_\z�0�������0bp��C�<���=�l~u��5_s�A_,�lގ��%Ƹ(���;(��P��3�o�9+w�V�Ҳ�z�i}4�˫Af��ɫA�������zB 	Ν��>���I��m�1N�Om���볡y��	zZi
�B:�gw0q�e��7 ���br&Ϊ�{��P���-�4�?nؖG�X�6� ǜ�꣪&{ON3[k�\W-{(֘_9|��`� 9��B���C�:{���B�,5'��$��(�Au#�*+��,)WJ��l��¶��~�n�GIs#�{f�G��~�ރ� ���Ec�������X���7qH�j�ѼI��+|x����23�)��D��>�}Ӿ�� �ZK<8@q�%������ M�/��x���(���>�v�.Cm-gx{Hjyܮ��X0�k1!�����IL�6'�rY�.���a����
���8%���>;�*�� ���0a�ZX/�o�ϫ�r�TQu�s���O��k�!��#�!QFȅ�ύˇ� hAs��9���9^kU�u��L?C��K��Ó_�o�El1���>`�bX󼋀=SPK�,�h�Q�����~����Ҩx��7����k	���)LMB��R8���{�,�9{���]g�%�*����E>^$������$��o��*���ɭ��/���;��#�/�ܷݠÃ���R"��N�í�;ߣ'*�ZGm�k�ƚ��/e&����i]�=����Q�k�՟D�B>8�&�2�%��X�uM�F�������g�t^��'n��Y�׬�x���G�����MX�Ur�Fb{��ɒ"zr�4��A�P,YHY0:g���
�0g+s�����d���u�e���q�8�]������ma�2`�p����姢��͛��v7Ph���9��h������""��5U�@��D7x��Z����C:�H�)��ɺ�a6����>(�&�l����Bzw�x]N&e��Y5V �
�S���̤�O��u/�UR
�C�m}�%�&R�S���B�����*Q[n�5�G��V�V޲pR�;���Bp��q�}��h�e�ԙ"���g{�# d0���FzI��\�d��м2Q�N�s�t�0� Q�?7�&�*���I�ݒ��!�)cy�"�OLYP�IEKV��+͕?�Ջ/�Z�����vj{<���\|T��D��3@��I�.����}L� �`���1��
k[���Cz�0 �ƥ�8'�4�u��j~[�/ȧ��O&�=Mu�8'�t���D��e��z�.�N.^!`օ���p��0`nܘ�\�u��s"U��M�s8I��;�q�ܥd�E��ȟ�l�J�Z�	 +c"̨�^��/ۂͼ�or�՗�~w�8:2I2���(.WŠX�ݧ��T�yכ��AT�d"t��9���;�|P���CkJm��A&��?��fb#Y:[S�CҐ�.wS&���!`����-�$�Q�ά� �D]�9t����>�Rf�I	j�����'�]kpOBB��Z�Q�I��d&=�!����	�-�ޟ!쀤'�Q��b��I��,j��{-�b,�l[�)� a�
�S�cq��
����Kx!���B�S�[�/����9��Y�{�.�u{����Lo��|�5Y�����`��8E�Tk�!yA�7����P�(�w��BA
�r��/��";�&B���O�Z�����T�l8�h:�(�8kШ[�^��X�T�;,ݗq��f��-q�X��C��(�����&�{6�y<rT-�(i�A4�f��\>�ulP���0@�Jo�R!4����j:b�o��rFP@o��c�������Aq�8�����C��`��AS�Ћ���{uKԄ��
kn�V�lF~���lrĻ|��"����p?kD��GM^g;��0�Sc�*U]������
��?�!~o1S񳠢�܊�b褹�?�5��q�+<E����Lq��t�{���bcL�N~�Ú�+�g�ڗ4^-��t�z�����d��Y�Ic�T�CB�L{p�y����L��qB��;����}�t�=�,�,r Ѷ�>�pu����38��A����E���j��T��yGX�Ot���4���/o`�����hr�Ez�{͛����58	ǶAV�i	��z���Xv�����M>t5�qRn����}3�a�}8�n��
�cպ�1�=�ܚ�]���F�	�d���&@0j9�q��f6D�������оe��Q9��7��bY�3�aWl�N�m�m}9����Ë� ��ܜ��)6��Gp��C�)8�)��2
G<7F��F4�}�S�?��<ZU��d�F�3nE�i�=&&����
�&�]�D��(�� XR�1eM����N��,���!]��o8�՜\���.�_cR+d�Ōa��r���l����H�����ա`qv��I�x@��|��%K���`��zT5y��Cy�g��x�G�sjaʤ@��ĺ�~m�=�id6M6!<��3�Bn�{Ӷ�X�Z� N��h�4�R�;�_S�V,��7��;!�qw`cY�*(�X�a|���U��_�d'^Y�s�5���P	&�+�� Gq������g%JY{hH=h]m�8S����M���ф׶)û!��R��.�Z\
a��ԍ�:r�4_HG�w�Џ�=<Hr�x���PGGxc�h��x�2PY�B�~̅�>��p��q#p��;V��Z�f�tz����P2�NP�q�B��^����nYZ3��n�X�j����$e�k'��!���:��"}x�Ű�'$܁��Vl����x��&�Y��Tɺ]�d����f��/U�+ۖ���e������Tj�Cտo˲���W�Ѧ.�W�HUͱ�s-���C=���;�9����9��bF#90��
v��n��`x{Ҍ��B'��8^����2}��0>4ӊ��!b���ϧz,w���
��珩����غZU��ە���J"����^�\�uw��At�����G*��4;��K��Ԯة,m� ��6$��f�M�Q���Y�.QJ_�т��2�r�����e�2TjQ������L��Mie�Pz�&,,̼τ�+8��/�P�o�d�(�/(/�n�vГ����ù}��q3��5*�2Ć�cQ�1}a���-i���A�����:�d˶ ��������:e�T뼷ERuj2�q��iI�gT��=�� ޘ���J�gQ9�{�U�7����W�	b���?��W���0^/�0�y�՟2 !��t-��g�*|:�u���?	��w���WqkKG�����y�W6rtL;B�.:��ѽ2bf1�s����&`��*�)]�V���O}�)�����Hm.��^�� ��)#��g��"�鑧}����,��.���N��-5���q}�0��K��P>���|��w��p�D䟞��6��2%u6΄a}��NB�Ɇ����:3�D�����mNI9�a1�om�ܱ�.:�\��g�a��/eŬ\R�-�1Cr�?}=�L��Q�B�����~�χӍ�4��B�x��� �U��U�^�r����;g�۰rP�oΟ���!�|eqL��C�	�Q��6.��=�Fj�dv�dN���4�W�nR�N�A	�!�ց]�F����D��+,���(����ix���|y����ٲ��2��� FF/�$.��οkd^uxwo��N��K;D�E��rI_hi������(��n���Ӑ�ڨ��l��%�P�k�j���C��B9����v������;��yY�������+�6����}���-�$U�Ѫ��r��n~O�נ)��|�A�V�P�6,������\mM_�ANRN�ኔ���D�d:B].%�cV�ɖ��!�U@"(9ɟ<0U�WZ?���sO��rwt>�?3�ػ��F$��d�~����Z���OD�/:ZB��'<��m�W�B`CG��J�ge���[i�d��t-Kc�C$G���d��Q��#���5i�x���m��Y��&��n����>�e� YK��;��+�0��^!���Ԟ	r����Q^a�|.���IZQF�N�YZ(�C�i'@E^AS<�?9������\��7�W�:¸i��(t~a\�/6R����颕����v+|����y[��o��z^�/���G1��/��n,ŭ�~g���a��.����\���j��}�r}���v�B|ָn1���|Uξ�"S�����\�u��yh��L��[�~��ǎ	K��'���oS+����M�U��I��ņ!��bEW��$�_-5d[�����bm�r/@�AO�TZ�!y�_c@e;��ԋ�iL,֝����7z-
t��ۂc\�祮S��ъ���S&Ə���H�_ȄQܪw�Z;�t�ֽ~���a?2u�UL���\������S�wj�F5!K��+j��`N�^V����Z������D�m%?�m��;�m��Mc�s���K,�ґ�v+!w��_���_v�>�d܊�l�"��+e���"+o):B�������ńf�����2����p�U�8{G�=�����2>.F٬{5��o-��cA���1 F���,�k�d���TL].��MHV�.�����4w��%����ˤ[H�*��"c2����[S�J��E�u�"n +S�v;SK��=,����i�����ѝ��c:����L^�1g��4scc�W�nM+�B�0P"��Z.d�ls����?��ʱ�w��na%�2��>���C;�}��7�z����8��ȣQ��:B���I�1�Cr;o�"A�"nZAE\�ƷMۚ�ږ'�nY˨9�/��܇�Z�4m?�%�,ޱ<q���&�*|M |���g,�9|�¶k�� m�l��T9���m�p���4�#��fH�j5h�l�n���l�2���9�#�*}�
�hnV�K����qN�un(JGY�8-�z̍gyG*���Hk!.�s%�'<��G�l���õ��n�MD׋�,t]��Ҵ�`�<S�!�m��y�ϋ�a�
�A�
��"�o=9�H����b��fz'a���J�����H��e�{�=�zȌ)� ����+Q8Pv��p�q��[����)���w�r�![�0zdv��ˀ'�;�%w2����*�!�v~PA�	P�+�Iq�@�2lb���5柦�s:��4A�ه���i�ϕ�{� 0�>h��Ab7i.^x�iX�i:��&�&C����m��s�atzl�u����J_B%�,�H���&�8�ԱN���={�*W��F:�#�\�?��&�oO�3&��n�9�h�9h�s�՛�$� N���dj�������-����������d�_��C�F�.� ؤ8��m��਀57�j�" �u��u�xh���0�C
b�4	�!q:Atؾ��F� &�F�p�&��^���w��;nb��}�tl�Dn�o������((�ıqSӃ0ǢS�ni_�(B"���?e8{AW\���� b��#�۟�(Y�	���LRm��v3�^}	�v�,�N���8��<A����h��ٱ�����w�L�
Xn�اbv<II�I���;�v�����\�<�=�o�K<�X�M*��ӥ���΄�V�HӼ�R%B�9��s	U�w�Q �]S5:<:c۷�p�5ظ��qIΒ(较$)�+��n����.ǉZ��tP�aR�=�\���W��m~ 2QMʾ���o{ϓ���(s��������������sՑ��L@���ˊf��g��Ԏ:�=��B{㻫��ӧ�[�����8.�y����K��=b������E38��s2�14?�]=lYX�z˼:|�2�y\�w�m!<MFE`+�E�>r6�evt4�g�v�{��S�v~h�P�R�;��^���"�����1p�X2}��5��ྊMl�����5*��l�6��%�ˇ2�y�%�죥��Z�@�������]��=��;E�Tt��� �m��&�D�w�Z��v����x6�e5�loTD��2�Ըɱ@���QC;o��� �5c�:�%k�F�"��/��H�5���1ub����v[_���ĝJ]n�tgr6M�D�Km�K��9St�d�,z_>x|�ԙ��Ύ7����g\rY�?��"]j�ƿ,m�A;�H;_.F�tխ��a����ط/n������A/7���@�&����7S����i���k��)M��W�	��^����W��\�fS&n�yn�߶۱���x�����3�6���X��-���������=���DY9���u����=����ȫ�i���j��ǧ���r�l'�����l��h��BSlq��� yW��c1��G}F���.N��4-`�N_4�ո�4=#륵������`��̬�������k��ܹ���b�V>���!~�\�t?�8��u,�A_�l�$��������6�=#]�n��)��bJ	�G(�������!8�U��b���h��S%�}	\�M��u]{����@�^�bj(�Cb�3 �1�|����_�]��
�b=��m�����Gi76���/L �n�"'b 2��>u���������i�?�"C�W�sR��ۤq����ӈ��p$��T#Af�K��G�me7C�Q��
�B��`ٲ��|��c�0��~�[6�0�7w(�(6��ʩ*���6���NcA?d|v�Q�NA���5 �����Wrf�1�ʤ�t[W�u���cM�B),�[tn R���tp���Ꙑ:,=�Ȳ~lp�f�d���B9�Q�^�d%�����5��=Ը�>`h-���A3�U����q�KcK�s��א�8Jk8F0�e�~;�����{�m�A�	��QN���Ic:�m҈ˍB�ȉ�DU���"�K6���
gbȷKן�-/�k���f7N�^>%%�_i�Mx}ˌI�MvM?=J�vC5JP&ɢ9gǧ�yD��LCME�P�9 ���k[�z/�z��%���.�<#�B�zRA��u_h��^GT�;� y����EiI=Q�o��X�u���|<�՜ ���.�m�#�07��J�99���oѳǳY3���nX�i�p.ն����kJ��#�*�v%~g�B�s�b�\�hC����z!B�LL[7.?���Lǅ/���bx�${\���P�V4�)/����
�B�|UA��
�� u�o:�?�>C�0��9���:/�O��=�eʵ=��5b��i&�{0<��gE���[��0�ND�Ȉ
?	g�L��/�����[I��5�u�A}��:�a%�.6�����RY/=d�1�*�=A��d�AJ
��V��e�<o�ҷ��P����n^�fe��;�aꤼ��n ��!���b 錡�)�|Hç
���۴wM�����X�a�)�u*/�!�w�����Nǖ�?��ߜ�k�#��w�Q'�L��1ʍo�{�[jEz�h9%ˈQ"R��왜���,�Y<�L�N�kp"���z^�ɻD�sU��k�?�ԫC�YY��(F[ƪ���@1������L�~�}hh��}G�{�>p�6�������q-7[��BH߂�����Su��N!"Mo������m���Wm\*I�(�Z��ȆTS�1��m������/��Py��paN�e��_Akl�I�"O�*�g�':����+9���{5 ��)-7l���6$�X�� �|��z��kڸX��dmZ�yvC!�_��c�^�C���+ٷK(�Ƽӕ߰?�hP�����{�-\MP��z�y�M��=�U�9���}����Ñ�(}B����u��XN��+
l�ˣ0���ϊ�O�)p���*�g�:ڄ��G&5��lU@�Û42�I���ܚ&�>4�x�3�����:;{%B�E϶moZ��[�-�w��D����q#�Q����z���-�g�]�2kM�:UX��,���$�:G0Iҝ�]Z�j�!141��R�lk�DfVx�{>��ã�C!��"t*�	�a<���06��
AP?e���'-�B�BDQ�����- ��4��r�Ao~�V28�5��s�ȵ|Gy�(q����^W��P���.&�frNa��5_J���q��hܞ;!��t�tp�]�O�+��	�H\�FNg$�d�VO�ʘ2�>l�û�G�4	�d�&J~�>n��_�h9P�����m����@_HZ�?��(���� 8��v>T�}W{��Y �$?t��옽-�va�Jw���6��&~����`��)2C���z?l�eZ��E#��F�p��tE�ꕏ�7����u[p�@���Z�lp3�F��s7���ܖ|�p�J���6̋����J�7Q�5_��q:К9C��z�Uׁ�fV1\~��������ȞہeccK�H�Ȁ}d����r�s$�Ě���w:z&�B�����]�}k�(gEpm����B�i�K��»F�Iy��cu�1��(B�	�ł\��QS�P	�H��O�
��vv�+�G�Cj���ȧ��;(��Z;5n���C�)[A��SB�{<`�������k:�ܐ����a��ag^���	cf�sn�h�FpQ�(�憳6�"���.�=��s�wr���z�Wo�y�D�a�U�2���4"Ox���ȧ�u��`ع���T-�saK��I���w5:��2ӣ�X��xjx�o�}��h���*�H��,j�N	��Gs}�dJi��z\��`!��"��#��Ð��1�*�q� �l�j��?V�ĮR�6@�c��M��Pc���g���w��_�S�g�	��'m�H��~.�`PK����R �+W(�.���Io��u�jvl7�m72�gE�'d(Bo+L��O3d���w���F+����Q�,j�P�y���"�'F 2�yz�	�e�����rT{m����3W� x�+ݡ!g&�^gRV=S߹i�V欀`>��ȧ�j��K�����ΧуfJ�<�Q�;��H�߂Kl�Y#�J�4�l1M�UqGD��ʢh���Ðt��y�� MՀ�Mҧ�xͣL��
s����%�m�li�f�
�́d�>��vz�]/���aK�(n��jz ݯ;��N^?�D��=C�7I�����>G���ye�9��oR���)��WݏP�S�Sz��gɥ*��/J����</X�_O� c�=e��M:u�"2�﷬�6C!�[4r�6����6�bxMF�!E鴇9[3����0:q3Ke���X�wR���E�)��f�ص�~����q���U�_cTI�C���y��"����Nmqjr�@Bχ)7� S�� �'�����\v/�w�h�VqI3_ǂ�(j/�u%��˖��T��3.����sMu��׍�A�ȇ�4>����� �T�=��)�e�K�K\��L�<h�P���I�u��C��<gF�GM�
����{�����A�{!����E�HnF�5�i| �����S�u�-)�y���ɿ�;B��`t�VJ����@^�J��e��Qa���V9v��gؿ��m);o:Jԣn�s���?q��� ;�p�`-���:o�
]4딄4-њ��|B����!S5m�j?4υ|Ck����[Rr���&S�[7��F��'S���>[h�y�}�x��X���(�י}�_!��S(z~���/X1hc}JG\z4��Zzh��]��OK ��nL#�yD/+K(��!RTw����g\�~h��4"s��-��Z��{�NT��~"a{�Q�}����N�EV:ŗ=Ӝ$f�5�S1���M�,�l�B�>���dJ�O EoUo����`�v溄8�7Me�P�*�^mIZ�B�X6;<rue���ɝWt{��kqb�	�	H�q�%׭*UPa\q�Dk G�����o�������xK�Yj���M8e���R���V��}X�>S��������C?�>�9;����(����P�?��4:`˘�*"�g>�
U�͍b-aݻ�!�k��L�wpx�b�9��3���������*D�g����/nf��[*F��(��V��X:�>>�&e��Vo�h�!�J�f{���*���|���);|�@m�N2���jn�%��V�!��#ǋ�,SFkt<��z
�������ҭ-&�W&*�J�L"�XL��8�sO)��F*c�-�Y�J.�������W~���?�����4�):a�A�w���K��r2$�v�zHݦ]�X�̾^5||�^,��.�����>�$�c���Գ�F�T��D}݉~l�_˓�k?sk�	>�9���Hb�p*��~_�a��<�e]EJ��0'�Rs��N�O�Lx��f�WHCo�H���c:��D���Z��P,�P�Y\�;%Mt��`�#����a{Ҽ���w+j��䑈�/�`<)v�Q�-!?.E��8��OW�pd�}�ݒd�r!\K�
���n�c�J�v2���%��Q�o�숾��Br�㟖��@�׹�Ur��0�"XElJ�b��GR�]S�u�?�h��L��M�Ky���)�p���;�D<�0=q~���n�g��
0�=^�-x2��0���yEj��Fщ�P��3�(k��qc�$B_�t3
V� y��&H�pyW��+�n_��2I�y�?1B>�X���:��
�:�� " Tfwdɚ#��'c�Ut�"�u��+Z���)j�3't9S_W����x��|5������fv��q'���U�m�k|��{�-�ю�.�H
w�~.D^����!P]�N�+/Ol/Gy�E{�D�!��G� �eP}y]�5�F��p���/�؟��x.TC���>>!���ւ��'zm����*�xِ.�L3V�����?�[�� Y�bǑ��RO-nFG���U���0�ɶW�o�d�p�Q�3	�A�5��Bl���Ɛ�������]�46,���]U��q�^"5t�l,Hq��<�4�ں>��m?�I.Ȭ���}ȿ:@�X"z�{�Bϖ�a�L�A�?k�����N�8+[w���@������Ùϰ�"XQ/��[�C��/�=�W��{�?U�J���(����j�I��U�"�=�)F��g�_�Ј���\�C��<گ�����(G>T�e�)��\V��;6�x3f�(>�ᙾ�%�~]�z>�����Q�u�1iøw��������;/��8����K��ٺ��Ǘ�byf�r�:H
����4�6���¦)�ς��qv�N�;�j���ɺ-O���Ӌ�&|b ߈��ΐ�q��L�o�}��;NCf�k�'RӳH�OOW�L}NI#�P�H=\�[R���)����1:�ݝ�>����g���L��sǦ���	�ǳ���&���q�|�*"|BT<.>D����㽽8o�ЫA��m�mJ4����w�d/;����m$RE�����2mȗ��4������}���@t�*��BEp D4�Ʃu�!B�Bތ^xN�OѭaѸ�+�����9�k{�Ż�����ѩ��[s'�Lɷ�&�Ro9��8�6O��M*�0P��@��;گ���D0����	�L0�5gIC��]��/�	4#�r���>sqd�������6{��j�	�|q�{r-�;*Ŷ���H�A!KC����d�ŹÀ�J�����8�V�4���z��	KESU� �i���~KR&+���|������@LxgU�o�z�o�Bd5F��MCU;���S?��j;+�$��ѫ��&H���Y[�����<,��:dA��R��ث[��]`��>g�M���ȑ�=v�����V6���?��-���-`�q��@����sQU�g)�J��"�i�ĥ��	O�`:��V���7����A��|&�6�]j9��`�114=��� ��śԸ�)[��.�Q��G���4`X��m��A	�Ӗ��@�L֮�="�sIw�i�a(��udJ�zH������m_���M���;�C��S�'ȽĘ��{�@G�U%M�����o�!���#� �Y��M����*�y�T��;٢�3�̝YS��	Dr�NN8@l�Sa��|��l���$ϋU���E\?F�O�$[$�q����Ș���W�O�;��DM
��/=ZO�������Uv�Ȩ���HZR���%؛�&�� �T�6�S�a�i�e����`z@���I�Ɇ�{Z�<�W��|��>Ũ���~�ֺ��c�Y��("�HL�N@���$ԭ��D�.UM�1E�>D���C?E̠Y5��Y�x⪷qC�rJ=�'�]	�F��H
zV��C�2J��f?����"ĥ�}[h��c�q��F��l\'1�J��9Ò镇"�	�hV/$d����ôe�o=F�����5Hf%Y���J�` ����` ��Ir�.i;RM���`"l6?\�&�6�h�d��	�|^��]�V���q���6��	�x��"��Q���� C1�	�$���/iudt p���j+�="�-�is�m���f�Yߩ��85@\,�e[n����-�Ya��-V�Qe�>�r]P!v�)I6�!8D��h�L��[Ê�$����GE�Y��{�R뤧�yH��uQ)n9� �[UMzu�U,K��9�Hn��ͺ�M�����1+Q>��OCwl�v'"*M�X�<�#�`��h>�.QΚ$p�Ɓ��J��yF����G�o#1ud!�4~B��9��F�z�v�s�5VgS��C��{������?�m��lBRH#T���[��f��c�����?Q�r��u{��B11���}��Ui1)������~���cs�+�+?݂��
`"j���p����L�����������[�`�	|KO��Pt&�\�i ��(aa�	ǳ!I9�s��g��b��d;��C'4W�"s���\�ϸ��l�;㬟�R�Ai�$�b��3�@��K&�r9����=��|��f��~�>o����@C���P��<��`j?�bp�	3{�5���tV�QO��@|�NT]9��{�)����6��)mѤ%1r#r4,�9��]��ܰ����hb��[飸O����!8/�<)�oR�k���ȿ_�>Z#�R��,,T�n��=� �/`�B
 4��@X�jLH�F�d¤75��}6�;C<k�_)���/rѮ�C���<���{f��M�	�/i��M��-�7M`C��)�]x����#�6�ĸ@#�l�W'�M��e�_���*�L4-�V���i*����{K��˹SƳ1-��5�T��,�'��A֮��OE�Ũ�m�vPm9�\B�^M�z,y�:��,U��`��� ��.�[�^�%���_�h&f�!��ɸЏ r��0	ژ�->�Ǿ�8��fll��	��<�����|�@7o�q5Grr6:���YO_�๘�{v,��ۯ�	�f��(�H�V�2� ���ko*�S(Ӈd�F1{�l$?a�������tN���_,��Q��}�:�S��7�aTg�X�w���}e�P��L�>��(m�����MgЕrG���A��v��E)-�>W׎k��;����%����E�wiCT�YK�]��_��u�,��V�q��;H�RC�k����CB;�X��w ��x��� �@{�#g>X��]Bn��Z�]LEh����.Ca��} @ӡ�@���;$�S\l���
�VJZ�*�"â���[l,3Q7 ����� @��l-e<�1��ѧX4ܬ��3���h��Ž�j��W�Bc�XQ-1k�P��M�����X̡ ����=�i�	��q\��Gaҫɘ��_qXF�U*;m�أ#�3n��	m5��uN3L�E�T���U�Ǹ�y�U���N��V���ʹG�C�$�Sd�����xb������3�b?�e-\O�rW)���,����V�"!Vkn�f|��Cm`�ՏP�1[N�.{ ^��{�fx�H=+9��;��4���z�ካ?s����G[6��u!]��QR�!�"p��'^
���(o
1��G�����M�#����͇
�_�����M)���B.��C<3�M��1n�H��.O�f�(h��z�x7���)~a Z*cHr����6 �G,�<ٵM�!3D򽊔�Ä�:�U�*U p֪<��aEQ�[ ����@3���ܹN�w=���G�1�Q-}~�h� "��
l�#|D� ��<_�`ɐ:��c��*�3ճ]o[4�H�_��l�5�0M!�q��6N���޴F�	����ֵ����7�1�����}�����:��j����}�:ƹݽ��,L�*��������%]y��*/��b�>�4V���ɾܥ��DuV�	A�L�˷*O4f��J4�5��+.0�2��tv`���\��ـHR ��8I1���2E�ږ���y�@�DS�� `md��<��w��&ZMI�E��,�=Z�u�|	?M� fLP P?�Ѧ���3�J�=�"pCv)���ҥ��Y|߬E���9$��"�<����@I���x�������=�˩8<���:�U� %��l+��&҉o�ݘN��TzRկ�4��%R
w< �S �!F�	����}�.�q����w/���M��.*&�EWܸ�w6j���e���Tۿ$(��TX���{ӫ�K��C2d�(-����a���C��C�@\���!k��O�t�q�R�tFJ]xh�;�(�ܡ�����}W���.)����~�^�2h��;��o�_�ovGS���`�/#��u=$U_p �ng��(�8�mKO���1b~f�&U�w�-���A�ɑ����嚟r$�TW��=j�I�fˉ��L�~W��q4V���.�)獜}��~�}>�j��8EF�R�]�p��6q����ܧ��o�ɗ�Dϔwa��g1}���D��Е�I7�O"�J�Y���<춈�n��*��Ƌ*`� ��:sw�^�@/FXcR��.����[��x���R���F��@+�+J>���+0�zW��7)A�l�69��8������sK�q��P��r�s\;ךj����rC=�c\6or;}F��3�:��Y�t������S���e��� �7��-�":��ώ��IBM��D��N�nm;KíPw;Z�T��y�����>m���J�?۔zM6Vv]6d?\~ ZlF�=k���P=�K�)����	� i��@��@+ﭽ�����F��o�"�£��"�P�f�6��@6]k��ow �ak�%9:Q�V��s�/�l{�"�&*e],�8�*�q��P�1����^yi �u�/���;~5a�Ĕ�>��l���( ��X�R�p;�x�[�-CGj�eG�άՠ8�l�\Y6���QN�m�_>��5���O���\���7E�
�H�A���Z��[�U{-�zF��^\r\�<��	'o��i2�~�6%�pV'�JGp�^�A(�;��l���1��9,Em�B4��K�	u�3M?+?�T賑-h���2�%T.F`��?O����.�̓���B���<�d���e�2e�%#���e�+���)�?�P���j��+���ݲ�_��J�|�r�N�ԃp
g�4X��H@��4���Lb�������,�',j�CwpA�ǉ���qv%�ie�-�fh����g7��y�@���D|��tѴ�7B[�|7c��c�JJ��z��l�qˑA~�}{���3����+�2�f���?VV�� �3�z +�m֛�~h/e3G0�	ܦ���{Nj�4jb����SH������C@�\����d1R����u�<����J i��Y�|h��XǍ� ����c��.ݖ:�Qd(�p㇖u� ����G���ʖ��H���v/0w�2�x�~���Q�G�vqNP����O�}�S4�%R����;�^Exy:T���CJ�w}A����,]���+���%���B�,��@���D��#yMDJ�2E��bܘ��b�3�Č���>Tm�%�mXQVcۤ��5�~�^ۈ�dm���I��LȢ�Q|ئ�|��|��pp{��)�}51lh!3ȊU�h�M���Z�;��(�\�M�gH#�b6�Um���WR|.��~�D�my��8�0��w��U��6��uc����6i�D
C=���H����+-���������v�=61���̊��W�m�P�iH]nW�X�ͅ�R�&�B:�R��=�ip}����$��Mn�A"���3Y�ڻP ���mAPV�} ���O��B<�����Y��&d�/��[E�����	,� =ʑN�	�fq�T�w;��v.�Bv�A�h�d$G���O^G��5������pr�G��!�c�K��৕�r� �3��fT%��u=��֣E�6 �8r��p6���+�uA�������tD�8��M�U��3����@���V,,����6*r�"|��A���${����C�V��7T�tˆ�RnPQ?Bׇ��>�B	 �h��H��D1ɋSǦI�V�E2Վ��j���3�Ax`�� �~�����c�{�M��LR1�[�R���)'yc��s~�������.�ץ���Kp]�i��f@U� ){����S�%���4&�*�,k�m�1y4^}:�.�^`�� 3�8��9��[�4���i<�sO������Y�f6Nk�l�ĵ�Lf��r��A5� 1��vX҅2�UY��_ �a�~߾���"WV��!�����V$C�����H�8���]Mx�:^=�$r�,� �8U�szo����4Q��xK�qB�<H�����+
*M�B�+��\f��*\c���QNB�N<��*��o�Q/�Ͷ�z��80d������	&��%����I[z�$�{7d�W��&nfx�LA�5�OO��3j�� �tR ��pQ�C�.���2%��"�#=�&T9X�!�G�����RR2��G��e�433&>��l�)oy���?�0ݳ�ɉ�:RC/~�Gk����A�P�;� >Ba��NB�o]�U@S�Xbm��A/��ó���st~��,�~�o�^M���gp�ya��ܚ�jr�4}���_Eb���mָ��k����< ;���*�`�Vm����~&�F��b������/��`i�# C
7H��f���@�~<�d0!˚a�H�����K�}`q��r�|���9���6	��Ɋk3g�F��;fas�Ơ�=���l����gS}F_�2ߞ��J`Ө�f�a>Y�Xo.A��i�
�����)�J@�`�ٛGY���zem�!�t$H��6��(V��f,}���+����:2�� ���ʥ	V|\>Rk��v��0��F���Qե+���/E,��� *�$]]ե�AQ ρ<u��t�z�.�U�{��pQ(	���Z�5$��2�%�(s�B �
iu�^	�ak� [��{�g�i������?���>�z_�`0>kc�>�k���>��膫������ތt��+�n�^�
f�T�8N�M}�2
3�5u�Ze�N��ͺ���FP�J�厛�gLLf4��2�Ŷ3p���`	x�'!z^p/�D@���O�^'{�A6�d-e~�V:L�$�W����_������c$��!t����~�����1/Y^Uc�`h���4�֑C���?�s����1L�k�B' �N��ţpX��XBߘ���jOn��g��R�T%;�_U\w�k�Hi���h ��u�حY�ꚽ�U$��fͧ.ֿn����%���?�¬�6����閕MJ��/�:��e�R��i��7@u3�§�7&�%Կ9;q��P�F��H�~D���jCC�/��"-/s;3�E�� e���s�
�4�2HF�