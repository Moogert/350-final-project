��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g������*���Li�ĉ�3���R�\��0}��N��i�b�QO3s��N��㐝p�W ��Kl]���BI숹�(�a$����=ZA��Z��<e�TrRd���t�o#��K7�QX3��O���� eT�2j�Ŝ�5�| ҭ��\���I$��Ng��^�i�cۣ
,�P\��B:�CN� z���� ��hc��GB	:b�[�5Rf���il��.Q��</4X <�Z*�Zv[Sr�w�P�����˘��C��\&�η��zR��bA�AE�Y�w��\�7¿ȣ���p�A
 I�!�C�^�@��r�>��+�5I�Y>?�A�����x)��a&U.�2����]L��^��Ȇ�{L�I4"���$���$�+�<ĥ�$�?LM`!��U6I��"�<�S�e�{܅��V���r��N����{���NdG����ğ\r;�ې<ɞ�iB�]�Gy�h��1����S�|�Qf��:�=����f;+�*_g��~0���N
�Z��9��ZUĔ���C�س�IBT�}O��֕�ϖߧ��B�{�ԗ5�9�幵?�.���U��}!GR�!=k�??l���@��M���U��_68_�Z�t���^x婋^�=)f}x,-~��Δ�p�a\e8#h��J٠6�]����ղ����y'Tp/vT8BQ���4 �� �ȱi��ʳ�q:Kи,K6�y4E�oHn�YS��l�����������A��5&QY���\y�G���b�z�������6y<�B��iIZ�?Հ��X0���dx*�,�Ÿ �bb��K��
��p���@vC�v�Tu��Ю�Ӎ�)�5���T�#�1|(&*���^V%�=&����D>��G��V��*c�����T�шy�9C̓wW-�\��)b&�w�,k$�]՘���
k:+������E�7Y��0�zo0>Ƈ�E1�S�������|��#���&��Qn�C1�iw�t�U<@��ܾCU�Ej���L�!��@^.&;M ��)�qBg\{N�%�������p9���/#��\�ު�5<j�u}^����^>*��"X�����)g
�xcmhz/�s") _��ӃLz<f4���<<#H��w�`ƚ�^�r��V����X��5�1\g?�@��N-�
��j2|����5�/���s�<� �w���]��`�]�V9d(�p�12��D��Ê��`�g^����N#xF�B�C�T��yc\� 14v���[����4*������E)q�41J��TC&^�*I��� �D;fz�?W&��?$�X,8��F)�bJ�������jʔ�hʤ�ݩm�L�S6妖�	�>��?���G�βU�[
��)�m�����C_�����M�q��9��7��o�" �抢�ɕ8�JE��؀jz�b�3���X%ř�U�v&e
A�5%k��A��Z���9�]0|��أs۩Yv�	 2B�3ǰ��.2��X���`fxq9.��*����eq���%c��^��i��$*��	"��N����^���E<����
`:��t����<���aΜuz��~[���\tA�?x�O�]�չ�M�FB�>܁!KR�P^����82���Y�P�=���mĳo3�Fh���V�g���i�+)�L*rh:󎦊HDYh �T��M��	_o�`�0dTB�y�`���<����:�Pc>V�J�~&{<2����10�1福)���޷�I���ҕp9���	�q�|�߿*-�q����9W��>InTN��k##_5�����D[�ޖ��� Lf�V�T�Kg��#W�w����J���s�y��r��f�9�W�1k}?-`��Bͫ<�0#��X��Sj&�&��� AL<���3+Pӥ��4�c���p�T��c�����j�ն�3I*��f��Ȥ؈�T}訏J����Q^\�y!f�]� �>뤳*g��$��h<O�f��jJڣ?f�*�Ӊ��bԆ���	\cOM��!&=񘥮�!b���7ex�I�l�;�8�iX):��Gĭ%���� Bf���H9ʹ��d]���!���k�c���d,5R��8��\�aN�1�"�؀�o������wH�򈍱��1�*ܨ�ny{7�4;�/pz� 1��ǕU��fn��.�g�� 1Ë�=j�-xe�c\z��k������6���ti���#��W*��"TP��e+E��*�ڽC.���^�:�wS����l�~�Z���Å�0�aUu*#�����~���-ҎO�n��ղ��?����	����B�1�
W2;�W�6֋�ͨ]�9��aug�z�+"1���b�W�0���<�W���:�	V���x�N��,��
����N'���uT��z��)xQ���ڛ/Ɏ~��_ƨ�jAUJܓ�zd�5I�|%�ۓo��Ы��Ϛ�1P.�JT=H ��Rٕ[P��$�������H���8�`�2�v��d+>�� �΃F�y��>gZv�<�(�����H�c��M�[�b��&$@%�}��5���Np9"(�s!F��S��A9�[7�!���}i�dz���u�.�0L(�-�T���l+tǥ9�΢Ԍ�XS��R����;_�t�IQ��=2ņ�S�ot�^���ɡ#{�_��s�ug������2ʳI!J�,S��=�����
�P#�͖i2�$��\�ƨC �͟�޷�h��6�J� ����]��8����~<�
T��$*p���7a#��@�Mwt���t#���1ƒ��Pl��-=�5l�<�9#3'C~TPF*��0���$(�xG�>wO����!m�}�{���B p�=e���2kT�"E���Z�� cܡ]�}�J!^N��V�6�f#Hd����Vi���0�T��lS��f�B��������G#��t��^P]!mԗ�y6~�;���ί]u��6K�ձ��Z�L_\G�k*4�R$�D��A;B��g	�N9����n�����7�PnN�����힒�%��,�W�|����� �2���
�\cN�����Қ�+鸝�sP!�|m[a?OE��܄�8oMhn����O �I��١������P1!$Y��C�t~��P���TCN�g��̦��|�!���js��\�6����Q����T�(�7;��=/���J�E	���yc� ٣7��?�:�E�ىKJ�-�	��
P�d�j�~�Ҳ.y�ٳ�x���ޯ��ϙ�!Ў{O�-d!��o���
٤)8���ǆEX������OOc�ā.����ql�������9�sP�Gg� �qw0�;����_�F�o��|���G���:ᓛ�2�t�+�V�����]�i��*?�w�]ߣ���8�Y�M�E��4�V3��oJM'�UA>��3gU'��XHo|�*��Q
�7�OI��¬��s;i[�U�#B���� �6U��X�̝kC���L:�E��p�b�t�<���U�\�E�![���_�G�ltuA
�k��w�D���G�juR��Ç���a_J�e�5:d6>~/әH��E3�K��^=�:y� W[�xh���`<�U)�%-6�,�n֤��0�/��.K�C_��.WWj����b��BDx��-~A�$���Q�*G��b�`�#B�-���IG�AV#�z9멼��@�2U�3��: ~p�_'�R�p�*R���>�i:!��HiУ~��126Rl�4|���<�R�w�a֙����η�����8�Q����
R�4b���iy5=v��{�B���W������x�3��.�O�7dTtHk��m9n�zz����]�k���9_�=�d���7.h��G[��~3�9�����wL�ٱd�_볦x��l��8�\�*:�L|`)F�yħ/3��}�݁�u��/vjS�^Vҳ�D2<�q�<�n��UF�T�Q�.��/9rz�1���|�-��aT־��\���w>�2����>�i{*b��
#姓��IU�w�i+s��f�+}�Zj��y~ͦ���Zu�-�&�Bw=�jW��� ���:��!��z����GS�Y��?Y���8����K�]�(��Ĩ��5:��RǦ�X�����4br2vY�F��{(��u����B ��G�[P1+ۉ�(�yN|j^X��#WAP�c|p��5n_U��g��)<D�PO^�gF�(�6#uuw���8Gs�w���ц�/��� ҟ�WOv�fF"v�:���*=�w`"�R l^?�N;�҈��p]MV�i��84�)���\V�S��:�S�_�ُ��>��4��6W�
�e��� �8�g��iJ�2��L|q+�)M�5m��S��g�R}�Z(�5TQ�A�|���-�Y�mE^�ۥ|��q붭ʽ^���ƴ�����naL���G-�A�M �AIQhխ�~���_��-yY�" g^zABP7u3��lUc|����ϞY���/�!��f<S�:Z��e�|	��\��~q�4:<�s{���ϯD�G]2J�rW!՜pS�|��U+sJ5��z�@��H��AC�m�:�o���j�����B_�ebj�F����'R���<*��3_˽�'�n��j|j�$T*q#B�}����*��MN��)���[-�j&�~��P�X���?��{�|K�ż*˹0rb����8��t��AL�z7K۫������j�mPwj�Q \�<�v=V�s^�s�)�|e�t�	f3��E���WŰPf�ڗlOK��H����\4Q<)�/����I�eP���Th�ͦZ�-��BPD�_B�ˇY4f"��f�;Hŏf���Ȉ�qe�{�V�'
w�M������xI��Vg�U��e-���T�ʯ[�W���C~�Xε���aw�mp�x�^���r�����1EET�ר�W�_����\�׃����I��>d��g��[(�#��մ���� U�Q@[zb���=QģTk�!O��L�̂��n��p:�>�� ���-އ���b����2ˌ;�J��U.��r�Y"�nexA��\/���:��o���`K~!(���m�&i�@Fq�#`n��eE�"�c	UZ�o�s��>u0�RX��;���v�؏���������A*��\p{��p���K(-�`����o#4�F
�����#i�z_[���:.��w7PҝCI���x��Vq��%��y4Ϊ�l.K0O�R<:�j�DL���K�`8�z���s�N����3%�e�l�����`�^Ņ	�k'�D�q��i���H�մmZ��h���Z�����5���Fs�(�׉RW�-y/#���yI%��ztɁ-�C!���etB�'�W/0�X4�N�K�h���4jY"US����ZP��'�d\';����}f��rJ3�*��f��;NV��gC��<T��,0�����|���u֡��V���
/�	Uu���#w� �S#�&W�"�+�����\0��Yet���=�K��.F!O%L�M��u�'��c���Ā�%�/�HJ�f]q���y���S���E'����a�"�<��M�u=�ӡ�����W��ޗ�6�0��!BH�6��p��b7NT�l0C��$1��;� O���#���r<F�Sz��cVZ�_��B귪,�d7�S8|y�����]@�:��x[9��A¦��{7lf�à�F�Ga5H��*�;"��vNE&�=L�uN�o�띓`,�J�Cy"��΋4(��b��,G�a��0k��[i��T�w7�ĹT�oA���=~0p����ɏ�`,S���|�O�sޣ�Μ��j(0ˎ��'���}1p��ܩ�+ӂ�<0M����6��-��u�82��Ef�����\�V,����N��q%�k_��[w��ʮ~�N�E�9.�2�'���������7[d�#y0;��������m[�}����=�.��3	���
��[��D凒�I(�c� ���>��:��!�,4"x+���-�|�V���Lk>ʠ�Ǡz1�r���Z�0����{�&�J�{��Kb:����]H۝���YM��F	�o�!&��B<�����縉��S��u�lb���.�l��}��3��.ַ(lE�i�H�_��H�Rc����W�Z�F�e��jf��d~��,�vv�}U�p�T��#�P�n
(R�
֤�TR�:��6�=�>hqy=�h�i ��t�����(J<q��-!Q���CDc+^��j�m�Jwi����nќ��Q���ne$�ùv����f攥r������̕	�N\�E�mP�L��SM鉁>�<��m^e��M�N����F�Z��YExv�Ҿ� +���oaQ�eډ�>�cӎ�ub^��2��YJ��%_���)<9�ؙ�i	����e��J�������V��I&ؼ)�@zbA��p��~<�Z���"_R�+aX�U]�T�� ���n��N[`-��#�����I�a��__@�:�h�Q�3.�S�c/��}���w���^���oіi.�A��oD �N;��,|����x�.��Q̬L�����L ��^�F�Z{�#�Ibn��b�	o��� S��Z)��5WNa8x՞袧�D�sǃ�d��bG+�	����D��s�a�[�\��1NTqp/������]OoV������� �G7�E�����d�5/FVZ�<�+���f�J-X�$���l�3^�J��Ca�4�ݒOﲬ�}l1������kГܶУ���:`��i䗏�t�X����V7�Ij���B�ݮ�F�\� (+Vb������Na�F��䌤�j:G���3��L��T`tQ����/�=�_�`�j=P���=/��|r8�,��)0��/���"��PO�֊��a�V�������ý{��l{�2��z���A줙r-� ����x!&(�G�I�L$>���鏈��u���3B�i,'*���D(W0.M{��"�̐�c>ҋ,�k���"�ۦ�*��`�[~ҿK�ϡ�`��X���5	h����x���j����2�`> 67 	[ņ�E��cU�K6��0{���gߵ-�Ap}�2����jǹM�����d�`t�[G�#���S��N�΢�-H��«r�ԉ�Ӗ�@B�[!yyV���v����N��*1II����φ4�tA�*��n��r%q˝�շ�/�B���6��\�K4��X*zIT@*�$��	Ӽک����]ER�Q�5��w�[��@>B��a�\h%@G�2'`L�Q�#r��:Y�d� �fz�`�rL��L�e9��e��Q�ܞ}v�1L[�ތ����������d�+�}�J,m^O��F��ʁA��&��M��Iz���bjn|�T�5���9%�D���G2�S� X;h�	5��($N!��/�O�����!o#��Z[�	�:�i�@͔����)�@F��D�	�3�Qz��~��8A�_u7��J�8�.� �W�˛|O�����Rʾ�+\q�D,�;��K+����!�hWW�99�(�����i0yDO��d��X�/~m�oJ%�����Z��H��♒�ī��AM���Bx֯=�WC|�L��e�����
EC�F�ͅ���Ɗ���'�)/�I������EQ9��� ?�]m�_��p���5�(�o�jd�s�:�"�U)8t�,3�@�䌖GG��������z��d{���Iz��*�.q8����6YO-���c�x
?�Y�9Z���]��{U@� �RD��:���L��?��inq=�ǹZ]g����(/vÜv�:g��D��<	r)��I��	I��$���}�In�.T���Ʋ뵜�6�7��2��zV{=eT�8G����{�J}�*��RV���tÔA����]B�(�ZF'�"�C�E_���?��y�H��Nץ@�R���� ���������.X��\tZGķ"�p��.���}��d����Uk�z-�F�L�1E����i�l���^~	�S��� �cb@f�(x[�}��'��"��*�f^�'���[�/��([�*M��VJ!٬w�F��;S�x_>{S��C% 5�O���s\4 Zss��Ow��u䘆��Mt�'�;G]R>[X������Yy���k�zS�Ӯ�%n;Ɵ|GP�����(gm��8-f+n��S�*j$j��_�
Z��/��$�2�d�K���D�������E�r��j�N4�w���x­n֡5�����8��$���8�����D�3����sP���c~8��͊vK�4�Ly=h�;��9R;�މr��U�ݤ��g7��J^B������BQ�ה�}��ɇ�7�Zb''�:n-��`��G�gN>�##3�@���0���
#>�Sg|2B�y�jg����q�dI���(���7ɍ�=�����vm��8��E���J�Qi���P��}p$��]Pu����=�#��j�㦅WG�:on�>8�a��'�(�x$j�l��4��ʁ�Q,���O$���}j��"?�G�h传�����$�)"�0i*��?az�sL���Z��AZ�%���� �n*2�8S+ ����i�/��0ՎTϴu_�����U���4pM�/�Z4>V�i�욉/�9�B�[��D�mH�d�����k4�����i�$�g�~�=�%�7��%���ⷲ�*]�R�R��dNt��le]�a������&F����@���=�$0!������cQ�p�WNS^nc�f^��Ɵ6���P�l�||���Dse�K���{T��|���r?��߰�J�!����P�z�Lv����}�l��괸�"`��[4��]�R}t Q��ا;��ZF�!�a>ы��
|��Y$���<X��L��`�5��X2	/峓�B�������I�Z���ȹ�3'i����+�Ҳɭ�T�����\�12x�p���0�z�f�j�A���(.7�{�v�Q���qw`x`1X�taGe�D��C_�P�}��=����*�J��D�2�Յ�o2�L*�n�}�^sI����R����d�$�?�o�	�a\��b<'���o[�#� :����R�E2�IF��j��]�������I_��ÒC�F���D��)OR��b&�@��	vʺ�<��Y������RR�	#%�j�yg��H��Y�g=z�����M��J[N�\�J�F�<�G#�"����]�%�e��m�P��G�\V�r���þ�Ô>N�4����k;�����i���ɰul]M�{HAMR�����)Գ�YM	K��ݍW8���g}���w?E�T�*l����_)M�C�1�*N��z5�ɿ��%Š�^A�Mj˪ЊУ�ǹ�L�����7V]�3c.�Uu@0fՈo���wS/V��n��"��L���9��J�l����r�.�.�\�W�t�4?����baS��������Y)�0�^���/egB[��d���T�59�w����ϳ�z_��ų��5-�C 94)%Q��;�ve���]�or�O�� ]v<zM(�XE�e%����%��o	,��)�?���1�����G5q���Ye'O�B��ߨ� 	���`&T�X�G��|�x�U0
_GK��]�X�� q�2�k�V!��C�r��B����2��@H�Fc�ī2jT��7f�R�u�
��(ş�H��"��à}��N��c4���@�AN[�q(��˚��+��<��m(���K�zu�25F��^�aL��k=hb�}�ߩq�=8B�H�k̒r��`�����:�z^�@	Ls�	jM"�yi猵:bb�/^���Ç��u`��A(�}2�C�na1������
��o!8G�|FyJ2�
"�Th�.�͉���ٝ�(������#���q~���b�Lg9��»������\$�� bw���Ԁ�%*Ӎ�Ҳ��β�T�C�l��8hQ��>���Ư~9�F�{��=��X#x�(�CG��G��T�3�w,t���0��	����۵���ux�66U������a��aH/�Ni_ueͨS�k�(�@q�,X}�%f���R���8��^�CO�E�G� �U ��T���e�_�'R�4��Q���q��Æ�ut\�ޫ����<�O�p�SLr�Y�_^J�<���ee!UΔ"x�f�sH$��*2%4�(�6]Dg���F�G��v�r�sAV�0���%��N���uteA�[�P7��r��}�5�6t<8�pLm���y��X0�1��x�$��ڞ��$ �Z=lC;��@�N��ϖ��D܀��m�>��Z�;J��d���	�3�
b��K��f��I-��h���y+�X�6�W�t=c"�u�'#�������w��]G�!��[F�$�f%�mש�c����C�"��_�5#Cs~��D7Y+u�'��ڨ���8�~)�` 	!G�J�Tz�N�<��>��o�B`��N}>��&�("�l?�F�+ Iƺ�7Xf�ݑ��U�tX�%f���"m���g6��M`�Wr�X��R�p(MxFK���wڌ0��Y"��EDb:����G�:U6g�+��@��P���=���K��	��D-���l�|�NJ>�"qc%Z(F�ѷ �kN5\7����oc��~,Y������u�:˻��b�·X���~k��خ����\$㊯;P��t�2�E W�����އ��d����y	Z/{�N�5�c�W6�e�s��������<Y\�Rb`dPT����){��g���һ��b���c|-����ʰ�X��}D��$��GO���o��V��%��q����b��C���2�`����B1#�tf5^HD�9��۞g��ی�~Trh�	?-=X
M���)�������.U�o"��d��_�Olz��ʠ����S[b�3��㉻AR�}.5�6^�Y���o�WRo�(�C�b����]+�Vs@V�%����]�(�D���\ �JJj�m��U�/��l��X�pF��/&G��IY4�P��i����:��� ���w�r�'�.��˖��I7����X��ӭ���,	vt �]�j�����z63�5��z�׽���+o�_5y��I��m��i[<w������i�F���9ʔy�Fj�ud"�D���ll&]��x?˃�j�0~�U���� M1�Z섈VCZ�Ϥ8ɸrZwM�_���$�h�V4ny{" F"a�$}Vܻ�r�S��e�����h�(`F:
����!i$~H����A��yYE�$��c��cH=���g���6g�bG}f~b9%��%��E���52#���|?�8 e�+��/8m0�m7�[�c��X}x�;�*X�+��gJP�)�����JA<rl�E3�Yx'���o�~�[�������h���f��m��Mk��b:���K����(�%Vs�*�a:|S?A�_1��$yF�|ɸ*=�7UX1�v��kaȥ1���w2˟	O����~�Ds���Y�V�dG~�FD6)W����x��\�e�*�����0`������Q���t�/:"ݭ�T�ş ĘD��>Wx�K?S�28��2���*گ��hB�Î�����g����<M�>��r���+���7`lm��$���Z7�;u���N�\ԾY=��r�5!fN��q�46���\������ⅶ��|r�p��V4i��E���_>ڣT����sZ&����:kj�v&+�BAOm�6E� >�Q8�n�/>S�w��#��=X�����ڜR�TBT����0�7��9y0�ne�l_g��`�����a�g:<Z�R*�����TL�߇{�ŉ��h�p@��$<I3}�U�q�|�BmUtS�f�Ħ�ٞާhEk�_�`S��A"�pc�X51��ðٶqQ<[:WH����-s���&Vz4lN�XN�̣������Q�0�X���ɼGq�~FM*|��|.ͶX�z_����#��4bD"�#л��U�|�y��rmni�E�:�^o @�ރu-����N�rYLn
�>!?E������'�t��'�/�9;f������=��7n�Z䊴�`y�s���)���i����YR�(��^jf̊]��~DÐ�{9��8�+�Č<��N�/5y�յ��
�;2�8",Y��kK�z�}=Ca���Eux���TIU�[T��b���f�o�߶R_�(�ϲ�%���=|f�؜.�Y�?���Q��˜|[=	4�q\jHp�[O} �V���c��0kӬQ@�h�c@����v���8����-��͢׆��䒖bT/9��H3�7H7��?C#k��2 g$�G�vE���q{璩��Q�gQ�U����d�m�5�-�x��s�F!�uP��s�eӭｑ4�
H��Mq��o³��yIͦIi3����%�r���n?�~F�1-�%���E�*I3T��J���9�֐�Ft�)3�� ��<���'�y� �;p41���y������&ҕ��x�8�W
�u�K9NM�XY�ԫ����M.o��"=�Q2uxd�T��>)�Q?Ü�zfA�W�hn�D�I��nӝ5����|��qoQ����ǃ��Ҩ]�G�U�X�I���mE�_��SYn��W���*W3.?[*�,
</�l��L,�9E�&7B�\��z����[$�jTnJ
���I/Y��7�ԍs�G���?H����ɶ���ٌ#��m��K�����z�� �m8=�L���$d��Bg�*,�\*���I����xG��k'�d���e���yToI�T�Y)���)��^��gM����,x��o��G3�p��lද���o�� +sx����׷�PY�%1�&�^K�x���q%k�h��ڟ���_� �&R����E���Ӳ���������ϩn.T�c�k�*�2^i�7M�~A�5P�Me���'������f_�r�O���(E�}��F�ڡ�w��f��Un�(��Lwnt{���0�Vz,%������V�<�VCb�c{��m��>��w��2Ǫ�!RH���Qp�Fmq����ia�M���ڮ�ˬ?=�W��8XV�ԻXK�W�0%:��ÆS��0��̒|5T��Ce*0�A}������G�����]��U�*�$/��.s��`#�'8܃V���F{y��w�f�V�/��E��@�؞����/.8�*�z��(�}Uo#ܲ�U�46�F���9T���w��	�)A�� ���Oa/g�]y<��@W���U��y�Ul}�hC����b�ǤN'�N^��RE�����{��S�-+>󐙛*�-���Ј�[�t��yeןdp��4�l�����I`��4|o��=�:ǔࢪ^&����՟��P�T}�QDIo�����É:��Zd�b!p%�#K�~��_�4�'�">j�t �}�j�hD�������R��@��	����F�ڎ�a��uL}�VM��e��Az��ݩS׎�i��k��[�����m��I4�L
a{�m�M��F@.~��"����;��qFMZ@���J��࿅�k��v�<�����\�eǍI��<� Uk��T~�0��E\.�cOgv��u�)��d���<)d��lOXTM�����ZK����+"�6��H�d��\��X1��#Lx"A�Ĝ��S��7�����ܐ�-l	�d���X��O��R6�aln�hw�Xl7�[-@L.?��*Ϲ72A&܍��;_x9=�P��ح2 N^S�P�[W�Y$�ʇ :W@�����\v�����@���%�]���ǵ��g"��C�#W�X��J�'1�ZW�n��.O�/P&����_�/�-�vJ��t!�{��(�=�.3y�=��)��+������J��U��?�%��,��É�h˛1���B��<��;>�� �eARC�����zF\�'@���iz�"���Y�n~M�c����a�we����̡o�>�VO��Al�=�����}���P�ʊ�1#��V�����S��*�x�hP1�6Cc�Z���$�����b�Ë�ʜp��L����$�s?�'8]�Ŷ����Xi᪞�:�H�z���0��- ��P����j�]6{��8D�	���<=�4�w�v+e�|SF=���r���9cOu�D�����g���y�(��^��垧�����o�x�GQL`&e�BF>��4P�u��ſ��.QK}(C�:��#� � 0�>��!g*�at��8�y��C��.B�3�K�����h�S��g�ܔ�7��g�	�a�02�p^���7���k���ɥG�:�+-=6�Ț�dlJ�Q��}�m���>��!��]I
�Lp�Uі�|�M ��E�T`Q�ķ ��[j�x����W�j��T��*�]Ŀ��IC
G���K!�����Rz͘��s�^���CR+ձ�C�I7�ᚋ�^M��M��?���l����5�������[��%�[� jE=�k^_�m�]m����:���̾�6����B��-�=�a�'����٧o#����aЄ�����%Y��7A��É����d��g�J�V�殜s/C*ٶZ�<�>x�K1W�31K���;�iVj=n��?�xR��%�y�Ib�}y�8}]f=4wQ֠�ke'�8�WV�t8L�&��F�t_c(�p��0J�p�[��{u���9�����=��חo�ha qi�Ep!��6>S�,�.ԐZ��p� q�üp���]�Y��enO'�1r���>���Ɵb"s��PVV�~���;/k����Y���T4�Y[o�\O]w�'n���u@��ʍR��`-<�'�X����j((��)��L�;�"�I�ߐW:^ons(�9i|��#���lZ����2?��S*_���h�� 4�e���K;wiY$����FXڎ��֎-\�����cvJ���:-�:ݬ��6B66���{E�̅U�l�A������^9}.�q�)�v��AF��*������\����t����WI�A�?���8����u221��d�ۤ�M�ǌ`:Vp)(�r��lj�G摉0�48�_����k1�*�% ��!H7���饄��`�k��P�E ���[�a��>R�S���oh��b��
cMk��&�>��cf��G�
ɹ��&4�	�P�u6��9� G�
(��[�\+T�+�t�[�gke�4����V���'� �#E��AZ����	���1]�V��)Si�g��:t���Zm��}�-��2�����U���NNe^�Rb>�����H�I����\�43`�Ą��J�$�>���U(
��Tq5���_������^�M�O(�b�5���Xц6SJ���Ō��U<��
7}:	��{�'���jR��S.U+6�{��v>��G�@j�r��5�f���P�v�_X�8I���ƾ'Q�����L�AY0V�DEm6��\���V���s�gAY���H0���@�W0R�(x*74yS�8	��7���!8c��;&���"�d�y��h2�B�����*d�ܘ��г��� $Z�`�\� &�	0��e�0�6��=Ϙ����Մ�?b�t�	ꔗ��.�{�J�=�QOU��Ѵj�\��K�&!��*K59Ny3���=۱���(�&���^q��� &��;���)�L���z���� �?�٥Z��D��SH�ݦF̞�:���d��6s�P����P(3pÇs��3����nMu�Z �PT�
���ū`<x#+��h�Z�9{��1s����R>KЃ��b��h8�|h��W4=�X-u��K�YK����Z>���:%��.�p�đ 4�@eВ�B�<���V.��V�1t��RFFf�����N���4�<7���Q��UN�Hd�&k��1r�-��p�&˽kq�������x���ٵ�2|�~���9��%$��;��~���3.)	�^@
2^�N��������T��b ��'�pE�h�p��]�3�M�:�/+��]{ʺ_�M��<��d������- P���x�ڒ���?$����N�b]i�qd�G���zH�:��~����\׎<�^��7$�?Cu�v#�?0��z������u�S�zr@͟»�?�R񅤅�����,r�FC�4��T(��sT�!&>�33R4pD��*p��yI\d$��5z�c�[�9#�Ԓu��4�j�9�Zx�,��ԏ����2<�V�%�]k�f]]�I������NR�s�,��cg>���Gj�ѳ�#�~�����k�SY����7�c�Ac1Nn���n4/r�*�B� �[�oL���].%*_�O���E�ۻ� �1��L9���#,��Ah��k��Z�bS����A�?'~��)��K�&�O!�I�����f` 7����:صA �u�I,����e:����`qи-��| :'����~Lhb� _ے���쟅��� ^E{�xI4e��bE��t?����z�A�f4i���W79_h#5":1�M/� u��-n/w�'�o*z�C3��ܶ;��V)TV�N=�^[K���1��y���nF���D�77`������Җ�R����2�1��I� �Ц@�\|�Ǚ�kQ/��6�c��2=/�÷�>���l-#����v����W#�f��}�\Ը�Z|���yg�9D�3&��:��;|��S6�\r6�5)	v�Pa"�渏H����Ȋ�)'MP �׉�ꌃ1`��5�
$;�nH�J!��jĪw�Q��-��h�OD+��]�yln�������@i
GA�C�E'Rm����a�i\�*�>Y����p���_��N���z�$,0*�tS�ƭ�ԍ�{�L�>�3�B�4e]��xo�4L�K�(E<�IiD�>�	�m-�1@���:;�>�[c	>����%�I��#[�a �;�G���t&�룩m���nE	��i��RQ�����Ci�P[Q��D�Cjـsc�3���bT|J/��b>L����'�2Hk���ZRax�{E�Ե��j���F�K�Ge������B�*R��2�Ĺ���͌zh9�`v�
����r�~@6��;3Ю�Y�F������(�b�9���r��C1����H-���Q��8�����4�-F�~��Eo$H�U��F���CV;��P	���`k� ��o�Ub�m"|�3/yP�w�c�J�U��	��ix�)w�B�t��%s�Wl?��PučUo!p�፠�n�j��mF�t�#�*ơ���3c���{�{�a\��={��T�g��T�-�U�y��砬�\nkm]+[�-dK�^}{}��x�6ⶂ���葬��J�&nrmqV�\!s6v���l�cwy)����g>��b�����~�n��F[z~y*�,6��5�l��	M�c���օ�מ�{tJ���$�TEc~�go����f>�?�`>+�g��wm�i<j?{�	�aܔFÍ<��#XU����3��j��C�-ˢ�n�����Ik΍$��JK'���E��C�5驻�Һ��0fU	R+���̵;}F]�e����Q��ǆ��@V�/��N�ٷ�+$Qx��*�Ŭ�K����k�ʘʓ)��/�3T��c��w�^*֬�x L�bm���C��v졪�u�)��3L�я:�8�u��]Ω}�5�Z���F鋥�!����%8Vg�n���v\;���3R:Q�`F�4��8�5c�"1��qпrzQ&���5_H1�ڃ��g���e���a+����c����*Z��/�r����-�5��#|��y���'�7��*�*���)�	��Q|�0R3�$���e���(my*~�A�����l���\��PD��2�n@WbLv(��U���m�"�n��#��}���r��]s`���9L ����i���3<h�?�־����:���9x�`ɔ�|�?��
p*-A <���;��7��t7�������)e�3o�/�+��º#�޼٭����/��7�}��,5�!����uQUz���O/T�a��&�����+w�~3�']��4H��9�3�2Ǚ��2�Q�-��_A�Q&�qu�����O"�0��uo�b���汲p���ar�����(v�G�;vX�,�Ni5w'v�1%�G�ٚ���k#����-R.r����V'"_F���m�7A�
�_Ea�5}$ �U����|�͌���Q1*bd�S�tJ3`��Jto#2Jʕ��tb�#I�*@X�ƌ�~ ݱBV��f�&�Y?����m���@�����|�Q��W�^�=�l�̑�|�9&�E�v���M�<��ͬ�(cC��a'[��i���`�o�7a�ii�\�c�>A�ȯ'i�W֓T��9�4������'�RZQ�W/CbR)����^���������g������	�zJ4�;D�d�eu��
�w�V� ��=���}v7c�M"I�+5ɳXD/�~8������$�PF�(�SH���2��Up�"�3�I����m����:}&O�6��H�ɿ5֞�v��]�xh��� �:]M??�3/��C�O%Iu����ɚ;Ij��ͬ�Yy�ӌ�ש��ѪZIڳ��_�h� �=	�X�[d�����7@��Y�w����v�)Gm]��ы\� 7!܀�~��{?��O�2�a99�m(�t:MW��v��T���p�?c��c)��3��B��T~o-�� ��֘zg%Gt���!��2Ȯ�C��g4�sjS�g��S�� ep^澒��hW���a��u���h���b�r��FA����\�=`�޹�� "ŋm`1V�k�ĕ�dS��щ�{��
 �N��CL
��j*�Y8�ԖNg�;�S<�� ny�bT�k,�Z�� 2�Gy/�A&���kF/q�>�AtTv�<���\8��`�w� ������%��7Zu�GN!8l�i�~��j��p�
�\�R�����N/�}q��Jw���x���IZ�c6�<mU+�0O�oM��A�S��|���k۝�O���5���?�.{=J^d��ހHO���8�gJ�K� �~�~[�v�Ֆ�%��4�6�Zp�=LZd���D�/0��k���B�NT,ai�+�1F�:�m��n��A�~.&L�yit�Z(.�W)�?����w�?En�u���A� $5f�@����.�B����E��Ac+?U�T�C����	�K-s��`��)�q+P�v��!u�/�T�FO���y�҇w��\S���]Om��	��C-!�҈��
�c�Qآ�iE��!�N�~���K�vyԓn2R��^$M���~���U��.	xǰW�$��<Ui/�k?���Av�db��k�|?��m�9U-5,{N�d��xi�|�ޟ�a#��W&E&��R6��W�与�m�3l�� �Gޭ�z�y��Ӎ�M��Z:�;p��0l,Ƃ@��B�.������Ve�։T��i�t��H�_&Sc�I]�g�%�f+	�qQ��Ά��|��-x�Ta(���3��BF��S�<<�̟��{SX C�ܞ��3MK6r�I��}�JpY��9E�ؤ�WT-7t:�)�C4U�4?ݥ�_��0��F���T9�B�������za����;YF��� �>]P�N�Ur��`;�ϑ �-�O�+�i�I=��(�I���#���WX�Hc�H}6*-�M��UD�A�˅A@d�� e�/��х�J�>ǫv�J�~G�WC��) ��?9�c���@�gbc��9!��,vN�%^>ZQ7�\x�n�N��|8K��ć�:BS+)H5Q*��Fw;����eP.Y[�bJ��K�Za޻1�?��@Î���)�%�C45�9[i�(5b�;A�������LV��C�5N�^|TTlc-�c����8� gB -�g��+mn�3��i����뢌�4ž?�b���Kx�e0���TA�~9P\[�IGkX�&�K�g�ߛ4�Dو?'�8��-ay/���.���l	�@�@;����2�_�4�Q��{V�ZZ�H3J֘ҙ�/Nz2�E�*�O��c
$$ni�5�4!��y�����dfo��l�p�y�N�˻�\Ͱ�7S+�`}���܌X_D�U��Q���d�ql��`�OײX_A耎�z8|�����-�F��2�Jlq�<8r6��l�ۊ�$y��̈́��*��):7�b��?7
1Z�a+P=�4�j��J_v�V��%Yeu�a�@���v�k�8�sfC�j/&�� s}�'�Mn�\x�
")s`���!�)�D!�~;�P�\��s��UE����7�=�ֆ_-��	��5x�E�Y+���(�M9��������K�f)��<��,�����x����xHz��mPX��j����7I�1�V5#�s�/j�������$x�﫲��f*��2V�1�@��	B���A/���s�&�o~���+�.�ϑ�tȪc!sǣ��6u�FoL����w�I���R��YjS�1.[n�ە��O�8��-���(�I��~��U@��2kCY�>��~����?��� ��%܆�m�`58�i���o:�nv6џя��^�S�������uV��3��l��G�{L<+�S��Б�<7o�M���M��).!�gD��9pH��c�$HYR�k��։�j� ����L#o]C��R1�>g=��p�������޼�����E��C?�
a}u�yO���7˙���i*-��9Y�-��)^��< �"{ӣ���Gv_.�6����@QDr7�7�@��O�yVZ�g���@�EM���0�6�x�#Pg����cX�j� +6���3��@�����l�L@�'�;���p#��t̸��3;
��S���w��D��S�ծ� �&%ܜ��{�G�ieP���BB��+; gk�4_�X�K��BR�u�PG��-!9Jɞ��c��'�٦a�l���N�`�+R��6�D1-�����c?����]�f���>e��	��M��~���B���]E�q�Bt]��PQ^�x��`������~2���:	�R��_����
4
ݢ޺# j'�b�>|A�և�/0G��m�Ĭ#�^�@�b��d.�p�t�cYC����t�������{IC}Ls�f}۵�y�ܿy�/L�Zf�e/��3������\}iz��N����`�a�*0���*�0�Ta�"�\[���G���sv+j�jǷ�����,������2M���%[`aX����1��D�<G�B=�ZG��#^���D_X,X��aa`�l'�����zx�?���w�H�T8 !J�T�>�b(xd�?{<�^l�o2�A2F�(MTg ���k�,=����(\��4��[�  ���J��d���9F׳ֱ�&L2���Tl��rĽ�7��p�(M�������$�N�����x�Iu���TX����������Z��" �p�ר<��E(��H�����3>9��L�_�7wW����o��nr�W�C����C��6�Wps�\��P���&�Z�|ӕ�������P0k��B���gH]u�3"[^sf�tZ����o�4�IP���Tz$����^7�r�k>�Wx�e�6�5����ʌ�(N.�pJ���
���)��t���@�p�ES� �Ɩa5�����5��p���{�
�Yd50US:.�������OeQz��cE�Af(߲P�w���]��#�5�<���b��ԅj�<�ADW����xX�p�m��nS:�hX�,ܧ��!��ܐ�ʼ�m��='�����wGs������!�`>���4بi��:ѻ��ƄB�uhUD�����)v�g�����3?�q�2�@�wKɠ�&z=�} ��NED
X�#�}f������	�@�71���*���(��m|s���i������ZBS����̴8�R��A�d����`j�����~Ʈ7�R�7�^��$k˷l[CLo��JӢ��j-2�n�P�EJj�a֢L��]lh�����!\�C��]� �b��;�:�O>��.E(s�x��=c��8o�Ț�	��H[̎+����`�n��=>s��P��[�2����߻��]uL��goCj:dd���\�a�J.��<1.a<=�� $�\�γ������X��`u��x�Ѻv���Tt�wC/(���<҆�m1g*���p�v����=6�3SX��.�g?Њ8���<9��V�X��@�����Z���.��[��X�>�>�����>���S)�UBPx;6����g�*l~�BS�.�A/�q�핑:��B�����ݭ��@����T�������
�&�z�|eT�uW�G�t�s��!����!��/�H~t�(�#�l�[�}��*�Z�dz�T�W?���D�5(6b�����ƪ0��њ�g��q��^��F.�^��7J�,z����݆�_~�(��n���fuF-�Z����x�`�wZ
������e��a�l.]���1��}���EDV���0jHc����Cm�����|�;�(�}م�主
@�c�f{�!�YuZ8K�/�`�F=��=����7<�S%��es���~��@l-
;��B�*u_ZW]�W�Nw�嗤���D`���M��49�%N#��X�1Z%�C�&�]��![P�d��<r|j��:q/�l�N*��S��BU�a�O�݂0|�	�ً�ѹP`���=��̈�!N��Oy�a!ܕ�,H�l��Ć���+3~�~����=�K^����Av�D��[A@�ԑ�{�L��V�5˹>�e �̩o��V��uc��x#��ݳ��&�Ф�Vr��In����q�Y���9��]�