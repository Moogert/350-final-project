-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hu7pT5nIqNcsSYGGM97gGa1qQuxHD0dWYWqKVQpnlvbN2PbohxoTmDYdWYscHW4oJ95iik//0WSE
DbImWelHXLmWQHerwCcqoqIdqcmv6zDDwOe6kjIXF6mM6YmELXYDtXLapqiyvv3Aom5Mpbp78RrX
PyHLOANM2X4eFInwd77I1lrpdfD17cHRm+cXW/bvRUe1K2wsukC5JiVz3ZV9gyfObIOPY8+uhhZ1
WxIMFd3165wL0gnR196pWSiIhEbkebDaOkH71OLatk1SQpvm5vEpp2dCr+H4xLUtJjw59jQzpVsl
IDz0nQziz1y7Pa5dYprrwC5Dw+j8QxZXN7GsjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
5/q4I2n1fFl385UdjXk0lx6oxfS+8njytyQM8e64t+m2J5scb3lWi9VSBbWKmh/oO6GVsolMvVZT
MJ+pMY5UT6fMLVm3Cmy4XSKppy6Y0OSl3Zkulmp75xpuMYH3FBTm14l6LCx/xQq5VpQrcj34OFvx
FZkGucCB4TmCXgJ8TCEF/dMMvxt5vk6q36XzDvE6x5Q9e+AdaYjco9vQHmu7awcJhcI8SxZnqjsN
UtR/NAy03+5ibwOhLXONgpbVi4J8foXtJ6LIJ/GTJxNc7lPDSChLFQjOqOK30lVifB95JRT8Kekt
RBgxHK0iTR+HlUE98XeU9aMW0d/kOIXEBbiplbjffCwHOp9dd5AY2WUNa58mMtARpeABgVpl9gii
C8L1nvTsNjcrfLi7hXugfIApc5C+pU0kcc65ERrRaZzboJaZpkaEjkjqAo+XzdE01uxZrkavj95n
IsoBBNKWRhi14gd1CBE5lPHr9eiK9B8IvFo6T8UqvVURIhP7s2g/gUwn1Yg4gZWtNsVm5n5+8DB0
37L6EerZzetaTCGc+vjm/G7cnez/8rZzT3gFTckYoiOzyrzzI1PJIYA0TD/mMj75s0cYiLvPGQc5
yMiOGFUUppAugrvuf9cMu4HcTD2MRWWLfX2Hb2XG41JTAVz9Nh1wrrk1grWLTD+fVGZsGLeUHNn1
hQ6tkHq9ZrUNEpnVZEOuRCDNi6RO1pdrSvHf9w2NJIkYJtJQrQr4Ysm7vBwH/5yqu0QPMV4ab/Oo
sBkIWgWyjyJ8A/BENNMJYvb23jqg+CLQWgLc98jEERPqzxR+2nA8RbS+O2F1kOdvYVH/Ox8+4R0P
f+BUs+FdPSE43zURm/fumu9Kk6SnsUB5p3jxDtvQmFRtkY8EL3TcaSqJpfzJb8WjEarAYWyKUWxW
ZPHI9J3DDbmdplsHNQo5MDRGGCo1ft3l8yLmqE/1k9Cu9D3w6b4IY9W5eD2M55WVir8JF5ve/p/O
bXSxEWslyh92Io48aStLskjq0ki9obPnJgkrZTjwJh2dxf5+sSNHzih6KJyYlVX/SFnHCihusuvj
CvmRRtobznCrGWWmOHejwnqILzKLGxlx9xfxF1huD349uLkb/ts4sBTY3EqjtO3EHlFHez5ADviK
fewe3P3aoxUwuEvhO2JfxuDltFGwueLk5eVxAeuD4NRbKNVR41JoWgPR244WGIZzkYUWen657Zqr
PyFOV+4wSEhfVIwFv/OjnomZCrkp4Xu4STX3YHfVtIO4W52zsNOdC5UeVY7N9owsUWK+ZoquFuQC
U+z3C+hoZTjmWfC5eevsE7ak2WuM2fN9HiR8/d8Lu2TtMHrJY3bVdhS6dooQR+W3n46DgdUTQFXn
f9aHG96f66Sh/UejfWSnoqdSYGc8XRlnrydbrCQW11dt3r/F1mpxC8XAt/Lzb75J6A7kFlYkLqOu
b9oUeK/UeLN/RHyWBZaBBc71d3O6mmiblf3oGdKESKC/TCpnw9EB0XZaZDLGedPQLR1vXtlgXHhK
EX5yi+S+gDt6iW+Qd1tQlsqx4tIzBZw2Jx95G5t/Z9QjKwGV++C5DD2lGK9rIMPZcEAlQhm1gwSe
0zdzx2iQNPfBPsuUfCIFWjz5HE9/DvSe0N2kjCfgRCz2B3pVGT7V8qIRqfOW2AnoUMW/dpBiCv1Q
rhDTcSSkaGBhZ7SDVjomMwO1wfOOpluVsgMQ+SBnCslKebSenZGvBm4TPOlO+eqCypnMbG3cEc/c
Pc/sbKEik6hDFT2ZtLYv0t11jhA/0mKS2GNVikyBCnDAtFpAYFRoEy8eMiMGw0uvMN4lusTbh+JK
y1a5p8G2oRl048IEuleYxIFIlFe64KOwOGAJ7NkCQaO4GlQy9rF+DL2KEb1+6l1yUki11BVneuJV
E6ui7FVpk2miYdV8/1cerMZiBen5Sb3tWOqUqx8wU5xsz5BacIWHso86dzczP5/97Q19LdfdHCIA
hYzvnDNoBawfJkCa3EYVC4Lbzz5gBVx4oWXvIPRvA48uCk12/HeZJqzfSIDH7BtohqkZ+JG49yvR
rCBoxtMspjxxIWivQ4lds77fYkpisIxOSxbkl2Voa8865unrnN+tUmDXJuG+Sp5ZdBe8aXmWyQjr
Y25+a7bKADdwes3vHlESu1JWGHGGQtNyzvlZYlmt3h8X8pH5nNOgPffeT3aCancAKl/MPnJQQ8DT
+zksTrOieum/YcsOM3VjWcZjfabEz7bwlzatIoGzM19oUdLEKi1jy509iALpFhLmwA556ZGf7vle
foYjff3oI6d4fhuG6vWM1BLp6hv3YaKwfG0pWuwun0XtRINxpmWXBZttqWkI9GgCREZdFM6VL6DA
rhou9CHrAkyNsBT1MggEcVu07U57HNjP8k+Xfhz0oVC0HID7CpVgJpHkwzpdoYo0tBggQQWZmOxc
0mFKGtYTwbvtAnKMM9PaK0QVtE1beQ1ywExpzsM+YaSBTdDAG/PxAlIljNXvGpMCoZITlTEzf9JQ
vM00SWqpSXKQ2dVZYulvcqzv82t7GjBlscap1kmiB8yXRQ2gCkpDuEN65+OmynJ/NZUs7W+HDEBw
gtCjmlRQXIPEs7XMVOtmXs5fHRoQJa2T49+rOxeYoL146Rc5uxdkGI7crUgWqV0l/e1SPW//9Siz
//PnJRkuh+ZmCLni7jxVXaWXO2X8J+zJghUszYfqLLEVX6Q35JLttLv8MKJexFYWGwwhP4vGpohA
HHPDgmdPtKC4s7vu449ywoO0b3qWJ+asqNWoyxz1LP4mAulkH2m/2UEWlGQhLyrwixmVfbafE7gH
DjWfexudC6FtCCXcZpmPBAorIC408n+ftWliH9knNBNOWYRm+SaBCqtqveRSKfqgR0qVuhgTEAZe
okBTsTF9Bl00BAmXJHbY1BxiX0+R7aiofVxc5TtxVHXDVGfJtyNTgkL5o5yy28wTlAJ2MiwPwI7n
UWat/J1qU13+VKrkPk2JX+4I5XWfn0/fNWyq7Z0wkwO2hPoUXs8XjpK7sbuiDHzH+kr5ZI8d8opc
5yCraU3kDpbJBxfbXzo7pGW1R4sPztc03uW4GLuI3RZ83qKy1ZIREXfqNoCJHmGw/8+/sI7/XmVo
u8ug4oFfi3c1waUrEAtNep25RDG5iMsTd+DG26cvq8VeUfg0uzBgxjimFm51AL6Lyy38FCPwEMNu
DhNVDfGHsz4LS56ut10QMO/h1kzfE8CFix2BBsVpUrR6egfXLs+oyJDI8ZYluPiukJUwc4GIhkcp
Tltt4a6GyCnSWnPZv8ZEjmQT1/59hawql38iS2/1oRon/wQ/8/dndT8F4Z8ujt/TKQqu0ro0GuM8
Va9kWoBbEzPGbUUXBilfVqwNJ/rhC4KnxqFFXYzy5ZYWgnahnOtALlinhLH7fZOmvGVNL129ZSjP
FwWhwhsDXhPtYPE18qVrPLPi218Jy056dOWYSh8VcVdlRG7YXDfTlDZWhk7pinDt6pL5w1UDDtaf
WPi4jml1S+YTJvAlvvBHzJGVKu5CsrIP5zAb4LHRtIXp61rN8i2IJne2Dd7/x+GbK//moYsbW30W
/PNEkncx4h7UW/n4cmYn0a6YknHZTMM6ri6l2tQKkJolSAwPsuOWVy1+Eakdx0NuGPiBDrQnJZXY
6H12+nQHdqEsBKFBnxW3PxhYq06LbWG5x7qJ/jck79s8RjTJW/jsIRv3NqmV9MDrEcLqIjKEqQKD
vVAktPJAvAXHdODWUKAeBUWF2fLQUgarXoyBEzM8dAexlGredzu/MqjCsGLupgLWc+PBG1b0qSe1
zfAXHGJbSNktlpagzBUbyh6aZwfjRgOIygaxY2K+t0vjFzPKMSY2NawCHnZswtEJw4idkotNaAhG
1bLWNRQmMyuoWLBdZsG0oHVCgij0IjcNEWuEPg3UzKdgYc7Xb7wtcVvgS/N6E0ZsCARg4gVqZhcU
oApOBQusipqn3X3gZ30Y0+HhgLyMc+/e5KOntIpzVNsjuVUqC7Y6BTTx8zNljK4eftBTohtmAJsq
t1hPjVnj3d7Ar8NXxTvsivtPr78A0ZKvLclu6LUYnYysdH4UilIQdMSiJQahcez1Yqswmz0uV7LL
pAARg3p6mQZznhjrGOphLSCGIe8XC4GAeyuuubZYhXxIKuvhHcMhoR3yzrTavIzMcjOw/Vw33YkS
Qa2zpd6bxWLft6XGUzOegtx10w4ahlekzGZoAM8nNfo+GJsQ9zHdv5ze+yC2lUy+3xGcHEsxYUp6
gp1AHxnjIeU4CuozPypa92Z8lw4VTnwcQz8CDwa4iRX3icduJpPso/QJkOvVEJzV8HEjU5oCR8bm
2aIicG8ZdAuM9N72qfjQ4phfXPaeaIlZKmHRTXp+4KmOm6bX8yv/ragwTK+urrFovzbQdwClSJvz
pivUYOWyN2jkCt2ICbKHq0agoHCn4I9oMAwT8PIl+TIJcGbCEvirJYfuFhUSx83xdzxt13iWrQ0T
/R1715sdPse0j50i/j20QeWOJkhQqJVPZNu9+orUX2ELI8NuGV3+zamaqPq7rW6v2WR4l5LxYFG3
Fg8FrczgMzbbhluqGzSpgR16/ySY1s0TRCTqhNxz0UI7mdAV/fBilnr3YfSvkpR1PLQejlX1P3dw
Qufv23W1OYRZ4AW7xk64UobhlRcTh4q2k06V3FqM6JIu8zmZCGCAAApuKGxpXxax7RrIZkpbWqF3
W/0FaZMF+wcL/8lFAjzkzw0wM63DZqrflcdZHW1AjzSSbGjce8nGtD9zpOZqpgWDlsy/lTwkqjZ0
bL5DIdohvWNcWZbo3P92ifgT/Zh9TzHWctmbJhePuzTGWniDrFYHPlMehUH23CdznJSKmOTfQbp0
RdGZrrc3Rpbw9IVBJO6EAYEhkfh7nsqKfRt+EdTDPZUPRge8v8RG7hG6aQQ0H5ejhxwUDQAMnNea
b2KDOc1gM8vI3kWxwpCNoy+Wy6yMHqMOQzyPNrjyXn0phYIBzTVZjyaIj/KXc4J04V9bQvIaHG3Q
9lkH5ij2ldIWNkAUZrXUEywuQSREY9sLJsrxFIud2zxF/JwxCE3BLp9uenzLwe+2zrA0xnyzKMTB
im+sVO5/9ZefZch5WsyY+OcdBVXfZo6rbV+WTvdqpUqDoGm/luiinVwsdJGlA3s5MSB1f7aY5sMV
WeDXgEVOqFVoVVhH/MrZ+cTIsxc0sNmAmhlLGp+155lNd6mMw7G9OCVBnTU3/DKNJj7mcSqzIgrN
MdQIa8HO34IGsz+SBXt44zpz7/t5wwMOl0dhRAyljQVlmZrsKpRcx1qALYKPEgEsBXyhiKK3VAb/
X2YVukXxQ/vSUTvanOJeevH7W9WTELCxOlNi8FgfVY8hjwCQe1I4s0lWh9r9vQ9xj7vpo3w5YOdJ
Q9xJUWCE9iIoJ2gwKnRAgP14xRqF5QfJ+ibTxT/BoFHF0lBw36k88Kw3Yd/uaWlrQbTknjcTkh0f
06jDRDrl0x9Lp22o79ic0lBhsAnJkKags+JzsPqsHxBd3kVjORoiOkduZfa6Nhnh13/3HyMqBTaN
hI4bq/pfkVNQz5EfjZpoKudd+1IiJGgXcQQtVzcLHBcPLtMM/CYP/UCe6qYnY4LhVIyU9bOaUv8r
Iqq3XVuFklrRunOoIMNcQiPYoyz8A1n+UhlgqlpOZlVOV8Nv5uA7c9VI91sBIA7Ki4PhXY79RmR3
U35YHIUtYzLTjiLlYyahIWzfJA5usVipddq/WFpbAOtT1Rd41o2r7Ku5sQdMdZPatbdyFXjVULK+
4OiSdvlZXeOeHvFQeblxV7xuYgqdH2EOOPHdhK1r8hhq+Wq63ZCZW1sndsr18Yv19l9myki5FFKp
ZJbqPjvTE3GcdSSXEHHXwXL5Q1l1JS4GNT+OV/e/j3R5JnD7L9JFr4StVjTKIFjw+YHPNHBTmFxq
1o1VaLN34cd7Pc5lI+NYlOrAXJj3cZBlO0TtMewNYmBZiJ80hi5xkZPU8iLqWfx5AeyVCi+TBqk3
S5bTiCwNxPnb4vjg9UFOjNTo7kpWmePi5ftIAPxRrbK0xPmSnt33mJjfRp67rAWlmo4JV8GeHwMo
28pcuMwUNY9/AmEcsSUBxk9sC+BcNuVa+xbj3gXWuO0opZ7Z5g/W03FMXX6N+YO9/ZSoGL6x4VXY
OzPhmsgLob13l1vDInEQoHxavfwYTocRUYxk/zFtLUUQCDZh1rEv5JtUkEbX8lNe7ANXNZsejg2+
KUYiNLlmAIV03kA+4qXXhgD2fD+IJT3g3+wsFIobCgss2FIS55EGiBJxsxYI74af23/IZie44klV
5mgC65yEq3Gea0Cilc7tsGMdwdCx8bR6J3kZeuj8q8ITjTLkJ3jpM536sfzeAfEF1VwqXUDqVENs
vlKR4jXs7H01eKzahLBqID0SI3jaOdlVmRbW2f/3wtbF2ofzGnbRKkyOQA3OkySf/sH6rBjJlSJq
18QysFQyhWpP4wmB8F2gpEO0f43LEaiTIiOmKczNKeTSbqjaP9y+XXCLKGJPBshBkZ6BAj09i7Bv
gukdPZqoFVEOv8SpZHgaKlZeJ9LgQ7hxPvHjJfFp+evO6V5SVd6Rs2EHpl0uMj6Jd4khAzPEMJvQ
2HzB0B9XLmJsrdANgUgPwezcYxRQX//+EAJ6I9SfMUiDH4iqcZEOPTOhkdLg8+knoTpQ3nNBPy9Q
BM/gxclTv9aBz0scuSY0ha6ZwoEN18fMsmN7Tua0WOzJS2HuWtp5q4NmaF2H6LSXUp/cKlueVoql
v25DDeNsTS9+iVkSyq8e8CX+Wk3Dr83Jy3JWb+9Kf94Z6ChB0liTuVZVjeWbWRaqz+KM0PiPKzKt
8zytN7zbxhDeZx7UhTKx/ZSj+wjt1QzcnJi0Yjn1e/fC+JdnOh0jqDxO19ZQnGYOExD6BIqXNFuV
1hDQ/q9G4thyxN4j6ivIgF4iLrSzrKQk7IiggdVClWas6JeOChPfLnoWedNoKoBIXyAPiW5Vmy80
DCNx6BuqO9XRyu08Dc6QY33pZS2fXryd/bziGsqLo0BCFG4GBh9FXVWyb4UUuqAmQWVqCo0AAQ96
lKAunMcbT7uAoETewKVnpooaYqKQF7DuDoSQcfcc73uDlS5oXvWB0EniouLubhoDI+7FqME1UuWQ
FIH8IxKHlHC/5gSr13Pj5nVBi/ScSFvxl7EpUm4/KddZNBYykc4j+eQqV6QCYe7WUsvuZJmR7o1a
JBXHCplTQae/DtpObQLFNv2XAdEFXILJmQ9F+DhoV8kQUqkjcicxBwJ0kBp08onJ6ss7KVtVU2Wn
jQzAYoDHwWBjTbvXrEA3bKgK3OYnMhoiVDu4OlhSB3JDeCu8wpGgMwUZGMSht18qUmnabacKiz2w
RhzSQa12/Dpy3N+2N0JXhsiWIKftr5Nr0Lfa0uL1NEt24B3mUvmM1hByxpT/o9ALMARrncjIJwL4
rX8Jxss6Boj/m7aTYdJAves3wvSvkE3FYu2vpCWhMqOliWpbayBD5Ag/euYU7dhjXD/jx9sbeH0Z
cqSqPHcvVbULOxF9EocNkowtX3KcngiVgmPxe6iNdc76pJZLLnGGAItQJlcD0yDOgYOlUxWyiLzl
ReKLY/Wqjn4vQl3LaUpc0CrSQoknBdaEJ1iTxPXI3NNtKUfII63NW6kdq1j1Pii84xjADBGrlc/4
anWbMSbP8wfAACYYpQ0DRC5P8Ufr6XLSk/aNQD9LzDl4QNtcCHQ0dcDFxYbt3ioYcjulnWTCgkH+
adDmXVTUngNHKHr24GtV/1u8jjua8gYDd+NGi/Qm3LnGx6sq9iWjHJ6fhG63g9pGA6lOfGyws5pD
GdHFAo76NEjvrMVefiwKhzrsxj0wNVJgeV+GhKR1rknOyIE6bHU487V2PnM9XB8K3NrTL95UE35q
f7rnJSfGx2DZp7UMcy5yuShIjEfvAzohHvnoaE2i0GuTKYaw1OgufRlWllxUDrjNoqb8lx8K0vp0
9UZK/ydyASieRJkaEx95EGOkOSEYE3DLZrxdNi8uh5xNb1sPAhysNmFFDz8cjKqI+4vI0maSiCZG
UqkGw6Jgp8rh4x3L2a1LXF0o5hcgwfz1TmHHJSu+fGh6qR0zx7fJO+0ae0HBU7g9TpwERCN8r6wZ
Rdk5KIz2scnAdtRBsuiMq5HytXGw02bVKQWpiQ8/FAK38GzFLsWqBSrM0K7qlSoJsZbqHVf7VOpn
VvXk/N2HMhXE5IwiU3SOYxksCAAl5X4zUOFsw8QAjeLp4427wTc10SNUnMBYockhAMSzQ9Rva9x7
jxeLYnAc+HYsGxzK2ntfOupDB9w1d9nT8pc1ILSS+7UzfiIOiCVWrg18ZA==
`protect end_protected
