��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�?u+οGݐ�>J�,��:.���;�g�m�k<�.��eG��>��Hۑj��k���Q���-V�h�KV��f�e�${��Dw��M��ڟZ�$���6ov�d���߷c�CӞ�2�����!)DO����^�����Н��T��3��{���3妄��|�*�!�n���멼��� �H��#Z�4kȴ����$���V�yJs��G�ע�!�S0}������fp@O���]��=Y��o�P�=�uę�>c��}8��!g�z�rr���jv��8 ����DXhCQan���������$u�1A��o�{DF���\�)j�`� �c��ˣ%B0���[2'�xr�@Y�it�1h�D�~E�ı��������nK�5e>�oKt�2���Ѡ;(F;�Y��ǈ^���cQ��m�+`���B�9�*1V�G2�_�&;���C��]#籋_�
�QD�kǠ�j��&�T~�����w#`i������j}JB@�M51�EH��WC�~�Q�J�8P�GmF�?��X��8@��5��
��ꓽ3�	z3ԕ"l��;��Ж�E�Gڠ��A��9�Ԕ���	�Q/l|	���e�~`)	�<�T�-�������C���`-��c��,�AE�kR6m�)J�$�SW�����5N ���3R��6jgQ�!�� �M&5�GZ�Cm�Ժ���T>D-\|�F�?����<$uL�3���uT+7����4.�Vqu#�3�񲎦~���	�� /w�����)��	�|�H#A�)�M1~ �R�r/��% C)����$�P����1�W�O5�ç��a'@z5	s�@>�yۺ��- �Fv���)�������EW *x�&��8���s��jI��uNZ���J_עd�H��DPc�Jԁ]Fn�ͯ�M�@fk+�dџ�׫8ǾQ�Oa\��Bņ��g��jj;�֔A7��I�.��#�b0�F�������Q���_�����F�x[xC���\��q��>?.u|�h�J5���b��<#	��q3��b�����"����z4��:)�ծ������gU(�E�x0c�����s�`�����E�$R�^۶ᦘ/\���|_ю��{�u,|�:H�9�Ǧܓ!*{�)4�������,�u�m�Q�v�gb�뉦��iqb�~�ݛ��^Q�/��@��d_��ӦaXQ+��e����	N+ѩ��z�����d-;���8� ?�/����o�ʏ���cM2X�bG�G��ݙoI��q�K-p���\n�]�[��9R�����pO��s�a���4��4�0X�;�u����p���m��j5�>���@�.��e��__EY�$
���̣As!Ԏǆ$�+AG���^��+�<G����G����.�:A�	ֆ����3c~HIEO Uz�CyK}!fa$��_�U7d��Бy�:�}��p6_[���	�v@��9�s2˙ψ�r6:R��lQ	t_<��I��;���}xG=�6����@�r�$�v�2*�޶ �Ӗ�OQM/��?��yl�y�N�!���&��[߯����8��w.ĨQ@�(Lv�o�h�У���M}�3������
��R	��'��Я���\ҵ�`�vY����Ư�F� �K�m`u^\B���A�D��>�
�79��kT[qK%bj��~�b˒W����鴻�gѱ:�V�p��ͨC1 =�����Q�����2�?�c%u���A��1n�UӴA���k�v�˧D�@�+�W��&2�(�Ǖ� 㾔������"R��B�0��5��^�Ahp�`�4bNb�>E�Pxfb��Q�``e��}�m�RC�X�892q��8g�9A�N��^��f	��:�#�n4a���Wdv�m�����*�R���mӿ84����V�Г^Zj�	�W7�xN�,��95����Y���#t��G�I��'�a��,�4o�$�iN��.[׋ 9�؜��t:zm�˿��2մ��X�A'QCH��Ds��L��DG(������ӎ��hy���n���h�dd����c������D�4er�F��*�dwrX��V�:[iWw��K�w�n7`��S�;-z��7�*�f�Pȯ�N��['D�v��D�ơA����+h�E9�_!/ ��=�n�^3)�n&�/��]>vқ��W����&��v��X.%�S�m!2R���@Is���U�*�CfЃ��^\��Va��ܵ�̍џ�Vw�.("�����'��Ze�I�v�/h��l̔:H����R�M���A���?z5NE��S�tŁ��u�����ώ�ϧ��A��ݓ���1��_��E���Rd�cVi�0����u�*(�����q���D�9��D��6�o?P"2���sn�\s�%/a�	a��#�#�.T�5��eɁ��XaA��{�;/�����4��( �M��[r"hd.助��~�!VY[x�ۚZ&ƴo�P?��N��D9\�Z=w�faԾ��;~�;��%�Ýw�s��s�� {�ւ1�)n�}OP�k��z�(�V%[���x��DL�;��i�����#�� �{ti�k!N�fG�I"�b�𮳸����2��پU�B�>sq�Z^6�B��B��?�����񡴧�m����{��k�kV�h)]��W�W��y��0<1?��FB_O��&?;���#�6Fc筝+֩5|����ɞ�U1tzwr�4�
"1$vb�in��R~\)Ob��6-���a�[�yOz3it�O�j�`��HJNl�sr����R�at1oea���ͪ�_�c$���`+۳E%�&��(�OF�dΝ�%0�?�=)_4�>wL�S_{�`g�$��Dn!4�����-<�cJe(;GK�p$��:�|gT���wĄ,_*��ؓ�*�(�2.�8e�S�(:���}���U<�CM&w�b�qX������#R$�Лv��2[2Q*��"�w��JD�4�&f����Q�#���WE�����%�rs��]�VG�H]�nOy�0�-7���l㣳�u���u0f��)��Io�P/ș�>cGà8�C2�X]{�ĸ�������+b���(ү�?y�z~���W���b�˱�$�:
i'4!A�R�YTY`c����ws�!d�gӿw����� �Ȯ���.��5�_��ƭ���Q�~��2�d�as�ƫ�e�л��Q�/Ι�����?��Tf�jҟ4����A}Ř_!�қ@�M�F����R��&,��u�,���I�.~ި闝3J�%���B��dV1����D�a}GG2Bo�e�G�C�	�Raod�Caa��\6�e|G��:��\9-�X|2,����Ζ���T��9*T���+#�D���ƪ��!�)&�kw�z��w��Ƞ^��C���]���2�3�f�a�ɫ�ɻm�%o��ǯ��E��! �ʰ�3�k���O.�����ּ�W��l|��C�,�8�9�E�������Dk��U_T;aD̛�d84R�p���{�j�8HZ��A�M�T�Ye�!������I�)�=�@���`�u�w��	>��|�)�"U{s�RѺuۇz�u
#t����NzYO�TS���fA���4K��R�� �}��Y�w�
��������B:� ���oV��(g|FB�MR'7�4Fd��2��Sc���x>5�X�>�řR����9��C�}C�a ^�Ⱥ�|Ϊ��-�fE:�r/�c����%���l�9�>�QnB�v�nל�b
�]Ы z�zY�di�0vA��'a�k�s�$�ʪ��wK
�����3�`����ރD��7�w:Մ���ĉ�5j�b��z>��D�	d�n�8��������s�VI�����w?�L<�����6J�N���{T�ERp�|���d�Yz$S�tJ�s�U$�I���� ���,�q�01zo��"ax>5��[Iu��b9jb�V8jB�:>��'(f��BD��+�=��CA��KLA� u����b���x,v���=�!0s7V_o����S�e�u�eA�Vd�{��;�v�Y���*1��̨	 k�B2q�;�*R����j�H�G�>0��yE)��C���bڬ�`�/
j9K��9\ZB�M��>v|;��X����}j��6�իY̧����qu����[k�>f�v�#�6Ή�'���&J$����O&����'j�P��D�0���FlG�2��eiJ�l��@����:J��[o����wm��z���3s�L2M��R�|,>$�U��"??�#��9T+�:˹�0�x���E��O��;�N*���Y��Ч��+�*|�d�ܗ��H�]�`O�.;���PA�{.��F��6���Nݤ�3\�Q?�5�~ᧆ���b|�z����3�P��?d6�|g�u�翡�-�Ӄ��]PPj>���u�K_�tt�w��?zB)��VJ��@�T�q�����vjE>���n��r���5���:����|�bT��O׿�#NIJf�����B�F�@k�,6���B|��`3a��An"��)� w�H,k��2b��G!��hM�J�JQ7=��ǿ!e����.hz���������~���n����8�wx���n��R��L�ߥ�i��Ii�զ��Q�<�%{�Z��v��;X���L���Ե�O����>���f"q(�{'kɾ%����>wݧQ<���l����_��k�l�Ѳ�@S����Ma�IM���	�&��u�z��w�C�S�8�1�4L��fB��0�z�,`Y���b��g%5$��f.�~�=��"�1���rD񜷾��g/G�kc��%�<��I�O�zi�o�Q��-e��~����%3Ʌ k���*h\ieke��Q�&�w�B� �3��x���V�]��mfP�ގmC)*_v��K�����_�DiI�.��85̴��v]�i��� ���U%d��i ��՛)�Y���}[�����L��0#�Q9Ð�~��n��8]#]��_� ��(��_OL�/ތ��x1 5�&K�Ӧ�'��o�b�!6��(R����Cߖ�0ik�v���0�f�ɢ�����H}$w{�G���A�������o��ni%��.�5!eY��w�H�_sU��KtS��9��-��[�?���Ȃ��mx9&2Y4I�) �����!Ҙ��j����`f*
��MA��\f��[ ��J�p�s��P�_�軯����6Q��iX��\ K<S'��ݕ�i�Ԡ �@�,�u�W�w��2�:�$�vnB��q���y�g�Y�e�<`"��q���)Pc�>��!o*���&G�����^�jPG]����ˍ�Ϛ�T�o_)L�[�{N��� �G����*.����}�T)j!9u���^.iP��)z:��-�&E�g1(��.��9�U�W=R�FT�g˽���_=vɣ�W�ZlN
W���	7z_�>��XL�/����-k]x>ƥ4�d�|I�����G�n�T�Y)@���\����A[�)t2��geUx��1@�Kq��#�6C@U��M}��3��|�3(���{+h��ͤ���y)�x߿Y��aK˘���jgZ���+����ַf��T�lRS�>�	��4��ό���8T�aỎ׾W�d@��WFzo�+�s+֛�ƶ�M�ʳ��*y�}kx���2���)}���PyJ2w�}7�G� $rxG�ݫ�Q�(W� �0��G���3b�=X�	݊��"���w*��%��r��\Dwc���I�{/��2��3@������U��@0($��mE�o�fxP��;��ȱ��V^
���K�r}�>��t]��ࡹ�	�LO߻��!iS���4U��^t�����pdnKJaD���p�+�OP�vĦ�5Q
^�t!��W�;W�mLޣ�T8��h���dާK�ѻd�����Ylg,AK�����=�~T�T�s�wnQ�5@���~[�U��KKe�#F�hҸEo�a�Y��a�j��VJ�Q��|�5*l&&o�x�q,9_F��2����E�t��Р}�[� �yvJ)�@@��W�&\`�L>Jc4g괌��3焵!���vن	"I�Jݹu��"�ss^�KT���}��͍C-��yY5���&�����DF�{�<����B�k4���%?�2L��L�����ɴ��n|X��,yN�v�w�����>��'+��B\-0���
R�6�$�����$��&�V �\�&E�����Sq r�;S�Z�v.���"�nRf�8��*�1��gc�V.�{|��l����:&�£���i]&A����θ�'ٞ>��	oRVg���#�Nd���:�!�3X��B3�����j[#b1�cs�Q.3|�h�^��3�z����t����[(�Y`��^1�}���!x�*�տ7��i���}�-��3�	Z�c*O�1o���$�.$�o�I�ƶ� �!!��O�P�1����7[�;S?Di��D6�e�yi�ߝ\V2]��z��qwo,���[����)ѳ��|)~qi;�:��~ƑO���#G�㶿�GX@.i�)7G!��B�y���X�'�W�u�=��]7�M�H���Y?���^��Ӫ�����Lw(���1
�J��T��+�`�Y�H7v4y��U+_D[���Lq-oHÊd��;�yU~�5���)g&��6�J0���gNnd�XϾ�%X�J�\RlԤ������0���BBH�������"�n��ɦ����:���oF��H�E�yʕXU0K���\H:�-��d^'7�H���x<�uϪ�8���]%��:~��]���x�RT��������5����6�յ���f#���\��+<��kZ���]<3�*<j��0�m�֘�#�S�<CP�'�ݭ]я���� ܞ�n�2�X;�Hr]�Y}ꨇdq�QC<���S�0]�|���x�5�f+: ��گ+3��vU�8h��E��Nȴ��:�\Z����n50���J����U]������/�QgP[���
~5~���2�);X�d�����.`�EsR�M֔U���~Am��0^Q_2^a�K�E������,����!�J�9�����FV6�yR�&Ϥa�;�8�ع�hn����l�JB9)~��d0p%Ti���ˬ��:f@���Lw���g��X���^�Qx��t��H����*�3)&�������6��"V���f���׮�~p��طU����Jrި�����:�|	�B򽡛�����C<[��cΑ����DR$���-�,i�~ꤲ�|��^�:\~�h븊��`��'V2R�858�6�2̭����{>ЮE��N�.���%��S���	k�Hz�-����E)nώ�@<ٯ� ;��}����|��ΐ1Xx7VL� \&�P�����ש+���u�q�c����? �E�vm�fh:�l)eM�fwe�C�^s<3C�@��.�R��b&a`Ԝ���b<�+/�����0Ǭ(N�v��duY���RGo�15�&���Q�F)$G� �z����"&)��!V<��T��b���&T^��JL��:��.��|/v���-h�-�7^��5kjE_/���Ϸ��&[Vms2Q�Ik�TnA"`0=�� �~PW�	jk� ��S��� �YM��@1`��:-`�������KۀIм��Cl&� �2��ꮙ�� J�Wo��e�4v+���;\�z�~S@C��'ݡ����>����-f�%nv��y�^в�d0
�""�G,A	%c�U�kf}L�&��qD<��/��<�2�X���{ׅckΆ�Z���N{�	�4�釁LE���pL�ɢ#�3߶p�(]4�`k�o1;���L�G��Z��P�j� ��&�Y�x�"�O�!�_ OQ,U758�l��sM�b\fK(��E��fp�=���91� �/T�9��c��yM^�D|:��P|�x62_���7����%��u��8A��U�F���)й!z�M�dd+��V7�UfT��O���&+>"ӼpqOp�PFqO64� �y/ՙ���t���(�X�٥r�^�^��#O�)�V� �S���V�RgT�i2�9����ˌ�n�:����X���bïv>�,����7C&eַƒ�/rLP� ��`?������/#�N�q���$���`�5gV��v�Z0�Lb��r0��/�M5��T͵������q"'�r'��S��T�/Yx����:�bo��C�DM�ߴ����^�*�
x�!�^'oY�P�@�t��Rv�ڍt�٧s(V޸��Vy�O�`^�a��U�y�m���P�����	-�����y"l���	~��1}dW�Ųa�����$7�Ff�����wh�eMtO�T����)��tF��9�z�u��d��3�ٽ�K�.Y�2c�ԩE�J����zA�Ѓ^�୧�_��QN�4�T)�"��T��s���օ�j�^�A�<�i��	��7�tM����M([g��[�����[*8�w+Hy���Y��i��D����%��Lisi]a��M8�	�Uɚ_f���xW)A��Md�z�B:���-p��!�Qc�G!{���S�b�qq�= ���!u����edi����x.v�GyD;�%��n��п�)	�e���x�	�R���&�0�2��չKϰ��2X�\��S���EFt�e�;�iHȝ}�����ve�C�$zVx��7z��?�q?��"w�e�q�Ǫ3:�,��SI>z0*�ơ�<S�z��t�C\|���-Y��kP�*��yM���c:��)�ޣnX�J@Ct~�CHI��������y3��
�d)TC�� ؄�pF��N���*15Z�j�����H��n�xM괾Wd��|y�p�9jQ}�ip�X���Dv�k�����'��΢?�]ctk��30ɪG&���^0�`C�USt<#�x��+���dq�y���a��:����!GH$��Xo�̭������g%Yk��L�7]ǐ�h,εF������[�J'�J���҄�y��� �e�n8\����y���#o�t�;;K1��,C�;rV�ꌘJ#@��oe�_�v.?_#XK���^��C_���.j��#���4�C�;[{���{�T���l�"W�Jǡ����wG���������ȃhIK���<T06�����7ʳ�N�h�<:��׳�q�Qy5�#�W��yz�ޣ�1���{��<���(�t�&��$�&�u���.��
#�Qn���6i/1@o)|B���ak�ǃ:��M�L!�8��8�PkI~�́x˵����:�g,t����侁*C@�-p��yH�+?�?�t+-q���6Ѷlbf�Y͙��� �6�3���IW!�!�O.�ǆ�ad�X��W��Gz���j���&��M-�Y]xHU��C�h�$v���ŤK{��8�V��>��?�:��b�<��򡼆6�d�(o6�j��Oa����dX���lmF�$"�)�HOt;������+�A��Z�Q�P6����d�㓬W�����sP1sa�ـ��G�s�ܙ*�=4�_b?|�3c0�U9[0w�3΂�Dp2�gO��|�>� �u�s�)���߫�F}�U�8Y^�ۍ���d�CR�5�`�ǐ�%�8Nh[��9�]x�S���~�.�L�;��BR���@q���^��q�:�Ps*�)�w�8���h�L!������a1z���1 ���W��P��}�Ov�J�7p������l޺ ��!�4��<�O)����C��8W%�Ew�Z4��D���ΑH�]������S.�+����E�Z��8�զ����wr�YBg�8�J��? �쵴�ށ`6̹B��m�Wʪ�0�W~�7z�;�t{�6o`�������VUu�z�2p.�"@�8	�o��xyz�?ypU�L�U���D�ޮGt'@�i��;a�ešDBa�A�:$����e�B,dKwR� �]�GZ��4����uk�N����$Z�x���*N���#��1���j <����ϔ)k��8���5�[�������p��)����q�jr_��0s�y���4�5�[���G�eoM����X8���[$�"ɷUVb�:]�`�b��GkZ�:2?�s-���G���c�$^��B����9E҆\=*�fAY	���E*�z���rU�E���N>�z�8�2R�kѲM�����3��!T�[Id�.҅u���C��q�/��Y��4ʅ(�/'4B���]A���t
A�f�߸"���D%�~\H�}�/�Y��<|��Kt���D�j`�B H踒gѻ�ِ���68��	�?e��,R�GR ��(V)K���Vo��7��Ǽ(�@�d�j7pبlE�g��T��|NYױ�G"	��e%;��m�oq�1��B��-H|~�|[	�K�@���2�w�[�/ہ��,t�xt���.ѣLt$"���dĪ�����W�i�%�d��27�
�~�.@�DD��`h�V�#(���F����G]O�c��k��TH��Z7�,}�D��1�>_���v�� |��@�*!�2�����'��_7T	����~����S�w��^n��!���t���%�Zj��{�p�ٗ��Vt#J
^�j,{��PT(�@c�#v������<m�����Os\���?��3�����y$cG���t��D�Է[�T�܋t��:�� �"2���b�bh
�{��q����^A7~���۬X+�Fa'��-����y�ˎ��1u�#����Td��$����a7N�Q�?�FmTy[������LF�P�\��?C��Ȅ��n|ٗ&>��6#�op��l��R��� �H4�&Y��������)�C
�』^����({<�q��{�ѯ�]3����ȉ�t,1�����IR�e�IŮ���	^?ETM��������_�Hދ���3Ve�w�M'鉑�����N�I�1O��uT[��Iw�)�uj"E��`[iu]���HϽ� d� �ל��1��@ ki�΋1�@�
��a�w�Bvg��M��@r�m�I�x����5�NN{�'�OGT�s������	F�s'�U7���F#�\g��������$ʝ�,�0E�t��q�!*�6ݺ�"�Z�B���T��:lU��3"��b��,�cSn,�F}���j/[Ŀa�b��/(����DZ�td/]�3qGecK6���p� L�,ޏ�,Kxc+:�f���X��[�Kqa=��ϡ%�i�1�d4%g���ɲs���(I5o<���U�� 3��du�"���5�f٩*��2�#4��`�'N�o=];���)�����n�{�Z���f�5�����f���u���q�<�2���/2Vm�{GB�\(�_�9ڑBJ�rЊ�Po��>���!�{ꟗe�Ɇw�z��nV';�~�7S�c��P«�X�y��X��yQq;��#)�)@��ح]�������˃��jA�¬�iu�4��9S��;�1ف4]��|��|p8h�h{�H�U�\��6�;>`{;�"ǭ��+��(!R����tjD��s��W�OA���{��y3�4K-�C������>o�)��T�vE��ףH�b�;p2���	��k������N�t�Kw������ga�l&W�ݏ�P<��OB}	@��d1q��k�ѥ�3W��0>�O�ZqGǗ{�����7�R9�_��4G��+�ˀk�3o&���i��\2�S�M[/�>`'����[j��F6�;�l�_
�_�/ADM$�di���C绑��m/�8��I;YU���;
8I�B4]x�Vr�S���8d�T�����c��j�s2��]CҬ]�ԃ��u�9�:ںs��4��ɍRǬ{�U�gIR�����}�@�{���-?�;$���&p�`��h�IP`H�W%H�ugO� Ai2�%����?�=zQ�R~�8i�2@uH��lhL��ձ����^�U.���V4�?6$���f�疛��'�}�#�ƭm�V~Y4����Ϭ�[�#0N��ŭD��-]�u�R�����v6�W5�/[��,�;������ j�\+.z�����%��D�&��P��E���߁����w�c��K�A������w��Ik,+�"/;<�J�9�Ƽ���G��-�l�p�ã��O�} ~�fE'v��tƕ;���LS�Ru��-H`ۧ��%�c�"�U�����3��7�/��j$��O��Dd��rY�
9?N�Ӌ�ל����(
�uPiW��Y+�1U?�V��&��Y%��O�� O��ەO���?�)������R�$c0�C�/x��L�ѽ���\(�e2��dHk a}�����:�� U� �D*4��V���U«_>�)-�{Ǭ:a��X��{��~lyY��������|���M�d�)� O���z��N�^����ڇ�l�T2��~e�(�w��2WM�׾�*ρ�b�[`�: H������ޑ�E�s�0��w��J[����6C��G�����̻�	?^-��,�tFVԤ%�n�G�8�k�P�.�z:m��>�FV����G�Cԛ5��k�t�r�ݷ6��RwKHޝ�K��{I��ٷ��ׯ���_q���Lϱ/��ˉ6�}��z@��Ė,ٰ���U�G@�Og������AeU�4�rg��p�s9���X�<�O���� qF�!ۑ��{o|Wb'�؍'G�$т��nj3����;�W	��� 3n�ӂ�P� ��C��գ�d|<m͙�3�i�ڍuz�V/�(��I|�׷��o���������e�r��:��	i�*b�nn-��J���Klu��q�?��!XџR��C�0xY��@Z�rxX?����JK�&&�е%#>-aO;b�T�$Hx�V)`�����������V�+l \Y�pt*";w6Rо�E|σ�Qѳ<�g���|"��#x8��~�r)��BvwJjI I��վ)��f� �/����H��KT����Qڭ�?��u:-���3,M��:/(p`ۍ��$�׌oim�Ƽ�ߝGD� �=�^�^O�tz�e�,�0+ ��0��B-�H�;
�f�ܖ�Xp@lU��μ�
�$��6ZOi*`g��HO�v괝���n�BfA1Pp���cOb�<,��,�э�RG�lL��q��!���c��i��@�1X��CA����������?Z�)�q�;M��pyW*RG�zw�4V\���J�Q-)L6wR
��%��!�5c=�K,��?�}o�8�p�a�_��{��S��?K�4���G���0�5�!�ޑ�\ɗ���hu�%������X>���y�P�:c��=�7�:I�_��6�7���D�	����%Ff��,c���2)~�K���XX��Ƥ#ؾ�`��j��.�N�m*;��ښ�Hz�%�\�+�^a��9�CR� ΄����8(����&K�1g�6E��/��3�q���O����K�m�_�"|���N������h	yjoqh���=Rh���쿡�d�^ғ��V��\Pj�|w�x���/�ã�˞�A�LL'��ew~t����tG�xН�Lqr�%�Pˡ& l�O���� `�L���I���ce�x�k��pks�6Z��'@�c���b���Y��/��s�<Pw��������r�Rw�Ed��J?,��y���:/4�>�	��
�RJ+csS������'[J���Tz�H�&RЋ��2 c������Vnj�����J/ƞ?8�у�<F��*t�o���7
�1�����) ������%f-�����?y}N��o�ǿ�=+�8�I���T�09J�ێ�$焍:s>����ƫ�4i��6e�'#���g6����@ÂW����1�����Ͻ���=(H�.h�l�N��c�=�.��U�G���\�$?m0������m�	���h��
����~&.X|6���Y5�]�[%�kk�w��w�w��u16f:MirUܬ%���e�|��gv1�`���o�0zy��$˭#Q��ʪ�(��.��٤9�Y
���brƌ������#5kt(e�sV��8����i��y�N�����pԳN�sŌ�b��J`sQ�Q{����`���Q�b~��ހ�1.��fx�N�4/ͭ��Wv5�,�wuxy�؋��Ȑ�(5^U%2�S���a�~9�(���.�ֳ�D�d�|�S��uk�Rd��*ʿ���'��'W�J`��S,L������
���	�C���o!��׺�aN�W�Bq]]{l.	nb|��=��΀�>�a���]f��'��K�g����0jz2n�H���{b��`�����G��ͮ�Ah�M\����F�߶S���t�;����i��j����'�"�">%;��MguEe��e��ꃓH ��s�����i �'�E!MLv �Z,fh%2_ұ˸��q�Q��[�E�b��A��/��G}e��ٽE��9}=��5ВUe8.�:5\:�l=F��s׭&gI�n�Ҩ!B���
�j�Jg�o���k���J���jhӝ���ܩ��t��z����M;�Ta=�ߡ��.(�������U��2Xg!���M�W�W/��/Ln��j����EeOi�gS,5�dA �K��J]��_�.�z�RI���h!\�#�N`�x��"��,���b5ٶk�=va�U9KދW�����Ն�*}�wb]Q�#e��#.��~G��4Ћ�f�	��[�v�鑪j��Kzl�d��QP@�a�zA�)`�Mߴ�ޘ��� �����`��>�@��K�#�u�}�A�g�9�p3�¦b'/NU,�~�3�yG�-���A�X�"�������K|1�NF�v��Χ�nݾTj�
#��=�3���*x�84�^?�O9��y��n����&{0�r1�޸����H]}+2ӗ�@�a�XE���*�	+ ^t��X�t�{}KqK_������J(�d��`h\��O�V����R�[�ָ���x#�[Z|�)�
7���-׭Bv�q�k�Z�EM�k��)�h�{ބ�yp����t��:XW��h�t�#�
���}�$FY�ăĭ�/7�����t��[�}� 3&�Ʌ�|b��V6~���,>�Bp�l�r|�8�[�f��~�>]x8Ԑ� �������>��+�wR�0�Pa��}�Wܧ���k�o�>��x4�=��L�c~b<�!|#�
���C80���:O�^P!]������B�j��`��Rd�ۇ��d� �Q�Ǝ�u^�*[[�X��8'+��6S	��I`����Rl�2�y���T)(ЭX/��A��A"��;{-!�i�cй�w�:m!sǃ��,	9>r�'	z�Z��|�o��&� �-�>�9`�R�55��Y��T��h��/�S���Aҏ.nB���c�th�9	Wtd����Dκ�`��<.�@X�E����C�U�u��]�NE��kr��
Lj<8��ޯ}ğS��M���'>��?��0�#�_�~����$�wm�eٚLD��mS�=�m���k� ���Ѽ+p����/C\UF �I@���D,�QU�����,���&��O ��a%�=;�]t�[�mCZ���D�ܵ���Ϫ��㿅�K���Ny�^ui`3T]��j��6a7�I.�{���egU	i(5���ҹ�§K��N3���A$r�z.T�2�I�YJJ0��꧱� ~g��b�Hw��!�43�_�O��G��{
BZ���~�c�(��vD$�ə��C���[X�(��,N�ͳ^�E(+��(��=m�#�&_T�\l��P���=cؓ��fu�ȧS��d�
��fÒ��>�!V���'�Y�"��[%,��;x�9��� hjl?��zb����c�st=v��]�?ƒ�Xg�f[��n�C�ud�F�>�2Z��eOY��&�n��@�O&y�
6���%=�o��
,��,<�������*�`k^a�����}|/�0�kC��Wˏx�54[j'�qb�蠩��Ȁ7��ё� ,�E�!<6��
a��ZTCL nMk��v��섢�D 
�|���u��'y�����J����>���_��oUi��%W7�uc�V� �Y%�j�&�u��`f��"�8�7%v���Џ�/�A�)CʬyJ�rFI.�H�L�j���&1v���pY�%�	X��U���« �Z�G�K����p����,��2��`��R�9�Y7���p�%f[�ؑ�.f��0�*�'�I�N��RP���� t!!�.$&8Z6p�T�>�����ե�&�F�m�Xܹo_@8'2Cb
�|�Z�C4L1s��N�'P 
�g��g��FTS	MS��n)xr�sJ(|�` I*�%Zy�	�j�xR�i��:�c\��M�	8��JLQ'�9{@T*����q{˒��WL}�H_��\���j��2o�yA��O62葟.��r{Uy�V��`�g���騗ЋҰm� !�!���GD�gG���-��Tt��_s���F&��)�uM��Ym'��'��o���qC�F�IZ
L�&1oдv|�j`���~��@�^���2�
�	���,�'o.����g��>�&CkD4��E���l`����Byͻb��އv�Yh����(/�~?��o_����ޒ�(s#�oc���6]Ó�a�NW<����I%���
��\"�Kn�D�Fq!	�V.����*%�C����-�@ӓ�Z��j&Ss�����b��_Z�FH]X��R��)(&X��̴�?,��9p����+=`���/�s$*�bB&	.5Ș_�Vmq��dA��2�J#2����ܙw�&�.��L�����2��`oU�r][c���mPE��&eCìn�������*y��XA������lB�2W���Rg������� �� ��Bxb��?P<b|?���D�_��5�e�vB�_�Ԕ��>k(7θ�o���
Q�m7K�J�-��?�[i)?B6P�(���D
��UŞ���s5�!S3��Wyv�M���G�|�ï͟ߤ�y��yk���Qӓ��7__�A��`����-��A@�
M^�� ˙v;B�(���=G��re���7�v\�H���"[
O������.	��3Q�[|ƌ�H9� �e�4aºI���q�j���/ŷ��������}�^X�����My�� ���JL�]�w- c��	�Y��>��]��j5�8N�������iw� 5���H�����+�FwM�Em�ߘ��|eu���ܥ� f2���d�x�W���`+=vp�w�(�w*h%ܻ(DM?�a��K����J��Ai�;�D!�>_�ɉmx�R�T0�-L������c��L�_��=�1gd�ܦ��d���V<��!�h�}|7��mb/�3<kL�/�����4��	׍$�����J�4��t�Y��)�'t� �%��T�p�������BÅP���a~����@i�[�2�xL�GGq�.YS<9��K�q���\)�PjG`*d	�8�wP	�����OP��8�~�YЗ�%̏m��T� �r�b/YT����%�����ڦr#a�]׆٪����iߛHU�>�j�(# �]�T{�ַ�/�n�*��qM��lis�55sʢ|�����%��X�������c�5�4�a�n��:����9���wn��uP�U2��^h�y	;_�W@��s�l~���N��[Y+QȒɷ���d+�rbQ�yE�_:m(a��Z�߉^sUق�6��	��Gک���,����͊��C��ː�:j^i<��x=\W���6L���@.K�Y�_�����KY ���S�yv�[��9�6�����<��AI�o�V��?�Q,9=iaz��y���ߖ��(�#�����t$��lU@��'���U�e`d��ߓ)M:&�Dj�U m}ȣ�_�3;�[�-�M�;3Ey��)ؾ"@Q�d>�O-|Z�HC�B�=��kf�ء�ׄw&P�{�ʕ[+��˻=�v�{�ֆ��[ŋ�{k��s�������Bp�zv�� �	i�$
����`�9�Gk"��yG8�>��֪-���7�?.�jG,������W@Mu�M��{��j�`5G���9J�Tܕ��.4hJ��C6B�h�I���"A�I��M�	�.gf��2���{^X�Ee��������́���G2��B��A���v�|I}�O�<"6�G�>=�~�u�0H�#�Z�����