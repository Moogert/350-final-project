-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YZFhzvLnac7LowKyvpgt7XNPoAJR15TwcB0WXKvIm0vFS0AIoC+B0QOEX/hN3ArbaZepjQrwY2aM
tmj/BJuYwHM4J45LhGyvd0wmvCpoCZplr71JEvGcVSkeuBFTJg8dCLNjqxjB2EijtPDXE/RO1ve2
Ti9qOi1jeuwu8J6EboQtqhfGcDvPpNvXub+dmgPPKzuvkrH7VVtnX6V+Dz8zGQyxkG2P4OsZHYQG
ExSgcXtaqwu+mMxFVZbw6bESH64QbHULuLMnQE5SpEZNnjcj7i8y9kNi5zjXdQOvHUQZgS+FVddd
uDcgOqB0q2Y6q+QyaWoAA9ISYBgomuA3TiOK5w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6800)
`protect data_block
eSkf/YLOdrJZfuaapz9tk0NFJqez/7fgFSCCIYA1dDLFNRMvmc7nRfH9K0jjQqJrILxwH0lnB2dt
B9McilDu6Pjv6nJD4jPC63N7Qf1Sos3q7p94SbojRLRdUFxxLU7FVT7N/QWVPsvpmsGYffEvWxYG
ajVDJSb8Kt6E9R6bRFTdqSGm1lsYVXf7maoQmL3bv2N03sP2GzayRH+mIxnDqQQl98M8nEOaErjX
s5PSHERWQzVUiEnzFzb8h+QBCbOMrxdUEUPu5nkgxlOpJRR/qJkAHGvZuw8WCm3WtHsZQiRG6ZDI
11ho4byivef1Bi1EFiQ3AhGHHBsUMuwV2k2K02vQIldPItjS0mWqnbM1H+Qcgql3btAJzNJykbhW
93H5CfnWYeqP52zNB/CmJS8f2BjFsCYvgMsvKL+/T498yh5btWp/IR/LhgdfZcX1nrUwS78ZpJqv
XmoYwQ1klHrSGCKyJlbpm4K8hL6SOYmWuzLsNOqr91UIIhyJfCPuAWTJBEbHtMXf0yiuxgRQnKCN
vNLnyM76HokQ8qZozZ64dzeyYmo0rkQqN2rHqLZ9MkMi1pEs9ALosqvFy5fLqH1BE+Y9RNNAGIg5
vAF4/8/oCXeZU1/Znn4ckq6ix6/dDigWX3qPSZhHxNB+CXZZIbI1LoUSKnZHc2OS7eREewQrpIk7
aZPQYH5h7ru9DgJS6V2YlVOck9CXgYGKf8vg20dwhYa2FNr0loPR33Jesq5lJvBT/jigPA7/Gvcs
wSk8a8MZ/OvYXV21KiA62qc88WglQ1tahvybB4o+tdk442Cy3VYjurdYILQBQUZktYBWvHAblqmc
LTnQ6rNNYG0podOpe/fDzw8qb3iXfsN5tZjVmpATXlEB8e0vMreBLehtsz0CiQSjjfshql+bzham
nqUi3DZhm7Mn6nprM3GUiwFSHdBRofR5NKJcj4RsmxQsxQ1ZOfqJWb9wNmNTxoDAhlVCWOJcy+AG
CaehPX9fwgboRGprCr59nr39/XwaECCGT+q1NWBpe0O1qo/QVg7zqpCDlkyzXVe7ykCa6TzMNZh5
WKuNTOT8Knu36CsEn0nY3ltJCDGo/Sjf5ZJg/NewlYOoCZUJVBPpPoZ7LiOvNT0Qk3P10O4g5Dic
gwXbRJ92Iei/apEXclA7XpIbcX1iVm+ElWn123+D072UhPXV1BnZErQyq3r7DBBeLp/64vY/ML2n
F9w182TTHWvjYXVpquWKcnmkSCdLC5kCicUqlS4vmdN9aIOrFg5JtFyptFkyIeGpXdgXiEbXxiL7
G5HMQKmi86B489axHf/CeEtDYUAulCpEHv1bN6Rr2f2m77oMJ8jM9BaWpGy7aZGKWq1Du6WL1TS7
IBQqE25B05sUS+BTOhbS1yy5vfCGV8z0KmL01it98rllPHFb1FKLiBgYlJwcvrnvSmi3VUKCc92B
Jz4yxWp1aUSPJN8FASDpzKxUqerrzujPOQ/DsU97JKYyIjLsSMKvJiPDhFVuHfCWfJGb0tToHaPb
VuLSCLTPo7R8xfd8HoHYUqLZWcuCZ1GXZ5RhgTTi+20kui6L7/fwsHB/TBK1h8G55i05xzRlqmJD
grSBD3JdbThDCBh9j6in2EGLNq7YP+furh1hQwKHh3ZjZxyQ7NE/+r2GDOZsNaRncZ8dMnO2cCqU
RbI1cNyQ52FsUFaQrG0/L1Vo8zAEZPNzkynVmNK4vz3r/1OW7N4TiTm/VCxD8GIzqlnzT8lUvumF
xaNBZmBlPWL7xG1vpXKYErpmsB/hzmaRyWczdsiEtEaAaGeEvznsi3W8WME1vIEb+OIgadeV667i
AzGAv4QZFxEljpajnwPTfATfeObCklzfeeoku4kTusUQrtQN8LrOOGRSUB+m+k+oXoetWu9arGKB
MCXIlfWGq4S3Wo22IARZJ9xIDQWtx+bDsU+YZsBDtvYvN6wpKjetNa5j4t7qbNUDqc9za3ZEyjOI
wyZGd8wr0MuCnvP7cOLaohgmyRdCY3kYtmWEUWUIwIcrZOWlgI5KGFShJdc+K9/rvkD2JXeJdvOR
sHcG9CLJ5cagz9FKAS7+MmkWuLlltWNFUxiXGcI4WOJgsAaSLToxBkQXgQYdCLPtkYaomNWjFZQo
jlJCwnlrJvkfftfS2wxUC7NqK5j7lA4iPNrsHX/c5KrFQdCDKN0PRwnVuUb0GN1IkS/dvugojAqN
/W+2oR1z65VIKJucewOPqVmbo+DmXrkh9XgDYkIjqUfYg426duzRr4DfjB4I4TR1vYFze7V8wb7f
wqy0Ly1N/JwLowfjAlZrnGjE0hsAQYLhIIsEW9iI3MAgQAmVR3YKm0EHnreAx7hBSIsu6MInT3j/
ccsE0FYF2fC9ocZvKcY/+Jo8P5tGmn5zbJMbOKa1+wvxTgeFqG8W/fHXm47gBHMBBb/BFG6H1XW9
cll/d7mAY8wZ8lfiRcbOBZfw5EuxEeRhIXDPj24gAMFmo5ggwYYUNvcGqMmfgf5gnfD1oN0ViJ1q
XKTogD//rUGj/ARC4TCIQ5+8FUCyMKk7bN5L/eI8mJ1AIgANavtdZTWRKQg66+Vxh0fDaTW+5TPa
OQPXMuwQvpqFITBNtkES4qFV/Tm7yAwCaD6TkhRjCWdOvx3plgT9nnpPNTKnAbzzD7luUrG/HzFG
uvVoCvRbL9yd8pWhbGw2En/FXSzJmrKUFdGb8n+1YIZBFVdclxe+Ej4lkxmhJV6KJu8VcOANJK+s
2ssRWTwuyhDeQg2z3kvgUXcO3GiTs5/rMnChRrZY0D8m//3WckAoLb8qT33QuX5s0glIb1iJTkes
dutfr3TzZ2G/dE4w0MGLW90I/fDf7gF/JEQFg23uVoMjCJltogxCPeQ+b9GDAcEm71kMGAwBx8Ke
LCVRkjTbUymBqhhSNdAln23ejOVQHIrXSyjeukMANHa4FVLLKaVdQRXaPgphWNsx31+Ur0Wt6tiJ
ZhnoXlXCku/DjWD04D7vu3cukE9KvNZ5XmnuRftUo0/JyxVrtXZCuzamf6P4/DUmUsqOYc+V9IQO
DFJbX41QpBIXLLdaftoNKeHnDoY2a3r8CLlVmKiLSsztfUKvyzIuu1fnk4IwfOI02LzdMXKu+jRc
sM1CWMj4vFhkW4pWSXEhGa6AozhrOaFw/CNH88V4MAFRpqtUzbA/N1duLU+MccX2WW2VBvIPLOT+
ohc3o2hIM663G6O5giV6hhTdKkOj+MuSEOtooUQyojLtkV0Nz0gSE/f1k9GzUBTS47lEGaxxQPMi
/wtxAO8wgLJe4x34szldXtHx4Qwi+XnDbRLZr1AeGLzu71PmyOKFYFH9HlHhA4RurbWPA+4K0GXd
mPpp26PcGw0G/6AfJ69JwviEJg3/vXRd5JwGyFubyXnAD//ceg4mvnRkz5JxBYj3AwISuVRFzi6t
ukNzD0UNc4lX99H/5EUeVipPIk4NPJD+0Azdt3DJcxITX5V2A1U8Dxmue+FxU6tiJGggZgRA5s7E
+gKGetMP2B8vzBT89hx/kel9s+6X+nN0sXIXqU5j7VsKCY6sKFobT6OAnRsFDhsGn3ARK+D8KGRc
aWb1fpOKLcg9gaxY7yeCOKS7sm2iej9ROFfgWsY535K/5tehupTsD2O0Fdi2Sv/pWaiUivxD6OpY
vDJ02A6AdbfRFqaMK1ebPL2tFPv0tyXHvQqHu4BceUWFTGG0bSwIiY6p6QJBvzNlFSo0oyGC4WDi
gAfnf1S0ReC3VPvCS5OB6Fdb0YeIiUf9n3GfmIYMG3SnOuNus+YuiVp+/I3afkNj9kUSYkVtUJPl
KuxsIP6lh3dP+P6Qpf5pr8pYBDUKetTLwos+4Fd5xrPfE11zWKXjUGCDpRgLW47GveJ3Z0lkiqHS
afJyw0ypF98FT6SvjMzSyENojHIdxULWUiABQtbt8b1W6ucaYHYk2pjJYMbItVOHivRPrKR/QXEr
Vhg5hzjV3vh0d3zU2SjtljSYAHKyNESxGUIdUokb+h71RquglYHiWAVqIDPpCsbWiQKNXLNCHhkd
vD6t+Ta9CtLRvTa0lvRDbzX6l5q8PMVSxQylWxpMFQNy3Nq1NnDyCNztp/jmhnkHwNSZJDmOs16D
85pqfGhayv2e87NMkzLqxrRC+9MYGQDr8KiCHYFu+2LmgcWXUgsQqeKL5k0X5xpqujoFdvH3Kx+8
ju8po29jvpnfYnZ/trjbF11D7lYSvR1UPNmEX2is/qpy6En0tc2nZwW6H0FF88gwjbiuJI58VC0D
qpMP9jYKXRJSE8AsgVfg3HHmjjxJQYyq2W2Ml2XHd0uw3Osk2zfQzteqWqDWt8iGvbCtyZii3gV6
u8+Wm89oAusJTzZVYVQeL/kAiunWQrCBiA5yjPKRzJeWKWxpCyLtR8Rtm+wz4vzXH194NvlD/zla
4qXYJbneP3P6A43ptshzS4okV2l1Cs5KoICdupFbKXHP/9kbhnPGVjX342yps8uDfH1CH1FG+VwJ
9rD6QDVN3tT10QxAoaSWgKbriQdUaFzUQRfrfbBXbb+76uyzEXrIHhjLXs9Lo3zGI2D/uvmmBtOl
OjWUrHNHWtea67OhuaF3zHIfyzfiJsg4EhfaUSNxVdD2j0MBu+a68EDlYNjM/EYsGKWdkdRCAmyb
whZEoAKcVT/K5waKfEvsdCLqfgRXt10yhYlmoXYxCDUnx7pyS4eHHIxO7q88qvYAbYlLCEyUawVj
URmygmC89Ui2bqLudjhK00dRe+pMRDMEzQi1upcyvIE2FBi8nTWwnBsM6gL3NcWamHS2QE/JFAug
LBNSUlV64R5yiWusx6hYSletdpXjTElPSzZquRFBSFKvmk6T60B8q9BzLDc7eeELHY3cCaa2pKp4
OVCJMCmCh//N2iqfQZOIKnI+Qxn1+iieMUv84oMLdU01Hg+qFd6tfnIJP3zcdLkDJp4D+vVB3dWk
ohUbzthMwyr+X7//wmn3LQinXi2uQm8tFOMc0HI08UAp1VD5TGz17nWPls029aNQJgioHlhpuLGG
WFYTP8TYU0akwFhsApVYGvqzNODgVj+tbsF8+b0DUq1JqSetnriKZ7b9+gs/kgt0FC7QXkijJFPW
zJXo86o8AYZyLXi+ne6GI6jWUCe77cTc+jUt1FzRgdx1RIuf/6OdrxxZ/l2owu9JhCe78h/8dCLZ
QPNSkdVw8Re6RURXc5k8wOVe9LzohMCiq+ZiYjRrYwkUjs+T07DO0MLF8KnL6Lw/Y6IgvjgH4RGI
OuCgyyJeoV+n2l8G7bI/+juEJeYsVjDg3dfM8ZI7i24coXKPU++VN50oXCW+aS+1gkBbgXsXBgpd
hKcvMtp+XwzIsepw3Sm0HImzPY12gxY47Pgxq+ijOYLNjHscPpp3X1mNla/D6/WRAqVgWmhRBbKt
UsQoDRO3QgeMb1IiObp/+mPRolLTUtTTkPIK6ErV9t3MWlX+VzeVEUOxq/3dgpBR+fUw2vby2hnF
xugYHhNkQugf93zpw1d77MPEabX/uiYGs0qXiTfyn/pii1/QHEvkI2nDjW4YbvKRkINTydLmIrqv
DLrpNLNdD4yG74lLsEgHYC8oNBDahjPhnUnVQEX6altRfLUSnFYIKdj9+QqxUkDtHb2VNimoUMy/
kFSZ58DUc0yiy2639nUBx0uOTvPXVLaheJQavqC3ms36RjjR5iP0OSeTRywa7H1gM6LwEmTMplZB
McwMwLtfAWBNZ+4V3yhDULLNoUpKwMoMOdVgePRkP39nAhk6LD8WKd2DvAuvjHUApoTwTHwm+N8o
OM3I9mhpLtNKBs1JmOkDXGiUZc2Vj0Fc7UpXVLN3hkoiU0FAD4kOt2wUYTQWtP/vJVLMTM6P5A0u
rfPAfoy7Ngoecmd5x/kKtShzQNigsoL3wScmlamZn4tYCctmUIkTQFptra2hdzONPa0aDSIHfopc
bhufhHk7MBOpgccDOMQsk8pmm/MgbZJ1NYrFkX0iQ1R08gDPRNKgCfJViPSyiuKcE+xA1P+AUp/w
ghg9lkP2A2F3Z+XTRXJJ79Am/PQeIzbL9pExHQjUeXVnr6HRuS2EvCiyq4f0Xy2xYwcEldc3QPkd
3TJGORkdBOOAougOpPpEq1Y4ZAccTSvNnbCe3aEGQL/CVGJ/fvewmTiIjLFOmJ2RUoVOEoH11Tiw
HyrzzvayNOae6oRNpPTJzUKafg9pn5kmnBEg5BLE7JptpRPbra4SNHl6i3q+xGRp5frh9eAwmWXH
pJA5UTwhWLzZcd5mRLYWovwgUVO4KEWjUSjvnzqb7vg4iig0TKHV1mpyZXbvKGWuSO92j481uJfr
8Q10BpGZ/ncZ4YbrkhlS1kTw7NLrgPAX9+Zdff1Z0XrVBeWFIVCzIviLmgu0xxErCT7epcPj0Szw
u4nYv1nvGwIAlX6n0mc7oUltCDPWeAUko4KKSKKz+7tcE+/8a2WdhMTT4EfcTYS7GY+MdUQl97HT
lBsUhW6bGvHGM+NdVTKLqNl3xYfWZB7V891BSmuxyCYa4oaY4qVgcM6s/kXm17UbOksbEdnvujKa
sSwpSrtmr6n3tFvaeFTZqY3oryCNhAOoSfG7LleX3hwNugJdLpWifZw/74E0jdL7oGOCGLraG30G
gEdLPgTsRXukWJsGJ7pf7Hjc+w2AR6lJwtUDvNdgoellLHNRhyz+LX36rFSePmZjpG5DQ1J7LtaJ
wPkdUemH8SYa0fUPB6wdLCabBV0+FNOyW4hvnGkZnNxedSTkpRW/1KXD0KqoOkP3CvvuW/KzSmw/
oidpjCPwNUNDdgQr6VYG102N3grGWFZoD2FMh+83JScOToWKU+f9kN3Vhm64zBG+NTakqWMydwAf
yXyxTGC/c5YVK1B7oEA/enPrw2ZPQ1xhRlEHEviWIcWRxWCNxVFidPNniM1YjoaV4VKs9c5qDdTT
xHujYpG4sMtvKHuMO4dL4L1IHhUFAqqiAOT5CpDmnk7OeA3PTm4Fp2ef2BHaPVWEP59LSUs2P+s3
aqkn70QlNBe4GtCPUrpWH3fNIwIX3irgVQJAFVJS4+GvJgqAQwa2mETPzjeRTJ4AyfujsVr2y6Ik
ZfhebbKpTATEICohq51OeExsbFiFW6mpRmw7R6rzqGnwIgqQOnbgBzieKl+swWd0oinKtO+NLhhS
s2+dnMcjjcMLWxX+TTLkeZ5fJNdwZ6VFo9NCNYQNgXD5Z6ZzLdE0hEsPfvaOTLM5CPB9UNh/rGAR
6xN+bQgRXqtSdPR7ed+BBhF4odvNvcxvD/TOAbAcxJVSDTxxtUMBlIZOxTxha4e2Q11g/i9NPPD4
xbpPqc/mbDnZnNSa3SBaE0IvmHfDsta56NyL6KXBOmfBW8nOSqq9aRkx9gh4qAFhMjF9kUYCUUFr
6SfcnZkg2zAN5pSSIS+vbaS7y9hX4uMcNRGxOCEVwq7fRG9bJsQ08BTktJ4gL+e9G+y5aW5Z7uX0
4pB7cCy1YjTUi/Wp6xefZg76IG6p7N7ZGthywS9pwC5ThhE0o5x9Y70ALvrWsoEUOOsCFTtu4Td9
UGVnZS3Dz3DTeJx/sBTXgUOt9LFMNDa3ftL12zspiXPmqfv+OzTFLbAjk5uv0A0hVjAaZJlHNTeo
Zih2XWHG6QzJi3OxjU3XBpDSp3FiA5SLj8tAXTGqG1VfLFFTmgNviu4C20JrW1uj8D8JRYIoN78a
SEkwYuI4b46WiKMx+b0fsBVF4XWuu/XD0SlFgxQ6CTiv/BI6UBg8t62mqYB43G8CAdX6MmMENEPW
sW/dvtu9AyjVH3kvlefO+BBVYNVlbVsIf8Y2eQ0L5vZCPs4nxsRl7QhlYwohqwS6i4oPHeKsOZM7
qIjn8fzxEPp9p8c3mErDBH2Qh2SzC3d16poJw4kbT1btNRSfuFiTGxS3ZBPot5YkhJYbz+oggCjI
IKbwIJ2WjkCHNXsPVYkkEYW7dW1j0TEMXJUUnejsaqBY9KUw08Scqkgd7E5NM5DpDzzBBTKl1U+e
gfLZDNIeMbDlp+hD6NVGo92ujm5XIy+ffdQzgHwPi6tYzVHLbzxWDWpyDLTi2KJCfWP98X0lmIpk
Z0nypW+Uh8l6166b/lMH3aydsMEtRZs/ZWbXSMKeYh0+VPNgecCMlA3tcadsKMHDON5r613qfTUw
sBULRLW4onyqeNFyxhf/W3xT2tffhCNUenIDAXWN7dfWUAsABRfbn5Co9M15+5KbfnYEk78mrnUl
+LxfpakDNlTQf5niRf2j+QMj9zZCN/PhEB2sium6334n9O/Iypfpwcx4mtmiHUWBKaOAVlRni4m9
8aREYqoGrziQzLkLUjSFj0bXfHMtRiNChcQELvGUa859oou/Kltg5YMbPCGWbQhwYhcIBaQaEqEy
EcOQQFpNg8TXKEIgd7Z7rzi24/zAsoDj6WQoQakglD+Uzr9/T9CZ4BiAOIFfuJDfOLbI6yx4gh02
baNwu9fRFD9dBnCUWkwWlDMzkKVc8wOlA3MsFasxAre50DHIeiHNIWuWYAIKkSpPjpwl2giwNYVK
JFQOSmoTJVo/i9QyIQ2GpkLy5z5QDaVakbERsQiZe0Pils9zDfZkV90Xad8/gkA5/1cd3jx1xp87
q0UN9j5W8gijDlL67XStOQkyVq5FnSJHFMXKjIXgYGxOCfl5YYggRT+Kq89xNL4vDk4n9OVw+mbe
LWmtY6C078J23zdd1ZkJiL/gASKt6LpVlq7PJU31wP7PFs16nvvngwN9QwlXo2lsXFVDg2fp4Zvq
Agugd6eWN6YgEuhkHMspjHLygqKpePxBAyRsfCF1icYRkIC81LsDjXT2a25cQKdNqh4w6rdsTtaN
bSUFCosmtMhBZvUs9aHJnHvhvML1HJlwkNcGJVWAt0iRLrKLTbReUqdEwuSVyE0xB8sGdrQFine1
As2AZWK93YCfjb6eU83Es+1Qs6ZAeqQRLhV6MACWZKcZZyQvsMhovQmAMkWYAR2VnP2LSnTwdbUB
bV8xzOAgqEjLZ+Yaz76NV9WbOJfbd0S9LlQ5a9O5JmpkZ/toRDLKRijeRgdESbHJga4kFKlrasiB
3ONjhZheXK9qu1mZ2LXHQY0=
`protect end_protected
