��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g�҃�f	��m�T���ƌ��"�C#~������VMb#�X�f�����|b���e���rQs��~����2����؋��&���K��٣�M�*�h��9�1��̻����d5!`�S�o����@Η�I�]���<N�����%F����0�8k<��~$��~!~��dV�Tm���s�@����Zl�U|{G�-?ҡ�(�K�ll9:߷dW��'!��ܗ��W��w�#W�q��ܬ���ݓ��Qy(%8jZ��{5�k.X*g���zۿ�@��S�k�!��������e;�����l9�&�V�����(�0mJo"PE������טf/1ه;�3���/���~3�S���8)�c�+�kO��p�4�Gu��k��gĖ��Ŧ矯��)��(�Y	��q�����<V�'*�o�����eD��b��6&�����Y�� �G(�g3|����]�a3v���t�\/¿�4��4��܃�G�_U'W�1�ަ%��K-7���Bz�ծ��@������#�VTRK�{6p�U7:T�k�
:"�!
ER�0X�R2�$ �X�̇
�6r@_�j��舂jU��㯓����Ê�/"HWC@�w3%\f���b�u`z��D�z�iH��m�OJ����,�O�1�����Itn9+Y�J�m2t�ᦺ�LOaLc+)������$���Z(�ߗ$_�l��:���>駗���cv���8L���tS}M0a<�d�0��#�B#ݪa��z���b�q�V�H�o @H֔	��#�}���?c}�O)�x�J \���鍍�F�f�[Ef��I�?�z��N�PS6 ���������N�	,5a"��5��dB"�V8����a��&�Z�,�?�*��`ظW�fD�qi0Y(S��̧�7��=�«�9��������O%9��+䓈�h�`M�,����I���C��� �00��m5+�Y`��r<1\{/r[��թ�
p)(��7�~0�ɏ��m�ڛ������C�]ũ���b�앨���#�y�%-i�$kKȧT�:ue��n7Ɯi��~�k��~]��t�2$vM;,��M�����xW��^�1�� ݵ-�8ըiFO%&ލ��'ǥ��܌6��m���Ϫӌ����p��+���Y1|��c�����?з�i�UH?�_{Zԃ�oI�a<ä���huXI����JSp�������t����%(��˝�,��I*`e��S����B�)d�d'IN& ���@#l�ɟӯ��>���K�*�-�r�������/Y49�w��e��s������Z���R׋��ٖ�Jfa*���M<���Xp�@�1 �;�X�,?,Q'�9~|ܙ��I@�g ���.!�����y��x�x{��.r�	��D5С�p<�����<��?-q'���{hN���:ԔߝV���NI��H#r�����n�5�b�������=5A���}�V�tΙ����Ϛ}�>�<�5ِ������Z5Q��� ���3Ѹ_|��å�}�3�22"h��UŴ�R�^�M�sI�I�n	"�a�C$�UEh�#_�\��F��P O8�ɻ��Y�f��;1ݨ~�H�ӑ� �����R�|��th�p+ܫ@�;yƛ��@�E1�e��RBH�lt��🳞���s�J�GEQ,.��=Lt1�w�RO��gЯ�w�~�aٰ�ɵ1����&;
#6q�����T?�i���JBq�g�%��&TW����{F�s� �%h�C
����qy��<pW���=V_��b�f'�V��������;�/��Kч���4��Ʈ*�ֻDL��z���4;W�f2r��\k�z�I,b��-���U�KN4K��D�w����PE��-�\��JB���Y�^�0M����}�e�|7�jX��;���)�=�0<�@�����lF ��X�`�8�q�:��R<�~�h��aE��be�(A��ν�`�V�m8��O�)��F}����ji�惡��1�����"�ķ���+I�fسJ>�6�����TW�z��^G�t�����Uu�]�6!��mh�R�~�pX�4f������uF��'k#�s_f�6K8��<㕸����Y�Y�@7�'f�����diC��\+.9�Ӎ!�uh�6��_
��(j>�Ƣ�3q3�At3r���i� �?��������G7��{����[�zG�m�+1����}c�_��چ:$�S�7�:�"�WU�%q̱�[hz��9�2]�M\�&�
�5gY���(\����b��`�p�0�xt����u�h5�E��k�x����uŘj'[�������P�l����V}EY,�PX��}C4�h�nN#��`'�^���G���ǫ����'�ێ}�C��^��\�҆����2�n��oP'38z�b��- �����m��1�����!��_���� �뫕��C�7ŅȡxW���!�p�`�?m��7��
�f���U���8��"��T/���&�C7��	Ҋ����(Sf�$����)��K��*�ݲd�	�Cg�IT���޵�������3�(�l87�~�t��9`׷d�ߡ���ZXѫBL��i�!��@L�4�������$$C!���?������u��;�Maֲ�5
��a���B׺���#�M��@p�n�3��^v��ԁ�W�d�8��i����W��70�.�����f0��Z}=]��h587K�Zly���_Sd%�vv�Y۳�|u�ɬ�{:���l9_>��^����ЩF���\,�[>��[�4�A4j)�H%��z`՟��Xt���{��������}�[:N}��؎�]MS�H�#�C4����Pȼߔ-���5<-]�_f���jEyi	�+trFA`^�QZ�)��]2��С�
	gu��3�})���y�7FY�R��i];d����U�S<'��;�S��%���!�Ioz\^��Ӈ;���풛��K,{+���;*"�*6UB��ஙc�aq�gWe)O�VGj�bJEU�> :���V�M7���T'}�h~�	���:f�e;�Ar���5Q��ş�3����!�|Q���,-SKh�k6�#��{Y�
`��
��\�C���iz����C�t��#,������\��g`��`�(�o�Y!��Y�?J �j{���� �I�G�$�/�r���7���>m�9�i�L������E�㮦�; ��5�11&��5�~ѷ��9saqvƺXɬ��Qu;u0@U]�S�9�o�x/��<�֜յC��Z�g�E~��#Q�SU��\�3����X2�����ō���,_�qt�uɷ!8P�!�p&?,�����\�#�"?�>�������i��OQ
����3}��%����w��ބPܦ{�e���oSN�Z	E"s|#�l�ly��k)X~;�C����{D�V��_�>�{�:B-ԣ��@RPΒ]}�N����q��KK���&yV�Q|խh#��,��C�(�o�e\16�B����-��;N6�x�(��-=/�.��[��rJ��eo�<*Dǫ0�3ֶ���J�7&9$�ׯ`�L�����fӠ���g�/,s<���L�	�Aoe�$�9TCͱ	�u�Q�kD�b:�h����a����Ae��T�$��6D��0�o%d%�z���.�=L��/�f@�w��(q�t����Y��1=J��j���4a<Wct��om0c�l%'��M���$&8��B$D4$�¶�Q���x|��Y��8�t�oK��ծ <�얎
�Q�-�Fp���x^��Ef/ِ6�Q"^�2,]�i�)tE��!!~�@
�.�u�U!�;'�����U��|�����J)��e��N�`�a�"/TE�iR��}�W�Tǌ)n#�[�>5>ɻpu�#Ą+C^�H�8;��&,;@��,v��*4'R��{���sȤ�9�+�u��>.����O�sy�d���!�<��=�C@����;3�S�kF�cPοR ��EN���[My�hW%��#����azEc �,ϸaJ95?q}�?A
�C쏥-n��D��h�r3���.��#��?�������,�\õSR>�d�d�)�7*z�e~Fs��m5���R�=L$p<���������VO����Lh���'���a�ph�׸k�݅��:YR�|���9�-�̍_��v��r|,\�aIZI/�X.�MH�(�ֱa�c1!<?D)� }*T�=	�� �۽�-1g�F�<�	ʜ y%�[�\�]�_�'�_�$Mt�0`����,M�Jǃ��aZG`����h4^Y({���Mc,��m��_�^Kl({p",s��¹+��� ���F�ι1��:-�r��VӀ��1�1�j;����Pr�#[%4}��]ݚ5��9���;]���|��=�����ݯ�2g���p�P�N�I�^rk���声��+��i�D����@F��ƃ�O&�E�k�y�Nuf��ԅl�|��t�[e�����F���9�w˚^���m�P;�;�@oh�>�U���������B�H�I
�UX<�qP&������.Xj�k-�a{P��N8� \�q
�@K�c�a���O��IŤ��+q�U�V�gM��$
r���#aR������^����[i;S�y-�cf%E���*}\��m�U|�M� U�̋�6�z|���CI�&�7ԩo� 	��P]����d�'�0G���[IXR��(�gR��˧��8�Z��io|u��8q��`�7I}��#3+>�G)�T�Cų'�fK��Q�JtV��u֮��6��3�̛�?�9"�O�*�9��w[:���=�r���`T�h��Y��'X]mNU&����aEE�Ӱ�w�T���?���K*b"�)ίF�Q$$��?DaʊO��@I��f���ġi���}�js�>�Ϡ���w�x��*�4��v���P3%?�wIʒ����v3�}�ش��~��ؚ�j�N�C��{`�@�D^p8�{^ݸ���%��G����"�w�h�}`DҖM[���ߢN2�۱�1�P:J
Qޜ�d��Cqڶ�"k�L��������;R*fk�?�>y�
���3���E�
(\�+d޿��2
��B?`ͬT���w�d�{3%����цv���t������p������wz!��Z��iq���������[��l�9��cLĢP��?��x�f��'��t�e~M����2���Ȼ�@ai�Zx�E�0��>鞵_�;*�=p�� �ᨂ�z>�M�S�z�d�Ϫ�ָ��vH$��Q���c��*��f�̞��#_��c�&'Q��3�+sQԒQ�z#W�� {���t��Ԁ�QY����#'�k�T4���Q�Tlh�|�Sm�Hc�/���W> A�	8T���@��|k ��:�~Z%�|�D5!�i�6� @��0p�!}�؆"p�"� ���l�R��it����`��z��U�S��� &��x��,$�sל�C���i�ɢ!��,�	�- <�1� /�ޟdm;/���m��;şFk��@��Mi�D���-�&�I{��;x�
�E�>uv�ַ�@AAM�_!6~�U������%����e�`^kEw嗴�����R�I�ݥ��)}=��K��"i	'b���$�3��`gfJ�nU�%���^����^-L�f
i�
�h\졒���wxNz���P�w���?�o�J�4-���;��-W��'o��]§�����&��X*B������G�b���.�F1 HKi+8��b�cG�H�"��=�C�g�ܷ}���3����XM�n��H�bX����[0�)��.�������K��rDd�z� I�Piw b�CNřq�O���/�YҜ�!^�� |ҏaǍ}������:^��<w���#�N�j���՜J<\�-È�b���n���9��sfao�"P��W\��դ�dWͤ.����������Fet�j��׷,��U�Zw���*�6�$�oC��6Km�)�T1�RP��O��'��6ے,��T��&�P�Ÿ���W��Y����H�N���x�^�I(^�+(Y"߀]'Z�p�����=�rt��϶R�����ۻ4ɖ�s��J�� _^z��Z��X|�o���������kD���ʹ�{m��6 ��>�/O�uO6Vop=�-(�i��'�c0�ش���)�Μ$4�Q�b�Qi&�	���֣�8$���͒��ͪ��at:0?x�X�=U.%|}�eE��i�)�%��E�7��a������|����^ф��S�p�ֵ�cC�rt�dz�h�w"�4#�j.M ��_�GD���4G���1%k�B�Ek�
�o�w�$�x���)���"'B��l���.ܼh��P3,wdry��K���(��Ke����Ƶ姿�-��
a�� �~�J5�7�(�P�J����L��a�_���dӑ�oI֋���'�iq6t>	 ����x3M"������3��~D@|F�^���}r�=|*"N&a+ W���^�Z�����!��^C��}c~Y��^/xm��g~(O��=/@�>Ֆ������Ag�zw��i^v
 ��8�u��r�~��}ډ,���o��T~�&�QC�F�q�a�iE�o��r-�_�#i�|����E�i���(��廣�5"�xK$�fs��\��s����¾��ɂ��"��oE�J-��̂�<���)��d�����$�g�8��4�**���A|��6"Ќ�>�p[��"����&����Գ~��v[����L����u���~ޚ_`T�{�$�	���@D�&�k@u8�H�D��v^���N�W����������sN���0z@q	E$�W�Е����ʾ��ʦ���9�5W�1 j8d��nd>B>v�D��'�\���Ēg�(�/?4U���M��=^2I�JN�G��Y�
�bM�U�c�XJq����9��M/�.Y�;\�L�eED�7���B�8>��)���$"ZÐ���x�✕����s�˥�s]�D�����4���w��#�8D�SU�Ɔ=B�aH>����Ѥ�pX��c��V͈Ź�����hc�����7)���H7*H�T�Y�S$So�2���uӋsu[�5�C4���ʗ�6�#'��_$?7`c˔}�h���rƯS�B%�
�r	�~��]�V���p:�������"��օ�Q�^�e͔��������k-;����_��t<��1i�t*_h�`z�� b䄀k�Bt�Iy�N@]��E��,�'�`�W�Y5/�^�r_�B����VWy4��@��n�zH��vrrp0��|����sS�.�{��ƅ�6�4�n��k���8W�M��%�}��}v���s�T[u*V5	���o���+�:W��sMw��OI�
Sҩse&7��!"PYT��'�~��.%9�[
�K�#��dɲ�g��`=�F��s�bh��A��(�3�DW_�!���l/���jNk%��;ru�A�g�"
Aa'~ѷ������!��!����4�(,V.�IͅV�K)�*�D��LT[P-D��\������s^y����:U|i�^��k���@�U��f>۫�wK�{���G�/�%)��W�;����.}R\�pc5t�q���Y��J�x<����� �L�jx��9\3��ےIq��ɹ�0'��D�e��,i����Z���(	�i���َr_A�$LGx��3�ܑ�ʱk�+�l�;6����fy����V7C�B���ډ}�>F$**j(G����l� %'��� PJ� �0�(�*�������PC���#�n�q���6��v�~�%d����K�m?��!J'��4?7�e�����g����z��?B�:�`e8�_a�8u�Z$�y��g�hڻ�Gt7& ��l�Ö�4�:bI����|D���D\�F�7O������ġ ;D��0 g��A��i�����-|'p$�Kh��W�'۟;�2��y�����@]�'Y�x�Z�̠����JS�q{#V����eU (�'�w�Z������m�V�[&�c�|)�%��?�0�iS󪯅ॽn�YO��0�� �Y"8���֝���-��ro��i1��s��7tۆCV	�v������P���2�?d9� ���y+�_�g$��2<ڮ`h@(�� L�;$ɺ^��\t��X4�	�Q'(w'ٗy�c��v�y�<�_����w��������jI�?��� �4͚���>l�-B�|�-D�����z���� �Qm =P�&S�j�d^�ݙB?oBza3>Q�
^~�����+�_�Dhu�,�VnO�u���.N�3Z����4>v���9t:�u��%�W5Po]��t:���G��9�\
A�!6F{Y��1�mi�rGd�j��R]�Fp��U��p�22<����oeH�ŪP�ᗰ��@����@Ǭ����Av6��!g�Μ�jJ�d��f�8��0~KXD����z�XV**�$�L���ӹ풨��4�k�R���+!�ۂWe��#^ZfR�pZ9�ƹ����*�:���&A�~]k�J���Ep�@�жBT��u��6�~$����)�T��DAa�Ś�Мp�� �]v��~��J��=m$K1����vͅJ�r�Z���;W�Y�<	H��F;�T�)xuj���>]���ܺ.`�}��Pm�Й��t8*<|î����-Z���eu�!�l%^�*���f�s����y<}zZ��+\bt3 2�A�Zm�6z���¯�@~�u2L��;���b�/#�oI�\_�k*#�{�{�@gu��!=��ؘ��=:T���ݾv��V�<�͓��z�	���{/, %����=�+�ZIERE��&4����s{��I�/8���}E����o�ƞe��U}
޿��J'p�)l`w~N����A��F�[K�z�]/<qLv{�(��4�J�L�*���QK����t�?F�+X�z�*����0lӫ��\G�����u�� ��f����^I��x0�6����?��2r~.X
�V#�p^�(3�m*�ǵ��q%�v�|� �C����%Z�oh��O�D��J�S�h������ѭ5u��]�����f����h�l���V5nE�H���Dd?D�=Ҫ*}���p���j���p�w�HOD��)�_��(��էK��/��z���)�'����A>�d+���TUV�Ȍ,6U��ĭiy�X/��-*��׎iTsq���<ʽ��r��ܼ�ZM�'2���"Ч.Hz��F}>;e���ᄺ)]�2r˿���F;H`ؘ#)�N���8��Z�R����cRCh�%0��qvf��	��F����e ���ڈ�co���H�+�����	�/��W�W*�s�i_oK����3Vw���;��_N���PdΪ9�
h�^��b�tH��q��� ���M��V���DОw�iS�9?W����T�1_�8��1-���B�I߫L���=�^�UH���X�1[F������nNۅ���ϳ�
Ap��Y0���D���EX�Ka#���T2Dֲ�kU�z�ʄ޽�lХNN+E�L� ��'�jXZ�B�լ��KZ�7�x��|},s8{��.�ҿD)�bG���\�/Ò��H�<�-M�D
4�=��4�t��~~şэF|kţ#x{�6��YA�<6YJ��,�e�*ٹ�e�	g{�MBڻ�ܟ���g��d	g�0���	�F���oΉa�֠�U�_�V3��4׌����xv��甬]�>���$X^�����Z�5�i��ͺtK"��*ZB�]1�)�+�� l��c�[/s�y�������k�_����O�eq�e��{��rǞ%����YSC�yH%*4��MC�!
kf $�<,;���:'(咞�Rｯ�� ��r����
~���F�MBO\�*�u������X!���n�bW��+��`>�8��"򻀋�Z8�{��_�����7���X����-���(B�VՆa;���M�*�&F�C��3�����K���Ɲ��E ��Y�@P�����}�S��d؇�r�������9��	��R�R�e�+�?Y^(�
a��źor��(�_5^NVW�n�k�X��]cj�|�i7Q� ����2�8�IN�x
N,?�Q�俩MvE3��t|1�PS�'; �9�WAL�'�6��F�|M�jƍ��������<�a�Xp���3;P)M��2n�n�ePD���u���X�1�:�ZN��%��VG�53V�h�B6,��?����-&U���[������n@���R��A�l�8.�/�ivC�T�CK�zn��i>Ů���L�@:Y5�%\c�%"�-X�.x�2�3��_)Bg�{�7���E�<�_����I�3.1l7���h��5{@�7���5������y�/�j��������j���@$��P��/:�� Ղ���tv�V7s$�����t;a���Ψ�vql���X��;:�[�j��nJN�I��Wk���2 Xw�!H�8��zaϏT��K���b瓲�ݜ���_6��$�D���>n�:�,�z��!W3��9�C>Nجʟ]l'!o�y|���I  �99 �T[�u�(L(��lF�f�	�7{��o��5ԩgs�l���ٙ�N��FY%VЂ&�Nm�7�M���H��3��(ج%τ���2�&��`�%�9'˶c���T����+�%	l�����r��q(���"Iz �.V=����֙h���V��"'�Da�h+)+���,�f�_�^�ɘW�̥��˙:+��Gi��R��u������~��-�!\�V�8'���19�����*�{o��Y`�V$��Q�d�7�gpnt4ϳyt2���:����\o��f�c;���R5Բ_"�f[�<V)�1MtܗEQ9�m<
,iNp��G�;��'��E��Ո<�(��ې.O��A�"�� WyR���9 ��%a�_P�S(� ���e���B�q�� fic�6� �h-h�_�i���9z��,aC��8F�����铐�mTC��iǑze�|�t��+������T��`�IC��E�׏/]ه_0��Kvo�����h���:�a��$�L�����o&�]���|J�C{£E�v�b�$@�Ѫba���'M��XQ��O���o�BX<7���t#4[=�"���F$�8��vd��PzCޕl�I�z�)SΈ�+��x�ܷ,�6�����Ү:�=�� �,�:�B�����|u��i�r��)Y��oi�	!1���S�f�5���­]��7�>���#O��F�q�݇9ũeg
 P��!�Ƣ���zO�1~��b�|RR��w���v��1K��,����c=`�S,���"�>@v�GC��o�d��P���+��>�/��.c�YK����YK�(�f�̬�d>�����ç�2�"4�����U��/��3��yK
ҕ�� K��&y܎��/�7�`�v�,"���k��v��Ӊ�$�iEN���4B�AleJ�|�~����T(�o��r���|�*��<��'�U�P����@��3�۳hN�	�@� 2d��5k��ba;����Z�I'�j��%>4�KeH R�Q���J
ģ��g��N��ǾP�Fad��R���MU�4q}��.�	|��E�*[���nW���/�"w�����򤚿��D�:0����p���CD�W9ƕ;��������Z!!ip`a_s�8���j�=s\�.��'N9�j�<�zI~�Vg���ߪ���ȡ�F���׀��i�=2��H�z���6�����i
���$�C0���0a�K��s�� �*V���`��D�3}��\�W��D��� �°W�Vn����g��� �φ��xN� 쯦��C��������v�W�p�h9��s��t?��e�30��/�zaORDĿT �v��4�\��|M�F��F������Y�?��,!`|�y��������46
����� `]��|���D?�6[� ̳Oǔ�z�4o'T'ivr�ixD����ki�d����7AsĐ7Ϥ ��L����`s�̫б��%*)Jz�3`�:Y��[��1W�!f�ŗ.H���� �Z��׭q�Ԟ���hAw�8w��Ĭ��m��C��\;b<R�j���
�ӷ�/��	@�Tg����m�o���ɖ��Z_B��8n!^I����8��(���f��EDx��}�)�����//M/&*o��b��n|��o���� e�3{$�M\���M��ñ��F�1���:�Fi�,����^1�,��	�y[X¡�P�����&��wBrP�+ jȳ7��Qϼv��8�)��j� �̉��]�P06�u���������'�z�ɐ^X[b�R��-U��=z��1�r�#4�A��I�=c�N	�h��r�M��_���t��XFU��aEi�ף�G6����Mfd):X�㔃����O�g��H�D��r�"�����`���$׎Z技e�^��ݎ�.�FrK�ʓe�|�_m��t ]���'��,�c\0������1���.��7��=���D�U�3����.oq�b�V,ǁ L�u	�uF�9�����p*�����i�}�P��R��K{����f�����\��Dam��a��j��Ws\,�����Ɗ'�VD�1 �s�t��F���H_��>Oj�3z��	�:�C,\�g�$T������d��Qb�h�kʚ�6�ʚ"�a[���q�D��sw,�58cl��P���f�x��\a��C=j���д��m��a
�|9g�p�� 2tX �t��$�%F��Ϸ^�S�`�]��e�ھOV�B�,��"|ë� ��1զ����.��x���T���v�>x��i߃�����W(�E���1"��*J�W[�I�����0�=�f��a8Ă/��q���O�)2P+�*"�)ĭ"w�2��.*yEU������=<����l�����ޏy��[���6<�\K�iT�E0T�9�?~Z�e��߬��XN&���G�i;����jf����}�n[�	�
��v������:��L��ߨ��6��TAT�G�>K�`�Ƭ�.�g��[\c$|h5}�=i�O�0�M���y�or�]A#��V�Y�"��I��[��ح�w{GY�Ic��ǱQ�B�r�õm�~�9�ޔj�����6�]����~$��� -�7J,�V��An��}��d���jI"d�G3��ꆦPat
��V8
��M�����;��̈4���)6F�Uje90=�sQ�K1F���/Z���Jx���E��sL޷,c)�g��&q�2x�����O3��lNL��W[��L�ɝ��r�	S�v���>v\��U��W�-1*�eQ����}���������/���J��Ex�5��%�����z���H��/���jy
���Zb����?�%e��W��7���p�x|a��jwSyb��T�L� T4Ũ'L�G)�x��˨\$g�:���Xͪ!OI�OB�M�s����9s�b����O�a�`�%Ⱊ�����_���^�ޱ���r�F��!l�9J��\
��\��O����D�y��-�_���̦�M��������_��Jd���IF[��_`['ǜ��njF����:�L9�ْ#J�6bo�w%�l	��Rr(�|���D�
���2rӂt�C�k[������t
��;����%/%oC>�x 	���'m�$(�d�ha<���_(�9"'�� �|�#:�H�����ih\&��}�?�a�o��L��q��llVDy�����ya��ZSp��!���r�V�92�����|Z�I:C�hWlR���b<��+X��t�p9�r��h�2���P�_��Lǃπr��>�9,�!�WΟ��I/�ꎔ(�����t���LJ�J;���jM��fIFy������ǁ�H@�]~S{ߟ��=���#���W'�a��������9-��!p��8�o�7���O��^H�������"w2�3��1y�`RW�v�����=8���ª�#N���ќLS����BJ���]$��#E��(��������֬���d ���<ݙ�A�L���.�J����H(��\N����(��4�?.�`}�f
?]M��zWPl}ֿC¤e��8���;��_B�ݪy����߻cyB��k-�4��>�P
5�:9�`�lh��� a�)���/�8H��Z�,�9�?�ERI�9%n�}��!���Ëp��!��o�z�j�.�h%�/�cej_�%O>Ԝŝu�����L�k̇��pl�}�+�QUi�����e�p�/�����]n�E�Ѿ�T<�M���Xuº���%����w�	�[;��+S7�3zVu�$���k�1� vb���� )�]l��Q��"���*s�*��I�	1Ϫ1��z>5�� %�'Kݾ��g��.�J�P����H^Ff"x�cxݞc������uC>� +�)iNa���h��b^t�����U&٫�~��	=NK���r!/%�t��+�-#�̖�#m��tz������<N�W��F���n�o�Ru��D�,�G�����6�f���T���;H�̨)^2��݅����ݩ�-J��^tB��X���>3�����P��'UN��y�	��.�ݪ�0���y_����]	rq�w���#���o��(�*����{�C�Y�ĝ�c�el?(y���/��r�h�Ztm�v�L��0�-��s!9a��֤�Bd[�2��:�%9�O&��oiT�FP�px�t�a�Pc���z�&��`�0[��\������̓�\�%G��ү��`�="��t�dO���}�HF��ǰ˹R�4{RAF����Q�S�$��'JPH����k2 ���i&;T���Z)w6��B�@����ɟ1f���/@����B(y��q!�|F(�j1W�ו�E��4��\1i?��&r�TIv��P��Q�̕k�����)o�a��x�u�u!v��3��~9u�������>L��@��X�8�i��Dחg4kUEȍP��D��q���.Ǆrxr��/>�����w�k�n���F�8-��	�)�Se��B�Q���j	�t]v����˭���(J��+��`	�>�!X�R7���+�O}ݵ�\�H��[{1s(i|��]��7P�M	αmn](_h�+}>
�2���c<��]>,vL�a��Ճ�#�-
9Y$��݁fUc�_]�p:^��3������s^��9��ma���������2t&�#D0�sP�;z�������!\�U\"�;݇�i��Xp:���+�Y�R�ֲG�%;�z���c�ע>(�j,�(���o&��N��� �ZY�0���]T6�Ń?�}�ݯ^�����JZ3��7�l�����7v�{��Um:�п���ks�����~r	{*�/v�|�լ'�xNg�q��Xr�|��<���/2䰆19���5��f�0����[1�%�n|ϗ!kع��`�`>� �8���g�5G�v��&�Z���_�ik�io�8�Δ����Å��
&ךb� �Z�/���ĦA�ѣ�[�����yۏ>�o�s`f3Z�m���=� ���fx�������K�0�1ej��T��W5��T��z�+[���[���lJ�4��K�_�7O�0`Ԫ�{Nwc��
B 01<b�u��y��:�M�Qy��9M���+I�`Y6y`�4���kM�1siR���n�W>8�lJ��θ�*-�I���5t~WE�<nD���\h�[�-`��4�/Ƨ3�����:F>���6��9^X��z�����C����Ym(��1�D�+[��V�~:mX %eOX>��M]�$�K�|�S�W�����8�ʀ���IzRb: Q�2 @���^j�������'�d��	1S�����y('*�������s���8���KAH��+� ��� 4��?�ە�d�%D�b�3� ����U`�,+wx|xO�)E�V�5ƶ@_^Yx��ً��%��B�-�)nOy�9�%^�y2(R�;�{=��X��4iLfMi��#J���&c���{���=]�~���Na
<��kF���9@��G[�_ǀ#�q�6X4&��-F+?F5CA��KNgy�mfk��y��OY��T}9"0��IG�}/�ͱ�,a����ow<��~�ɂ����cO�q^z�{H����N�my@9���݀��nn��,F��~�o��q*R/�ڼ譝�q,�v�m;�/s�@^?M������QI�5�r<�3��ի��	�*��]~��*{W ��:w�ʁ�1���jY���(��(La��d�mȬϙ]�kix�YNŶ�)��+�h\��h����$��y�e�+ *������G�x7�4��rJqk4b�B���L[��=�@Q�r�G�OHFb�`�A����-А�fݚQ$^/5�V��وx7S��e�n�PI��t�~�gL�P Fk����4���]��`�ƔM��f�q��|Ͷ�{*4��=č�#!碇��M�a��Tj�&��"Q7k�E�0�����c�j����oO?�g�>!	7
)rf�i�]�7K�,����)���&���N���lE���/�]�?�rv�U�0�p�NA�&��:~�u4�9�]XD1��3�j��Z餳@;��*(�CL�,Ul��������+�\/U	�4	� s5�z����o��B���� WZ���ǵjƥ5@d�2k�H!trSp���]��;o3��-,)��Χ���(jL��n���34�����8�w1}�KtHs�9nsn�o9���@3�ِ�f^�1������~T��󱁳�<�M���x/wv�+�I"�A��}i"��yP�9o��6sO�&�<��x�eJ���F�#ص\	g�VB6��p�����v��FWd@ô0)�)���Lr\aڀO�~D��xA|u��]X	O}��-sr���}����p������֫5a�;Vn2�U�\NT�T�������� #D���A�z�>�_�)�����&r}D8[�\Q;�R[	bCì�U���/E4�,ګ���N]~�#�l����P-��� �H��}6fJIr��1�Fo#;\��,0x
4ה����U|̀��kb��,��-���IdA=J��?�pn�3$ztv�U������7-���7���qѸd����l�`/��x�t?��Rn�!��\����bf ���6�t���r��}�p�7�V�O����Q�<n
0��/�#����"wK�j�W{RM,�$k���ƄO���Z2Gd̂��#���fvK̂�T���tHF}E.��ON;� �-�`T�-,s���R���� �&�л{��1!�,z���Bfa�Ii�8�$���Ȳ��DB*����9��I#�D.���Z~�7r�Gݴ����:��t�]����@���Zfx���ɹ�2(��:�w����aZ
w덯�_�V��j�R_�ar���ʤ!$W�z���9��8������!�)��B�g��ˮ��z�o�v@+%�-��()��߉�� ��h�-��|!8��E����+Mp��L���yٸO%�Ǽ��b4M�H�~���N.���v���i]]t�&�7=�6Wd�d�V-ro��M���m�.f�/3�9��H�����[� �_!�T�(�����vh'���a�7'�Y�6���ʗ}���a�;�o�"%~{�.���?�b�p|�o�h|/�:�Г��㛩~�P�D�
���,^��[�����ϔ[՚Àqw��U���8m(��A��:����v���6�N��VW�D"~���Z2[�"�H�o"���ml�2���E�����ܺ|���^uA�C��(N[9���m,�)$0���W�>�_gab/6Ϗ<&9;E�·R�W�vo�o#xy.И���@�Ł�#�yy~�c����:�<
�'�(T�8T�]��qM|�i��K�d!~�qƬsre-ϙ��C�Nqi��Jdr��
��g�,�?Ô-�!�AX5^C��ݜ� ߟ}0݇'Z)��}fU�@e�ɡ<��@N��;�G�c�[IP��n��1�9$�UI)o^��z��A�Z�	c��Ouъ"u�(�>9.��#!�X틵OV�֨?�5iS?�:v�`Ԇ#�d��+��.:!��vc�%-p����A`�ʂ�B7MA��XN�d̪��]����DjT���7����Ah���N�k� ���A�~#XO�t���Ji��%*3��r$�r�9���v98*Z��l�?zݍ�>��9�� =]�H���&T�c}��1�$:!J�h+Nn��	+%���>�:�}v��-�Ƿ+�{9oV��!}�K�=���|�R�h�Q
@q~^|N2>�S*\�Ϯ�FOH�o�Z4�g>�9o�qr���My�Y��4K�޼���J[��x���
_�#�/�HQ�B�0��|m} ��!1%n��7����AFн����9r��rz�l[�;|b�&5h�����o�o��^�dKfs2r6%1��V!�A�����R�?��4��U}17Յ�������P
��/PNYt�-�E��lG�U�s��ڸ�;\��me#X�^�����I�n��d��WF�0A�	v�!j^�6.!�A�渤CO��d1�&�>�Lr�"�%�� N�d�FE�� ���:�����k>��N���H�x���("�P[Z��x6�j��g7�ˌyrc	�:��&aE��	��ӂ3�x�bY{�Zoh�8�%)��aӄz������]���0�pɪ*i�˜��K���c$oi1�ۑ_�7Td��hƸh� �6�9$i˂B�ׂQ�N�_�2�@���@�M��v[w��~��L�"�#�ԅKĆ>r��I*������ i(v�]��(#@�͂H
�B`��%>9u��������Y���F<庪*�u��\�{�̈́�Q�Q��Ȳ!Q�<��d,�~Lȕ}�kQ��w$�t�a�w]�:���+Xwy8SGǚ&#�V�B�V���fj�l�+~=q0ކn\f�)Z��w��LYgu���&�W�NA$�-`Ҫ��7o��*���D-�`��	��A(R)*˿X�~�zC�6¹�&*��ݣ?&����줰�K��v"Ɖۖ�g�z�a�!0;}@��]���^��|l-3�7�q��a}�@�]a
j���6q�DJ���v�}[�ij��Ąe�	L���ڿe(V���B�Xj�}������E�j8�Y;��2#���[g2��D�4�fk~g����Pn��"���v�P�2�������e���#̜I� ���	7���	&`��Zc7�
�=��,c=zJի�mY��z=��Z��E���p���ĂI�p��Qp�o���L���2�k$e��P�#��w���r$�=�.�D[$<����MfZ7Q ^� ����W��'��\p�ۋ����ӷ	Ӥ�D/�I_FzyA�?A�A���d�c&�S���6�<�~�N�K����}�^��C~ѻu�/ז`qnL������K��-�Y�TF���ڡ��r��h���Gю	�����6lN.��(N#>^DGy,�#������`h fiú�X��I�����v��-}g�<��]6�c�U��8�&{�,���������w�i�<)H�������0�{T��q�I<�������D5����%棪=�LX��%�l��nm����������|�s����gA�_
�G���[0cl��`'&��<�6'���S����c��e�*G��]�:�&���HS�u���p�7P���������t�nY#GL��j�e�
���c_��3���.1ق�J=�}:��|���o��p���T��;>���-8:���rq�+<X(\?e�
�;8�;C��9�5O�����[���a�}R�B�8ڝ~��N���ڞ���PKS��X�o����bR��X��t�U,��sɑ��%�IM�Ҿ��"og�w́���~��o�ҿ�SK#]7`���1����9�L.칦�
����(��E;���H`�bH��������l?qf�ԧ�@��+��*��o�G��&�������9��/U�	-
����Yr����Ok�GYa��MBj��W�v�q�$fU���pz���W?��ZΔ�Q�F���vef���ām���h��qc��B�PQS���X��& �w:��Qb`8���ʚ˳��%� �$~<��cNL�!�t�h�N��ӭ7�l��dTӴ=�y�����b�4�D~�<�4�P<X���V	S'+�9� ��o𻓰;O�p��/u�7������ p�u����N����6G��/�ܾ��q��ۿ�*�D�PE_E��M��2Cp�T,�P!q�1�=�]i�gQlNL�N��R�c�)�����ir��<�赩2�#b�t�<=�˵0O���Ξ���4�M�1�k�����??��`\B��[�m4���k欺'�`��_ٺ����:΢��Q�ɔ�;�El��ь(����}�5��oݨ���bG�	U+��z��Da���G�����w�F�͗��o��Q%G�m!H�>JyW�XӃh�'�E��7����ȇ�=����.���	r����D�r�1���R~<�nH��XC.2�����JY�C�BwÀm2J�a ��N�������&���s�G�2��"�	�9t�p�-����������0��#v�1z ���w, �7{H�����a�'���=����Ǎ_zI�)p�jP�3g|�>*d�d�1�op����J�9�[�3J��˲zA =�������� ��":��(Cr0�?�خ���u:���5��H�����\nS����,�wI��eHa^܂�

��H��Fz�������mfܙS��W�F��M��M��k��5����*��843� �����Q�m�a��������>���a�w*��exm�\���i�r/ױ�l�RVI]jq�d��xg���9��ĸ���'ŕ�_�Dۦ��U3�;�
�?����j��P���ӵ�^2���'�ښa�Y�G��Vz�kO����%�N��Z(��y���:.����,gZp�}~KSt�G�7n�V�}��T�H��Cn����r����-vC
C5~!Q	A��O��x3g]\)�D@�����P��v�~=�	����_�P0�ȋrb��E*���c,!��WR<sf���)�\0m���M��A�^��G�C��v~��#�w.ZO�@�EKl��(��J��sҘ_@M���b9J,��?&Ќ��X�ui;~wv�4�!���q89��tB�t�G��2>t�&K7����C�f�ix��vB�,�
�kȄ��4�Q*�����	@u.~����Q�4�h���C������׻B��x������Q���j�5�up�����aƗ�K����$�"����*�C�J�?ٵ�}!��`)�z Y� �N6����2��[��m�%�ّ���?r20r�.��a���2�����E�(ۜ�SA�Qh4Dx���R!V�ٯ�Zzc���l6ǧ��7B�U��8���`5�>5��`�9��^��o�^��A#�p&��b.Ա^5Q�(�
���bGk64%�S���$ٹV��o����[O��]�m������ԕ\am΄�J��_��W�#�l!�X�>z�8����`�3d��\FM����	�mh��M������)9�}�=�;��I9�|k�4�T�5'#4Z`�\��&�M�l#��P��0.�W'p T!_��#�^ܷ(���_i/,x"`6�x�
��'O�Vz��p0��	ԇ/���4��Y��ۂtv~�D˚&� �s~��� �' ׈���B�yՔ�7�wt�W�A��0`>�o�doxSH�wk�,x�s�i25�`|H�����mk��c��u�8�������fM%�Ẅ$�l�/Z�#b1�g9�~���iU}>���X��ۦ)��y�',��:�?Њ2���Q��x��V^>q�Y&yj~0CE?p$��f3���woAL�gT��<@K��j��7�����m��JȰ����F��L=?�߷B��bh�X���Sä#�bxɘ:��V��bܖhe\�g�#����LHH�K�4x���X�	!,�&S�^���E��Ѯ�{��e�j��=Tr��*��f����%N�#������\���bod�m]���El�����ͩ�!�����z���BF��jo��^ž��3���Z��Ǳ��o�.h�W����X�d[��h+�7��Ft�&ݗ:���e�U��&'FH���?�s�c��{��
���(�%#J����k�A%�����{=���j]�Ȫh��I<�y �R�����C���^�Y��>��"z�0p�3��n��-��\�mʫ�ߧ*�����vC���P����FU'Z�8 .�E q��@�?����˚߱��b��a
XS�{'ɹ*O"�}y�}BiwW���U�(4�$�%� �g��a�]/g/��.\,T���3ڨ��Ѓ����q��J�j�j�m@��u�a�����f�ܧ�G1�T����G�,������CI�����&�n������q��9%p�8��z�M��'����ą���Xܟ�]Y���X3�H�o�,��q���䌟J�\�Y?��Κ*@Nk�J���
�>L��ݑg��-�~ �{��m�^�i<����܊4���ϔ��(�3<�K@߇
��H��~d���Jj�S�MY
wQx��\67�PD�r�j[�M=Y�ɚ��s@#s[%Ul�cF'9��"	��5���
a��K�Tw��Œ�a.$9,������%���h�.��R�����0�p���ςf/#Ҵ��'�j����W�7Wi��~o0�I�_��0��J�y��A���Z���*e����b��^ʫw\۳.sQ%6��IN�T\���۪��H���pKBŵ��E��6Ce�<���?W���7�"���`�"�������V�=9#�934I
�
��8�K���{2pcB�Β��Sp0����F�X����>�=�����|�v�z"�8�m>4@�v9Vq�܇�D���{L#(��9����tGuc���A$+��T@�l8���Ku�t=��F�%Ug��m��,m@[�nQǬ�F�sb�Pp~vn.��Ld��]��I �]M�Ȥ��Q�A9��& ��M���z���@��1J(�F����\�;t����G�	��7���Ix.���NP@Pj�ԭ�2	`]�]�������&�st!��	�}�JY���*�SԲ���ۮ��w�`W�_P�c4	�`������xD�>�����\�y<p� &� ��� z/�'^F�����>���s
"�.�l�C ��$&�B'2w��my/��H҈��鹘=�8p�Թ_����og��8����k����j��O
�}tGr$E�����O�$Ģ��&A���K�j��,4�ԓ�:UFK�F{9]8fpc��2�t��r�~�	�$]�U�#�����*�#n�VcmMN˽[�T\�$u���"�֗�O�Wb�tjh��IZ� Iى!�ai*�ۮ�%U{��F�	"�]��z�b(:������"����c�<��(��6�w��b��)�lj0ri6lX�����1����'��ޙ*פ̧|w�Yƹ���?�I��D��lN�+��pF�|�=Hi��YQ�T��]�	�[`VG-��D
�IVQwh�^q���N���Ǵ	�`؋���}��o��j�9�3��YjL#�_F�����b9�r�A���x�._��C�T�U����,>q�$�g �'-�����$�ķ9S���ku�gc���*��3IT�h\C��'Epă�g�A�b]�pD6�}�/!�j�G�:�]��?�Y�.�cmo�!���5�ؑm�p�b��/@�Vnl�}��qЧaa�6O!�g��d��|>�h��=5��ԓ�vF7{�]���}9g�����Ru_��&u�lH�Y��
(��9�3�K[k��?ƅ��k��uh��-�8E�-4T>Q�mDqE�x|{�֎�u���V�� ��~*=������&��V���4��Ǝ2R
O�Nb78�y���[f�;}��L�U�r��j�
�����սU/��8�u� ���ʮ�>�*ƣk�=Q�"�dֺ��)z="�Q^.c�f?)���H��-E�lI�e�J��8�l{Kk��$�~,�r��iw��}U���)�Y]z��:*sڞd���[]�Z�"Sð��Y�.zpOl�y̸.드���!x:�RT�݃��b�g�3/���Q�@$\X5�����ႋ����A��z�+��)�I�W���	қZ��g�8���կf����f�鄕}с������Z�屮�zd��ó_J��z�$ݩy>zeak���^.<�Ӯ햖ؠw�����d8&�,��A@��e�Ȅ�'I�Q
<�nm�R��g����Ij���U5=��1[.���^,�^QԯuPџ��m+�1����(�H�btN� ��9*�.s�q�`~����q��5���s+K^�:��~��S�%ǘ����Ⱥh�e�."�� =�@��UNC��P�WC�����2�+ƹn��ap�����}���d��^������XλI�M�@�z]Ly9��$p����;��CYì�Vז��@�ךeD����i�,����a\�Yv[)g����Er�}��H:ح���Ϸ<'��M'Z�="�O�OM��\�ֶ���Ӑ�<F}���F��9$�y!����tl�V�	�^��}�]�h	~��چ��eZ�q&���@�d��&ġZV�o&���Ô����[+�G��W�qjvz���Ph҃�*+K��J0ܛ�;(a���.u�Nqi09�Er�׻�.��#3���H�~[Q婎��#�a^�����wM��{O�:�+�'q¤��bE��P�R�C��K:��;�r���z�i39i�8*�ۤ�دL�ϵ�ʜ���;�]�<�Ϥ�[vfwQN����"�����,_fT'��+`^Q�k}@+���1��:��.���t��Q��ZȠm,��LOi�Z�A�08i?��T`(�˄�ЋB~�;�1�.�����'yX���i��?��z?�z�u>�,^�DS�jH��b?�c��}�$/NE[gt�S(G{��<�w�X+2��$&Z}�{��J�K�5e7�т��o�ƚ������5T�uـ@V�E%��Y�ve���3ɿ-��܍�^�>�f�/+��E���X�\0>4�F/�~dIQ�j7h��x�Rh�_G}�|�L7(���ߔ�V���~ҁ�p=⣶L	�%�͑W�[4�N�8��Q ��=����	n~1fs&�/2�%�����EN]<��0��g�$� �U~��:~t$.��=F(L��l
�w;[�����B��-��I��Gqu���,�J��+~S�� g��SJ)�P��sVm��������ۗF/wʜG.�.��sZ���\�;���*ά/QE �i�������y���w��>�����/���Y�!�#n t\(��u��t������kI\�!�W����$c��/l��Mfm��.�F���
be�lj8�M~,_�!�f ���O�B�@j�O� ¨��T=���
���� �*b����~�Շ�� ����7�n��E��6��0!f&y��~G�/�������Xc;�/{�J�^N�ݪ;*�f��4`^����>l�SωM���4H��L��JrňV��:y)3�z�����VH&E���+VI[P��<�f'B���kd��eL��>������_�0.�핢)�s>X��m#+�f��\+Mw7�ާ�V;?襩�����1?�Wƭ�k�S��f�7��k?���I�a>����6�X[gH�Es*��!{�tA��c�b���,9>]%$$�Z�ou�'�֟m8��'�3k����Q�ݴ
�e�;.c��Ork"���Y���	�$ei������=�4Ll��qd<�X�n�=�#^+���iqWDf����dʻ�
��8��b3��Qx�K�ek�O��C��EO%t�q�E���^�W�ܿT%�ml�.>1��P��X���G|;}�Jئx�O\b%���Y��g�������$�ݏ� �N��&���h�2p����/���d�f��.��C\�Q�|Ŭ^���%/�t����� |,�&y�@�{ ��jH�1#D��D^'f��l���X��R�Q"�?��Я�a� L�څ�1T
�OE� �+�$�HS/�?b���Kѭ��Y7�,�!�n�ťfG������Nr�9�O��d�, �v��
�����u���+-��1?ȅv���-�.�3����|z��A�O���}��ВT�A��"lk�]�2R��R�	�Gm�Z��%�v,�����PQ~�yO�a���8~O )J�&�P����Pϰ�E'�O�P/oX���"g$�ٙ�����nۦ~���O l#m�����,8�L������r�u؝�`d���-z�6�lH���n2�8)�	!�a�㦰/#/uB�W3�l���������� ��O�C�  �?�$h���|d�l�Ӽ���ǐ�����W��T�W-��!��s�I�@�:�Z��h��#P�툺Ց4#�VȰ����Eiz���5(��6�WqFBC�U��B02����L�>�;������e������N���fY'DqHQ�G��A�l��!�U��
Չ��,�i�̹D}��Υ���o����О1̙�dO@l��M�D�,������$���J���ӛф�\�[+½K�%��O<x��Q�x��b�xzY+D�� +����l�WS�`�Ӵ����e�����|��x������m��;
vG���Ă��\h~+�-H�[��I�%\sP����X睯:�B�3��D`A˺�78!�s�Q���<&F��7$RF�8S�Ԡ���i�q8�ʬ���h��@X�=��$8}�z�#V�lbFb���e�a�=�~�΋�β��G�j:��53�h��6,D�?K�+�^y�/�9�y��PC�����]��s�� �k�eV���1Έ�eԾ�ژ�#� ��
*����&Vp�G[��T�4J�j��x�ҕ�zR>�z�1�]�y��{F�E�&k6*6nn�����#R�L��pG�d �c��mO�zbz�^� �窞�9-�5��2���y�k�\"�����&ջ��~&�2/���]��ms��1�����7nឹX	��q\��薮�����X9�K��%�&#�T���q�c�'�����h�A]��C+�q�g�%������ ~���d�������)E�\��Fh�Y<M�����5���IQ{o�VǕ7@����K�8?�@%ܜ�7�\���G^��<��Ɏ�p9ot��K��6L�����	��Y�qgZw���Ì�v��qo)��Q��b�  �ݢ�m�틬z�.�v��b� �|�9��/�䙠�}��f�[�j�u��h�,'�*�#<�4�ר[�'0+�O��y�)��Ҟ�&\����i��o�j�OJ�i�9�GQ��Տ?�Ӹ�U��p��FP1�����s���1w,E��`K�����#b�4	�ɀ����;LNի�1��BpY����NpO�T�#��}j��57�&�R�}�����7�x�P�C�4�E+>�kCC�gW��������n>�q[m�:K�\R�K�����"/:�)ݦI���Ӈ�	�b��N�R	��PB�S�0�����&���=��F���}�����J�~���nD�I,����;,����S��s���@������ܖ�����I�G��C��z���d��G�՝��^�}�����p�<k)�#吥:�����~Pگ�44�^�g!�q!�t8�O[�s`Ϳ�� ��sj�KaW|�A7]\U����h��A(�&b��m�`��K���d}�'�S�_�-�
��U�9�ɃE���{'r8�E�^?Ep/�܅FN��π%����S�G;D�ɶ;��.>��V;��tq�i�.���F�	��z��h�-��m����c�,��~���ێ��c�m2&R��'��<S,�dH
��tV�BK�ʰ�	K�W��� 2��8�n��|zy���S��T��n�������ep F�?Q�?N�;�<]d0�� �Kp4*޽�#A��2t�� �hIj%��=}*�0x�\���u��~P����(8��-H�uq$[6�X�:�)��{Q����}������up�a���b7�(·@��@UR���m���UU�~��}ç���f���%m�1#��w�&H~����ƣ��F��P�*�/�xdV#ck��J�tE��&i*���+�"w�F��=��D�@�Řls���`�A����n���e����"�I5h�*c�=�e�3.����S�0޶ZL%<���C�Px[��J��`�����2���Z1�Ҹ�ia�C�+�[Kr���vz��T�|�2N��
��3ī����n��/[��N��쳒^�1�[R{%Y��=���#�_! �p�f��0eT.|�J� �9�I�"������Q��.�2��L��G����j��Ư�vڀKb��v���(<�L��?ِR�  '�*�aW��E��D2|�ž|M�duL�YZ�$�"L��LT�}}�oP��Q3�*d������~�)?Y�"����u�ϻ���}���:Ce�Ê��]�%�kF~kVb�mFH��2`6)޴�	?k��|p������:���H��$g2���<^���Lb�
�w� 5{qY{m]�3UC��N��V#nfn`\;��71�����W)�����$�&���q����Ɯ����u��MQ�az�T/%w��&2(m�T]:��#�o��H�n�����}�ś庿�z���I���S�<��`�Mm�Oc�a֕o4�>[�/g���[JH��L��K�`y�������n%���F�?�Ut�K��Vj��O�&����6�D4�.��!����4�M*�h6��K덪�Y�ˤ��cMfub`�.?�6��#M�(p0�W�k����)\�df�1W�u5�"C֕���d��2Qg����n�����UY��
��65����3������a-�V'�*����\�)F�e-�����g�����16�n�[>�zO�uȿJ�5������\�:��RU��N������g��o��&�.Wz�M�؍�-�G9�(�'"�7@�s�WR�~U�������ݯoհ�6r���D��w���$���?�Z�hYp�G(�/����$S��'�!�P���vscF�`o�دҳZ�k-��7�x�/�GK�"N�-���ƕ\�f�ߒNT�JN�j�ټr��`QM��nT�<üui��(s�b��#�8,�Ĕ��{�>Q�Ą�c�y�i��F�$�M�MࡵΓ��Ǖ��k��H��z�5�_2�s�<�"�8�!���*㞯@�c����͍�"���ˠ�bF�b�]��	wV0��Zz6/�T#Ծ��m&��|�r}_����~Mb	c6D;Ɩ�Bs֊��=t�ַf^���j��(��B�Bk���8�����R��D1�E`�c�m/Y5$|_$��� 8˫�O�@��?��t�)��UrA�p�2�(]=�P�lK!�A����D�Z,�V�!J�w�
O�y�紣�x���{��bb�?�v��C�w�Md�̪�����x���M|��4�ܶC ��W�: ��H��Q�b�q��AFukH����2 ���(��Z�pY2��[l�r��Q�@�|=���� p:�P�p�f�A!�K��x��ucAY�|�T�M!��1�����44��R��[uo�_sM.�/���l�Ӻ��SH$��K��]��]h��.�����n��NrOX�,��eܮo���X+�4��/���ծ��:P�gryL.=�R���`�^d�zd�׫hd������#wn��(��]G���J]����5�g�Pt:�H�V2��H�{XSܭS��, ��vťo���9��rT@���b	��L�_}m��8r(��b���\�}%�mC~�մoɧG#0:�
�sN���g�Mm3:fA�Fz�ǀ��D��`K Θ��<O��V�m�Po�&�,�H��l���^�^�g(>�σ��:c����r-�8B(�e��uȍ+�6nKQ����%3	(�o,�0��t���OZ��>�U�ڭ�_���E����7�?�Mp��h�p���RO]�߃��8��	o��2K�z���z�
�{F���¿�,0x�C���Q�ګ�b ��T��Qч^��8��Gт���
.���z���Ѧ��O��Z$���N����y����9ET"��s��D��!p�+9o��"ᭋr1ĭ9����h��ĸ�x�I��rZ����$ԩ��[>��0#E �.�xx���5
	*��1t���Ӣ!�ʴ x��k����`�у�}O:5���[�,��U�y<s$Bb�fb��fk+�&���a*j�բ�G���1ߦ
��V0/�(��vP�~Wҭ���s�)�'���l��V��b�\���psEz�!��囿�H��h�Q*�;l�a�@}؉nK˼��'ϰ�cv��X�!��|r�l��Gc°�|�oP�0�pp�P�zkr�YlUL��Tݵ�6�u���fەf�]�����U�f�r1���&�ŬU�&h!n�/24��XJ@|i]�p�	�7s��!`R�w� ����v���R���������DU�>�p��)��d�S����N��#ڃ���}Rq��++�˸G�j�����5Nص��^*d#�,Ŀk�LH��|���縀�7�JX�~;��^���7��7�QP7��c��'�T�t�fԾ<�Ƥ��4 j9z�sV�&�<�]��(�1f�#�`;�=�`w���|E�ʄ+�c: O�tJ6��6�~:M��qho2�M%S�XR�6�l�ؿ�@�26?��������`8��b)�6�^
����"Z�l��=�M@�r�d�:F<�Zp��><����J��Ē#C�o&����b`xT%�bn����k{I/qElO�����
��,G>����h�6�3W\i�0 �
��'M^�x�A��3Ķɲ�r�\�� ��Q���Э��hdV����a�At'Rͮ����$N����.�<��n����(�ڨ�7),�ؒ)K��{%�Ѡ�����R#�	����[���nt�$Asd>˪�ΰ�M����T�� �(��@bS�Y���� .Oϣ�xuV�'cs'�;8 ��v�}R��\�p�|�^J�u����b�7�f�VJ���f0AA��}Fi��΄���hp�x�R��,� 	U}2�h*	�k5��n� #�� ��g_wޣ7]���WcE�M�d=��֞�m�(�gcǛ�O��H�d�a�m�4��D?P,�$�d�{ ��L� %A$L�p��ϩ�Ճ��(��E������c7��e�zP� ����P��C���^��vh�X�B���r
=eT}�#,)L��M��e�DI��?���+���9Xہ}ܸe�@��;e9��g0�D{(���bt��+����B�ܖ߅�qC�H��I��H4�*�������9v5��o|qL�e�S�#�M/ї�4���#
 ��A���x��vO����Zc��A�����D��E��P������c[2aY��b6<Ѱ
�$~���QtGȇ
v�G+F�ެS~�_Ӣ��8���)p��X,��c�g	��Ε`�FXw���V#�,�56��N�h�Q�*:&���P�&��͉g^�BS�&�v�h�	�R~E�-g�K��
e��:;�ŕ�f�Ԓs�1��m@�S�7l�E��3a�t�o��99e�<_�E�8-x9mK���D��^f���Q�w���� O#1y2c5[ ꭵ��&E����|g�X���E�'B�������ſ�i�Ԉ�;�Pd��}p���g�P=7�ZA���ԡe�����%<��D�F�g�y_���,S����%�|������������}��p��+�I+�U���
Ფ���s�ԁ<`�\�W�]h�c�4��ME��>�@��IA��
�����W@}�Fn��� �n�.25������]�/3�d��;{��	Tlƚ`�L��tt�p0�N0Y����|��J��g����Ԗ8%;�W7Y�O�k�ȍ]�8���|���
����PU�;���E�X��P
��x:�o��a��?xP���xN��%N��_j1e8��=>_��q	���J�f̶uc�k�B/M՞��Pa�UIE���=�����$5��n~G�B33U�)�!���QJ���ݣbۊk�Ѭ`v?��"]�yfܨO�D
lk@��L]�d�*�qL�w��E��ÞեR
�Bf��]�U�L��T�r������!�zޑ���M5b���m)Ǝ�����hX��Cb��?���������IL��*��b^gO������ƿAH#������G���i��Ҧ/�e���	��� +�M�B0ZZ��9�2N���'�TY�A�̠Z��U�"_�B�='�P��Y��������9�����Id��?GZ%E�4/�P�!�����X�L#��ҨَqQ\�o=K�["���o�s� _B���� �B��0�(�GiE=4��GNR��iN���n����;o�&�bQ 2�Kyp}�#��m�f���0�ZO,!򴋌=/	����=Ј��6j�l�B-��r�hv�:=!6̳`?�L��Y�]pk�X�p|y���8%}�C��%]�>-�����%�{�Ӭ�����O�X���|!:H���La8�٤�Y�k��s�!M�z�I��`�c���j��4���h������J6��-��&D�O�Þ���9��L44�tp(�óWv��!�Xq�ld���6�a\�r�)O"��\���c]���Dn.��'�D�aZ�YB���D�L1]F�I����v�x���8���V��m��s?�r��ƶ�����ޣ��62�4����7J\���)A��Oy���Zj-�����y���-M�`o&��g�Ǹ\���7PM:!�E"0�#�C�+��Ӭ�@��z���a��c�ùM1[��I��&���ɔ��|�@Q��=< N�q{MO�EN�M���<�SQ�����U��iK9^;���yO���~�|ˏ��a q��Q���f�w�͡���4���t���0#�?�Ӈ 5����D����Th`9n���&"~md\��K�h,§��v"ID1h_ܰ�.�u����P�Ώ"��<�ۑ�Crk ]*1]b�+������R3$��j]�֦�FkÐ��R�	�tW"ly�&e���oe �VY�p��Lq�f<�����{��{E��/�$btDi�`���hQ4��|'�A
ۮYw�8׏
\}t�j�$�X)��Sw�rc���E���z��.�@��!)�pv�����{<�V�DH+jy�:�(�2�$,0&I�<���h܊���,�� AU�@�e�4��K�/+5~���_�@���@�i��ai�?��9;1�X_�+ֽ#�]$��mw�ݥ&wTUq��DH���΀��e�⾭!�b�������5VmM��
��Lv>�h��ӄ�3��n�b3�%���%�r�j!�L���P 9Nlɔ�gc}��,	}�\ ו�p�p���E>�?̕6��)8k����g��1�~,�<��X�B���
4�����V�^W�(�B�E�0X��]���X$��"�!7���4.�����(QM�E��x���$�J�7!r$L���Ḵ`%�M�5�V�eă<4K@�$ ��x���R������+��>/�f��^���{��`�n�_B���bV��i�-�����o�m�):�F�f݇��D����]M�)��Ĕ�O�e1$��ö�c�j�u�V/���(j+��eIܻ���c��O��-���Vf)�C��Id�-�?$o���Doo!�H"��\O�H�	�B�jM�/�sB��S�$�Y;���� �w�����%��&|��/��v��w]0a �����R�DU���0.8��_0�E:���!�.w��k�&d�o0�gɏlFE�)@���u.����o�6w�� 9͠��k_��a(`9��t�w�ȳ�o[>�b*(�	�2,����m�x=0�S�s�h>c$�>}݇7'��Wj�T�Q�'5��z'��(�<a[��_���[N�3	���|��S �Ȳ���M(6�ft���3��O�Pg�{�檈4��o��x�╜�l�,���@�;��-��7!&��3qO���*l��5l�T��#���KoFι�� E�=�a�i(]�����Z�]�-�H_�s�sM��U��f4}�'r5���"��=]F#Ro D�j&�'��{<\�*
��G� ��3�5q��ֺ��)<ʔ̲�� -��W(u�^P�`�>B5v��nOs��eY��)߼�؍>R�b �8`�������i���bm���|lĥ�k�>Ԇ.pD}�*�x�}O����q���Y����e�B�s%�#��G]�A3uџ�U���1��9�8�}^L�q��]�Y��7����äј�ꔯ�%	���!�	֏\a���c;��Bc�:�1
�6�"j�����4���/����N����L	��U`*��Q�z�w��|��,LV-^sР 䜧�]k�
G����{���]2�)!{�e�~A�B֪?g@����L�}
��*�v����3�q�K�j����C5��,����3Et�j6�pc����r���8S��[�v��
@�Z;埠�qց>����� ������IcW�-�i��`F�]E�h�54��kk��'ha��R�@@Ƅ����р�ԏt��pv׆��A�m�'�uF���Sy+��*'?u�Vc��ª���5D6��Xi�f����1�\���M���]�1\�o��%�2
a�%,ۋõ��sr�%����4zm�d�*�;�o�U�(���W��g��߽�y���2c�X`!�䉠�A(\A"��%��������pp�X��0�e�B���netom��G 1N�q$LG�*�x.C�1ݭ�a�yT����M�����	�'P��cie���l�.��2����r줥��o�fGhSw
�H�kH޲������q�VFm|�O����%�`����m��Q=��~���-mFb����X������L/�"5_1,�(�����Ah)� � ik��Gj��b8�GƁm?w~G��*��@�0hT����Pl^z��g�k�N����Ւ �EAoI�(�����$^��rQS�����)zz���q�Iͨu3�L��b�H�����M�Ç�o��8Ra�A�j���w��w�o�ت�&Y�A�2��R+����
�I�x����s:Uv��aE�E+<$���$���v�����aj��$�q2X�q(��W���i�_cO��O���b@����"��;���=�-!.X��J�V���&Z�B��ob83����Ud,�i��DY&�CM�`�:�"Z�*��I9H�����v� ys�5��b[�[lv@�#ǥf@�����[ �1f���`*�����7Y�-���B7\���o��`H��0S�)�8
���D#h1�-$U+�b/�M��H��a��Ԍ2MN9�Q-	5�J�])8�� �0������3�I��X"����Q��C�AKQn"󕽲���7��� \?*x� ܸ�OwO�vǵ� ,\5y���K2u�?�.`�ET��@������U�k�~�!8�dAy��#�q�^�M�`�Y��]���P�0���+}SLҼ��(^ȝ�~X�^3�_���z�f'�Λ�3�C�/��lB�(���52���7ro<�m���z`D+_;A�@F��+m7g�\_��A���Y1����qA�F_�#����;WnY��׼MT��6̖�%n��&�� 
��r��0�=R���]�X�GMe�_��_(eQY9$_����f�s��tU��w�������6�m��hp�_��^��`7��'�	6B�I�i�{�h�m�����ě.VhQ��=�G7��{@��C�|-�YRԌM^̤K!���H�Ro=�_�7�4�\�i����e�02�"Z�nWq�i��6�P\���h5U��_��#���X�<����� +ܱ�M7K��p����\��#<���GўͿ�.&�W��_Ա�u�^Y�h?A�V��VwZ� \wΆ�Nn����H���2�<� :j^� ��R ��9L��Z�B�Hj�K�v9_����}Ǝ����)Jn�{~ �.O�b��Σ�g���ҿ���|p��?��z9/��흨�8{����$;�Ff���muL-"#���L�ڸ6�z��W0�k�1��e��B��o$��S|J��[�޹0Y��ȅt@��4��&�<�6�b5p��ܟ������{��Yb�N{�n�2�"o'oK��H)_-Jog�="�]"3ȁj�H�� f �q>�T���y׈��w2Q�0ݮ[Y���s��E��t�n��o�*�n@NƗ�,g��L�Ⱦb�;�)�'�9�"o��.˚b��щ�֔8��[��ɢ}�`lLJ^۷?A�l:����=�o����!��� La<	��G��l[[_S[��]�+.��,/�e�����
y�t����Gq�)HkR�i����aG�ܷ2wt�+�gE�76��UcX�)����d/%x���r"Hv�y���V==U���:�bʛb�΋�r��H%����,�hΨdd�Z,����Ip�P�98�eH�>�j0m�?�87˴�9��{ۀu��\�ѫ'cG�����q����q[��~�+@J��>+'l����T@V�/Nw/Pd��8&�E��,Bș*�2�	�$�d���&*�.*���ũ���ں�z�!3"�N��e_�pۮ���aA���w��r�8�-O7�#V���,"���~�m5�d�0�q7� ̈́؜��;b��t���)�h�=x���Fﱵ^��?X��H.�q%���԰�P�&Z��K��O�^�-��,/knj;P����^���=�	k��*���Y!+�j�2\Cf�B���<c�N��'K���s�^<U!��P�����́JnǛ;�2�=�AuR��y*fn�@sB��*<eo�X��q�[�d�HkV�q�����Dp�z��QZ��uPMT�\������^�C^�C]!H�gMT2ͭ+�L�S�^:9�S%3U~F�$u ���|(�a.
�����5X�
M�]a�-?��O�n���[[�U;����M�8�-eW5$��(Ŀ�:'05=g|��Z��5���F�i ��c5aO����xzӲ����M��O��J��� ����L'n¥B��H��f�h�--�K_\�b���
c�嘯bʟGӣ?~��F���������Y�R'NB�h��b�����@�=�E΋�H(��g�N����'1�Ϯ� �e̪W�Ĳw�:��w3+�(o�
@�3^t8Vg��s��
_�,����#1�]��{��$��yiEZy���-;�]����E�aՋ�gj�֥��Q�� ���Z�~R�^lgX9�����l�v����y,�`#Q�,i�4.�p	�����Mٛ�3~�/�*��x2�S��Slq#�H���j��{=����r����h�qP� ���2r����is��%�h���k��)�t���'�v��}�*�$���_Y0���KP�j��ZT��M_���3���P+ Y�b)�p�!ؽ���k��(E;'w~�� ��a�n�|D��H�&;�}?�~�@�xr-�j���)���/���."|� �l�0�ݖ��������f �e�wI	�1�$A���O�2P|���IB��g� Ƥ.t���NN�JA���Ƕ"�$D��v��n.%�v�-9D4��@?���F�瘿�$C}z,Iy6�K�c�(|b}�Pv ��zn�<�b��I��9x�nòGv�S���(�!��6`�U���O�sf��I�J�_�JH��ݧׅD����"ƎCQj�w�YW(+(�^ �1����2��d#���klykV�Ŏᅼ(I��)be;;��y�����9�3�̼2]����[�I0h��0ҷ�h�[��7�D�gm�kq��֩���ڦi�_'������ɄV�Q� �� ��y���<ܧ��������n+~^��Y�I��`�W|����`�9����Z>7{୻_�8�����Dr?-+���2� K���_�>֒��+�(��C�P����Ũp�o[�8�V�n�
���t�`c�u/"�����HN�E�	�d��:��`� ����bС�a��|��	���1����nB�:L���o��鷉�o@���G9�Ll+�?ٰ���L������,�`H�߯+���č�&�V�G�1���1H<食�f���3��+S�f
�����r	Wz1��>�'"I�rw�}j�26it�'���椄�d��%��'t�n�qٷ�~*���a��~~���Q�~l�M��#vsn���2��3�`]&��:��*x jQ��ݓ:&���UK5�\�{9�
^pwxE�p-Xi���Ϫ,мӾ6����M�?sџ��c����*M��q�^� hCq�ʪUI�4�a���	3!o;�D*�Ѱ���K�ݲ�����5�A `����޺����11/)#��cW@�c�x��J������=��3��E0�BR?^����x���LR /u��&%+h+yu���ʨ@bC���,�6`7P� �b2�6R�C�H��c޳n���.<�5D~��t����i.c�I*{��,�#�9q��9jk I1ٲ��I(�k�� X9�V��G��Y�j�/TI���pB�®:�>��W��B���jHiH6Ĺ��_��u?�u��:����h�>=��3��W�y�8ANդ��f�eMͷ���y��I�3Y�ìC��8�0�y���%��,�lPk���%)28�����H�'����QhX��r�B��3�{��[��_�D��)��t���P����[�{S;��LUrf=[�^�F�"�O�K�)�e��ȵ���|�����.N7�tO6��dv�7��(���ep`�_�/�Y��*�5��+�O�ߞ�rZ�e憺1׳�����C��e�X0��1Q,���`��F�mR�'R$VR�����Ⱦ�qJ=E��3�=ݓ{��a]���������yaK���z��np9d�@P�m�F!��isfD�F��@�W'|� D^��ϵ�D���,�|s\1D��BXw(^�8��cdUzo�(2O��?=#��a����G0i����H�Cu9V��;��  �Ë����f�./u��P����eO6Ȅ˭�>BɳM}?�%G|���Z�?6q��pwF����*���X����d3����~�g&|tEܓOZ/��4�@������Z[ڴs`B��o����M�;$"p#�����Cw�J��=�zt��=�2[O��Ɔe: \&8��B�����̢��"���ą���8�'��ɠ�	�Ԛ#��a���mm2:W{X	3��b.6|�WW!İՀ�]&��ޱŒ@�1��*3�D��֓���Fl�9�O\GF@@��8�ƵZݮ�(M�_����!x����;X��3�����OB��Q?2Y{�6o�I�+�=az4ϝ�Plz����}:{�.����C����Y�̊��i�k��������_��������+�lɝ�6n�q����ۧ�DhY[�u���R�	]�х�ev���Ӯ4�/�}�_��iJ����W��j��d�BO�YN���?��m<ƥ��/�Tl�;5ꕄrm��M(a$���U��GE�L;>8��z��K���5c�	�O0f҃�m�2�c��o�Mj�K��� +�jD$�F�$H�di���Wh�{�/*&�e�[�Z���/�IŸX��G� {�g~tC"�:U�kOp]��FҦ��H[Q41�*ī��N�E���m��p���Y�]�:&9c������o��w��3�`���~��4õykhy̆%fl�U�O�@���;s�b�LQ��Ek��[����$�G�����lX�%-����9�5ѝ����0��TN��y��	�����|���:�	�2�-���U\sy�Ńx��1���[� ӏ���qbz��-ݪX�W?��h��Uz�p4Õ��Ӭs����vi��y���Zߘ*H׈�{	��1�F��n�cB�z�m�=bС�3����M��m2+�hH��#B,\�����Q�����၀��qd∱co�3���u���}��dG|��r�����(�gCr����4��j�J�gZ�*�o�a����v�&��,��10cc4_��@>1_�S�,4)�ӹ�G����Ƹ]�����l3Q��g#���C����P*	��x�W5���*��J�}�f�_Ym�Y@���L}�tmt��8��?S�X/�*�넅Ur��)h�/�K&<��ыv�ޕ�#�.���3�~��]��?E�ֶV��͛pn��'�i9����%�����b��|�Vˉ����~��/!ҟI [��@z�A��;冖�Sp*���bto	�/��n1b�.���P8��Tw�탓�y\����@F ��@w2��n���'2�2,_����5E��6F�_�VE�&Mچq�����C?��t}����ܠN3X����t�Mە.?�;_��E*�t���c:I�ң�^@R�O�}1egH��Dw�8��{'��$>�=@nKm^�D(@�,h�{�-�� s���I�[xה�i&<�����ͨbp�̪��M��3*�`��Y�[�$��)�5 ��b��Mں��#Jʎ7 \�kгU��Ab�^�:k/l�\q|�v�h�����ƜY�E]2���!�C�:���և!���`8�[����0������������P�,(k*Sc��}���%���~A� �zE�H��h^�߫>�lkW��c����^�8�߶�|.��j1>[��\���g��vQ	{���fJ){T�#wIJh�#2Q:�����իE?�y3s��H�\�gm���?����i��V[�9+�TzZ��RYd���I�
�>oA�."����poׄ����X����:bC������I�jw0.����Ot��@�]ɏK$��j��g����?<|GFQ�'����U�:p�!�G��$�`}�������ye?i5��e�e7���W�:��\�b��#e�M�� +��٩�E��`k�d��x�p���mp�"���i'�1�e�&ɦY���P09�<D,Y��Y+3Q']��mQIZ@lUq��JQ�{��ݺԲR��h�|�8���D�ϒ� c¥r/��@7ɔ����f�EBke���+/�]e�����gM[#�d�
<�<�i��fQ�]����f���R(�.N9 Gkiߦ�2Lvz���������h�N��$h��) �7c������ˉ��!��k2]�j�m1�%�2�-i�����GqS��LDQ��z<����;�� ��/��<��G��s�y�3ݬ��/d��5�R
ן�ӆ/����S��)���2A�<{/t;������ϵ��� �3���ܬ�i��[Z{�Ԭܺa�á�g��%�I�.f��t�s_��p#m��=^�G��ki3m��W+l~�-�(������ ��f��_��W��}>�K4���9ko}-T#��̬5��'�; ���RB�G����3�n^p �60Z�8I��
����W=$L�PӼ���H�e'��,/�(�R5TJ�WbGN/HUb[��p_+����t��rF.h�z�Fj��������.�)�+M��V��w{T�z/�O�)n=�{ֻt��M��Fn�t�.�Ҡ�������
�6�Ǭ>v}H�.͊Wᮌ1���t����>��b��˒�S�����:/a]Sm�0�wp���#�V�
W6ܟ,�A�����(��)�s &%k<����0��z���+���H��Gg�H�Ф�(�Q0ș�4��ћ>i��&)U�D�f���l��-�	<����k��T7�.�����^�x\ω��X����`��5VU���c�׭��q�i[
m���Yν[�� )mEC�f�_����C���Ͼ;�k��g���n ���Tb�Nhz�������4���|]�Ħ�ǋ�a&�J!]W^�m�PG"oR�~�~J_�?nj.G��]>̫��n�K�)2[}�w.�=1�9Ȅ[� ��:��w�h?�ɩ���EQ=�����Y��1c��b��*b[ƪ2X�y��|�
Q�[+���G3GA�j،�_��F�g�{�ҍյ���RQKb�Z/�v�J��i�ԫ�C�����>�'Ή�%����|C^q�]��YѤH�E��ˣe�XQJ���D
7X�(�H�I����ew �Z`2�H�܁3�_W���;�1���T3F@�§dw��-m�K��k��Q��7z��D��&j*)T��2��>]QR�^�����w�;;�����n�T��dI_i��Ls�w�cՠ(�q&��'x���d�DD4{�	��AQV}�G����"4u��X'(=_@��=���3T��e��0S^n	�E���k���Xl�"4qj-]�6
&+q��N\�����$�"Mj�u`c(f���t���>Px�<J�h����<Fo���5>�<��<�V�mN!�$_��d�_�X5�?�>�x�[����6d��<�C�$E���6�7
�-�LM�o��p�7��v��#b��&�<�r�⣼����B�����ce��� ���h�(h�����ӓ+�Yhy�e=��y��|��D�f��u�����,JfO��EC��u(f�1�N_<�ɴF�Q�fe}
'����<��b�0��t��i��(��m�|�� !r��'�ہ����1�\e�,)�qB�,
}T��t�����<�z�؄^����vn�9+3�+�e&>ދ<�|]��3ܕ�ԝ��]�oe̞r�`��=zy��t��E�z��ŋ��o6��\l�-�}�P~���N���(��a��a��w�M��5$�7���WuT���s�_�4�O������?�]���V��੡Z`	JSZ�o*i����p�r9é����r8l��Ih�	T>�:�U%də���c�B�
�M/�S�up�����s��pT5�V�P"S\��������	�,�ݔ�-k��>!�	�߷��g�o��l ��Y?��
�EѢ3��k�FS�`O�m/�#&+����,c�����	n&�N����9�i&���+E���s�W��d̰�s���'�cT����W�d>Fk,���C�&�z�G}!P�'�L�J��xo����ӂsK=G���Prn��f�C� �p�=*�;������v�Y��u.�
i���ɡ���Y-���,b@�ZB-��(.I2`��9f�`������@�Ј8�Ҋ�D^Z�k�4��yo�5��e��%�l�1�ؼEf�(g��R�Q������S }\U寑��,4���S���)|6�]���j�dj� ���⺕�)��f%�%0W�@R�����5��鼶���u��S��O�±�#zt%��Ҭ'Ӹk-P�098MJy�,�� $ǈ�"����wo��%vQ��~G�q��R�;f0��[��Y��5I�&XJT
ϫ0Z������M��]���m]��/���j�Ibq��p�yl
�Ճ�]p91K(��Tr 佒yB��1��}�w�U�D&_ � �kd�	v���3�Iq�Ϥ�j��H �)b�!/r����+�9���v�g�"�+�����O�ӾvxpƱ��[®y���m^/�~yJ��_�2���&��ǃO�RS�l�#�;:M��Ջ�DC*���[�;*_��)g怿�7�,������p�塔���yu<�8�^�;�)�!��a?�C<�ᩁ��H�J�`e&��#X���64��3���®���*�Fi�B�������2�.g�@^=��w�;3˷�G��Ɣ��ӽ�=��+Ri��oT�sqa���ڷ��'��z6ꤽ��ܰW���w��
7�����KS"�Xb}�$j�s�MWS�)a����톘!���©�^c��Rs�!���Iw�-�Irkoa��,�g�qw&�!	G@���u��]�T�����#��~��O_�>/Ԅ!�S9Y�8fD��C�%:�qE�����<,�j���TpNUh����q���&�c�*��-@�����q!��(�jcd)�V&C�x]�+�/�D}��S����t=%�XVMHLt��Wc� ���^��~^��	(R�7P��f��@J���eDTee�*V���T`��黀�^�_��� ,�R��������q� ū�?{�
�P�^�6Y3.b��}U�(����c�r�ej0C������sq�Xwȣ�� .S<�֢.��\%,���/ٳh��]���6e�vA�P�g��.�a-�|�v�^��/A�au��L��fT��H�B��t���F�}��UeM��A�RB�r�S�rӗ�5�R�����'��A��f�$�ă[|�����!�l�m���`2t��Mlh���m�E��B�~�oğZI\K��'B��̸�R�I)j����q#�b��g'gTWa��$��ǞNf��^�}�B��y���r�\m��6���9��J�p!��H82ډ^$�1�1��4kSI��zc6S)L�p8�*'TL|$G���/j����Tá4��cX�M�_]H�g,�+#H-{[�0{\Ez�/��﫡�6��^��5�/w����1�9�e�'�}
����?����%5��MP`$nTD��=H���P�������Ns����/��(������N7`*ȥ��y2q��������3z
A[��Q�E_K���umӢ�D�f��8�ݐ :�ԢLmD蛢�w���o!��!���<�}/ៜr���u�>��d�����%D�\H��{_G�ݩa�V������p)�i�٪���r����K��/��C��`��Smt*Zp%b���X��ʤ �c��ٲ�*��4$�m������8e�Em	=p ?�D�ҪF�>y���Dեuð�P<h�u���H���˱��7���f��ݴ����\5��rt��T+��g�� F��^�ZA��/����W���{�)ә	��2��UC�@&���c�?85����s(bMC�fiB#�Sf���7+/�,M�2ݼ:;f�hF���8rS;q�¡=�׫(���/#a��*�����{��+��΀B����w�ωn{ș�Rms�3RS�Xc�w{9%<,h��]B�M�(W��PB���0cU���qy.��L��"т��prnH��s)/�V1ۢVOQw2q�[�ØHw]!�^n�>޵_�X�6�EŻxz��ty��6�Cы[MEmO�n?�
�����͸Pn��i�j��;t�t����!��/v����A�ɽv�o1�TE�n���(M�6cmi�N_�� ����"N�?M�v��@�;�V�����g��L��u1+� *'B�.� �k*z����"��p�gR�9�Qp��S���cd]֞&rn�@�x��Z����1׬@=�4<�V�r'��$��u�CB���V-�~mL=��	�t��V���"o7~cD���t���'�$��T��&.�����mܸ����{�U�)�_����.��I������hGDԚ��JF��F�S�3-OZ����m3m&�ɟ8k����[-->tTau�B�2�t���Ee//���ϧP�s�"&���-������S+T��cd�i���[幽|ĸ;�yີ
SP�%ў�De��,�W�ى�ζ�r�ڧΪ�R��� ��3�W�X���M;�"%��f��`_>+$�/��S����U�\�qY�s�A�K��ǫ��n_̈́�k��&M_���+���q��	� 7�:;�ܶ,�\{��E� ��Au�Xk �L[=QOL�F@���<���24_���.�vK1`s��
!Wɞ���,�J��r�m?�A�l�5~�e3g���5����#� ��˒�>B�Tz-�����1�ܬ���L��@"��	h��C��8�4���1I�O��_ _pg�t�����:��W[����7Oy��B�����g�'43�r^��1X�|�Nd�v�&F�ث6*OR�E����[.��+!2$�����^q@��l_ba����sE1��6�.Q���@����QVy?]�u�@S\Z� QsQ��x���D<28���z���f��!b�o������6�w�ѩ�$`�D�q�]bu��5C��:ﰾ�?�~�0E�k�ތcT�#O�}���V�B�ɂ-�8�H	�I�u�2�i���	��'��ņ��ox^�� �)�(��B���fGѣ��[\���r�N��SM9���[I7�i����߈����*�!��'��U~�gۺ��wǠE]���/~7��hq(0Wf`��0؈�`�i4R1(��s&�I�����c�]��P�Y0TN4��-+Jċ�������:�Mv�jү���(r���|���G���A(�����=�}ߣ��v1>��a3�C1WV��9C�R[��kN7��:8�9еu�r
�����8�>����+x<Q�Y��ԧ����)W�zs���[�*�7YL����|� �����[��ܵ�V-t��6�AKl)��T�S.k��w������ڹ��l{n�S��s�i�柖C���͊��i��|_�� �Y�o�*݋`K�v�f�.�Z�ձ����E��N�!�9�9�|_=�_VI�	~lEd�cr,�? T��ϝ���������G��\�� ��}��ëׁQ.�h���]����� "Z�B���(@e%��1�b	�g���̗�����C�sc���I>����;X�2�n�36Tڡ��bZ¢�@�zٗvǊZ�����0�e0YI��z�8�c$l.8�L���z��n��W����V���y��['<Ru*9}�(���D�� e$�g��(�6�3����?{�x�r�6�]��C?���XNr�׮ۊ�}�IHK�dԢ�����ǗNr=������W��H��_��!Nc-�7j�dp6�xd�'	���8�&�,����������H�*��%����D�=� ���2�6BF�_X9C��V���<s\׻B���S/dV�/n��S���7�Л�@�w��n��P^ӊ ���#�u�I^���=�����>AC�9�g[t�NXjV�&\���O��~��#u���Z�@�nwm���y�7
�s�l�c:�S��F���E�Ë�<�m�u8�+������xҪ^w�?���Ү�A��>���oZ�t2;&�i*h-�8g���)�U#� O�X޲@�����"���CK�
������r=s)���N�B�RE��3�h�Le��Im�%Qi��zI%�⑕�~i^�ȝ������ѳ���jD���7ѱ]�r?���۴��0���c�9v(��UZ��J�s�e��=�����=�ϱ�ިq;�TO2�jF|^�5���(܋Sm`
�Y���)�����C$̔���Ǚj��A��@��� 9Qd*��E�K;�已��XX<�Q�q�9���`��e<��l̖YSe����-����V+)�mE����R>�Y�.���}>��䠨��x[1x� Ŵ�U*|h�Z ]�-���s��5އ8�7"4�[/���>���O���  x��]+>���,k)��w�͈�S�S!E�,)�Ek<vL�-���]a�A~Tf�,�(�uӟ�d��]�IyJ���vZr��t]�^FQ3�4$^A�Q����J����X�|Ժ�͂�5W,I��X��ҭ�k�y��W�45��7���'��owWj�+O�DM���;�h�28�{*ͨ�b>K��$g�wD1� �끉�S��}7)�Fē~��f�&,�ٟl�U{Ǩg=����Zl����6�S���L�7�|����Z��U�DE|�ݤ�e.��yANt]ō�e&����pF�nT6&��a�e�k��p[,��zʎ��׏b�ߩ8Xw��~��ꂻ�	/��0��('J_^����NsO0��K|���;{Վ�Z��UF��3-3ɳ�yА'�ZH)�����f�1!˝Q�>��� �6��lP�>w���K'�t���V�@dt��v����+�ٕ�qZyIx`^N�pg�%A��fr��]ā�ԀJ�9�Y�����w��iz�4���K�c����l�L$��@%�&4��!����E�l.�ߘj�}�,���0N��ӡy3f�� ��2Z��O#�jMܞ��%�[Q̉aONQ\�0_���[;����:�E�c�D3��]
�]Tu�D���h�3A@]; [aN�8"Ҿ�"�mc39ߴ9�I�����:jU쟁O�^��ޝu�@1��+�B���ގ6��K�|�~ �b�b��Υ�H
|�4E �?Z��J������͑�,��?�L�=x��7���z\�g�tC)�u!�1���c��YM�.��;�2B�#8
�X|E�.`�� i���*@l�q�����QQ��"�$2Z+6r�����V�Ʒ��}<�#��e�^�&�=G�"���Z�4�w��*��?r��ie�Ԏ�NQ���<d�ך�(�[����Te�����R���)�V�dk����9cQ��#�&hO���S˕s�iwB�K��Hva���>�D@��\�6�� P���A#���ʌ؈$���̧�g�4����˃�P�S���𬇶@q�wPBcj�I��-��w6�P� cN�{�8�#[�"�q���*Q��p��]�� ��AĆǋos Im������ �����y簐��.�sc���y}o�d�כ0���v~%2g>�>���4.ʗbP�V��A������Qx�
��8��6��)"�O�-����6H�l7De��."Y�P�Ù������zV)/����B:φ�L�9��}п�:A��;��H�o	O��L{s��\`���P���35�6��/�ݐ��ֈ˼��|6�]XN�EL0���6�Nɖ�%%����/p;6qDFD���UF� @F�m z�:c�w"e�2�-����g{�*�v�4x_n�	�Q�lA(�t�i�a^7M�qi]I)�'���5}b6�$�ߏ�b7��oɖϋ`�؟�]T�;U� �|�@$�ւ=JaL1��C
{��[c�-Wڎ��~}���G� �q�ʓ[wj4�0B8�7��z����lus4���ZU��iňIa6O�q�㷶��͕���ͽ+���g��:*%O�Q�{~r.ky��^T�[��}���������b��� �#x�{��@�N�份�P�����^�~
�b=�m1W�/T��<�wl���}�|����lP�P{���Y��I�#F�ͱ����E+i	����')���s�LpM�7�y���s*���d���Bş7g�옄1h#�J��4.G����o�J��j5�<���&��;�1�7Cw�_NN�A��D�9�Q���D��(���	��Fh��L�K��������dc��9��}��W蒓ٵ��&������ҙ�����(���i��.)J[�uM��/E���y�Ҿ�ۦڅ�"�1��4i���ԩ3�ƬP�2�a_C|I�1AH"Y��7�?�˛�E˸xQ��}ϥw ݧ�z���^4,��p_q��ёT:ҵV����w9l�c��i��R�Գ��$v#��
(��1U�	��ڣN����L�ڠ�oJ�]��C�0��-�U� ����e��*̭8�p|#A�B�G��6��֖IZdK��ʰ����ʭ	%j(�j�@�[����?=)?�핞]O��������п�x�җU9�qrL�2Ί��맷�����[����`n��?��>fP�ˌ��V7%�A��Qb~�
����|�В��X����koO�Ӻh��aUS,H�~ӥo{�/6��]8��g�r���;B��j������bT��Sz����:uW$p���u\h`�ĩT�ă��ul�#����1ݒ�l�j��<Ky��XL�� ³�/f���~�l��8�?S怢��{U��k��)K�p�t�����m��n��u4N*"D��鳹se��Ղz�~��e!���rta�S���/*^�x�$��<(�7
zݸ��Q��0�W��S��*�㻏�ʟ�/�k�k��%%���<$8�q��,�%�e����1�7�",�B��Y[;�Am��f�|�Z��J��$��w�jp\�a�B�޾�$�*t�S%>Ť����-g�
ut#�Í{{?S��Ύ7-4e��N����RPA�!@��)�|\+��RL=y�q�<��`S&��ˠ���v������Bs�3a*��N�j��aŜ��B���T�`|���J@�M�v%�����:�L��T��[4�6B��r�@��2C��I�"��A:�.�r���rd=w2%3E�����d����y�����y�,���\W�!;�m�������\�.�������G��bV���>�]QԤ͢�
����l�Yu���,�%��`�����끱%AZ�}s����aq�Z8�/�"�LG캃��sd��P�J|ޢ�0�b���(��I+{,���$�����
8?�4I-�R���������X��O�p��r�����i�g�:�s�ה�����5l��FL+�������6�⁕� H??:۱��n�8����[-#ڰI�[WR�w��6>�����e�83E�ɲ��?}!|��L*�Q��J���Yc̗������f�����L��uh Jx��!���Ǎ����Ps���M�%��!�����ť�D��?���`^�.O:i�"��Ϻ/�|���㹮Igl�bƕs�VHv�0Q�i���C}��ڦy��3Z��}6�r��P�(�N���u�e��9�j<Ϣ�~<�#���罜O:��_7���y�u�줁۪5JH�d�rC}��b�q��3U`[�9�g<�P�Re�G�FS/���5�d���*�n=�E=s�T�c`SRi���D��0Cܲ�#d~��yO>[�� ᅌ�$v:�l���T���@w �3�P�A�#�X�c���t ��f�%^5(��?@�,_� ;� �(-��g����՗���m�Kuq0qx'�kB��}��o��%�����"�S/�}��p$�N	����տ	<1�OVy�OM�?*�k�,H�p���/�ڵ>��T�rUx�A�j�����4_��Ɋڡ�ɜ��:r=k_9�#S�GV�ɸ���/���9(�q\��m��Jic@�l�1o�1q�h�{v��{�f�C�1`ͼ�����_K<�@򯤔Dj�˝�d$��L]ա.rjT򢟺[�����=7x:T���!�*���@�N��= ���`n���R}�	�+�Ϩ ��kJdw�ik�Q�1ԟIҽ�+�'�0���Qg����,L�F�?��cD7�L��[4i�n]B/�z���T��L�Ij�
I㧓*��eh�/��#�ۢZ���dĐ��3��/��ޛ���S�B �o�F{�����\�ļ����`;�{�hEQ �z��)8��֓5g�p��Pww�X�">�L��`��
�ַ7�V|R�?�����L�=�Ѓ_! �Q���>i�����]6tn���xy�䴋�#���� �5��{���M�*�\U���9���-����f��Kc�H�2:D.�:ԓN?sq�@���i�V)l�������:�RN/W]���;R�x5gX�pll��yW4�z�\��&V�(̆������]K�ŢKH�i��`/n�p�'ܥ���֑H��)�c?*%;3]����C�S=(�%��$T����fmW�C=���YZM�h���!�e-�' ���eͭ�lg������3؛��� ���?����'��!%�h����<IӔc��A�$<0Zf�L��ă�=��y vEoyp_��.��1�yG|=mM�b��^��/�}��Ш�s\��-cYh�d�@\��2]@ͭ��:��׬"a3�Ro���g�Z��a
�4(쮥��2i�d9�����pg^h��bK��N�$���e����"��8�:]HJ��(�!�)�U6��I��Xo�W�3N�/l*���L�7n�����Qa���5��.Z��J��:VJ������%
�ŭ�T�$���P�
�*%������x�a�tu���5�R1�ى�W})6�fH�ğY�J�=��Ա���2C�
���a��T��6c`�������)�o���r��+�[�*�)��u���64RP��op��3��}��i�[����x�sh^�8�X��[K٣ ��&�����5�n�BE���EC�8�b������լe����{����W�q�8>���ݏ��`ŪV�˔��sl��M��VOo���I��lû�~��q/�ѡ�=��b{���eXkN'�=���ވA��hc|������y���؇h�\��m�R:�Y�������p���B��ɂSZK'Q�� {C�٬f����#�d��t��Ku��J=����<�/�#�W�R�Μ-0�����ż�Ӯ݀ :8��n�~v��$����5���٩[7-.�Q��Ľ���$��ތuÉ��a�/�"�-�/�	"B!����؂�-��|@7��:;'�_���D	��65-X�X!K'��g����灹S��d�q1�����U�[�k7�CFɃ�7�y��h��b~�0�����1��q]b�9��d����eՐ��J�]U0��n�����ܧQ��_��66�n�ʩ���蓏�K�p��e��A��z���'�
���L.�y���U4�kci*�PX�7�N�Xf-�qN ?���Y28�׉.���ٳ
]_ 8m�ߣ�bn�?�X�sO��>w��%m�J�sA:@H��fs=*7�����@m�y����j�(ơ�:@5�3'�X�.~rs����>����\.��iqo[4��e�O�Pyy%���jl�n��'2�s�~<CG�+�S��A $��k�*3B~�>���R�Cf�w|��@�=��m�ۡ�N�D�OQ�=l�����������HYXRr=�^Ne�љ`<�TV�a:��Lq�˺T���0Dd'L�l������~���8>
,i�0668�NO���%�_ۍ�G)������g�7��[�
�q����)@<'��2k�(X��$ת,$�*z~�M|%�*>�,�wu�M�5�%0��a�u"�(P$�T�M�`�6e���D�z�$E$�/ob��Zx�@���.YA}J=�MqM�v7�	��_ �v}�g��Gٕ�6r6�X�����ƚ�,�0v���7-�e�E٤����5@�����J&E���pC�sU�*9W)|��9q�w��o�҂Y��/]�+�&�^������k��Y����#e�ު��!��,�up7�>�>39H�T!hlpv۬�-��ah�,�Zll�zT��x~e��rG����H�w<��Zn����#is��|�bF�򳜁ϰ�����;x:Y�8%\����f	P�vGK\���Τ���<I��+���`91L��|�zT� ����:�b?�w����U�a.
jP��]���2f��eﺊU�&J�y���Ly<��w^�Xt��y���,�V���Q���`�Uv����u}⥋� �wntKA��n��:ła��N����^-�ǫ�hsٜY:��@� �a��iI�Q�B�K�}�z�� �A2wP�q�/����S�u�
�2�xCx�H��Mx*Do�6Ȋ{+Nؑ=
Ǭ��h�Z�<�3Lߵ�Ǝr &��8.T&�Lˁ��X�W^�o%i�[�tq�
ǣAT�^dj>����u��~kkK��N���ݢ@�o��>����k��q7�
^ʱ;@eG�`y�,}��[�H:6(ݑd` =��6��h�y����}��#X7�ݝ����t�F�w�
�fБ��~M�[E]`�f�0	�j�v���w��+�n���~e�2�#_,���� ϔ�]��Ǟ���=|j3U�ɘ�p�6G{H0�%mBvtL�/L�x~�<�)0���5��B��Xz:�h@���E��]j��'�oT���i�I�'R�.��%�wQ؏@�,���0��5z#b7^$:��-Sj��^�fu�,�S������-渐�~����8�.� �CX�H���ގ�[���ƐǬ�W{�<�/+��(UK륞/.ba�8||�f��LY`j����JE����J��HX�W�S5�X�>)�Xl������ �?�=���������|F�ue�k\�-pW2o�4��AnH X&͸'Aa'�����h���4�+��6������h��Ǎ1�O	!�����:>#f�%f�>�UXJ�#�tq��v$p��Gl�ߠ{DI��9�V��C��B+g�Q@�����4aQ9�CAH�g1z�Jɭ��5{k�i�R�c4���'D���>���o�9�?�	)�Ll��ap,�#��G�q�p�IH�6�&N�c)!��"l�-�V����f�����h��&~� h��I:���{�m��-Q�7�1q��H����k�g�U�F,�i�=�����r��l^�1�eIj��Ձ�ĸD�tS/�f�zr$�O�vbq��N�6�q�6!.n�/����Ǹ�cR<B���AZF=83�U��~ʽҪ��+l�Ճ{B���p"�6a&�B7��*ei\�xyX�j�B�v��5��%�t$�sx_K��و���өI��Th�}�������UGv�+K��r_�J���#e;���z���a��1���mo'[,T2�,�$8ƚŸPЌ�xP���Z�������>,�����G�/-�;4V�*B��pK��T�W��@h�4���a�'Q/~r�U��O���$T�z?�*���l�����K�`��X��&�j������g�Z
F�n1�]�
�����&����,*��C8�kDU/E�z��Q(d��r^[ұ��%����r��V�w�AL~�!/��f��_bSD���R,BH%AG�&s��1|��:�Y Z��-��ot�|���&�n!}�<C&)����~��un�%k���@֦W�T�u|��$�m�t4�~3 �`P��M`c��ʥ�� V�Ql���߼�篔����JJD�{�� ���nop~�o�k�ȹj4�ј�#)�)kl��Y��|�.�U	1����f��3�iY�vEP�L6{�W�U�Ҕ5�ڡL��o��#uxC�(o�&3b��x�q���ʲ��e޳��E"�+��B�WMסmw2H*���QB�~��u>Xá��Z�A�,���Z\"�6�Ա��7g�*eZ�Y�$!v�e�/@_��`m���0rD{Z~��O�𛬹t�Ud�ed����ӈ�?^��Ř�ǡ��=�<c�~*����q@f��=*�ؑ���x"���۴Rz�P&��5�H�.���i3`/%��ScL-cѾ�
�|�t8�~
E�nH��%8v�a�W��me�,�[o�zj��ـO��6��𙁜q�K�X��Y`�oVA�M����.ޚ!TZ����}����e%��R��$����XDc�ڱ �S�S��
��f�̍���Nn�0մmҏ�Je�E՛M��&����x�_�3����L��&4)��"��W�4�f��xcw�x?�ޅe��Oye2����}S�'k�
��md���7�e�����; ��SμC��s�ՃU[n0:����f���s�j��G�a|c��F5�l�ڻu��;7z� ��� R����ɋ�`���%��)����{��N��Z��� p4��X�\��؍��
�a�.2n���[Y�C�<��XŲ�.�[tۼd�S�"ǅ�?�X�P�,�si�:G���r���:��2�r���!ͳ�"%`��p/&�T�:�`�̉me3����%�ZY7ZQxzDB�ݥ楫�0�a����)�(��g��U.)4�Cy�ُ"0Cqg�$J�%ͤ�X4��1E�%ڲ]]��oq��o�y�x��]�02˦��S��<�@�r�-�О^1��=5+)E3=檃��>�`�h�Ј���8����9�č��6XTJR�bn�[���݁��O\9zE0��h�6�ė�텪�[�=8��bu��k��l�z�R,q�Ri��?��+Q�{��˅���s�o3��}�
��̕g'-�S?��|N�]�<B�X8�����R�������%�8b[�H�M_��*]��̬����ߴ�/���0,�ҵ��a��=3���zְ�ei��:q���P� ~5�
u8'C��	���������|9���Q-P���RJ�h����E���A�k�����ėH�>H0��:���t�^���`� �>5Q���C�208p}���	h�϶q��90<I��2�)�ϳ\��@y�U��!� ��/5&� �fKG�LW�_�F?�&^�!�����GS�b�Le���@�172%�����'e#��w/���3�w���?z��M��͒\�,z����<�i؞g�I$�5i�|��>JG���C5
="�
6��l�*W�Og��9���5.��O�'����`��+n�Ri�}������'���XE�$wul�ꤏ �����2�`o�j.}�ɵm#��F����Y22�rǇ5����I!nՋ��"��R=����0Gj�Eʯf/c�6�����j����!�(�VA�U�W���I'�sY9~>)���y)��9,�'��������ᐑ���|naϜ���}!������"���0.�'�|��/��G����,>*�Ҷ�s�(K��ɼ�ϟ�j`�x�,L|'Lmm2��mE;a�
$� eU�"Z�`��Bκ��Q��"h_%�y�*��f��)$����A�RܒfA]=�|xBLݢ9-�%5}�5-��n�>̾�e�C8�-�rPh�ܗ�b�?k��

j�(���7I���\G�����&��!'蕟�Oa��у����V�RC���w��$�4<-���;=���'�0��T9 3L�C�>HW,I���э�g�����b�*D�"L�XDݿO��j_�r��:�.������ӹ��a?g�;I1�[��,x�+E"��ܴM|����1�60���x"Kc�����tC�^���Z?��x��Zx�2˄>ĳf0E��ߣ>t�,H��v�wEd�Z�B�����ʀ��,�jx�f�S�9-��yG��R��ʝ�4),��K�r�2-^��;�Oo��K6�V�,�[������gOx��6����+�#ɦց�^��X��J���3��\@س��t�=�ч�1��C?�!�?�T���&L����	\�շ@m|yw!���񼛓�or�{�K���U��dF��	;�uf^���F�e)a���8���������T>5��Ɏ��P[j�Fࠋ� ���&�j���\��6��ƀ��?� ���$dd,OK٢"�n)���L�39��,0���B���É��Q��� 	bҐ���L�����8�Y���+(ZKKD:�+��c���ۇ�xQ��#qP�9Y��d���6�����g嘰���o�1W>?�тkr._�[��+
�lԪH�Θ�==mm�����a�M�27*᎛!vp����$X��-AJ�KA@|�0rn{���,���9������ A�A��p6��K7�K��>߅��i����a�MC�1!4J���)� 6�95.�0ng� ^��п2�s&�!�&U���ڻ�֙; br[�bo�]�ۛH��Y�;ؼ�������:0���Y�[�����]%%Y�pK�G�ٙ��k�D�r�n�;�M��Wn�`+MSv�b3P�M�a�w��o-Ƭn��}�1�5^���T+m2�nVc���o�l���0�3W#�'��a�r��w @�߽b�K��'g]� �	���y����0��B'ofԾr�V�����.I�$0^Q�`�yC���ya���F�xuU����ߑF�=ECh0��[w�OŬY�v�-�B�f�Uv%+�<nl�-��T��#�)8��YgG�/W�u��^`r���ֲ�J�|3��abN���;�ۗ^CjN�3�!�d�4�7@	���<���5���Θ	���ϯj������R73�3�=-�b53i�_��M�|m�b�@t3�g�f#�APz�q�����)��c�ق0@j^�%'U��	�$�a�T����o�=1�-��o�*�*)��$ӧ������'t�ʵx�X<���I|#�q�O����WW%5I�Ӧ ��3�<Q�S����D1Q�'1��q�@�T���p�/�8�R۟�`�I��>�26-đ=mcJxv$<�J��+�8L�9��=\ ^��N�m�R�m��a�3��o�T�e�W�&��Ġ�ET�3��6޷
80Q����^/
>�������=~�D�U�W/γ{�,�A}eS/IIմ��F[�!MN|��x�r���P}�2�7H�Q�i��,o�.&�Y*D�H�%��!�rrDoI��=�V�l�r�@�#�Lܳ�ĥ�bv�:���?Y���IBŻ X"B��Q��3�i花4�Н�A)����}�]gT�~�A ]��1W��co���}�.�$&�L�����AX\Y_2����Ԫ��h�L�K*��7���^��5�"�ѷЕ�$�6�n����:��Ç�����t����#�p������#j��=y�[�Tpi,S�����,��ݠ�
�KF��\���.�b��-�ͽ�o��<5����v��c8��1H�_���-����#p���p��O�k��g�nj?=sj N�l�l�!�D���"AG�)�
l�y$�0��tبc֊��$�OOl��g:�Pi�M�.�i�4�xs������y��J']�6U��kC�jx�Q�5Jr8z�w� H��1	����/���L^�Sb�iu�o�H>��k2���U�~b�7��y{�<�d�~�x�i�l+��B�)��Xۭ��I�Z^�ݐ��Z,��V��Ӡ+"#yp�w̆!U��~�J�K��?h�F���2F*%[г�/�bԼ���i�ɴ.��5�j��ݡ�.hhe�9.p����1���� �q�$����8)�C�d��p	��.��3L���ixቱ�ǁR�ygQ�r~��@�L �;nD�+$NU�����Ѣ��>=Kq隬��qR��7�g0LS���Hx�@ejK<��v00������m�	�D�fAg�"�������Nd��W���?c;��0@���'�Hk���q=��.��Ԭ̄�to��Q�[F�hd̾6 ]��v��5NhsXO���eX�/*?#W�:D|�V\�į�X:�ֺ�6���e)r���%����b_�|0���{�k�bG.gUM��l7�f����/.C�Epq����`��F^J�\�%H�3�v�.leeK�)���Z���u��%��������;�/�.W�H�V�̴N�1\Y.�DNT�r7�� I23�X�\�[&}�̍�0�I�6!�����c� �4����>�z"c(k��7�f���S ��w��0�g��'����j�!DP��+�<�"qmv�j��7�f�	���/�р���2�R�����P�e���9^�#�c/�ҥ��^�` i��ѕE��+ZMK<}��EP�Y۽�sa���Ms\X��x0�?�� �e�%0��D��s���7��}��G�v|wbA�������r��ؤd>0�p�J��-�=L ���H�{���cMk�� }s�؅�_��j?Ҧ��$�K���¢ �.jʻ��(g��[ؼ�Vo�
�`�~����Ԋ�л��|Гy՘ц��?���>��k#C���9Q�\K8��~&�v��mȘ�"�_1�ܱxF�R8��^+Q���{f��kN��)3�'��W�qS�9|^V��tۢ�3���Z+��c�3�咷�s:��6�Z3���]�;��,h��(����9�Npl�V�3,'���%�me.����	y�������և�Z�oQI���3����5���)�>M��T���$��>��(��[����]�˚	 _��h�÷�G?6i+&���7S�fW�,������f0�����&�o. ��'��`m��'g5A�I��f&E'���l�U��D����kE���n�aуYc�_ 3�����E�#�D72*�ɨ����ӱ�މ��m0<����{��E��D<�+9�g�!Y6��F-E��{C�M<�H��Rd�$�µf?��`�y!j߶�K��Uˀ5|<ⱍ<���f�
��=BA��ȇ�X���Z ua\�5��չ���*F�� �)R��9"���P�:�����M�d�7�^y�+.	�����7�=��ö1��pS��$��&�c��w������&o�<j[�E~����E;��}��f�(� �`x���3˓uC��Vm��?����B�B�4�B�T��=<96�����UT�y{�=�3D+P�K�.N�(�=��f��	�&(�v!UJ�h��e�$L�����z�d� ����ѯܷP�0�.�C����@�Q?����g}����ߚ���$�~y�Ps�<� ɯG�_��n�Ҥ�ܻ�'�4�]��ϵ)՘E��K/�@�R������Jp�>`y�]G�a:i̇1�s�z7��� Z�"�/���U��H�.�j�������fȫy��չ+����j���Hvƒ\�~��v	v�>k"\,=�>dv4.$I
"�� ��B��)�͠��s�ƣ��b�޸�lF�~�k�5��I��XB����_*�t�TW�Ru�<D�(G�����&�!�ܸ�~�)Aj)�ʗ���S@�����,�u�j��D~��O���@g�v����T\8è�c��ڑ�k�<9U.�U����s)E�*T�#�-�NX�S�C߫��b��"0pp�e��D
�,��>ZQ�IgQ,l5�.�G�6�'�Z;����_^x�ƛ�2�k���o�}�������߼&v@��o��J�ӧ���rϙ���Xt�z�6��>iœ�V�S�D���~!Kd��<�%�U�+'�"�6���o�V��f����T���n������Ѱ�]wb%���Q���I����`�m��:�H?�]�S{t<w�o�h����{����v-�v&��CR��B;9�<�u��fq��i��z܂�k��KZ����	t�O#٥=RϨ�u����	�|m@{{���{:���nL��f���Z��%)2�$af�XS��>��3�Om�﯄o5TIL��K�E^����k�K ,��]����<i�m ��\���x�ek)�!�O�xm[�ULq��`���j�xZ�P�;�m����������Ө���ܰ��-����l=�_)\��~$i�}�wm�O�����3u�o������mB(1��V8aP��i�&B�Hrَ��O�F�4�_ҥZ8�,/�L״���z!��;��ӫ#%��L�6���M��KlP{7$�?��g㐤V���f-��l�dn(v7�x>�3>��	�a�����`|i��1e烅��iPYc��W�7�'��q�[�6i�++�����	��,����.&.%z���Lfp�U���o��'�+>��g�
�\�U��X�_Z��X4+uVV�s����ۈҔ�<q��N�m-�e�M��2@&w��+B����H��SY�C3��,^��u��q��L$ĥ'GgkL�EK�*#�O������xWN2�Ev���.j+ٴ7�೹��&�i7&��|L�j�y���W[O���!ݔ��5�ލj����?�ta�X��쇏�wp��Tb[괜��]Ħ��ZTFgSj�qٔ�ϟ\)��bO���7�f
�g���!�5�z��S��8n���nf��v.�@~�*�ɰC��laD�k[_-nd������H��֞�I���ץ�5ۡ�;' e'}��~����L��`bނ3�ă�w�����@��i��Z�������M�QV��?����Mw;ϳ�\�[�}��coC�l�ԘF=��g��u���O�~���X��a{��P�*-�B�I沫��J�G��T���=8��{�t~���ª�����l�/�ś7��Z_����I/�N$᤭ybf�N҅��L�$>"�Y������TcO��>a�?��A�Rk��(�9��V*Nd4�i�m�	��%l[�Z���fʝqn�aTzw��e�ᩁ�������t1�%%�jB��_�^�����RĺIO��P~k�=�W�,�ű�Ⱦ^O�O�Pr�?�k�|��u*r��TRq�3H�=�9���0%	�Y0학b�e�����> �,�AX���rh`W�'_�1�ȥ\�e8aU��#z�j���%�@._Z��;��K���M���uP��\Y?zK�A߿^�Bs�jy��[n��F� b�#�H�{9�w�g,�Ԕ�(JƝ�J�ߞ�D�����P�.�<'anEXU���Q�S�q��[��q�j��FpK�:��%���/ߋ�[���wװ"m���h�i< �Wʳ��(��2�,+�+y���b�)�o��ͧb�-��5�?W���X�J��`��_�̕π��,8�O g[Ш�V[py��Q��4�)lqi ��{�V��k|,�c�A]���sPEt�'�=?0�1ȱ]��9Y���Mˠ�*�#���M�pdB�v�hh�a��90�?��u�B��V�ʽg��)���.v��9֣���k���M��^/h�&���:���0�,]4�c����W��^�4;ǽ��_AN8c\����1v|��K�LKw�1+MJ��Tg�ˊ�0.�.��f��0�ת|�c����w������D3@�+���F9���4b��[^ �2��b���kQ��*��G�
j=��;˩��d�S��`�T��YW�6� N�u˅U����f�m�C6�&��N1t]Bē_�㦖o�q���>�Z��&�<",B�a�U���\���l'���v82�gP�䀋�
��~�L|RT�z��G�;���P�n�s5Q �l�-�:Z�+б#��������M~&�s�o]e���D�C�t��j�Y�U@��_˩��֡^��o]������xBz��b��V�pٍ8j��dF�O;�Q�Tl�#��M5��f*�Һ�:O����v�Z�E����&R�mv��@��nLp����������	CA4P����U�y�G'CJ�����������������Yf�*+`w7��Oƚ2&�M=����jdѻ���ů��u4`�N���R��6�mGl�����IN_+�ӭ��1�¶{D��2�|��僊��������I�n�11:4�p9.��G��0J.Y�����)4uh~#����U�ݯ������K�-����K�(�NE�qZT�3JB;���w�b�E��X�c>�p�9�a�R���ѻ�X�2�΢t����e"bS좂n�?�w.��rܖҭ�M#��&q$s:���C����ڋ:U�<�Y�R���E�ۍb�"R��By$ ����g"}���e��Q�d�]���4�-{-A��'���Ezw�wgW����,l��c��^G�nXoH� g�l~(>�L'���g?���_8�|8�m+uh�}:�/���&A:'e2�&-�+��ƫJ���c�5S�,��ZE�[D�(� ��"d���#g�9l�� ��\����uP�	�����I<�4¤���E����x�ib�J�\9��,��.�[Ӭ��Dʋ����(eF�s��u{��t'oF�sU��c4�R��	��e���| _�[��Ȣ�%�<Й\�r�job�έk�*:I��T�aRҫZL=����I�>!��	v�3�ٌ�M�M6���\��N#���4�2�h���~0��(�:2h��!����K�%���X ���k9eͥ�����a~�UENK����$@��'!�u*'�1��5>�'�0�<p�<<K�Ɛ�M��z�
��=�Y�r���x9=�;>r�28�7O���&=n����S�����X<�c]��	`�����`��E����*4g�!M��:�����D�39�1ͫ.�M�:�J}@#��L�+ݧ~x5�ًiV�XRtǮ���
_��������3�*T8�X��@3����6����ò�uӰ<��/���{WKw~�Ů|0���O5��@$�b�q4:h7Ѣ�ZZ߶��6I-��}�F��Z:tc��T((���[�9���m'�Yɪ�ܸ��4�O#tC�s��ܬ�{1��lHC�ʆ���z��QC�vhv�z���5�0pO ���&O@�-,w�J���v�T��`m,O�Y��������Dnl]NH��p9y�Lm��C+c�ry�Sܟo5n���T�Q yV�����MsFCgԨ�^�
.͒^�қF�W2j!��Ů�4&:1�)�� @i���r���d1����B���RD�óv�9L��ײ���ˤ/N�tΏr=x��\��9�k�' c�wj��R�'��%X\�~B�.��B9Y.�4�����g��a��4�9��u�}��V���-�<9�r �ݿ`����}��%��v�l1�ZD�k|�`�O��U�D|�:��!�v��&(x��6>X �,o��)�I#.����	��0_�Ѿʦ�ViMLҊ���N�C�#�E��|Mq�=J�90�F���%�011DU�(��w��8�@�%�$'����޻��~[U�������9
Y79���̝`�ˠ߄�&�(#A6 �jO����"����澏 �^I��P��@��חqOb.k}��>wf(�;:R���y3�x��=����/y�W&_?Bp^C���'��q�,�Фӫ�5뜪.��ăAlL\�uTL�����6�-��zѫ�A���ɴ��c�qa����x�<�ӿ�I%�h�Iy?A'?)�ܧ�R���
R0BK�)��b_�Ɖ�L��ܳ��ކ�U�Q�&q���N9�Q��pr	(Ҽ.�99H!����%e��x<�GC�M�vO�b�Q〇$�F��}%r�kps��kgҤ�l�Y����c��|�8�� f2~4��ö�T8*�(+BQ�4�5h�p7�B?�湎� ��|�0�/O���&���>e���}�e~��{��~1���e'�خh�QU&����F(�
�^����S[�Q3����gl
�
7�7��.6�@�d�Z:ގu8�&9������q�ܡ�7Y��*i	�jKswD�.�MH���,�_~W?a;��O�}����5�77-�e¾�y��HN�������f�����zj��w64�M��%Kj�D ����!���H?�4!i(뤉�7!�{���4���2�'�Ecc��*��㔘"+��Bt�N�̜��i-�5�41�`ҁ�6���o�qm]C�w�-uU��U#�,����:/2�/0tǬܾ�ן��@�+$�qo{���oQ�C���-�h������ȶ!�{�E�R�ף���%�	�����L!ϗ)��a�X�E�ڭnO�I�y�w��Y����2�w��M/8���р�fi������T�xP�U�M鵾#�]����6܀+(O悆�����Ds����f,�+3��`t����+�t�[=`92�3ֹ����q0�6��^p��� ׳i�0�@]�i��%���~���S�`AN^���j����/�CN��g�����9j�4Ot��Y�ٹ{v�O�#\#���)�UZ��8���u>�e�I��W���ձg��"�I�û&	�3n�i~��� ���Fs����+�,l8�N��/V��깈nKˈ��㉾�X�=��ԧ�,y�G�ЎQs<�~����ʢ�ٸ��#��d(��6>��ѯ��u��/u����?�����Q�"��Q		i;�TҢ��߱�ੳ�N�D̀�mZ�abg���>�M��S<�.	���p�g-��������v��-qi�a�N/�������UHy������&�5�u�:6���9৛?-&��ҋ?�.�8�X�K��Y�]�҄�����H�%G�ˢ�����R�q�ը�9�v}1g1�@��pjɳ� C��r�C�:k��{{ʗs��+�W��.�W�/B��x8O�C���+%A�w�
f�0�E\���D�x����hF��]A���ɕ�� ���F��Խ��:h7�8�N��p��	Ae)۳b奅ܫ��L3��ş�ЈN}�vv������b�V��[v��8T�>�BDr�!&�
d��t���,tI���1RR��2��(䚍�0B�}yU�bk�����"o[�f4��u��݀sV�Oj:D|�<�2J*����;�n��sKY|�sZ��.����|���d5k�1��|x+���cv�WK������Z���.a�Kc��c�G����I�X�YB�␩BL{���ee��[[i���,|�{.N��=$�t�֑��h��u ��b!�>�S>�Ƞp�/M�O�9s�zlՙJd��ɪ7#��	%�-��]u[[T�i����ӂh��+A�9V �EЩ&���w>]�"@ˁZ�:��}�ej=�ԯ3�Hn�b��NQ^eUߏng�$��2	Z�����֣r�`X��w[�����i.�3
�����]\�  if1`�D���d%�8PR�u��7�B�:��9�xdߛ��E	v��<���@ 	��ʂ��E��{��������6A�6��� ����5X���a�;��4]t��J�To������U�+�=O<rͳǟq+�̏ɿ�-�~9|�R��u�(��XP���)��K����9�#C��+��Dh��d,���CÇ��s�4�C*�%j�
!qq8���r��lٰx��mhi:�Ĳ��IR�8��dXwO�W=�?w�{2��w�����{�"�*�K��1E����љ��""V���H��ǲ�WP�y�V*Y6�4����h���]�BJ0�����-�0*�~�uТ0���G�q
���Gg���uU���i�.{�;�Jc[":ӵ��q���&�6g�e���{�9�w����l����濛�G��#0y1"�/סi�~��ۘ��`%��`�A��Z�0�F)�T,k%d�J��y8�plD��n_�?Ib< �gN��5���3�?��Lu�W�F����m>��S2�ݨ؞�i��S�<�b�=V?�@*��-�M���'�U�Tx��0�_��1)���>���#�Uq�ڧ5�%]�P"���s�u��;�pڸ�RƄ*q2�o�l��*0�&fd|u���F8�ODGB`3���2�w47�߽+��Z�T���l�������kN�c���ظ���\�a�aЩ��̢a�������	>h����:r�+uO�����nrm}$��Sط�c`Q���B�-3��r¢�^��p������$��,v�i�]�8V��8�X�2���`�HI8�}����a4�i�����ʋ��դ�������,[w��`A
��'���:�MSK75M��s���+{��m�&��>Z`
_��]�4xcK���B��[���q��Aw)t�z8L�N��g����o_j��-T'h`�����XYa�Hn��P#������L����.g��{]��C�^��31֍��^9<ʚ�������c.�����!3�~@7��{]�R�:a�gup�2߽U�* �છq��
>�WD����
�Gb�#�n?<�t��:�h�� �r}���U�k�?�];KJoJ���'y����]�Qgv�B��`���޳�8���P�'a(��q�6et����<�A+�ͿQ6��|I�4��(���+Nf�������*�Lr��Yxp0��
<�t����6d^��.GQ�<�ڛ� ���ϕN��)����v����������������Y��ABc�����Y,͕7NC�!��;/���8�^�9��ǝeU�����mX�Y�RA-��/#�o�����S��Uf���|�Q2���D��Y�������-b|TB�Ea"�ߛ�x,���{�-�L@G#�XKM����a|���A���j;.�^�K]?T5��c��b���S� �!F
��R�	�5���W�  ֟�Yj�ωH�[2���.�Q����.�J)�[Sޠ��t��@���.H�L��l��)D|����g/����ו..A �sg]�Yd_���\�Ab0�j�":���2h�..!#�!b�4H+�}Ha����D�5���b�0
ةKk��a���� �QJnZ��U^�8�5�X<����17`�u�z<�_�.>d�9y��6�­�8�7�u�cw��%Њ�@8���~MÙ9�k��jM��;�@�"GCk�Wv���k����vN.Zs5�R�/S��h	28��r+�`o`��4�m�`"��m�T�,h��x��������f�����qx����]ʹ����7q�]T�A��6<q�{�ɣ�_�?����VTX����ƸzZ�7�?2#�	�k�IV����,�F��Ԃ�W����a'xCQN߮\�Nn}S�+�V>����D��}.��p�`/�F����ٺ��U�,��1d�db�ئlh[���v!+!�M1q�w����0�0���	���.���PLгk�	��Zx�ұ�4�,.�#�1U��Xf0�������E����bc�N�|�s{�N����{�ᇜv�U�#	��M '�B�?q����2��5�R�ʁ}�d��&�G���[��Y�rJ��QTZE�\n�0�a��87�,?7�>��. ��� �L>�����`̇NQ<$�Q�v�w��p�HsiY4��F,�Bو@-����M�6~ f��>м��puJ��G&2��Q��G�X��4�ʳ7n�3��e?���V;�7��ZQ����8F/����
LЧ	$1����7��n"GжU	�_��;A��iCd^�؛��/BD���4OP��zg��bTС  w�C/z�q�u� �-,��Ɇ���bS9�٩�ǡ�3
baS�٢�(F�Q�ȋ?�<�'�����t(�FY�Y���*�[	��k%�'���^��Y�tH;�7���zD�������l�^{$�6��O �7����ڢ�������.�+��o�ؾ�N���'��2�`'7;��Nh�٧?tgN'�/Z�nk�j�_G�M��� q��~6(�
:l�1,Uy���	�|˽�\�M'�H�7)���&gx]\��¼���ķGJQ��ң~n�(���Pv՚�P�������60l �rM�h7������̃�@�0��W�/N��^�d�����T�GrX���|���[���	T��sD�
����e�/mΈ��/(�v蟶��r�c� �}�1`0��L��w��ǺwXY	��sM'������`�	AG��DDTs�
�����`���*bnr�3�[��cY�F�2c��R�E�\y������ �!�1���Cݐ$w�59e�\
K��=��v�X����㚼%����0.w�ùŖ�|�H��䣡#FWO�ld4`w�a�;�]�l'�F�,��BպU�?�\l�`����j�~m���bP]r��=���r
[����^��T��M	K)V_��:VH�*_�0
_����N,� � ����L�>��[f�'�!'Xi-�
 >7u,_}���ee[��	I����+����^e��7z�v�����D�;d��H��7aE mJ�ڲ�emK�8Z��ZN��SE-Sum�ˢ��	�δ��U�W��)�]7�k$��+X���_)j����I������
�~���#�0�@*|v!��k�z�މ���\4	�>0�<KC�/�!5��~�qi'�2�`���r�mY?� ���O���n�@]����8�;ӌ7ctN�}��V|����j���Ǆ�[�}�'��G�g�����z�v	�R{���]j͡�:���(�;��N�����Mʤ&I�Z�	&�5�L��<�"����a(}�̗b��V�^� <�h<� Y�����C:>�Ƒ�7a�a��ֲq��(��W6�*)hr�P�^��X$�@G���H���Y�|m�Sϳ����T��.`����Fq�E;���,��-r	ŉ�0^��+����ڦL��p�[�������S���0��x��"}u�fp<�i�ʗ��ȱ�z]�ֹ;-��-(8��M���Ζ�p|�&���6!K�ip�:ԕ'J�Z���2�E���sK>O\5M� �)�Q��V�r{w)�օ���6NjӈOU]1*y|�W�I~���0�߃	_������WD�Y��~��{v3-�@��u�e��!܄�kz�P��V��`�j�f�ʣ�g����Dd�o�Ϊ��" �޿����qD��٨k>��[���[�%�a; <�'&����Dk$DYd�IV�s�(�}9�(kA�~ʟ���.�����i�ģ`6�����E�_�]4�)Q4�/=��4��10��+��u���,��Ьbyw8Mt�m�ZA���҅��Cf(�nV*�u ���u�F)�q�Y��Z�/�K�0˞�!���W�Gr��Mḣ>"�����諆��g�0]�:ǼK���*O��TSkD�(L��	{@6�0M���r?4�fӡ���ě��t<V����h��=>eG
���*o�!X�����������I�E��+Y*����Ue�Bor�g �~�"K(R�%#�&��¶��ڀM�=4�
k�G�֢�䣣Z�����Yܶ�@�N�&�s�'� ���3r9󗨠���ʅ���8��[�{�g��vHz ]�@Z?!B!�����ir'��;i|���n�2/P�͕>K�]�U�c�Ǜ�8����9[�n�9K�M�*oԹ�
��wl��*倁��&�H7�p�a�����Rg���b��(gC����	�mI�:dȭ��hA�H�r�i�$-�C\'z��F���j�v�NVge��Q(�*>ӫ����}��diRu�e������.���"�P�R�Le�P��ا�3Pʦ~�:���`�l9Knö1%v�.����K-�t�t醙3���x�^���7��?i@bƫ(�쵫�{^(�O˴f/6���w�N�N���;�Z��9�P����k#�f���%���������5~V K� �X׎-p�ca�D�FmfZ��vw2H"1j���+��'���}Κ|�l=3y�5���p�>)������!���Hh�Z돕����� `�~�;n�&�9pK���>0��6Z����G��"	������Ւy���\M"9�0^)?��V�{ο�������V�o1ˊ�P�cb�
���>V'\եm	��߂�6���6}��jZ%Q����+q *6`���.L�'Ė��r��	i�s��5�Ȝbd����N�C��<<�x���Ml��^�����^���#cW~vfa�u(R�/�v��1��NY�b��BKz�2<��T'���\�`19T}ٌ�/D�~��ԟ�=7�3��n�KT�P'�ʃ��N?'MJ�?|��2�_'=���~��|��YN��q�����R������gϼń��,�/"�X�
��,��ﶠ��滅�&��<��욺7<�m5C�܂�⌵����n��V;�8������z����FxR~�S��J{M��0XW]B�j�hU�wߟ����"{�1X����|���+�i!�%�fEG���mXM�t�+{��ӬQ�ĀWFJC?1/I�@MZ����>Y��b�?A��Ϗc��Ʉ�[Jj��7N���M��������G�1��� z��( �bL��~ѽZp��C�>>j�U"��I6�V��߂�%'H+[�e��p!�����4��H����+����v�պ$�͉7)¶���*!��H`���& 5�4a�P�{�����j	���L��v%�}��<�Qv�M6����, m��T_��8B'�F�=%	i�.������$�C�d؀�3G��)�^<((�2*YOˊ�������c�Q	�B&/2n���p�􊅨�C�^����v��5j%�E�P2���ɘ�����A��N�z,I棐�Z��]�i�c9h��F��J������!��������H*���9��c�yÞ��k[PHi�4zRY��\�V~$���7��>�,`@��'��r=�3
��&�:N;s�����r�5�Ȟ�d�Ux{N�L0���%��^��~*�G��ǽ�mY�� �>v7�ԕ!t��b�s�#a㮆�H�ka��0Wò������H�pD�������ì�c+Y�[��3�K�Bhg
֔r7m�2���F(M[��vc�)��N_�gA.�0|�����}D��S$yخG	�	_��&w_u-F�ݺ�AZ$Г��p��'��c�QC��Oav٬�ެ���&u��7��� ᷄bY�|y�c_��5Dv�F�q���������L �n	.I`�%)GV�C���Rrao��9|���ދ������]��W����v�-�7�j�q������S 	�N���@ZC,Ed}�2�{�}��X��(\(�[�F�2T/ً��9ek8�߰1en����	0���<a���kZ����s�Ǌ�5���4�	����R�	�B_��Ȫ F����9{A�� ��o��V ��6æ��
	.¦�f�s=����A&�c�mt���Pb>��0I��u	xG���!j��H=�L�ӎ�����������Q@z��"��"T<����KG�Ϝ�#�-s#�<DN_�uRK���V���6a�ѭ��8Y�W�u���H��S� ������b�Z}�R��L�p�i�ƽw��6�n@[�r��Y���g=~�̉ <�B8H��nP$pЂ?�_�[�N�F.h���� 7�-L�*��yij�γC5��%�6j�f�S��r�P�ss4�R*bk�Vӳt�o+`ia����`253&��t�߼.,���c`%~��JǵGH�bȤ�^'�>�_���g�	����v�w#��)A������>�f�?6��5��:@�U��H���:/y��]y?��kT�bp��y��&���g�VW�t9zh��D9�=������
��SJB"G�x�{Q;�h9|�_��
���	=�{���G�n�:�zs�H�Vؾ�<ϛ�ډ��s�"7�4�4|6}}�W%����@��0��=��ӓ���^*b��R���J����N�i��7�����<�W*��?��J>���!E������JfP/��xf:Y7��(nτI�3�����a���BZ��RBh�	�-�J�ݚ�!��:1�)��s��^C�f��)J<��_Z<�	V&�$�O�K�Dv��m��d��2ʔ̽!�C��I�\�!� ,Y&w��?����o��}ce����dRo
n�ߔ���ce!�)�W���t�s����e���y�����3y�kRs]��V���'̴��[Ra@���=v�kб]��[ji�C���v�`�L)u�@A�_�l07�{T�8����Ns?i���B�.[�����1',#��T�X*د/��J�ܲ�r�Adw����I�t���L��
8뎜Jj E�T��hh��Z�F�JFq�u�(h�;��\!d$��Q�R@�Jo��\Ą��W�Oݑ�FE(�Ak �3��璱$���_8��Ԥ��J�p��u�.�"Ѽ��u*h��9uj�f���.9�K%�It����$xY�F6�/!A�7���O�p3~R���K*#��؆E��~�s�xp���~_���68�_e_��%�bO�C�|�.Qc?�ݕ��F�s��%ˉmO/�/3�Ƹҏ	��<�!z�ˈ7̗�C;���B�K�1��ٽ'uګ� � �4?�CUD�Mk��l��z�	�I��'XAM+<���~a�|���7�����BZ��+�ͧ�F��)�٧{`d���F������Ə^υ�FQ��YL낄�L}�֑�����9�����k��wpLJY���Y,4t4܄��	�6����p�|�QvWW'{��z�W��`�n=U
Lm����]��6?�͘�@���	�y�jd�]�fp.^��&>A�;�ҷ��E�m(��td[���B5����)C�@#��-w5�N���S��Y9a_���|�>����q�B�)1u����ڛ��L�f�{�[qSbDu����%�>tA�JWG�V�dQ����IL	LS�e��*�E+�?x��c�J��=�/�M�wd�u�,i`uꍏ�=)B	g�6���ﺅ�Z`r����G~�wn3��
�֓ ����Q�}��	��w7���96*�4���;W�x��R�3���+n85�uMRnW��Q���De	���}r��x"�I��)
t���Ծp,XT�^��6X+A�\r��W������ ֜��5Z+��}����I&��s�b���2����|\��&l�i(=�/��<�tT"��p��^�U8-	�P3<p���|�<ժ����O���\V┰�;�����X�.����v*H3: Pc�!)�0+�p���IUp5�b�c��)�y"�)*(���UN7�bS�C±%;��P�4�{\f*
�hN�o���eIv��F��Z����\t,���7��.��<<�J��dke&���q�t�-h��Q��s�k���K�`�,�2N<z���>���T+���4��p7B��c���*���d���*�R�I�\��;7��na���m���.(?�䑼Q�%����:�)���.!��~���u_��1��J��!�qbJ�Qi�3����J(��3Q��`���������s�iz�����׼��#t�U�{k�#���1����z}lAh�MJD�Rh f(8l ��5��ܗWg�)@�3��o��_�� X�����r�֛Z
}���Ku�N���%�f����J&�)�
k�3cm�ȶ��5a�b��gA8�Ψ{��'�f�W�ۇu������g%`0�zF�k�ў�rQʞ��+NQ19hS�{=���_O��q�Q���5�ј���2��-s���-�:m&�T��]����1H�r?/�ڹv��="��B��:5Jd��%�R��mC��C���$�'��9�&�qn�)�{�\��0��X�������-�5�g��Ǟ���s��@��[���^L�C�-���B�5��NP������^��?['�q9�+Ttc����$�H����%��o��)����q�ɖ& �z��;�~���*/�n0qVjj4�H�\p�Ss���f�(�F4��:J�/�7R,c(zi+��&��v�Z����e&g~b�D1�]�s_$x�~>|N�q�(��g���~ԁ��D�U_"	��,���"P�d�&K�,����Ye0�:��hN�#�Vb<_��Va)���U�V���"��W޽
�������u��^��S�!����0��l5�_Ď�#�n��cEAQ��e8V4�i+�kF�zge~Xz;r�hir)��f�q8��d���6�b�?���dUˊ�K���`g���da"B%C�t6­�z�jZcits��b����T��{u3S����*��7[�'u���YS�Q�hV�+��tڞw#D-��1m�I6�/���p�X�e]K�0�S��Q�� �u��C�{^Ғr;�Q�(I�N	@�%#E<1��y�J���B��ܩ.W�ݽ�����Z(F&�J�ʇ�7Foh*k9<=A�R@<%���_Sd��L/`�uz(��a����U�+Ǝ�֐ϒ�>��!�������řr2�<�X�3���<�i�m�b��|���a�hЄ�Hcdxu���T�C����H�	�Ąz����rņ�����Q%��f�G|0��q�8��Oc��vH��|�`[V�	w���9�����l�8�ho���#�M�Z��'�G�ˢ{�Sh���1gH1�o޽��
Q��S�2]�֯�ȍ/�]o�'��.�|Гģ�\�4��Y�fz������ʯK�,���\J��W�>G�V�|�'�&k�������f�s�;y��7���c2X��{�ӀF��Ɛ'E�u�n�ߡ��T̈́�p�o7qp*]��{Yk {����J�R�O��5=��z#���6�����NZ7���	����K5.s�:=~�B�lc'��t�g6���eɲ�I�K��-ug"���0%����*1x��O8��x�z4�B�K#�v�;6�Gc�R��T��5u�'�J��x��U��9=�&�⫠�q��,�pF���B
���tF����iT[E<Bh�`�F��b��� /DQ8gt!K+���)��E�}���GGC�n�u�p��"x=)L����z�^��R��Q̓���X�:�ҊeO�|��ử� �A��ۣ�5�yTgL����Ћ����9� �:9EMH"_ eH�l����-�H5���R��|T{)��l�(ˎ5���������*\��9����T���=cNx�>fZ̦BM[1���R8�:h^f�9%�iﯣz̖����-��d��c�����i��;�U%:c��g�F��_�S���0�Ȓѕ�"�8����H#�d�\��H�W���?�Y%I���������`�cc���E����<�Z��Lj�W�fP���f����&x�ǿ�ZU�:gqY���������̟����y�'K]��W��vᵪU�����vh]߱�OB�4i�[>HͶGU�V^�Ʈ�$>Cwe�q��w�q3�B�;��\�]��)Vo�No��ȶ.��X2?�wpm�u��̀��bRD�����Jl�ɼdw|�K�Ev��"�tsl��׃��ĕ��O��z5�R��Wyw�k�(i@�̍վ��vc�+�#�7�B�1Hc�a:�/c�rؐ�ά�������ի��j�_YR�/�.g��)���Cʭ�b��I���-���<+`��޴wM���a���R�̈́X��i��%�.���tj���1�^�Y�z��r&�G4���-���ЎK�[(�.B�&m��/D��-�#f��=0��+�Md��F��~f��aM3���;�`l��Y�Zp�a.�js����JD$k�9�F"E\1~�Q��~`֣6��kuE��
{-�WW����(�x qu�r�FNX�a�%Hৈ�O���E�sSۛ��� �O4Z�3����6��1�ǂ�z�LpU�a4���`�d���G���tG6�2�5TJ/1�����a�9[%a������N�u]7v�/$����N��	�����ǟ�'��n���O�8�@�R���o�K�ÓZ~c��:K�(aT�*͓����^����zS�v���s˱�MU�$A��̪�Vx���"r�J�)��b?�k�X����I-H|3���V���ɩ����am�.�d�`,^�s��I�����x[�I*I��H�:�
FD�?Xb��jO%��	u����-B��8�$ �NPo.g��Bw��d����Xs�������]O)G�>�9U���Y��E&���t�*P8���;�a+��������ꃋ�RA���Y����x����D�ݭKȉ�T;�o�gT��Ak�ػA|\-ѯ��{�\.� �쨖�����Nܳ�WqV�>�5���N�5Q?*l�~)p@Uû����(J�n�@d\� !�5W{I?������
ݘQ<	��VBv��7�F4�F�{PE��y�]�UjU:~ࡘ)�����&h�?Q�C�Io�L*�R�Q��U��A�q=��9�@v�p���r@�J����̊:�tr:���v�Q'���Jsk֚:���'�I���,֌�����k�4�Gd(��v�Hl��A�:���2��Hu���O��#=��.��o�7��=�J�-����?���(���p�{����@��G,����Jc�]���I\7�|"������p�F0 �5��]��	��/���#�uS����Tm�����'pu>�.�O	��;Gߪ{k�\�Y�5_�n"����&'�ć���Ǩ݀L���h�I^�U���Y�&����P��G���T%!�)�ϖ��,PWM��dd
$�����_\�ʧH΂(E�vA�mM�z+�d�K� ���P�٤l�&&�`ĦB�w�@�{�Y��%Oޢg] B:oF6[���E鸃/?�M���O������-�B��+���a��$�{Z�8��m��@��f9����|i�rʤ}1�t�v(^�:�x����J�NC�N�E95!�_R�a��.<�	I�͈�a���~�$��'�槠��;�e�z��Q��~r:�э�WG��vDoRy�3Ӏ���'eS|%}7Aٻ+�b�r�	���wϪ�|��#���0���e��߰�Q�DTy�@EW��|i׊ss�Z	�X=�m���Ϻ��/ȩ��N��^T}Ȥ���7�>Q����KB�hz���s������=���d�ʫ��/��=�j��rl�J��!����kj�FQ��tXR	*�a���'ڰV̾�^8�nK��3g1ᩍq{�ۅ����22���5�3:׉򚲕;^�<a`ù9��n��%�9��9��v�K�n�*H#�ժ`�#F6��<��'k,bǼٌ%$Y�:���oN
@F]�ӳ_I�e\<�E�(�'c�7�� �����ŉ�񺊕+Ѕn�*)�9�"9�B���d@?�~p��� �;O�d�iZ1|�����Am�p4�+�W+�E�ZQ���*�� �0�N��J��G�,�v[��`0n�В<V�3��e����o�>�-p̀�(�ٱ��N���Rl��4DXD�Z7��ͅ(���N48qK�M��,�g|t��l�^d����+�ժ]*��0Ic�A#pK�BW�����8���W��W���"�n^J�F�,�<4�}����� �}_�a&������sŲ�1.��t���YE-�����&��y׼� �
�\�(	�W���Ze �B��#�$��� Q�$�OA�
ձ��<bF���#3`�Q08��!��U��*P�ט�}����UҊ�R���B�S�9V�y���Hį7:��A�*hRJI�WY�?K�l��$W�ߤ����v%BǢ�T���'[	!���#��eR�&�C�J��C�'�ܪ���`�s���T�űvnl`��*-�DA3
��-#���;���e���#���%���:y��v���"$0�������"�n���*��ė<+�Ղ��]�ڎ���9�AX�Wm7(Ueaə=|Jb�FP~�K���;�~h��<�+��򣯾e܎z?'����9�d�?�kԟm���R�o�|oK�&�_p�x��,��:[�l]pSk&��*Qg�s�F��e��:�� :<��Zv�����{d���vI k�ɱ+��Lp��
�Z��o�&n�]�.䯐��PSJd�i]Z~��9�ᯕQ#�>�C��\AB�܍��V�]ǆ��Z�q�� =�4�9f>��̇7�3p3h��;��.�8Bd��W1(�� �S��%U��}��d�����5�1&fF�?�Y����w�E�ϼ�֐�f�74�x�g[���׹.�+7"D �ponwm�ڲ�x"=E��P1�[�x�+����E|��@��Ϭ����� �A�Q�w�[G7^�h�w\��/�&&�� I��h,�ϙls�^��SL)ܤ帢�ӉD`.�y��m�� *������7�j�1�P����2Ep�U�	�2���mX�oxC#-���*.���)��?&P^�P#��K�n�Q���ă�W�?&�(&��$��'���xqӁ��	�Όe�H�����*��8�:�?��}h�@EfW��[W�O	�T�,����:��n1��	��O��a�3����bJ�n�g�����|~�76�[���/]=� �#f�:��Kaȍ0�jKI�0oF;�V���~����xJ��O�d�g�C�xB�%�=�A�n���+>��r���R�%&Ո`~ox�욒�Uf���\��^pk��(�;̼�5�1k�Qw�%"*IS�+����g}���§Bc��(a-�@@�����$�~K$}9|(����i�i��>0K�79�4�����YcPam���<:+���hѫ��}�#�9�É�$�ţ�-��߱D�#sa���]�oJ�x~NXXR��DK�<�Ku�q�S��]�L�+wpb��
o�$�gb��]<�Oոz��]s�G�{Å�!��shm����L��_��X��,џ߬��'������M� ڟB��`;:�T���)��"�'-���a}�,���=+2A�z����n�������ӜW=��c�Nr8��Q���?�#\)��#�p� �]2l�?�q����>�	�ԆJ#	Vż�8�E�TY��?W1�%R�s��|���W���vz����t�ľ�> �1Ż�x��G��*L���a9/��Ǟ���m=�^X�ێ��5�ӊ. ���#��+���ײ��J��[�����3�(����#��������'����'oԠ?(\M��h�O���Y���|~��L��4獟��6�&���$�#!l:�tB0(����QڊFح�ȑcO��
�,�ڍ�@D�QtX�Z�ZJ���|AA�����'}��a�k��c��,���i`���Du#�=	�g������ѩ�0'	ģIk�-/����A�'��PV�WK��wt6UO�Y2}���v�[�^��~9��S����5���Y��K���lL�J���YQf�=����-)��)Q|���,f�r�v���N#�Z��D[]�H·�i�h�A���+���ʎ(�f��r&M�]簙
Z)��o|d6��}Z[�"i�4��4'�ʹ:� �-��*8��;,"N|��{���ʼv�'�����S	���o8/I��`�l�'�Þ�(�> P;�F6�p~ 6�[�G�5&;�q:���z�>���r���M��[�!��zP
�聭�_ۈ�#k-�BJ)���M�^��H�4l�V��K!3Ӛ%����0C@��d:��]��J��f�O��_y�d��!�l�p���T���|��n���Tc==�M�0� �Cƭ"�ّg�7S�P�ޢtw��D�L�9�"�������V1DN0
�̩�Rl��٪����Lj�+���y��|�t����|u ��EݏU�#���4Ѣ5�U�Ӧ}����&��O�ZtN>���Qlէea�j�KIP�����6���ͅu=��}C���a�f���(r�f�x�<����3'c���c�.�2Z{}U	0��r�L����ok���pRT�.��g���_:��l�M�TW`�O��&!���gP_�
$�\L�F���sۜ(�N0��E�x�mG!�<�1(dO���U}�{g%�]�v��+�9���f�?Ǖy�Xώ���4:j]�I9g����l/b�c������QH�H�"
_�f��S��ԛ�)y�,i~ ���`V|�'9xx��2�G`?B�z�����3��O��fJ @��8����x�Qc)̣� C+[፬B�O6�#�u��_%��f�s���Nq)�׳zm	�p��e�w�:�<�ǒ���w�6�ʆ��Y8�b�,��)E�_�|n�zAh�(���=OU��6]ڰ�]��~r�}8��n@W,�2�b�_M D��iw,�R΀Q����,�}}�<�g�q'����?�H5�9���-7�(f&F�Q�}�BHJ"�X��&gVf^7=����������H��һ܂�A