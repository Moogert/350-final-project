-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
t20jniB5tjPnj4WI8pQgrY62CU7yW0hNevkAy9wCwjFwGWtMjFEX1TcyVzWDLoc4XIucJRRHCYpJ
xLTB1lTT07ydsG4nB43cKxVrGkA3K2bPNTMKb0ydGkU5wdNUDD6B9suVv1h4Gf2fPeheuGNRmcSO
tPQeYUyLMzwtcRi03BatIjWzri74ggzQYzopGfu3W/miuydex1lWrUi4TXYheGuryX+i2ciF8rqY
WEsb5wyjZxtwjlQ6bZDCV4/k2UCh8u9Bx1GbEFGSml6zNxX3zxsQgrg8LGOXeEvo3jXtQOCuhZ6w
fLC0U2zNMaRRDGo4x0zU3Z5G/V8EWxyTQgvBsQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10272)
`protect data_block
iNlD9Hd74mBNlIZvrrn38MjfzsKLH6iqXxSEYeUGzmAIqTrMNmG68v2BSUwqEoUVfg+8AOSOeb/q
KvV7nOWZ4De5pERYOWzaVkL4hSh9sBPcDEwbncuUSvCLkyNRm2Fkpx3P6mMGtKZTRRhvt37BDkZu
pc9Vhtz/zEh1gwC/mtBij2Gvvu3RUYAXRKXU6h8mJrnFgQ7rRDazzFWtd9MnsMASZjlWYew+zLYM
yvMLjh8QMlTgbqMA/RjhluqHYCEtdwHeLtUhMuVlTJp1RrdgCM6FvYNRHL6Hu7czsSgcN0u27pAv
XMs5z6GyiKbdyE6EtXtt5EhKxf4BnxQ+tsODYql6iD2l6rkL/pSwVWScc4UDm1hTZ4qaa5PyJj5N
RFa/TUN1PPjEjZIsoRi/A8skrxdZL9s4kXyf/PPGQZz9xdXGGxgNOhywbrmu8jjz5uguMsGpOoX1
I/4n/dxnpuXKMZpo88JjFed6FSqrRnJTFG0IFtLa23g+D/cv/DDJy1ma8oz29V7tVfUAphx7FxOl
cjtSHVJFfQg0487nFNBPMHeaTZLcLhScI/H215X6e64zijmNH/tbrmRzMmxQfS4bvVeF7+MNAHLf
76BuzDIDzXs+U1rAYF/8xcfhEjPJur6QmduWWmFh0AdoSvR5cXIoh17VxDFIVM2H9R5MulQ9zBe+
7VQxh+YNjsRqXjxqwn33o0DMrw/6bjkqH+x65q6kYbZSqsYi6EOFhkXyc5HvpAa1gp/k0yEElnOg
8UmmG8E6Ta6M8Puv9gtHPN0RAX894G904vQ1FQHGgldtXDet9VlxWRyS4dYwVrmDav5+r0YSSKZH
TbTRBHrgSdzWSRvJuT6HeBWPFe+ro8VN1Ge6Pa0oF8mWUw0gxapKTZ+VT3o1d+jdXZz3+LHt+dBU
lkOgAKJkiFCwZ3grOam46iNrITLVgkq0vqqDPsm5qxhiJgeg/SDOaSa7ENUZDykb5Ous+D2MyilL
WjOO9NTKnrG5aN8Ehkb2OmIGl3HjgieH5IyjbCzg3C+pZCxIFqyITGrfA9uDPX5so+7KoSIaU9Wc
CGDoIK+diK4/R73EsZjQrnebkZoh6eOEv/3Al6QLYgYuuMHEragINQe2lEfmOyqLqh4RYfW5x+dM
j42ecX1NfJfQRWBJ/v6qzj727GfetB+wgfbAUGR/ArBmpJlUrcaYtIUADGs4S+ufnOHZRngLqT5P
9gbLrN2JIO1f+TuHEdce95AgRk/iT1BZ7lhOwpEdYSSeQMxYGdQE/Xkd1v3ORABynFQRC7qI3YvZ
UmUFzSJBAh92FkVG+UAgNKEN8B9ANaSrIgYk3SLAO9sK6+mAPys5Jxk3BWFIGNW+qOFhGvpdIvBu
Q34WgIan1w7c3oftEpnWrXyPjHUHOmkW2UmijMg4jTUaq/SglnZY9WV8OT+0cTIrx0o8aW7kGaxx
GiwCRuJeeH8MKbbiK8MhpchMEWTmiIWXFLw5U/sj/dIg+xIBOIwFoU8R2FxJdpYChxjj03rurnpp
Vp+kBwrDboRSoqJAt2IeU2v+FW49bd5HB+gMkio73bGN/Juq15Hf58Fxw/cmefc+Mb87mGHuB/l/
xhPYXjsWCgph4L3ncXONTtBwimtZyw6eIWJaavsiTDdPbH8NCm2wEKnbYNN+qxOF4DPr35rwCFcy
40HMCXEr/7yMFuUrG9aV5a6NJCGHjsZbpvSPNk2oKZAry/S3yrB3hV92FEzMb1VLcBUsXBBxXCM1
TTefl0r1K1dNPno2iDqMuVpbmRfH0KQvrz8y8tOIiHlCox+FLRcAt8Wn0lOGmD9YlsB7bE/LADVG
bzjCB1si1Ko3U46RwR2qnT6WDNEqYLGmKPbpM/oL6yee7Uot31PZLuPSpyBKeccIycmkbSEuRUz9
kBlBoodvBzT4cJtbsH/XH5Kuuv6400+CXiMvyg9O1GrWyyzdu/El3OcZSBk9a44JE3OAQrPMBUGt
/zmUr/gNp61v49IkDRC6dWgI9hOW/tySjSHpdVPtMkyoXhJFLHDWzrFO5ZsnkoNgcwsryOopXXpO
4+2JxJydWL3aUSv/rY1JP7neyJ9VKnwuOa9bcczwBliSJR+5c9qrtFt64UKFJas38xax5dV7DiNG
fl/9SjR9ciL+TT/WmPHfRpDNVbzOI2+0w5V/EsPD6a74sPBbhpR8YM6a7V5Od60sBTOXTnNiyuAw
vBodOrq81AiBz4/ajtJKkHvwwZg0LpHjM7BCpxISgF6MOqokni7omXi1EdYZ3KrULt6AHJcxF4EZ
xyIK1tOAaUP/k43rYhICUZYBagF0z/aaoL0Mk9ylpaWvQwYMm6ZUftBM7pU8rXp1XcEI/xi7xz1r
mdrYEmZv3v1vqZg8zFI+IUXJXuANuZQ6fuwk0WP2hK9BiB8rqvq2vKOLzFI6goyKuTx+MVX6KXDp
M4w7H8T2CDXIIYpxiksOWj7HxbgMpCaaeRMbZEZENFBbiYCZV3a7cEKquhys6TOrk4U6HXKDM+3f
DuBcIwFzgUvjsUQLwYVLXG02vnbKIyfueX8JGaQR4WjC1mlP6FL8lj+j/GbknkmW/m7aoQ+snz2Q
BqpxRu7vRS7Ta2O2so8ZGhJagZUd/R3J/AJBn9KRfJHH0no177BPdrSCnb+FUBNwFKUywaPPwcjA
ZLpHTbXgW00Es3u1HGBjQDd7ltB3euXRHtzyosjOp1+jbDgTVyXoq7aVRnV5Ne03DKQv17iLrXPt
V4wBfNni/m69+p3zluNKCWAB+rCZiZrqKyXCCQmePkBtgVQtKBqiXLWOk10KCR1D54/wJsh4zR2R
eWFhVQq8iI7iexUysBr6q2h/31cGu5WadFWetkeOsFj+Puw4AozUZHImhmUAAYoZ5tt/CsZD3Pcn
31qqGFwlzcCJMF9oGKIGmyCkq+5MpVsmJUHxZrSlZxZnel3nMnL76uiN/dv0XPQP43ToPN5I0jb2
STrHOH9AwSeXQm1Iwj43KYnePkwsQkFClb+YO2GpLpd33iZRSBjN6dS8PjXwQLzKEGd0UNmlopmw
glpU4xJkQCTuMkdchNjiTQpiLIuDBG+Vk5K+r+fehT6P1TkJocpxKCzvGQ8h67i2WidRVM8rM+Cm
vJql93DdjTXSwCkmySx6KV1ItuCMAdRfEsTj6HLJjw8SHBmbsdfMDrnIiqA2xQWvaMl6AcLa3yck
CYt3wtmrSks1I2PEhHWKUMliG6EzL0Lf6TolUOLw4rowv98m1vgflSE6aVYamsfiWu1AuSRJdR/w
9hjaqsnkEU3wNY2PF82RS/CWVmt1HXyyMeUfw9w2kTO37RYBXz1HBiesLBfhBES0WFPL/mYkBn3D
95mCwaTnWK2ck16vUuZrQp3b5Lw1nzSmrDx7qqWaEGra7wG5SbluBlIBZ6EMQRB6M2YD9QqeUpla
QO/7OwU3BUVY8amcMA5TSEdxLiUNggaf3JlHDi8TM4ROQEh+vZtrXEEwz4lzsc+S3jUyvsxN+P+/
SiBqRcqOj1nYNMPCgXvDZzC4eU2DKbqEkaQ/V1O8qYd5a5To0bfNgSILA55y7M6feIKkZFk90Zvy
qqI/cnomnqnUZhyjvoWM7XSsDRFk1+ooZiZb5lP5yibWdEUhQMGn3qfxdU8W3aWIVBrxsUHxUt3n
k7V14mSULn3VIqUJ7tyJFEb/9sIS6pHFABcM4YfDJJjYJGbUN4h+Mjp8M+OAG6adP6Ub37Ow2TAq
IpW9x/O0/A3XPd2R40MeU5KnppTAXXJQm22HSH8JaMtgru48QCnU9X4ULJYE3uzIOq2NboUZE+Ak
3w2+gjaDcIWAGdmok2fU8pkEF1e/xsET+0UDyXq5c7SHTRzgoiQESeyO+rR5K4shOaPpvr2fHvRy
ZkDl30fjVrFthr07Gu2ANDczTVTCP6mtFPPACnwI2bUycZqmjTzTtNbLbsiUKfPIiOrhHmfZmaLI
qwATJomC2qfIKa+evt6/tW6BR4IsCTo4517DudPLO8esbvfooGbsBw+WhU8cxlk9ooKXh6Q992C/
Te+mzogULbeDvBh6kvmFLyAOEEpc1mAP/HxEFrbgLHg6kCndoOP+SnbiGaiUYXJMZ7nrc5FX9Ito
sqsYL/FVzVlavAAJIk6XmW6HtN5q3UiO6ZLSLfQoHtd6VHmdcZNJ8ARcVAJPceNqqpdd7Y+aGdR+
oXdiO1iWeQi8JsSMr3aayzgnqGTl5ZyX04AXh5fyNs4jx93HCB9ApT4/fAwLEh7ewCT5a/5/zDA1
7TJ6wFkVC4agJhYTXXr7P0EaoDmwuurTVF2PDoeN5o4MdEx0CsBRkjJ8lz9vWdGO7OP/19yopG5T
xjSaJnRj2Rm7qM9pW8dBN62McVNNMqDSOcmpxngc3G66j9pU4IsybixEbJZwR1kcFMd9k4x9Cuva
+DCvJbFizRaFqcAiGE2s/0pkacoInFRLhjtwpOAtiP6IthyaWp0B77s96s/4BoauhfSeqI8JofTK
yQPHJtauV7TEF4A/M2vu+FJm0raYtJE+NaID/x1TiUh39D/cNXLz8Y9IBt4owvGLZpzjSStjUjKU
s9y29JneqMCSjS81kWmtnfStPwjZvsGkTA6xuzlnSGVpO+A6nEF+ibYTWBzrTAO9A+HsOVjik21Q
/hSvzFpkFGtOlQmeZ+jdtM1ipcvfdoVePr2SmMdfLUOC+sCKHnfHcWBLCSGh8ftqzhp/eYhdkxSr
ZoXTvAA1TPeecMx+rV0KR/Q8a6V1PdbUYRBS39E9S4NcESmA1qzcAtMVsPbAXJ3aurtWE90JZTvl
JMDxHcjISo8taMWS15ltqOZz5RSYIj4+CXo8biIsYuxhGcNPMj3wDpg+3OI99a49S/YJs1glwY/O
H+5pWcbY6uwO55W/JNRTEknFH06Q/pSOpan6NC0zCZu5UPUnRBLKIohPO9RjZDimrsnhclrlqaZF
Cu+8VXDNJ2ikVZoStsM6QLIb6N73Fwh9PlysJxtA0GEaL78nO/A/Y3cYS0C6Wk17Qvqbv32ljeMy
hczPJEX2zx3Fyl6p/t79GDw/if69/zpey8ox1ne4ahtd+eMhGz0uCQmch3+hVklu0btaHnWMEWlh
V53AlKfqT8FUpzy8NWa4YrF1Hrt0iLXsMTOuHjpC0Nau2ksSqQIj486VPS146M67M5SL86PzBMp5
rCQY1VE4xyRpZYK1DNxZGAJXqi8Mj077k29rt5e5lzAus/zNd1DAqdKM7nfjb4NZWrUjORSWK4NY
bTwRr9Zw8OTwLnHcMH0z7wUL4F/CyWTZVuLjUD1aSY2lxoSxJCC7ZxJDlojaG9DVIm4nYrGr96qw
3wMOZIbxB3PyzaE9QE7JgmP+m1v/jfMylO2ZeAU1JpT2hgwOYput/n/kCCswUjN2Vc8ZzIyyFMxi
m0cEcUrEE4ZXFEBH1cBFLa3GYUkcnGSHGWfkSHfagclddXgTNxTUy/884UTZnwtarAR0Lbt/QouI
1lpaIEAe0+8p/SyWyhtMMf9terI2yHmku1l2a2gEnDbQSUdB3z6CgZuLjUOtWwvYDHrZmzIm3H62
gVLDO7KLm4H3zu+GvRdTnAwZIo7UW2otAWs/OlougKtLXfPHZYkU2tEhhXwcHU3nv/5znWeo5DA4
sV/mFjyPzfklw79Y9px3v2CHpP1kYsr8p0QPrGPCpXmcqCmX0PfboDwWe9A8vYYb33h6sQp1uFyY
UmZhp3Y9IpVnGW+TqlAi0ZxnuefzNiEL/8CDmmdrPERuAGaaOMfduwp3oSb1fmBpYeC3Wg0gtoa3
zVmhT+LnGQQJjFQThnitFuKyobGwQdIthsNxlQOvt7ZTdg4IgJLBFeUppjH25ETJgicDVUdo8aI8
7jl67FXtDcYhRjnuyvmRohBWYy9JyGar/uNEF+yZQ+6b2qZd3aVmLtp6ej2kDQZ2IGvbRNYkaPOn
lVmB07isYGQx73PQsGEocNCMv64Q1i1jgeubx1wNGaavHC1IPxmvxJWpPJDsgnS4nJXOZhaFnl9S
LEbuecmohw6hCDQZGRnM2IvEbCAhMgdWo9kPST+XOrxNh+2gQwbqNvttlb88J/b8mHQvZaPX6KYa
RCu3vTrxE0FqLmP6y15+4bxAS+6MxK+YbdRs23f/buBi8Qc+8wUMvUTBZ6izKF1t2D+WL25MVGcK
ouAQIP0FrWCevQba24035XT6cSXLfwEJOHZL5m57SHpHv9Rr7VgCBs69M89+tqjBWFIuIZFGAThL
/LtZRAFGLLpqwuifv6m5hk8GXFdub9bk8mNKb16l6W5nAycXAq9mHrKzKi3c7xGRK3wBukz6iJKS
eHAkFJ7psqoxU150UAFJGQCS9ZmfjLyTlgzorMVWUYwlYsVMFbbzRWxDzR8Cn0X2uY6fMoEUxgpn
uM4AtkII0u8PkqJzD1jXL3ALK1uBJ6Qu+1oVjZBdY1bhKcrzCnkyLjFEeaPEfNd2QvvnrUqsIjuI
XV/wU2vMi3/HjPQiaI0DLjCZKcOeFm0Fkb6ZWZXH1nshOhxa/Wh0+NKsefy5Yncb+sod2vNJ53aP
TtOjV6704TUI9fCnYCHkH2v6fSkvzxZBy9Ut98+Ebm1Ttpjmal6qcbiffILDhmm0EtqAFOzIHR6O
rScL1rxQ3O8s+Kfw2d61+3A8Gw2rMV9lZb6wFm9ENGfCh1FhwnF/vLtafqpglcXe76NxqzdcVSYh
5wmRZVSQsp6OTahW2PTgGMMGVsP9g2cLaRjQE+5wmlmBo51l3mEhpHtp08p8/rSgcySxiW5XltQS
lMJdhrksdLUPnkAveyrvX3WRD1RGvPVf1BC1LE4oJmPxpguxXgryRzicEHPlM9eWC953syoQ+nyn
KaJ4z2OYRqZG01/qbts4ddA+uldTYCUEAr8vR1OUdHo9gDDtFJK8z4uzFadw/GprMW8qvKBUV1O0
oYEUd+wRiiCXuWuJM7ag7epoJHWXpaZYbhxZ7h88g14vivDulGLc+aTfIN5jTF/taZUD68spmv6D
CQ7Tjs59+3sQ9nZAP00K3ELdVV2Aw3I8/zb7QJbHxiQFo3SrmoHJXOxdDZ2qk/bYgQFNngyc5KS9
VS1stIMWTm/4DOvFP1iyGk95cq/bYMlZmujiWoD/Ox3hABM1vwdwESnY7JnNeQ8/LSmg5Bge4cfw
8pdaXqB75ehdweXqNkL6ibZ8moY/VxUgjWNR6gbxrYz7K2xs30KOyyQCPS6HryCriTUZE+fuHWBD
tf5eVvSIORfyZhgi4gdzxn+hwLjFwIF7CGgpQSsv7B+KL81e5c7usg8Wya8AVXM+rMQxLwy0gyyE
PD5NKNuEw/EOGaXmOGHUu1PKmHMsIC+iRlZwY3U5S1OWWO9dy5o/OqUwDZ97xN6iMaAKBRzqrTIs
HjtDzL5hdYGGcYSUSXqvGiY/kYZFU8keApC1KTAVP8/AfqPDaOsSUhbaOgOs1iNqAnnUWavTHJn7
HTDjOmL00TZaqnXViWytcD+cXczcixtn6nEPUJGtyQuIlcvUlQfAii7LPZYcewtOrusEQ6N3scx+
d/UJuY5g5IqrFsQLqjiuJC+jNNjCodmc5a9hIxixdgkOntrtj7/fTru+glhrDAW/Ti8L01iHNVMz
0Cl5frwHi0qmt9tBfI/MWls1f6oeYGy1R1gxq0coD6S5i/6aTHYUgrJzMKFDNpTMtsA1eJFjDfow
F353uPEge9i+6kjQKvxZKAuvqrtHSNdxKzsN1Mwx5dw86nJL3pPEb6TYmysH7xoqRAkM0KTcI/aE
21T2W+8Tfmv/zkAXBLS8JQ9niSDhXpvvx2LzhuodquBkEsdTfzTMEnlWgIMY6xSAe7w/aZlbuZTF
kzFi9Y3UvZZA/Wm4SJ/w2thGte3zfJM8nq+sWH3RlsytopG592FUfilM94BXhZNRVSfttxIHga/q
WHpVbW/9eno0zNBC7iIVbU+Cgx5ptaHpic5osh950YsXi7vSvjE1E6f1G1Mnd6UOeph71vJs0xa+
aSBqiMmdcI4Kq5SiUdMDLvmaPpgLiMMK4EmcaKplvNinSBSmYn6QOy8Z5c/0xVkW1qnOUFATiwZt
qi/8YlfMjhgFWgwm2msuh95ihHeO6X28jTKNupEC69mkZZhUeWD2d+q3gGW6UBZ4lgH5sesyfiLb
A/UQo3NY1mm0ZTMW5J2EkjGU/vyFO+u+lqzR7/DgYNHBjORmKQGQcpwUq/xmqMuypAp16PvOJxeZ
a04bpBlWMMMPy9kmabSG/W/NvyAFbi1XusS0kjC+00KiCt49Exam0EJXt15ZlgFVKNFg4GYi7BiB
mEoseacODR5ikGxc2lzmSfHlx4nLrOxnT6u399GzY1mXS6MFuyZA+W9EF7fMYizMxY9lZvxo8+ra
ExiZlOU0Wqn7gndTd1omSYu6x141jUYzAxw4VhvRkjYYQQsA6DqiGbKxi+orChwudAZ3uckZDrlp
7SegUo9IWKimzecuzFwj8e/vA/GExejVppMo1unN4bPfvrUJ6NZpRcgK2jdArRAzzA6SG4xuzSrb
APxe6xB81cY1lGZ3E2dMxLD7HfybUi7CbrA7Zhpiz2U6KrwHva0LSe+QNmhsNgO2HRSF+rHxB0fz
9yjn3pMxRkBDywf3kGDHD5licyIYx6nBNOwY9KA9XVDBu8kGXsXqcdHMkarfht73G4SL0EPJsd54
eQn/cWPulfSG6sIgJZ7kupmOPqeWaNk35jr9mUs7NCNdBhei6zcrof/vprP+5tIfL9IMViDQ3A3i
xLXPc1B6Omw43VgfvS0zTDpukINH+zJC77ZUCkvb4fPeuJlIgvAlvt+roGvzAWUgAIARSb9iWvI6
1QRESfbZ71HOyfJBvYaVblK3QhP27fa9WmbjYaPsn1ipi/9mD1qlf9FR+/Lvlksl10wim5eSnGTf
HdBTkeujzE/ckYyd1cQHmI0/UXIFLNjux2qPK2H2kjNDWJK2E3Pd0tnz8U5ifQFHkUyDvCNRRVm8
sjnDd105AB7q02teBm4MMT6GPhaK9IdhW9Bxt5KslCliF0FDxz0QWMsaxiTFxekDxsvPq7zJIgwp
eIElrvdrEUcS923ozNyOcq5AiBExUmcb60d6P3yVJN/oNceZ8q2ZFlajAUYyrPPDRrIRnKHa3ESn
TJJFIMxSO7xNIfz3Fr51LO5CfgCnU1vZk7GC63bvGXzL/EhJW7/3Q9tq6Php7SxCHGBTKchUwnA9
GlqQ70aCfTrsH39y2/py+GP94glEt/E+9GegxGwEh4sczQIYMLD5cGMV6NVTQsbJtXXWZUJP+rAF
i8lrxAlvzK5IEoab2dNyD4PSjzbjn2XuPTXWh8Tl9kTg+WJeFnuXd0WAA2IYB8qFi+tGpt7g96V1
x8bmEDhlZtiHk/afMgkqQCOLezXjGo5sQXHhCtgCbOPjx0ZNIGJAuQOlIqGOqONWRBSiPZFy6tdH
rSu5EPmnTT8G52kcpzEsaxdrFGVS+TbkhkVuItbyhvX1RzOaMTk3HDSvk94uNB6KNG7Yd/WXzrrV
fgnofGJbyJtyrYEjsQlSoU87mv8P6+aTe7remGiDZv0CWmMeqfsvINAncSsRSJLT2oPjEQ8kK0J8
/dNnQqPixAhX/pnE1pe63Bo0bTcIs24X1ozriKqK5bGsEqyN5ISZLFmLU4yiEV8qtqAAiVC/Ct27
ccHO1ZAI2D2TN7hxeeDjD41q8gy8jJSkfe/qbUK7H/fFPJ5pf18m1wQdouvCLsUG5KEVaowlQW95
PYkzBD0IDZ08TW2tpx7z10E9xbPM6W0kY2kOxxmYWtsOvagN+c+0evB63OOMNLiOLcuia3T8XG3w
K9zY0kDtaq+5ujn2r7w4zx7MqEC+f33zswwxFKcN8PjA7xnV81Jfbo6lJPKxbNyIeBnb1LzPB0fH
WJWpQWKvBG4jWGOFo6WV8bEAz6H+N1S5CFYvTNMvl6PQvx1NOyE5aDoWsIU4aroT6z9S/fv4I3kL
Sp492BXezic4K6g6u0dGrjT0aU/h08N8DdhgWOSC6DCuWqSw9PF8zvsi++CpWX4u3MFFRGQq15kd
8elq+9Iik/4G0ls4X4Xch5ijLPNduEKPcr9zneVa8Uxnj2Z8jU/oYJIqQLpB8ONK2TOfuhAa99Tx
u7lfYP8e381hpr9BE/wCjgEpd1pQ02Lx048NUEVkTmAnGzI0CGk/FfbnoMs9bj/IRCPDwZdlccre
Uh4KqaO3B6UEuSJWKsI6EZQ5s4F1kR4dOZvqr4UVOW8vamLiZpUKDucc96KxlS1tuh+13o9695gC
vaxJlggHb7JUVLnfEXeblk+0b0XMbOGcswyaY5GsQe2h3x2nhupwRchhTKTUcAvnXMLZaEXbsFjs
16E7S0h/7Q/ccdLqk/PEkfwIT7L9sHIu2zsA/qrU7t/pI8KhN83GSr6TgBdNPxd0iafcl7+AgvOC
Y797ZPjg3Leea8yPQ5NdXGzRfhJSaWaki6k06yY930sVNQV1Uyym/x25TArUnJS97ferRLskWkA+
eeJqx8YunOg/UuwNDAXzyqeuxcwvv06fyaY18CuHsnItp20R8M6x0Lr8Dv4d0BpKVJx6gkUA+hP/
b/ZUu0Y9QV3RzDPiS/yieQcfdREBVgbs/hHu1cJEw95VDqQywqDuxJ7HGv7M/thnaLklTXj+bEZa
PBECS8OJYYAy72EvS90Lawch47cLGmAWq53OSJFN5n5FU5aNHy1SU7rGDaNuBfUH/LZR/+CvMS8p
05S/sJ/ubPyT9pj9kRZn/VWHdZCR5S1cue3e7+5jim1ZV753FvtPA2ZxBTiq7yyiiAI5hIABmIKf
USdOp1mkWg9qVLokrn9q/KshzZLXY7HScn36onX15Ng1hFICCUgYDd3EgRr1r4O5+X1PtVaume1W
BI9r4Sh3LO742Fp2Sojdh8s7q2kbZNvIQ39BBQP13RUQ4Rt5rtPhIFz32AE8jOW1Ngrb6GFtne5e
PSeEaGp987OBgG0YhHJ3iS6xCjMZHED1VTk86ot9JZ5xFgIhi1ZLfYKbO6hPSEt6nXYnwLNL2XXE
wWoDu7vp6BKnG4BMGRnFZUjqppZFMv4hR5eRx+bEYPJcbG+TeO4jAAuWrerW9/MMw0S3UToudOqm
87y8UulQpcvIm5KA3DYMPDso8nftPAtie9MeFpcsOKMJ0MPR1PpDzXZqOQRGyKYu4yF8BVlvPFj9
mPfycYecXSLku8TrHUR7aZ/YyVz+d2iYrYw8wk/MKqTAdIStmYuFer2Bn1XU/C+d3WepzHtrOX1P
zJmj2vBZ1VWNE5kuXYYQb55+/D75aZp0id65X+4JArdiOU/XMrf8odVHac3666jDIw+vmj+iHkQN
2+9eyi+mWLv78JFOTeY9ih5g8/tsEKAsT41H35sXgtYOvDDFBynY3Z+QTafmJaxY5WHL0SJmL+Gr
1X5sEMYUQkdIwYXVW15j9jWjysErnSdmvghwuM4BrzWIfV4ColoIOknTOhsnPcDFR+48oz5MYDCy
AyKkFdOqKQHLQfU+ykZBuN+q7Ti+MzSN/+x+2ESzuiQo/GQUZ75S/ieP062IAFHvqGEu+ylioguK
G4n7ghE4KVnKJWf2b4s1vvoYYFqs84Wwzxyk2DmngXElc1jODKy/pcDX9+YY1wfeIRA6SHcygvNB
Kl/3ESuMgpMQqs0VyJsWmA7ncGTNx/oyWzpcnGxeUKpBXP2AMixhi84LD7mq7EyD+/Sv0zZe024U
jWMvy7MSLq+b9c7h626TCqI5QJIpGFjbGqk07bzEcXJxjqQJQh9Ins0wqpv5l92k6dIbjRS22w1k
qa+UOKCmEhx69XEPsBDcPm+W7RxzcTNBWMynywsZU7a+q90s1xNOV2KRiWLVnRJ509ZUeLQd1mkw
+LagdB4hq/1C4Lf8cx4kwhEJS9eD0ldrL52CZVlr27rnfcZjnsiaIujv/lq/EX+otG0LQAx5eo8s
Fuf93F69ry5et0vsCTm4/gaJp1eeu6hFwL75YEttCdggFgPvmDNpBB80bm89nJvOK9eDG7SmkbzI
QkUxqA/YVH4D2pHPMBCDIea0nC4emSIDQClF9ROqXqNmMLwiM2Icc9bc71u1S9pcKCk2OMVEJZZw
XZ924wfqGoEUGTytLqQq8QiaBZ1dUXPnDw/H06leYkjqOUS7t11e1W/I3tTOrUnm47P5EV39q7hC
2+B+Q9lsFLYW/f46wLcQ+DshEPMqq80uGQmUcxuO8XYrJM0A8BkqLKb8uMweJYOB5Il4AckPnqOE
8paUfQHTbRXKZ4PFEeJP4+QunPnfhdGhMq4xrKP6w+1aKpZYejl+qKmQZEUYAPpjkVBT7IYvqSHx
9OFLfp5pFyuRldoBgPT+6SZ+EzkV2sRbfvkOqP0SVmlhuxaLdkvDOSLGwhxbMcqRMs9NvMdeUOIa
J900xyz+KiUrqAxE5hqnPl0q3FV3v2xp+RbaS5rB9OVKKA0gZBS6Yy/ezvU/1SLo3dRX3djuDpVo
oiTaedNOML0QmL2VQWnIp4JNACJgt6Tivzq8PxbwFNA3EogGZ1ldrYgnp6p/HXaMa+yPVt+UTWbA
4AUDcVcJ7zk9fwqFyrqc7Vtggae27o9n3yenlcVmdMW17f3lXYBYHdqBk8h7xTMpySwYwLjOBK3j
oxMK1RtSNZaEHt1wyfOWrB6em0hH18W3c6El2dKBHGT7oy2McbQahVOnTIldqoXBcBzIhPb83wTg
mLMDwqUX10o92yHF8pFfUER2ASw9O13JOXCkJbWuMNv2MkzhoTNZig9j9KMiuwt5SHLTSe61PKDc
S6eLggUh4IutdvNrpI+CgbLQSlQrNgJ9eAUJ+MqlkxoZlehkJ2DCEW0Pv0xi+PakTmLfGDfQPHLt
NqcuiM/cvM0XUBEgtq8vuQ52xJxxEFmg6AGgLDLFVOysWQ0X0L16pL8lnV3TvPnnZiyCDGo2gPrX
gYE9d9MWiDNGZLJ3FQMJbV+zIGW0krx1md23OpkTInwB51Fs+M/0I0X/lgBr7sG0YfUCqYNTSeUK
fnvlOuCFrFS3h4abmzs1rLGDpqQXBh25DXnMKXSQzVSdfHlkaVs54Jz1eqJLSD1vS9wUZV+BDYU+
ws0KFOgLKT1rkbPfHrlkJHFBeVqxZYwFTuMwRdrTLuDRXw8E1uHhWvfg3ZXIl5LB/GOYo/q7MxBN
zkZR8pVC4rELB+nkWKbu0ql1yngzJeZCSuK8NI/ptb2ynN5nnuyGyzdeuclWv0L60IPVWiwZOHno
CvPuPhKEODrqczN7qpnY/L1oj54F0fW/VzqMSypLPsNIe57B/ctDbyQEY5zqi595tYaxfYT+mEMS
C/62tZpPGcRL4nxnFLrpaIP7rBAMSrT81wLd+r92pwYgPnyeZgcsLNjs711pL9zmZ2Txa/y/T13K
z9TrtYXzEvki3jSThXa7TdkKiTUdK2d7jqPVGHALFp2W3aUzjATlH6WJYeibOZA7Uprwmxc/9FGi
0JFlsjSJy4H3DFps/22gkPaEk8IBC6rB9E5U1V/8/KIbPEdznaw8jqZ6d8dY8GxmuFav7F31WjH9
CE8vF8+eICFqdshPi+goQ5nbD5a5uHvALhgAZP5JuxWdl/a8ioMtwOrBTfqgKvqlFJEFbnOusiOG
93beoXpBvC8KwzvNzS6sghyuLJmPcYbigh6i9DVyNWnrpxp/1rv4NZb1p8KrebOxN7zR0zk/Dqf8
RtJWd2O14coyRas/
`protect end_protected
