��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g�҃�f	��m�T���ƌ��"�C#~������VMb#�X�f�����|b���e���rQs��~����2����؋��&���K��٣�M�*�h��9�1��̻����d5!`�S�o����@Η�I�]���<N�����%F����0�8k<��~$��~!~��dV�Tm���s�@����Zl�U|{G�-?ҡ�(�K�ll9:߷dW��'!��ܗ��W��w�#W�q��ܬ���ݓ��Qy(%8jZ��{5�k.X*g���zۿ�@��S�k�!��������e;�����l9�&�V�����(�0mJo"PE���N��G-��,��4�y��]���]!��,��p�O�_��)�����`#��b*gxx�����x�[��Y�I������4��J^P�������X;�k���Q�Y��_7�O]>o,��(#�I4$I�$�@�~�Q_��C@e���k�ߡ���ܲ
k~K?�I1sUBmv\|��S��R�p�!ヘ��y�W�*�3�笺�2��!��!�^W֭�����������u�p�LF�#l��i��yT0�{��LN��3���6]��~��z�	�zJ<�2��τR��6��p�h���Y���W���ԲzɥFݔ.`R�̲��̆s��A*�A7�&�D`����*�7.B��C��~ M
��7��[X=�~F�3��p��Ao���T�B�P�#P@��`�^œ5�PB�3��s{g�T��	�U�ur�t9�;KHu��o<umi�xl��&;8�=4߮�������M�P<$<��VK���ш��=s:�`��'��d�0[r�v�Eo0e�'�*�V"��CM�ķ�k�5+�|�q�5g˙�/�f��IT ��� &9��]��O��җG�'1��Pݞ?�E�_����6�W���ݏ���~��B].�@���el��d�|�Op�� p�ٽ�ن�����~rp�)r�U`1�
��A����2im�Z#o�f!�涖�^��U5(s剋c�9�A_s�$�#+���m�������/�H��jL)���w�m���C��(���X1.B�Wؐi��;v5g���aŸ�ZE��)S�(|3IG��Zп�p�����bc%F�bX��F��a�5�J҂��8���o�dL)������д	�c�,�!>�qB�R=��4��s:�R��-@��(�?v�Iϥ� n@�ʅA����(z��$g�/�ğ:�P�&����TzZ��(\�W%B�����0o�H8�(W�gsav3����fg��]�Zޥ��gݤ]k������?"bQ4�3�A����e��	�ieՎ]!�E?/�H�MjI x�L| ǅ"ʬY��Gh����j,�v�M/�%\�>�k����֯[��&/�2�>�C��9� C�H�F�x^�ko�@�CòT�o��f���k�\�Ċ�Vp��L���Y�d��3Z�؝�ze�do�]Y����� F{~���>p8�9_�.-����_7�Cfh�0VS�*��_�!��˪�:Zw���#K���}t �^�xT��N��O�O��c�܊������_yE���jڮ�E°��L��\}��&�zcq����K
0�Li]�wU�dJG3�����\^T\%�,��*�u1�4W�g'�2l�4��T�R��%?�`��>J}�C3E�v2�VE�*�0��F���_]�:�=V��J��vC��HNwI��j��U@]?��-%���(tshi��D�WLm	_	p/�A�uX��k�8K��v���|-ꯒj�����i����s8e��|n��p����#eZ�RL�\Ѣ�B�`O��;%_GvB�F���X�'0�Ӝ�r�94(�Ź�1���y��a*�-O�3.�%��T���6F�
>���=����>��L�s%���|D�O�Ojy)���$��I�g�3.-�����8[aFunTh8�>ܶ���om��W=eqL[Cm�a�%�����F�]x��3��W�"m�����ƜnT�||S<�E�Sz�Y/ԝaAZ�8�gf>�}��V<
�����>%�6{�x�N���M<����ZW��ׅt�I�3��<mf_fa))�U�Y�'y��>)�-mW
8F�Gӯ�����Oˊ��������1���AG�h����Ka�!���}W�1V]�$�Oʧ̠��C���������W���9�gv�+���Ę4{��@> E��n�lg*R�D�Ɯ�$�l����b{��jb��4O�<�P�r�:�J�n�p��5�嚔�;k�>�a�ݳ�s��u�p�;��-��3R�ʥ-�X�8�"wi9g����Ǚ�	��T{K�nb��i����ݐ�
�<��)*�l s[ds_ϩ�RCf�ā�H�t��ܺ�2aNq5X����~S^�4G��c*�U8�z��NQM��1�f)$�0�P��(��z�ނ�d�Q�W�ߢ�Hq�~s�f?��92��o�$M�'�r��V���P���:\�q�ށL�X~S��Z��4��(��k����Fʋ���6��g�[��q�7���P���d�l\H�(��4���~�T�i���R�GK�˖���������t��;�z�5����%�qO�i,�w=/ɔ�p]Y��$��/�h�Q$�J�~-���!�ri��O��{��n�G|� N��f��$��*^��B�~�*�3XyWhE�gj]X}d07K�]m�*qZa�(�,q\����P:M*0(
�����6�P�B"�5R-�����x|f`gv��j���-��!�o���a�x�U)�Ŧ���g�e�`kCP�g�I���-%��?��Ya �v�v;�j�n�q��N{�wHJ�ٜ�7�?E
`c �;��zs����%�I�q�T��� ��꨻��x����y��?���d^}a�M��*��G�mH�L�nќ)�Kb/Ϙ�Kn��p�ݯKn�T�����<aI��٭�:K���i7�]؃�Ƒ�rhD+E\M`ى��# �x���
�<*��RS|&��K�� P8�Y�Y9����h�SL-�S�bCZ)B�O�iz��\`�e�ח-&epI��&�_��kR�q+#����^z���*�pl�R��g��L��G��5�7_5�g��j�KQ�x����0�!��U$��T�!V��6CP�4�-���}$�Byڡ�Q���x���k�_�q	yz-�]��>e��^_�cg�	]�k-���%L�'6��§����e_:�3Tq�	�W��]A��Kqg��"-���n�����rc��fB���-��;̜�ڲ��F������~?��2�P�R9WpK�B�P6��-jiR�gBlV��DI� %�?�8Q�V���߀X�z�%8�~�8��v��-��-�U� ��d�q;��8�&�ǄM��|�!����,�1��s�E�Q�Y��ҠG��Vi̡ʇ�![����=Bڙ�� 	�G�J_�=sz�3��y9y�� ]c�0�v�i�a0�x�#��u��+�s���`�������>!�cw��6�E��lo�w0ڻ�1'�;�E�(4���a&����:&�~IQ�e*;��ܛ sn�W��D/`�a��v�6���B���IO>,�Ғ,vv���!���ʛ\�f��C��<��n�P��2R1�e�e u	��.���t��W�\��W�SL����*rw����sdg7�Y(#�$}��}�ne�l(�[e�{>RY��e��Ks��$Tx�*�ױP|���I��-����(-��"���o��\e���?���H���|���5�~kʯ@8*Yk��l��~ z�/ϣb�_�J6;�p֨�>����e>�:��C�c�^�]d#�Վ�!|�B[똟nf���2L�}+�@����y$�A�j��-a_ 8k��W���E$���Pj�K��ߊ۬�S�F�a�Fz Z�e֯_�U���x�J���|��2�5�k�b�l����+��`�~�r��qр��JV/O~��
H�gƥ���]3����M��-SOW�ϣ�~�^�5"6nQ�P'W�U��5֤$��t�]J�]���}x��7���=0�;��K��"HM�-`�.��p�<
!�F���gNL�=o�BP	g���@0Sp9��Z��U^34��rѮ�Q�U�n�Nk��h@�oE�cB֋��8"( ���j��|�0��Y@�F7锸	~$Q��(E�Y ��<U�r	�e���u��|-�b{�nU2���L���U)���C�?ר�GN���d؞�üV�.�|Gd�nX ��	Ň�Wyu@L,Y�(�-
�[�tȶlb�W��Kh���F���zZܢm-���!��Q��9���y�j��?��>@���3�Q�4�_��BQ�ަ,Wq��*M��iw��L�G���9��Y�Í��d��������2��֋�<'�l�&�I��Wi[�j�Ĵ���dpH~o��ʙ�FIUa�"<ff�=�!�p��*J�|&
�48������">Gi���b[���?u��#�s�ʊ��� �\�V�2=e^�L�-={5:���)	M|`��&̕�5|"Anʋ�ɔ�6������_9�H�u�w�f#��g�����uX��GVN@
��z-���`��<[���=��^�7Q�r��g�-=g�*c-�� '��n	���GM��d`�Ɍ� _e��&�?���)�z��#����td����F��._NS�g�`�E����P�+��Դj|؆U���L��+z�-&ُK�j�%�4V !n(�V���9޸�>�d��H�ۗKG�,.h{ѐY��"�i,'+ap*΍R�>��y�Jyb~�a��}J��g���c+��B���!��F��^�
o�B���
��M��yE��e��CW<1tR�����[�W��6�d� +��C��RU�Iߤ3�����I��I����j����;��N���Kщ�::_$�P޹��"Y�v}���0<���I�[)�?"�,��w<)'<���?}�(�1f0���0���3�Cs�ڵ����F�ޯ_����u�dI)9jV8��z��^X���\��o2��z�����k�;�<���S����g��::jȁ�y����"_��n7\ɹ���&Ċz���|K�����ϭ��D�D��;�#N��)���%�]9DL�4�O=�+>�#_2�R�ߚى��څ���C��܍yY�45� 4�υ$��;�d�ݷ[*�^8���J(�J��L��pF|�g0I��ޜ�d�٠��~Eݹ��$UM6u�PY����'�zm�<)�F:��Kr4z�5FK���b��vs|%�E�w��$���,���dKs�q�5�X�`^��S��ƞA�_u7�Իʏ�Zv/^o�n��]�����H�e�Yʁ� zX�6�#T���#��#�Py{2=��b �E�<vVҮ��"�� �d�Gِ�\f����?fÜ������G�}H~$dg�P������=6Gn�aE>nt�WI/++�I�ǉaǸ#�<�>�a�SM���b�}\6��;����[�VH@�a��4�� ��Z��s���땧��_�����ɕƸn�m�j���'�/�����Up���][�m��������S���<A��l:��/�M ��Q�H>UǴs�1��2�!�xa������$ D��$��(pxO��%�����˧�RT�]�Fy��?./�k�$�r�iZ %�ω��OÆ�|� ���#�5���T`�$I��w�:�]����`�F��00��;���O�ǟ�?k�y��FrB �t?[��-�x���d}���ԺL��n���)w��] ��@u��r*�P3���w�dH�c����Gp:}����|ƶ=@X/�j�uR}VK�t��37B�ǭt�$�J���Ne���kM6_�/��]rQ�:�0�lS��J Qp
25u���o�{����tx��X*Z�S�����k����Vb=���U�c��w�h,U����!�,���{y��ǫ 0Z�p�C(WK�%]�{��>4�ϭuU�dVЍ�(�Q%��O��|�Ǆ$'m[�O�`(�B���IM#�b�����K�gi,$n;4��3G���U�*�~�۴̛�O/��azs����m®9e��(Ɇ��4�\n�R�0������!���0,pQ�:��3&�z��ڦ=�)�2b\#6�5�;	���#�B�KS#rGO����QOZ�B�@y���6�Ӳ����+�<W����q��H�УN����t]�޿��~gė�1�e���?�w�xS-^���ׄ��D���\7W��\�N���Qta��d��[E&�KX��{�H��U���h�҂�:�r��9l3�h�)��[�zu�{����:��N|�-#�y�}ꓭ߇�oy��p�ލ�
m�����8M��xɎ��RQf>1��J� Ύ@��m:?y���%��4��(
+̬�WTa��C�yc�]i��u�t�^F�NF���*�qxE(Z�煚QOO�W�e�n���҂�-���$��_[&�Z2g���3}�`�� ���r
�X��H�צ=L�mи�@�:�����͔H�2"y3w0�x�?��ٞU|{��S-�x�o*��:�a\��<�a�� h��5�#�VK����8�v;�%�&18_�����U	�W*Z5�F�S�k>�k�v�zƣ�o��I햼�
\�
2z�/yQ�ߒO�,����<���[w�+vB��O��+��M\.x��ON'�c�:�f^_�����߿�����
x��/�f��E�!��9|b�@������٤	�OC�h∔��7� 1�/�{���
U/��VK'�/U��G��\]����_E�3��O�=S
��o��_ _������'C���qK@���ryiT�M����\^*
�GH��}\�����/��}���5"0{� �s�o�j�1�_k%��m�Rfp�����eU�%�K��UH6D��m��v4� ~����A�`i�,rԼDP]����'S^�ُ2��TDP@;\�5Y"������{+��w��^���eo�h{��+����_�D�t�P�&:Z�ӆ ��z����X��N�Q3���'�U|,�r뚎�H�U������3#8�Y��*~�g���*��4+ �Z�6"�5I��@������ɔ��C�u	Ǩgx�d�5�4n'ΖW^U�|�Qm�DK�&��4���R�[��Fȟ��C��xi��_�ѓkDNyD�b���J��lE^E=g�A9�a�\|ݾ޹�Mꉕ�c��w�xY����̓@��w:�ϯ���z�I��S�!��6��TT	�qXq{8�=UD�<��x�fXTa� Q�8����HU��K�(Y+�ĜKn��| �~�EYDh�kmE�q#k�De���O�[�\�a�߇1�hSЩ��.�Ћ#]La��|��ƹ@�.�1�;��|u�PpY�%ʪ�h8W��P�iSm�������QI_Z�h��R��9A$}c���z	 hX0THɢ�y������ì%��{�� �����ug���~���D���4�':�<����m������&�=	��GU��v��B���\2���W�@������L��tX��S:��ׅ��
h4��ch����h���Bʎ9�������0���])+X=g(A�1��{�!4��KǬ��G��k�n-OM?�V�����.��\�0���8��0u�i��m#����]7lmⴇ�N�W��k:�I�#s�C8o��Ӛv��U9z�0j�'���î(�P��r*B
������-f)���kM����RT�>�? �H��<+�p�������A�L�vS�$��g:!�K�^�/�+��x���*
.1afA WR[�k�l�����`;�ǳo����<� �m�����V�п�HT��>��,a|�U.�2�3�M��搬�]��oGQ�Ǌ�v�(o{�*�4t���Aw�`�������>ܠ����\��H������7��%���$����l�K�A{9�0D)�Q,h��LYb�i[�[��.=��s��0��2Ԫ~C�^�qI��4���RneC�i��q�d�\0=a� �E����`�����9W&��V���BH�������8��p|(��{	�m�W�bPM���&�w�z^�,��3ZfH���_=��!#K���t#�(�X��+�'6��o�u/�!���}'�����ך��>4��T��-j� ~�46z �?� ���Y�����)D�����j�o)w�\WTb���[�"tڨ\��
\{��"��W�{����e{7�|�������}cؒ�QC������"�О#�9�<%2��:,�L�mY�~�k�Q��o)���"I	������{KXI�����5s�@9sմ�ڞ��6��`��#Cֱ�5��3Kʕ��1 m��Ɂy��"w��Q�=_��7x�M��&ۺ�T�LjF�"�`)t���߇���1 ���:�Rq0yF枊���B�/�
�էs������@t"hDz�9է/;Y�t����ޞ�iF�$%2��+�ȹ��衉W����.is>�
T��Ə�48��PPEI|�KZ���.aɿ���� -�mhM���c@=�����C���XA�����S�jާ�������1a5��vd6�;�)A���� �Wl��z\?�X Ln�M�\��la��Ȩ*O#�(���>���6��l�ǈ¨�K]*@Ζ���Eǯ?κ!���?��̝��BxOo�p��cP���U`�ޖ��
��稣�7p�X4y����u��;�`�7zq���hv�`c��=\5�b_�`T&�*���e���4<O'KW���J��x��Owj<�����DՇ1Dw���\[K��E�ڍg�զ�f��L��@{b.y�C֩j��(��](Y��ů�� �:5���(�Zv�����pn�:c���6v��C��-��aܰ�Ei�@};��:ZN��{F��B/l��&���6�WP:�np�LB��t�^�
T�\�tMmܧ�r�'	�7�_�����BC]���\�� b�x`�Ԕ���e��\ָk$^�Ӛ��߰b>	��A"�*���kvW��庭�s�ao�i�OV��D*�n�#�C1�מ�g+����f�\�%!!��̂� 0��o�_����v`K�IX�%]�P?p=C���[-a�UA��M�2'�Z:���sTs��G�UV�9��v �{ŋW�gp�HcG�W�t�	_�y�\rfZt�{β�-Ƽ�����{�#[�-�����?�V�Ih7/f�{ߌ�0�YzePɊNT�$��1���C6��5��mC�!���M��;i]����� ���w_Ħ��b�N��\�k��b2�i���(���z����F;�h�mjA|����=e����r2��Pˉǽ�5k���%��V�3���򒓕|=���hu�r�V99I��zw��1Ƹ��1{] M^�AEffq�@�pi�ޥ�S�s;�|
��X�?����=�UlP�� ^k�A}1���?���H�^�cО�#E ~�0!�(����QUe���`4EF;-�7�b���n�n��k��@�鱾Ǡ�������N�=uERQ4"�=�����2hw�
����T�5Y�%ɧ`Zfq��ċdW(�^�;��g�8
�de�1;���F8�R���^��Kn��O ������|�������i�J����S��[iԪ����_=i(�AT��S{� ��: ����F��
͟��#�J\emM��mE*�|3�:K���l%�H���R�h����+��[@gI��.��U���� �_V��EDyk����oc9o��ONʎN_!V�淾{i�74��a@�~�Ò36ԫ� ���fY�lU���G�	����N����o���+�zÀ^��hj�����X����"��{�/��RV�$载C����j3ŵPB�W�$ǉ�;��yd��G�aq��W!���iѥ�Oo�6pw���:Ç���.uB�
����ؗS鋜u'�����%�id ~��&�
��r��ME��/M��G�v|�'�/�r��{2P������5�����z��j祕&�bJg\�٧�w����c��f�V�5�X�n�Y@r�F��H��Amsu�"�ŦX�r�?��S�Q���m���l�E��wK�{<�m?=L���wu-��a(ٛ:�5A�`������<����'>h�m�(��K��<,2 zq��Ip�tE|�Ku�S��0��*>B�6�{3ƥ�
�/�$�Zow+�w��.�qñ���r��U�o������I~:�����1is�)f Ϳ4���K��Q/�V�R��n@EV=�.J�:#���E��3v�	{a�Ej�x92������o���ٚ,V7叇�i���0���p
 �jWwe��e,q�h�	��TG�����W`����nی��L綖���I+��и�eU��h�UX�<PSz`SR���H�󛟃9�$&�p�8 �,�B*r��~W���\�$�%C!���A�b�Qeh�%?���Ϧ��A�eq��RqSt����������G�#$J7xKY���?�� �(m�椫�:|$[�b�0��n��B\g��LDͱz\�˞� WQ9!N')!��\��ʌ.:�
�fI�p;�[�)�*0��V�Ȁ��߄M��x�HpȾ�stO��+*V�:���w�!e`?���(x-�0�!��v����"���#27�e���<�"����%�g�f�	��OV�ƌg���\�Ѥ�tt��6s=b�%F�':���!I|���?�+`W�)���M�SЌa�C_?h���+��ډ�yUkykC_�Đ�V����\�YϽ��� ��3�GkV�Cs�Ƌw��~�鋂���+�u�Ʊ$�8����!���Rʐ�SV�f���E�dk��Ei��$���p�t��@ێ�ޖ�$�y��#�7z�73��X"@��=>��?�%M4�D���I�2*��`� �^ִB���u��m���НNG�L�r�����	��҈ڑ�?��\���:n��!�=��pm�L��a�fB�$�q�z�6ȣ�a��I!�����)B�h�r��(�eOS��G�Jv/�,���2W���}�����}�pi�V�, M�O���\.ȑ�j�C����eT	#�]u���?���R��,r��[�K)?��u[)�@^o==�|˧h�sM��,A�'�a�� �l�����x��\Q?�?B>����y;/���`��������p���Кj�H&�/Z�-�O���,������Q	��1�h��G|��+9(��&��,�T�f�{�ZK ����P���#VXC��K�i����hR�u��Z�P[0g�;��i�HB\0��;[91�_��NQ�yG����~:Ә5�d6eV��l}�S
�+jٝgT}y��I�C6�"I#�uf?ʯ�*(N�E�u}�%���vV�Ĳ�1:Q���M���.[�R2�����%;�h(�PYd"κ�"���2��q':���^�""�9��ԏn��c젏~6;t����X\��c�b��|���n�%�4�Z�������X�(���IU5��{��f�'�QE�#y���O>wW�c��TvፘQǀ�߫�?ɧ��u���΀�r!"t���7JZ.3����گ֚�Tx�����|�>r&�-�`���I��БZkV�B�5q�E�ᇃ��`�!)C�3t�j��gT�"?�������'���@�a�G.W��R��+H���}���sv��Z��B���d#�'$�*�Z�=@��C?���suā���\3��f��3�Ѹ��HN�����dHT��t6���.s��n<����Nc)��ܪ�ݔ��Q��r��$�y_�;�?�}}H�Lw��/ͨ��K:�rh)R�Cꚹ�i5�}i¬�������aY%{i�z����zv�-*[jȒ�yΆØ�
���F��F
��Xh�!��2���]�V�.I�T�U��0�h$�Fo	Dxﯮ� cT��H���%�
Ij�]�h��e��\z��+�V�� _����>���|9��V+J��U2`��G�Y.&��^���X+E)dy�e�A������r�IÏ�]ќ���"��Ǧ�~c�.;���Dc�����yI73^.�g�O~��dD�+�jB��;�z=�)��ܜ,?5}�{�	o�#H���	�z�@CA��:W�Ǖ]F����M�
N�kp��Z�p[��J�J�� �b-k^�Lp�%C	���%M�}������<��Ps�O9>H���D��%�zSC�	�@�Q��=����LH��7����o7��o敞���^���pe��i��D���U����e J{/I�G6��!lu�%Z�w�w9
������U%�����,�a8��Bv�ܪ�쵽���}oN��q��2v��P���=�+�󶈧L�y�פE+����v-��A���bѳ����48y����2a���wɐ���yy]��L"����ӫ71к�o��K@�I�4~ȍ�-����������8�,�Э-ab]��Bڇ얷;8 ��E��!�"]����ˬ� ��|-]��I\r����c�00XG3:�|�yuS�0,��m�Xj���qj�@�k�Ms\Ej�;��k���A�u08;��m0��K����6�W�{�$�R�EH�`��{bѰ}8e���[U��C�eNd��)�����':a��~�� �/:{Wa�2�ުO���Nuр8�n�Q[\P���*F(.���<ϕQP�:�h��	D�\�ͼ��C��/aTd>|��/c�,�
��l�����x@�~=�����KJ��`�56�>���j�l'��[0�l��M��Y?�<�d!�0�����3N�"̽�x�ZIr�t����R�$�	b�k�p�ٿ$����__�3�D���:�����oe���BW�9X� Y��W�	H��c~�_u?��"�%i@lД(y�7"�Y�bzK��!����e�źEU�84Az��,1R�?�R�S����J�^�LǫQ�g3�B��PB5]�cN�t/�.��֛r�2*6B�,�6������ne4w�b�7�e2�vBU�ċ�+<����}?�~y�P=	ƃ�Q�*��B��N��_(rhus|���
���uhΈO{����{�A\����|��5���ߥJ��Px�k5�*�.�C�/������L�)^���BԄJ2^L�5��K�?H���"��о�)�n\48A}.�<7��w�tq�z'A�7c:/g���9�	�,.� K���8t��o�4���:��Y�'��%BJ�=+�e��g�X�� ��#k�2�ۥ	x�q�{Wy�6��z�`�r�Ef�H�q�o>:��ͼZ,���F�Y��sW|���i���|#rC��E!���Y������˘���]�)���K�G0 �8Z�ݴ3*�~U�OQ��"��n�y��a���muȷ�� �m��m���\�!����X���A2�%�����z9�\Z�}��ɍ�3/1?���8�E��ߟv�djn�|��� [@G���(�@'3�kX�I�Ze>"��f.�z"b�ݵׄ�1B.�f��%?F7#+��J�MK>���kr�\ ������DM����}�e�_�K���_B"9_��~ѩTq�	�� 9�e�{r�G���g�{r�C%ժ�H�ŮQ��de���nu�۵A0��� ��ǁ�(mq���h�ld�mL�\�z�膔�j<TΥ�̎��|�`��S*IK&������r���*�����fUA�»h�NeZ�������wԬ$<nmY�Z��u��`M���g��-ʍD��}'����R����}Z����ɭ~i��-��o_��÷;��2�a���}�#u��2D+Q�=��>pT��|?������9��x�~Z�IDC�+M�����Ѧ\q�zr��]��Jg�S������Y�&m�j����C� �ì��*��IP_v�ic�ʜ	V9{ϱﴶR� ~8�x���?�DC��BxOi��-��M�-���w�����Hc�g�U�k*���������k�E45h���0�(/b"�{�V������zGʪ��WwU�
ļU¬:̆	���-#�G[��2?@��i�3��m�8諥��iq�#����*&�"[1����:��E��g}�u���d>����ß����6΂UF�C?Ex��R%܆-Z5]�b�����W�0\T�N�D�����y�����㬝�x:�/l��k��,�u�E=h����+.���o8<�ӕUMs
�� �4�>�=�7�Eۅ������uk85EgV���g���n�K���]M�B�6&�f����o�m,��vV��:�D�}��E5M=
�T�Y�ƪ������-~+)�25d
"�X����mk�7*�)(�@��D�b�-���;$�<CϬL8�mT���t�e��|�Eur: �%��i���� ַq�&�6XgC����HJ���u�p1��������e��OCƲ2#������%�u��I�N�V��P��z��F�z�y�i7�&BZ��g����
8�)Ć� ;J��"	��l~g���Z*Y��>F�Ʋa}��u�I��jp�<��ٿ�]�n�eVYs͕�!�y�͸�γ4ٰ'^�"cek���kW���y����31�Ի�Ǵi���干��{�`�yc��lN��]�O꓃5�1P��D>��v�.P��<J<C�#���܀8�%���Q!4���1�4��m�my���[&WB�M!k��O�h*<�������d#bMTbOG�&�ί�a����n��p
Q����U�V�L(������0���r#�h���U:[���"��r��^�d��H^�c�W.��^݉�,���z�J�N;m�:Z���I�l���������A�nps-��Ʌ|*GqM��K|�_����l�KIx�B"1Y+�)��NM��+���B��;v!
�ܛ���TW}��< 2ð�"ʖށ\� �H�J޴~��O�]G9>y��L/��m}�S9萰أ�Q|��(�&���D�ñ6G�m���v���+��=��?�s�[�||�^\Rh��A�9�&��4�/�;��'co��H����t*b�4��[���}�&�SS���3�%t(>��:9<��zl���� �����6�lј�,l���KR=�胱=b�X��{i��8xꪮ�B���)hТ�ޘ�I$'��ʇq�E������*a��:��s���>�~��A0͉O;�k~�5��w�	�
/DN����+�gl�WQ�T��{��=-i�(�����%�p0ym�'o=�o�C���6O�?�{"]*F���	T��8t�A��q���a�}�
T�}#N���ޞi�h����G��XM��w1�[ē��-�h�J�aE5ſ�Pa9��+M�W��U�Nɲ߲�P;��t���9ӰJ�Y��cу�Ϧ���c�q�1������+���pZ�nl�|�Ow�j�십V�L��q�)Q��	�@^d��L��'�n���ʥ��V��Z6�{�[���%�Z��PǱ���o]�������b����f�Vi���IK���� Y���C�"�R�r=���$ͽ���]�<4�����s2G��|OK�*фd)�Eb�oIH����@�2�L�S<��6��֗R���[kNG��'�!%Ae��!�xvt<����If����Tc��*E���l��m���.�*����)��cnڎ�p7W��Cɾ���[j�p��T�П�5%��Ot�3c�B��SQ�.�%�����\d�:��V��E���V���)���Z&��&�K��$T���R�m6v\����4
�|[lx&���!^���ܠ�w�F�n�����n����U����m6~��$}��g̔�]�
���2���@���F�#�kɟ�c(���G�J�`��D7�]rzJɘr 0G���mT6� ����ؾ;��M�j�;H�8�/����c�We�aS��m�݆+��B@���sǴ�r�l�k?w���ɭb��=R���m�h۲��~ģ ��j{t�Y����N��(.rD�ѪP�e��,������E9>��P��.�k�,��g��́j��D�΁�,�<�W��7���T�$��p+�	~�\{����F������Tv�鉒^r�����3��LM��F�0��[���]�D+��8;��z�.9�?,>�-{��/E�_�f���#y�E,ú�p��ε����J+�}_�/#��޴:��4$���=@5����|�Nl��-�ވ��D���rG0H~��D��M��x��h�C.u�������(!�]�_�֚�;G�
���$����m�6q��"'�Mb���5x��8JCBTcn%+E�gv�p������~=��߱���Bc ��i���}fԃ��Q�&?]��H��:Ō����^bl-%l_����4� <���)�a`�f?�{��|Z�W-��4<�c�ohŞ�cx��*Q�A��9��B ���u�$+S�/����ܬ๲SO��X�KёKO�ѭ����q0�汊cA�X<���U���2�8�c9���ȢE���N���y��(?���KB������ʿ�S��t�%Fʪ(#R�2��=��
.9����V:TTY���ܝH툽MM�7��z#��O�F����{��;�1^2�Z6�6�����r{�=����Y5�:n׭^d�oX�\��"(���bTg��ڰ�mm��E8W�^�[����z�dQF7�W�v;�P?�E�b)���±��yƖ�04�AGcf��ڱ	v/��[�*����4���$��Ӹ�[b�1ّ ��8C��'�u���r{�3n�����c�X�������q�JgU�Uw���MCc��ŖW��.E����I�7��*b�5<Ȼ.���gZ�2�O엖,"�+:��<d��i���n��T1� ]5P�e?k�}�z�|n��:)W��-�3��@A��S�A��Ų�f'|<Pw{�{��o9��r9݄\�'q�U�fW'�����s �8��YR� �����E�Ȋ��Y|�:�����anr�1�84s#�z���n����rd����f������:�rR�1V�lK���
대�4۟�{���Ŷ]�n�imM�=���	�f��sp���v`x��(Œ��(hHo��������x�ϻ�+�� 6���"S� 7��N��'��+��t�n�ǹ���)!H�u�
�i4����������o/֯E�K7�@��sǏF� �>��
G��+�,���y�X�N��$����}��'���2Z �4��k�^�˞�`��.sH�~ ��l��sB
�u[Č��30+Ƣ�j�$������8OLC�E���c2q���1�C�[8ݼ����'��P���2��6��B�`�&�i�8�gZC�2�z��vcxJ��I`6�ݢvP�iz�m�/�)e�y�����	�����{��h�;ۃ�?䗇)�'�Z�i��X
��xsʲKW�y����4:�P��l�w�L]1l۸Vڥ�F�U����(^��a���\���s-�%���PSf�w���
i[Q�7" ������֛�2�ʘ�>���e�by%�x��Գ�r��8 �k�Ԝ��|�'haw'�Mn��5��H`���\�rК_���UQ�e�K��t�7a�l���($瘼:E9�x�C�r�GVg�d�c��.�Mu�-�$�{�����s�X���^ꦜig�ﵘX$�YS5��d������$�4��������|���Ȋ_!&���5�0�{��Y�K,'�Z)n+"���ߦOE��:3�6k�Zv�&Vu��E3J�ʚ�h�`��qc.�f�o��gr��.��@ \4uE++��.h]Ҫ>@'E�AK|����慠1��rM�Җp|bS${Ϛ0K�
4?��+#G�}�h����r�}���6�?4�yƐW�4~A�y��B��)e}I)H������A��P����5e�:��i�@PC�_�h�y��ro ����;t���%��x�.r�lZd^\��|F�f�z�EV��RL���n��n����a$3���8�Z)!����1h}��ڇ&��q�u�4R�

��m(NG�O��~�f�}�t=!S �6��-]HHߨS����mY���E3��M�-@(��T�ˏ)X��Q���9�ۇC`[�[z)��G���xB��E��I&vŴ"1�{$��$��겍�.(�ů��{��}���"�Z0��-�!^�.���yK,�~��� �Յl��\��0>CEJ�ֵ%�a./rKb$�:hQÔ���k�)e�ݾ��dz��H=�G�C<>7���A;d����������.��(�K�&�ʮ����|<)�u��3�i�.���!��i�~�o{m�ZZ^�Y�����kL9#�p�<f�o������vϋÜ8��4&� @�E�f���Ͷz�	c��v�9TL��8C�=���Ϙ+
�{k$%X��砷%�*6:�5�
W�<!���%%��1���p9'����s�����M��
+WF�
l��p��h�2��iJ���h��g�YsD�D����R��<���Eج�j�/���jq���A���U2o����G�q�����=��S�Ĩ����Y�${��}�z�ŧ�uяB�����,���4��v�̩�fl�+��P;�aEg��0���Z�G	��ٌ#_ܞ�"K'OxT�x��Ȯ��)���6F uv��a,"�Ű��P>%B�D�uEo�1�q�L%�Z�ivl�@Y^�L�,!��������^Y_r�~E^��a� F����P��QS�Y ٩�|��=}��͘��L��0F$�Y»��5$0�N�p������;~���7����]���~C.����$U5��8�fs�!Z/ۼ��wf5�tU�1�<�ngײ��F;.����h���zV�)���yZ����H� ��J15_�{_�_t&���&M`b�IA��=U��dd��> 1�@����Zå���B�g�߳���݋n�Z8c��񊈷uyn���%�m���*��mT��:��w-1#�`{nb��G����i�Ы^�)�t|������3����+�e���g���ֱ��n�`��2b�¡��HD��T}�tp��G�'�W%
��RV�����"���g4�l���K30�����,�����բ����=SXR�̈́�$[��3� �x��w�i,�F �M ��D�\���Tz�H��t�t9+�L����4>���蓴�Vz��yQ�ȓZne��V Ϊ���8:��Ĳ�f�߃k��*=PiW[��u$�Vf�����#�Trj������D����,{����-��+_�����qwC�6[S ��w�W[wj��K?^�w�s��B���L��wy��8�J�s��KGpƲ<d�T�J��f���3Ϋ�m�����m5�� �$d<�a�_\�g��$�h�	�R-�T�%���E���|E{��#c��N�s17/S�����Ja!ZMh�I�#H?~`Z���Y�4�B�o��`c�>	�d�2̱b���,EѽO�?�F��ۈ�S$	k�D��\�B�y�
�|Q��N�q����ϛG��~���c�l�t]|ܮ?����$���;��>�{�P�Eks\	��Dې���pob�<�Q��P��f�(�����:��φn�*��Xo�g͵�9�0
u{��M#����d�/:3�B��2���O��/���W�6Cfǁ�c!=ԢjW3}41�HU�nw��'ԗ*zV�·qW@�1F���ѐ�E�%���-y8ň���PT,����fV�yrN�0��Le�祘��=��X��NJ�%7Z�3�Ƅii�Bv.��a"���&`��_}��N�ԏ>ڔ^�]��r���{� �V�t1�%P7���o���;�8o��0T�C!�(���*R��pU�1A
�֢��F��u���Y�g�V~���J�{�:�Pe=�8u��x$i��r�U��s�Tq[���⠀�A��H��|U����"�c�m�a+�C��9f��5#�(����n���g�Mx=�< s�A�\轰���_�8vf<]���8�5$�YD�X��F�F�.(�⁥���s�M&��4��1�V�Ka5U�M�і]��-,�s�]�M�]�b��^ g����W��[8���i[_����D��<ց�aU�Gn�u�J;gz�.o9R|#>!^��<w�����/�ev�a�A�[�jŖɩ�y���_cG]V:6�����& �J3��c�TN�F��'A���0m6�⡱�i��u�厩�Ӯ�����	�g&K8o����D�Ji4m�{�l���C�4,��b���3���yZ�\����;5�W �����5���F�ƫ�o4�d���~�މ�ٝ����Өh�ľx>��h���b�qgY7vD�{���0�6��o(D[�rU������7��T�eVdDI��Kj�̂8�b����l'@�����g������� �G5�xľ��[f��k��~;��۝(�)�˚w5P�b�uB���/��9��~~��L�>��h(�D��| ����OhS�q��5O�w5�lhIdծ��m7aQ����o�A��(�C�v�d�z^oj��> �?�_Qb]�&1��ت �nݐY���i���n��ks��W$�y�աX"���Ar�QkpGN�
�Ox{���qki��8�-�iJ���Y� �i:���HjL��l�hg���>�d��l��8��lPj�|�B�4X�M���.�
�y�I�7�s�_^"U͋����I�V��H�`�� _w��u�s3�����eJ�]� Z������v��;-<��]���t� �vI�f�NB"�=�2yͻ6S^�D*>_���{,�$S�a��eAF���ä�	�2���1+�$ӧD/����Q��d|��ժ�G	P-�5KZ)=N�k�xL/wgfg[��2׸2̹f�� ������\������ ����c1��&���N`R��X� 6��ְ�{��)��.)�w&p]�)�6�T2��@��e����mJگs���W�I�n^�N�1r2�;���K�[l��?#�{7�1C��|�@�s���J����b�{�A�u��n�̮�,p��|_�o��-���7�Ǝ�2S� eDm��j�۴j��Zq�M��Zת뙃��f����^�K�tj#|�S�%�D�~cx�i��϶�`:�Q!Sf���(;�@�c��D�g"���+��1*�ʞߺ^I��POE|fq����Z!ю�8�E>&#/%�9�\9㦬���9[�(�+5��a&a֞x��R�{k*Z�9(�)�jr+�WBHGs���������n��p�����!��Wy�bd:�%�M�X�Z)J��e��N���-��#]��8��圇�٭������dE�-���8�6�uk�q�^Y9p��?�d;�voO�l�?�D./�Y�7Y�Z�	N��IZ�����HMWÑ�A�$<���T"F�8�۷oz���@p<YE9��?����4^�c��\j�h�w*P�m����B�n�V�He�Rz%����'8AԪ]p!ֿ�A5HP���*�яo�d��9(/D�⼶b�S���3�4ƨ.N=V��#B����k#�`>Z��_���o�ָ�}k���@ۂ�a�u��˼�Ju���7J�%�����tְrj�nP҆lv�I2�7�3��Yw$Hp���@���k.�Υ1�0l��	�[HQ����N-�� �͂��
��4,��nq
�w8��,i>��0���:�<$�	 ET�Q�>���w1H�R�D��pl5P�Q�!��?�ĩ$��/5a�0f�ց5�N��@p�f���g�O:v��[=�A���
䌴�B�/�8�1��w5��ď�KU_���jE�u���雮�2Ջ� ���V@ 84BG=�\u��30	Y#����}ݎ�l�=ɲV]wi?QK|����R�'f��y���D�p�
�x�6����u�c.�C�7s���}��p�e4М��^q�u�L�{?>]�` 0o��	fTKF�I1̑�R{3Xl1闟�!m���c��A%��%�;Ap�)<�#9Y�A�@���n�J�Tu�Hx��ҡXK� \]�.8���Y`ɽ�7�	y��ށ�ί�<���N�|{�&�on�Z/�΂aGqH��-Y��U�Mly�rɴi�%������ҧn
�LV�q_ޭ�@av�"v��T�� e������\����i땤�VV��}��ޱƙ((a{�N���s������㺗��0��0z?ۼ��\�D���+�¤�5���v�����6v؈Ƹ���9���+�Tݡ���ͺ-9��#Yƽ��|�RL��Y��?�aW���L} ��	,�
;�r,��&n�+tN�;�%<rD.!t���d�/�;���W셅��x��.�df$A����T	w���#S��c�$"/�I}�ݥ'�m��iH��û��E�"1_H=>��⛞�A�M���Ћ��>�u���qh�*4A�#޼g^�,V��b�1,���+�}����S�̽�~���b���.z��~������<���$d~�{W�#���e ިi����UD�p������X���7��̌���M�nߵ������A�f2'�����Spʎ썇�!�V,\��4���l�Y��g:%�1�N��u�����D)��3%.*�f�k
��B>��OQ-KS�� �^v�媘8�b�c�.W�!��?�)�@z�ɝ�	�ٶ8�J�T��b����l��w	�Ӓ<S!66Ԧ]��ޑp�,�&)଺���l��}ll�NV�^�?H���7��3��^�Hǩ|�~�P���7���oiO��������E�?�~���R#�_��8��h�6�{�����N�[��_�0�D���W&��*-����vWUS�����-�J���v>��6���nt�"s\v�F�El���E��~���Aُq�ǰ�)�4�����n	�p�`�y��An�߄��5�鳛�̬V�*xDQ��X��T����F�.eJkU���p~��|<ɕ,��w$�R8���=�1��\�Y�ۺ�):���C�)Xt�U�Q͍���H_��\���8�	n�Y����EV�_��`�s'g�R�����;��H~�eD���@��y:�JG[Ay3�Yh~|,��6dݎ7���2�u�S3l�/�����>wHI�tFi��C�EU��S?d��D)vAw���0����E'�hlu��깟T���ꓕ�m�Dy�� sf}�����E>�S�7[�+�[� ��C���nJ�n����< � ��H��g0[���"��;�H����ON�����Lj��j$�N�28kjy�#�ͪ�x�k�+�Ş�;+ �fs�ܧB듀��km�%H"ᘳm�2WeB��U��?��01V���!�oA3�}����i7_����I�S�+ ���6u�^f�Y-���6x��HDe�Y�C�!�9d��ei�5��>��:������s�Pǿ�^������ӖS�pǟNy?:�	���}1��v��!���D����Ւ��D%g�Dp��@"��nXi��E<�	�a]mW'��c��<r�iq|�Ӗ *ʥ�}���]Q&�
g��
|�L!M�̒�
ʭl�!��:�4��J�<W1M,n��~c�c�y�Ȍ��1�ch�,k�w>���)�&�ױ��cՋ[-4��Y+��N��uS
vR�� �l�
��?�G��#�ĝg[�����?��e:5=V��z� ����lh,�=��'c���m�&���_������gJaj�����.��z	��bMK�G1��x1U�y��R�,	���ț0�Ü²۩�ö�~g�S�<5���i@d��|["�H��e��Ri�Nv��΁e�O���f_K�DB11���%�5JZ��R�d�l'���_���Y����8ϒ�9��{��S:��
?c�>��*/tp��^2U1u����8��ѱ���
m9���M��_G��f�[,�1��I_�s_�������!%�~|_�Ĝs�c��fa?�O/j��Wݍ|��aג�r���O�3T�䌗dmj54�'r^q����ԙQKs�t�����8!�M�����5�?Nw�%!������Xe��o��M��4�%�4��b�)�|{
���i¼��F��@|zNh@�xci���Y>dg��U�<-��(��Q�د<�M�z�]�G�T7�����{��$-��I	T�$�w�z°L7�/�OA�v�|�3p�%�D���M��Śn�����M$�Sd*#og��6د�ct	�� +Q��iu���Zf�����ap#{�~B
� �����z� �V�̽R�{��Dc�����=��H����c>=��S-c}� ��M� M7F%�~K-��:b�De���3C;}�����u[���b��/�-\���u=�Qw2�^��_�����~[��'��j G������s;��B�-�L�k��)[g!Zs\�N
0�@k��a�d0|�Q��v�t~���X�J�x8�K��+��X���*�p��n(���6�Ç�����RِS56�=o}�?�'��b$x�}�6����|���u����qnlb���o??��ܿP�	߿]I5���!���c����1<״C�������6��a)�\�/S-�yoڄ���u���?8��g��<-�_&h���=�E7B�8oJK	��Ye«�]녕\�(;ͫI���h��E9���wz^��A�mJ�!�'�����\�9O� �k�ѤO}Qg)zQ� 6ꦁ��o��f������_��`��%iLO��E��:���jnYN�۟en�ׄ�\��B��S�PѝG�m�� �\ �E��}k�K~�4.�K��R�"�O���G��Vw˸5(��o�m�T|M}y��K�k��,ر�p�&��5/L;y��k��,W� ɖ+��Ek��FK˅�O�E4�2Р;,���&j��<xŪ?nnx[V]�/M�x�����8lp�y���bA��U�D���9)����J�nu3]R�e��UkG?����C͊[�D���� ����nl����V�VY�����"��}��F����ߌ����9q���zN˘�������YO�����P��2��(��dh�.(��0>��vp���y^0Ku��	.F4^�c3��x�?�A߾�͇FUI4& i�p���ƚ`��j��p�aw��t�8H�V�=�c����q�f��>��E��[
���a�ls�@�㣫��;��V[p����.lYy��J����� �p�{z� c��A����+^�C��z�/�Vٳ�\����^P���,�l�P�_�姝�*Ֆ��xC\���غ�H�Җt�:�Tğ�-�B`�w˅3�����o�G��;>3�$�`/����l��OJ�d)�w�@"�Ia������lS9p��Nd;t����!M�XD+�a�g����*k�����_�S��%H����'�L��W`���3�Ya����J�+~۾1.R��YK��o���Om^N/���ϲhԟRآ�������E+�����;�e�"���@!zy!�D�6�}�H���yKJ���mcC\IY��	6V]�g�b��,�!H��
���Pˣ�I�o��A¹1gL)��#��0��n�)1�Nτv'xA�U�J�X�[X��Ylת,���n;����D{j�#ZA�6��76b�+���эn"���l5��7V�6�UA���d�p[_�e�C�A� �(��}�׫!@H���gW>
�rݔ֢��� <�]6d���i��Z�)[h�wS��,��9ci����غ�Sg�ޜc���'�������6T ӧ-o]!�@lS�`w��q.�ylJ
^����y �б�/gjZ�����&#�k"Zw���`��f�T*&�"�@��x��c)"UCQ��� ��a�ц����drT���=��C����	�4_� ��sJz!���C #S=�ݻ�S��k)����Mױ��6�N�6�ha�S��mg���Fߒ�b �.����a��e�S�4�.�VUC~`^�"o��FS#�1>
���M�o�SV��qf2�C���W��5,ں� �_
�,���R�F�� �},��7܆�q������6OW=��܊�r>����^RMD8�a`�W���L��6�lqy�ԓ���J�U+F ��2D�~�s4����=@O-$
����=$nz��@��̍UG��8�d���t���1�ݐ� w3� 6c�u��=.�����7(ԫ�n���Rnfr���7��4>�����2�ЈLV���M��S!#��>�W+��RK��1�q@��� �3�G�p�
�D�����Ԁ�|�ʲ��p:�D��������� 9
K��W$���	� ��w���Sw��9I�T�~�H�����Qϐ�J@z�;И���8t�O��f����D�mwBG��!�֋eQ'��d(_5��e�U�	4����'��8Q%�a��q��iK��
d��!�5�a�[Ҥ���o�+M����,�m1n��r��H�8,��e�ݐt<!#���u�.G!�)Ϡҳ�����	,�B�^�b�T�l��7��M��������Du�EJz��3����hA������7� �Viٛ�H�pc��mVb�_��H��pX�h��Qې���2��M��[l���Ȏ��t]`#>YpTg�+~w0�7o�=}�=��:2O[MΚ<׆4� "� �j�y�,��LB���v9nU�^ ����	.�a�P��G4�`�w�*2>_l���s�zG�&Vy:?�ʰ��i�Fk�g��S�tP��bT<�1�˛_���95Th��4�;NUHWr8�N�|�>����9/�1Q�^�O�W{g>�"|������.s
ض�5�A�j�S�&�������J���M;@zߥ��g���K�fE�Y[���5��0<
�Ꮂ��s��E�/'j�ݞH
:�.o��9��d^�bC���џ+��@iyu���Ф٥�)>:�ҷ������6��*̂�]|������f�8eJ���sn�x��q�rr��=��>*MS�����@G���< �i2��tD�`�ubV:���q%ʎ�:�u82O��J]x��ż�$`V��o��v��ًy��AZ���2��3g2�e��V�/"��,�K�i]��A,w�):z�C�Q�Z2f�&<`�%�u�Xr8Ӻ���Z�lؔχx�@�Bqj�T?|Ōro^���T��z~��`ѣ��y̪6��V��V	���(Z9�O'�[�v	����o3oc�Q��d��e�v{[�'��R��L@��¾����$��E�q��`�,�m�B���pX��5L�6�1;�t��9���ɘ~��˯8�h|����/��2�>$p��_��U�E,�m��D%����1�ū-����Z�D������h�f��DG�GA�Y_x�et���E�����?�fO�����$��h�duԴ�k��s��8���hr یy�V�V�`�Ka�~�Dcz�bY�
-��Z�V2���V��$�c͕S{��fJw��F�[���,+��qq�$�����������p���F�Un�,�.|0rn2�cju�} �=<3r^/ �K�'�[�������pE�D3����L0w�VH���0C-��x�S� Z��W�s�gΌ��28�ϡ8�	��s��04�f�'�u���Ӓ����^|��*|�$�d@�jY/����n[�/������Y���*���f��/�!1��YC=WGr<������b~�:,�s+����iNC'*���m�tԺ��=�Ԩ��D�n��_n�轠m�կ#��|���H���hN+;���iNsW[��@�#�LY���Be���8ܯ0��Q�nݘ`Z��x�e>���V���*8�9�?���,]�[p���J����+��1i�M&����Aj�B��3�� 0��mXФ�;���~yO>�F�d�3#a�5�^����x���&_И4?o��)S`8T�l��%�	���yV�$Q��@_Ji�-�H}0S�%���I�)��Ɵ-k���=mt��h�ז'�����u~�V�[4���k�'gӖI
>Q,k��ߔ5��	b{����L�@�h�7-Vn]��/j/'�Yifa�
�����!�Ǆgj-��&�#�+>�͖����4pr��%��U�zoM�|���
��տ�O��4 l�ؖ���D���H�K�B´4iU'�Y��鴚��NZ�Zuke�U,�t��8�H�����j�q����d�c�J����W�Ľ�����W�C�IE���(٩0Z�U�=���`�O訾����x\��`y�5\���W��&�&.�#=��-�>�!�C?�$��W��Q�����~�Y��I�%{c�=���Հ��ֽ�<ҥ2nMR�BJ�X'�Iwu�ϥ�W�;��!�
dv$�i���X����=�R���{�_�o�~�¬��;!�� "��s���j��`/GAߚ}P�����^g5�p�Ok����v�9F���\��j�` �X�����ފAhē�
,GR�=1rBM�ԓ�� ���~s�2�&c�xtJ�Z�GUJ����0� ���^}����E�z�{��U��|�m49�/�����_���@$���Q�}�SS�8�z!�*��SBn��ZA�JZ��K��+�=;�p�Es�fɻ�M�n=��t��N���D$��S��x�5���f5_sH�)�V�e��7�lv��K�p9�����|����tX�4�rn/�Ch-9!d�Z�Ff��x�	��^a���
�>e���QY]�l}����9u� �w�{���O�<�e7��}C��J�� E`�SL�R;�"ovt��ȏʱ,@�N�q.��;�*�Tl���*����MTcdC��Ό��
e<��$f���Q��M���؎�L�ԑ�$����ewu[���zh���b�A����Ln�a�D7��:Uњ��1�V�a�N���9�&�b)i:���ί�O��&�i�����܅�Vo�<�I�&
��P�u��IT������
�{�0�f7|�GWG��4W���s+im��}�Z�MG�u{['ӿ�u�ր$��U�#M_v����R�	�¨�>�U��N�TX���+����E�>�8��L�3l��f� e�ܨjͺ8�sD!d:�
q��3nf)�
����`��<��d��z�<���'��cS�>��ժ
����fcU,��?W�����bC(��\=��d�{��D�@�η;�&�_�^$.��z]N��M�h��N<{�E̠8_�J�����5B�<t-Q����ٖ�����tȉ�(ʷ�UY�!�g"d�\�Az��|�hH�O�5"���R���33����H�Ht�è��]�۳s*f�.q+ӻ���۶JL�z���?0�Ԣ�c�h�������&�nN�{�g�Z���ǹ������9T1zU��YL�}��ZX���*n@Ю�=��+�F��ؤэc��	 pm�b�!W6����	����,��\� �P W�ܓ�0�_�].@�=/#���$l��۳W��1�Ztc����|[��0�D�=�V��h���\b�"'j���wP������z(��B�(Lx����荤�۸+Z0���>��n�����S�c�USX��Y	o9L���W����	-*bg�� +���y��(���Fg\��}��;�K���f� Q
�����?�d�
�fƃ���9Th�F_P�����F���~�.�����5�X�q�h�f�VYS��W�Z���k7ԅ�c���\����r��v8Ja����Rh���[l��6��������l�6��4����s�����V#�c� �2}*様�e��\�aa�'-^��%y� �l=D��b��q�:%��E S�JBX4X'���Fq��'t��m���/��Bp��v;f?�Vju���]N��s,��Ĉ,}6��ܯ_��h-{�Нړ������gV��u�aC�l#PR����m�d��w�IL�-�Q��/
��#��jQ��j��p�q���8}'�q��J�3�q{�S
��p.�ؑqi$g����=x��]��^�-L{�ND�H+gۂ�?��}T񊫕%��E�e��6��5UW�LA�m0�2��CV��F�"]��9�3��X�l{���F�^On��^����Z���ҷB=	F��2Rs��Ȕᚲ���U��#]7�"����t�k� �v+ʦ?z#G/J>��nP'���������|�H��Ԏ���dgEq�KLy��j6�sH��Zta�%�x��+[{�k	��ȥC��\�v�EQ�k�Z��;_f5i겥I���0�U5�%��E��&+��ҝ�m�.m,������v��a&Ɠ�)Ya��0�Ka����6e�l�Fu���:�I͍�O�X� 	�k�u�Ҽ��J1ɫ�"�e���zf��]���ǈG��y ��'�{q���\s����`\���&2W����G�Z�J�c�٘p�m�+�2T��mD�a(1��5�tP���J�%EW#=u� S�n 5�i��qQ<x�������n��/������qmu���j����j�N�l=L]Z���B�
�}VCb�5@�6��u���׏T;tars�[l��_i��t���J�%4�Z�����gGz߆�SO���-�j�C+u���y�e�ߏ`Pq���6�|(Ɵ���#��Ow��r3�ѹ}Y��ьT>ٗe�F=�bS��!�d�z���赘�y�L4&��,4)D���C}h�[����Z~32���{��?pV���#��¸�B�\{9~Ӹч���ɲ�afx��Ŕ|���'�HnV3bZ#��J�.���]˄$��������=x���_ �DaWbK&�.A�������Z����`8�����c����R��XGQ�Co���Y���x����Q��
`�1 Hrb%��ƆEʵ���n�|r���_ڻ�1���h��x ��}X^�p������B.�3z�cWڤҰ��$��Mo�K7�z�<�x\������)��;FzuH�2J�T���xw��Q��G	���I������7�PD�Y�������8/'�}�3ǵ˝<À^P'^�I�=��{w�_$���:�յs�n��(��j>9?I��H?��yN ��5�U�3�/O�A��4�$�`��hbd��n
�J��^��o�:�"u�[�V��_4�	�'���&,��n��]�����T��g����W�eZ뻳l/�-\E�t����G�s��Y�Ӥ&z�$'u1vJVÅǧ�3�`��	4F�w��-?�P��nJ�B��ς�M̗6'_qړ�vD��\���m��ڕG�e�=2-���5G�*��� WK��q�16�(��h��R4m���T�nIx�����V��w�uD;	���۳&���U{�h�Qk}B���tq)�ҞԈ��#����]�8"��=��f���e����7ז����̜�=���bVٚ�=g9s��|2�S������N�on������l���-�V�� ]�pd�J�!h�(A���sMXP�3f��+1��r;�#���;���I���@���mxA&I@2�=���B@8��1`$�q� ʩ���1�*Ko�0��m���v�ѵ�"vB�a���3ݐ��`ݢx�w[��Ꜧ0sպ�o��X���)?�~=v��� u3z%x��3Q�LBj�|_�A6�~�+�(�@2��v&?��2UiuK���:{,�M?ς�q��u��0*��e��A)��{����YC�A�+�D�0����%I���^��g�Q�c� �h�$U��� A���ޚ
⵰ǣ��a����⌘[4?�X �=J��*�Ar�ba��z��{a���G͢���I��P�ݚJ�]W��YVH�L�]��87<t������GI�}�1;x�G�p/mwIw�m~�������?�ӷ��H\
[4T�������/�!��鄎��� D2^�oK|�`�/0���_H�e@���}���Տr���扵j��l��S�8����S�8�ZH��蹿��1f���wb��f�����N���2YJ	O�WÂ��o�衵��U�\5n(�0���1l ��No�~��K�E{=��u��{>scA< ���t�1i��f��&��W�$U[A����(a=7K��2y� n������ޔd�Ǐx��8~�s���O�z@���$^��\
����50Ja����(�� i��!կ2@s>c��~Ė?ݗ�w�Վ�' ���!l�ż�G�u�Q�Y�t!����0�,��`1%RN��1���� ^9����cSn�SBr�L3�96��nE<��tQ\Fv*��ˢ�4X"L�Gd�+�#IN8;8X�`FUyzu���$�>�D���j��-�����?�� ���r��)��?W��Y���3?�e�_��f����H��}�V���k��(��D��� ͦR���`�~�^�Am�p�=��_�%ޘm�{)�TЫ��o垻غ���!�]M���/�F�%���w�om即�i�!�>C�p�艚Sj�K��5sG�>f�� ��t��o�ؿm�_1	6�$�n���J|Y>�F��v����w5�ǝ�����A��:�f':�5�<��t�S�羓�o�!qLyM����S�d�顆�6�j�Q��M� ��|uW�[�@)��b��%`�:�'@�����bke��[���$n:�/K���q��go�օb�����*������q�$�S?շ���g��	��d�:u�[�Oܖ�B��L���y[�JUK����t��/�2���;�dr;�~'�AU3%dDap�� ��7�=ݛK��9�V����Kp�%��uR#���w�d����&ۿ����9v&]�(!H�Ů4�
�{�w�2��ۍ�La>���LVo12�{����I*vT��6f4�����o�(KL�-aƫ�$&��~��Y
�l�W��q ��x���0�M���XT�/)�T�K�v#�[�X௘`�Ί}�3�n�UXN�+-�����|Fb��4�zX�˨+�$�0
>j�qk���Ƿ�#c7��Be�TQ/@{��r�pw�-���ECF	/#C�����#�'0"Q����{%I��@&`X�\����Y�����S��s�� �h4b^M��)�Y��fq�� '�ѯ�Ծ�w<�K��D6P�A��B�]�����B�z��7mR�H��_Mt�*f���(:��V�[5-��<���)�&RT6�ۏ ��.r��s."�;H��Է H�-��G�G�n�"zy|�VT����<jn�FAs1����ȓ�P��L6dd�ͤ�BЌl�kT�Z�6~�C�`;���۲C��������ÿ)o4�\��mBT]3ؒ��ҝ�e.R�m��7:��'�H��e��M3۾�߸k�W���
�oV?����RW���A��X�Ǒ�A�?�b��YͮL`f�3�-��k�H�/�o�}�ö�3}ٮ��u"��i���d�Kve{�O�T@׵�p!�7Go`�wQJ����ac7n%�0�87�2�* �v$���}����d�A��]�^MO\�l~�{��N^208�wa��o��2��7'F>� r����JfdLzt�ϭ�z�On+�������	P�Re��:��z7I�G��m���>���{
�m�q5#Hj�a荡K�EnTN�G�g���(
�R�ѴI��z�w�3˖�~�����쫭;�ht��$��3���/7��{��)�gX�VF������b�/ñ�]x�qe^c�9g�ué�u���g���<b���ħ(F�[`þ-��{K�G��y�j����w9��d��h�6�**���9�4||лJ�ou��m��?�Z�4$�PY��߰KÂ�F��*"�*�������&���Y���3BEps�'����BdU�!gPHU�|�.�r�w�bck�S�Q�@��ԝ�<x(غ���B8�96ԟB42S��0_`S
Ჳ]l�` b�
����18�ꔟ��a�1��JsT�l|���9�A�*<s*Z�wp;��;�\�*�߮��v&U>a����� �� |��6<��#�}���/��~�u�[��=�h�dP
�C�B��ߥ6`�ޟ���t�z^?�̓hS�򕦩Qg���4��H\���P��:����C2:�P�J���3�h���
��)�$Ԯ�l4��͜��{�&�!*��F��w�\�w�Z��؞G��Awd=s�c]����X9�WG��*!���-���v��jK>7!��R����a�8Y��PX�z��Fep�'�}:���8�����*I&E#����p�*�S���^������
���r������7,�԰�KΚ`��CuPR;����T����S�;
�-���؀\�M��YO0�,oV1�y�yi�B,���O�R"�q �����فĀ��g�7�+�&��
w#n�EtA
]u�;��"���l�i��׶�����m涞�--�J:�t/�a�6�)��2���j9�F�!�d����1���@%���0k��]<������#@[������rz��QU�8��>JK�uo����3�=� ,sD��i% �Բ�'�~s�����q8=��g�e�4MO#�_C~�O:�������&��ɞ2y>=���5-��һ��W�&�4I)���F-+��
�||��3�'4!�>�t��ʳ������e9�ů݅�_�Uo�K5�X���c���;�ћ�PA��`�� oZ�|�@
�n@\Q�31�b�̶�wBvw�qo,��"6� õ��b�qz�v��*�8��E�뛯f�ɒv �̭Za���AG�����3��_@ص�����	�t[����okJ���� �N �Z>�D;�%��$��p��{��^:�e�ʠd���[GE�[�yo_Ҹ����]����v���_ŰIu����O4u�Ǌ�� \T�G�͈�/���h���LU(��(__à<W���R/+8ld�
�~� p�G�"����R.���|�D�_Vf�-Q=a(��j�����};'���A������z��q�Z�v�ܸ	�J� �w��.j��@��^���Ш�}g��g_�qn��xA�z�1��&[�dag	3R�[��-��O��\c���'w.Z���d�����<6�ʚ�۾	z��@|��V��L��Q�w��F�c<
�o>�Bl|V�����!IS����7[�$cY�y��h�P=�rڠ.g�8��?���%뀳�|��ƫ�0�Ϳby1B�҈%�_���q$@�6r2��)r�M"��at�(<��^�|w!���f]$�{��Q��^O��^�w^I	@i�c��~h2J̗�Ďg5�}e����W���M3�֡�l���l�P�o@�G�ؒ�	n�oť۰��&e���v2Y�3HM����'6ND`�c< �s�-Y�]_x�>te:�������jo�'7��'|�z ]z+��^lf���|~֊_]�ݣ�ft0��EM�T���
4�>����)�W�I蒓ސ�E[N�E	[(�BU6�%*
��2��-�\~kHCc��_O�&�4�����ʉO�2� ����^��;��|u�6��Y���-��/�Q�
�� J���Z7{Xq/�a�<�p��`�[�P���P�5���glP#��і`U��Ľ��I�����ܔ #bK�`ݸ"�j8A �<5��U��]R!�&����q|��6���!�K�������mdx�N0�Gt�Q����z�����3��鑸y��H��8���� (qF�n*[/Ŝ4Ɯ �W�yӮ�|h�0^�|l.�D3�)(�3Tԟ.�5A"�+���v�p}h�u$��� ��e�5]s�p���E.�w	Dז�S�Xj2�ꍓ������]EsƠ��d'�rf��pF��m�Mz�9j�����s�{d�m���N��Iw~��U�ī��V���
l�')yU=$
 6�f������5�m3�'k8�:��0K��ŏ�`���^N*C� Oa��3�n�y����>�oH�Y�5���v���4�X5� �2��j�u��|�zdK/@�%�N��uCT<o�Q�����������vO߲��׸T�æ����[�lP!D9��;��쁗݊��9oo�D�'͸�}c}�H���i?Uҙ/�he��*[u�7�O`�
��, ����A:^��\(J ���������E��!#��XЯ�s�5���h)�Yo��⏣��'��Qq��W/�g�>�#��WV�n��8���i|����\����Y��"�������ܖ%���ؽI(h�hy$�ƪ��a T ���\մ�FF�a�V�93n,
r��{�l��b h���jOn��b��M����,���;j�����MK���z4M�lpc�W����g�逘|��Jz�V��=�y-����F�-}�>��S�����H23�U�ƻ�n��V�7ъ�~D�{�J�$(?�ELڶ(a�L�(�:��9��^��`]��d?��H멬��6�e�Gj�d�Lo���m���g*l���m�鋧�֕�tEU{xY��-��O���T��a�V�V�R�8ρ\�ˍ��������� %AdN>8��%�X���f����;1LG�p1b�I�U��6�Yw�@�p_9���cw6�
�w�㕟�����`��=1��*K
h�UVy;U�ŪZ�Ƀ!��[yα�f���]��Uu4�����!�gt#:����vb�9��b�Zb}-�8S�����}�`ڜ($}�U\&|��M� �NYd�g��CB�i\8y�6m򀓗�Q#:���qV�Ui����wXd����Q��uj���x0���~��� *�{�X,�9��Ӽ 5fJ�0��B�^è�"�F�;��\����Q�5�I�� �
�D ����HǮ�澨�}�l���SA]r�缴s/&@�6�DI�RQ�r���F�w0��P��\�V��m�N�~�#d��>w�g;��z+��ي�ץ|��2p~���vD�D������X�shՊ��xi�D�jŎ�H����]Ăŉ�6�K��+ǫ��[��WXB�TB�/��4��VZ��&B�N�M����8��_��
��Xbw&W:i����E�E��*b�m���oE�?��lz:�'|lhN���7<�`R�O��w}Mc�H��XN�MH��k�|���I��ȟ�/���/���|E߯����Zi����!��'�5��`镟��*XZ�M���3^t"�#����o��͏�0�9X;�BDO�b��"�F�:`ӭ�����W����3)#p��ɴ�7�аC�Q[�U��I�F�`�~(�HtS��N�k/�г�5+g�,��>w�>#���0��1э{�1�b�K�����v��t��]W$���������T�
�듺�~�\`
j=�J�OwW��׳�8����BtO�$�o`aG���$üJ[��>�\�3^�RB���Ա}UYag���A0�\|5�C�k��v�X1Y��|�
IJ�.�
[R�N�]�H��?e_��Ņ��o�ʦ�z~S�W��Ş��?|+��l#����PF:==���y� H�z2b�\aA>�oQ��K���5 ������H1Oj��=y�j)��$�*f>�v|�����?b1�L��Y����uu%�����鄹C�8$�"pn��B�1��{.P�8��V�"�2���?��D��Ε�d��3<�v��4T\(%a+Jޙ��a�	���|k� h�o�h;�kY�}6D��XZCf0��^B�Z<�`�t�ԝ��`JW�?��V���i�;�:�ZB(�oTj�a�����P�+Us�i���T�N���/��y�ߛ�g5��¢����
����ڑ=C���_�L��`������b�tIY�P�r���o����C�W!��]�A��bDV�b�oV��8X'vr��M+Aū�n� |�E96�U*�����`}
J\���I('E�Sk���%�/N�Z&nl�����gױY*�0��X�l95/!A.�p�R��X��*��rt���$�:%��q#��-8�¥d�O�[�b��P�T��}�sa�	��i�S�~��YA�1Uc_Y�N��5fڋO#sGX�`�jX�bj���������)��'�{]�!��ت�%?(�x�߁ᥞ�(R�/���zե_:�k!|�M9��[�ɱg�$R�/x���'X'�JB_��� p��m�7|����P����aM<�7<`C%����?�kqN�=��s��d����}��atz#y$�T�?-lTre;A���2&�2-��z)��M�ĥy��ջ
@�7�n+J�;utK�|IB�6����HH�b�5J,D�fO4�ҫ��2�n;l�i�d�Bn�U��	r6(���I`.)��7[v��ɩ3A��4�5%]�� �ydH*}��-�&���-�IDm��M���{��k|�B�.����69h�Z�����F�l�A>(-Ŧ��@���{@Z��;�\CC�%ǳ�T�T��EU�7�<�0�U�;��o4Ok��B;�Y%L�exŢ^p�Sa����2�P=h6Umh��������;v&�̨χo���_���_�V(@�(���{��������\Ծj���~/�ew�)�^��Z�)���Xg�a8*����^�|̡�)?��7�<[�a*�{��1�; ���vBj;�ٓ��K*'/K�+RD�B�2`� S�4/؞�Q����7n�H,#��b�-oyt������ AEQ(�l���hZa@Ay�^JGWVp�J�(+|t������қo�3ﶍ%|�-X�E_#�z�j\4��~�`3��*r���eK����%M`rlY��[zU^@q(��b�_7��H�-yl�$qD��|x�R��` ��1T��;β0���fpk `�BT�T�(PD `�!!�P�����"����pFIY�)���Od��s�#�c�?���	�B�gn谄p]U/�kq}�`����l�C�����h��6��h��YP����By�úHp��\�8��+|~��{HF)�jN7�íw��;����3���<Z����@ra�F�8�������Gc�Rڌ�p� S��=�vb^M�^�]e��͙D���	m�f�=��Z`p������7�FcA@��\��">�ħ��1}_���+��%*6�F֔-u��%�������~�5��潿o�I&)�F���>
]�_t�6�ʊ",p�?6�f�>��a�5#��}��>V�B+#�cӾi�5#E�T%m��H�7ZD�<@�}C�Z���?����u�iKß P�45�.䮩��w���9�|]%���r���8	����O��@C�d	{�Y�0bǴ�{�(��X!�m�0�Ǽ��!���)�d�l�[��66�G-��k�+������q�tj��N{���'���2�#����w`�̤���?��e����	�a��Jɻ'E�Q�TPB�д}"i�׏:du��Jɱ�U��ڢ�˖�tkp �l8X�5P�V���w�<:�%�ve��s+.`5O�v��'E.Փ�X�Et3Ɓ��;h�팺a�I��1A�����>�%`��[m�E�(l�2�[A(��1$O�BѨ|\�����=
�vc>�F�. �.~Ȗ�zP(PD��j`�j�.a�m�l�@�w�5 �~�^핎����Ō��Ab�z�Ģ��*1Ѱ׈�������x��]���3��Zt���s:�tpp�ˣ� 8��:����=��"�B�Ct�ߴ��������o�p��i8�����w;�x��K���[����w�R��!�_ �GPgD���*�O�'4;�9?}���߮�+б�u�k:cx޴	<�ͼ�7L��n$Z��zq �~5K\aYT~d� ���nڗ���!V�.4�qC>��� �n���5C�p���/�,P*Y�)��|q��x ���eb+�٣ݎ���ؔ���Hb��UK�f_��U�ߍ?���H���d�.��|�{�4j�\c�]��2k���7���U����$k�w�vg�r_�_l�QȓUB�d`�K��LN��H"���I�R<���]�/�>O��2<������c�X���v���U@�M	Qe��a�j� Զ��=��'@�����|���(lY�~uପ�CC�mC-m���u���n���\7�l��~�>�H��� �p���S��v�S�B;F�?�p�u������z�����5���3�G�A��tjMԷ�0�뇭�*�м���|��ʓ=-۷�F]Z�t¿2���e��06�P�mb�W}�]�)�F:�#"�/�V� �8SЪ?F,�.��0����}�x"A0 ,Ujk��&8�vbs����A���^�,0y�O��Zay����������;�<�&/L�K��I��q��{h��Ӏ�vkf0?ըt�(��zA��_�Ӥ0�d+nU��eߏ#�#"�2�-�W����͛l?���1��b;kC��,���>KE�\o	��ل&�C����s�#8ay�L⸈��u�Ho��ޥ�T��D�ů�գ�l�㫹� �["�
4?q�i�2�U.����&� �	g`\��#b�lv֏�cn�8�鳯��R̿��&�Y�����Q�(��)�T�TW�'�n��2�¢�F1=��d����&�LROT�tԜ]+pyȠ��v������A<U4u�Fr���V���F]�In�q�Y����OǷV%�Ε�5h)ʧ���xO�X��s�lt�",�ְp���Ԉ2E���/ ���$r	� ��s/l|kH����k��/���I�z/�X����K6G�7���[26��x����5���� ��\6�)��|V��g�Bq~��ri�t�IϠ�#S.� z�� ��&E'�ԭ~]�Y�o�Md;�
��ir\��,A��K�����qd,��:��Λ���Ҡ��[9т 6+���E�\���q���I�������Sr�g�)�ߋ�kӅr�N_��? �y�O27}LF��¿i|�'�>}Su�f����x��~��8�pQ��O����spt��(�w\�A��­E,��4�'��ufن�����>�U����	��ۛ�g*�-�,A
NO��:�����j����*W�!q$T����~ķ5�G3WK/�]���I��(�6)��H}����nC�'Z8�ȿa��v�"E� �ŧ{�m���=h��3�\�������%q�{4N�Ж�a7F�G�m�mh���v��	��HDN�S�կ�߂/�18�D���7�ж�6]L�[��ŀ��s3a|�5�����#�V��/��SCJץ�`�|���>�'?N�C@�
P!�\��G�;W+��W[�W0��B���}�����0���}�rE��H�G�>zsj�)�N�b�^�kIj:E~���yxI���"|�U�2}�T �p�|���w�bd�6��=#O^n|Ő����uBp���7������ ,i[h ��4����;�۶r	�Ӡ��ߋ�<ǒ�?i
���^wE�B�	�=t�����Q���õ�}o�R8
uyt7�5�pٯ)T�U��b�"�B5mu�vi���tj��(��wj�r���ϫ���]��UE9���;he�3�t&����l��f&9�����ljݼ��ȉ�MK�6ہ�g+J��.E-�"�ձ���^�teH-k��*�ѣ@�zi��������'C��^����u3�����s�"��>PoY���oJz���͠�6����r�	�cD��C���j3w]MK��f�a#��y�;Uk�ZF�eu<c�E��0;;|g��B^���,�Co�[�3a��t"��y��:��|�If >��uR���d��,��덟�˸P���O��3����U�R{cG�)���`�R�/�wf
�]2�qin���O�o�,�g�+Dќ�l��ҷ��]�E0-D$ �}KB�ɓ���>��Cgú6�P�yy\���p�lesu%������_� �#�ߎ�2<HwU��Hޥ[J���ߢ�9f�>�r�3J?���o��e��u�ڼ�Uk�-ȹ�z.븡���nDa��p��}f�����x�.�|;#���ꭣ�ݍ�~
t�ŗ�JX�EÝA*a��?�.�z���yb&��:Z�����[VՋo.R�'�|��4C��x5�fc�I��=�J�&jRLh��7J=��Di�X<����m8-c+C�Q�	}�\���I$��,�<�#4���C�@�Hq���'+ �r��2��W�;�/>�j";--���^?������ˉ���`�g�s Y�#'�bM��ע���&��!���`����Q�R�.�dT?Ӫ��*���($��D��x�7L�d�t���غ�jbz�ި�I+h��x<#׈�Jț���K9b�x�O���1��0 �HO'=r���<! ��)��V",t7�����Z sW�i�W��Vv.S�����y.:�9DXD$��
b�뵂�O�/������B݈4�EiQ���6�'0)�q[�&c��U9MlV���S�W���a{u*�z��L�QL5N�����q�����ȩ?��l��bc�����H���95]�6������{���,���R'�+1x��OIgu8��+z�x3o�#|�eh�������Y����d.3v�(]�Bq��r��\����<X>w�+mb�E��(H��']D%b	_���f��󠮉�4���\��p�Y�^�����͢OS��dH�pcS�1��^�"��6����Ӈ�Y�]F�pU��,�u�2��th7p9{�^J�������ob�U�N��
���I9���/��p�?h�/�&�х�)�e��S��)�ǧ9HG��j�^�L�沖i�kl�2�>���e���|���F-ܺ���!#��._KcY�=>l����z�P	[�n��=MM��L��߹[��H�ޠX��X�%#;�����/7IzO�/Ө��\���듣3,t#6�Kz������m��uh�J��$�[	��a�_Gt�;ߤ���[�;�ӷ[�c�h�+���8e�r̓���$r8ĕM nz=;�ޗH�x޺�R�����Qe��۾����	����l2�h�7���*~ �#�-��Y��	�v}�R_/��#]o��0.�H�W�&F��,�bo�bߔv���k��E��z.Iux�LE�R�1ZU�1����Q�v�2�J�$�c�xs��3��R�2*��-���َ��LA�_��SB�Y6��4a����N���&���UR�#���=�u:��&�] T(d�,�vF �|Ȼ!X=}� ��h;����K�G,R���"�.�R��衵�l�gf���3il�H4�^J�>�r^@[4�A�b�~���_*DU�} (�+�CΘ�`H��!�e�7c��^`��4 �6�6���5h�{#~-�ӏ���T/ӫ�Q+ ��)���`xm-#�^���w���eǡ��s�E��[���?�ò)|�p���fi�֔#�%H��R_��-��U��"iF�4�j����/�f)��hbӢ%��a�X�?k��&y�5��Vu�Yǁ��G����~�x�8��7U�z�ԓ4;�9WYW�E�`�[Y/`�<H�4�\����+��R ��*�4v^w�pL�=�l��
�~Au�LI��HG9#r��9��1isGs6��ߛۿ<�ޚ�>-�n`�����mc���2k����_뒉�����p�>��=���?MVk�j��/x���$��K_�~/� �y��qZ���22,���l��o�����1F'U����6'16�{]��6�ޥCV�ٯ�s'�KG�b���s��JZ�Sx��` "K�0�(�p�9�����}�q��$��CX�M�p�ɂ�|��к�A�mr�d�U�`�n���X��L��.R�Dz�x�KO'����E�	�����n-�V#9w	 �T�G�v���K�#bJ�8{b#:3��>�T!���A�Z��RJ��#�t��%�	��_:��_V��$�81>zĴ�:�[L�sH��!}u�����3^t/��e���
H��3�_��oL5��3����\�ต��s0Ϸe�ᔜx_�F�
��R���h�o6|-'_!�q7C��Yd\kf�7ھ�иS�[ 6�}���?Zڶɶ[<�J2U��q^���O��%U~,�SDH�	D�svg����;�&@��={p�:Q�Z�����٪��O��[5:����	^��.Ճ2���y�K zy�4����,A���H�KO����B�H|����C���D�N�a\�s��@��>��
��?8�	U�?�e����r?�=ʴr�vk�;.�(�k�s�OX��j7!kf�V�QpK<@y�-�E�Ӕ�L_��n�,��X&��⤛~�:�o�<�N;�7�$�f/jl\r\�Nkx���?�& ���#}�%�����r�^��٭�!T�#�3_�$mK�ѕ�m���Ӗ֩���\�p����sNF��w�eX0��u%��C/�G>����}.��[����e��j�z��<���� b��\_V�сb���qPԐ�٫k��� ����=pO�������0�)����A��tm�����I�+�SyB��V�w�E5���L����RG.���y9�U�5�~[F�WoD:픞-ǫ.�a��y�	
���i���/)H�)U�ѷ�?��ߑ�#։p�s@st�U�!>UXVѦ�Z�}�ʔ�7�1��R�S5�V1�hL�.&:��-[����x{���2'�벒�|�w�`'^3��Y��c�xZY��Q,���c���
>�����ϝ�/b�Ć���'687�k�u���ha�Gp���.���:�k�Jf�>;j-�,o#^�"?�8Z@aڿUjs��P��rf��0>�6��<�{tZ�aE��N���D��,�� �!)��·t����OH���zT�ūy{�{k�j����-���M�!)�>;|$|��H������^5��f�d���%�?*]3ΰ�%�˦h�IE���H;����KN�t*z�-�����W[hz��g�1���:�I��qi��P}%�/��	$����6Ti���,���wE��Wp�k�Z_ܳ�~��q��V� 6�ogX�� �����5i��$�P�x;߃' }��Q[���Q���	}���~}_(҉��z��:猪	N-�Y��@���\=�!���R�kd��e�k��!X�4#�Xn0%���E�:��)�3a^ɯI���_�A�ҫf�����逌
%9��L��jqQi��_/)�7@+*/?�V� �v�pUI��#����߼�\[�Z�V��Y�ލ\��7���09w�"l&gB�Q�G��~H�c3/uz���Q/#R8q����0;�慰֛x3���A4�����a�!�@q�_�h���ʌ�Ԩ�����W\'8l�jTT���%���� ��ι�f�y��;Wix:!�,ȢҦ�]�}�p����w9	k��������'x��&%��
L�K5>���P��z�(��TK^<�@*�=>����x苏����a#�S���3h���N�@⹼�a���8w]TGu��E ���\Y>��o@�	�P�j�H}�zwC6���׺�.���b��I	)��z�kU��ȃ�7a�G��ŷ�L��A��[�x�ӫW���_m����Lt5���:���$���=���S�;�_:�̮U��V9VuH�`�w3�t�>��"�0��\�ݯl��O���x�B�<�=v�〈�u&�Q��H}��7u�ɂ]�����&����G��ƚ�{��Xŉ�����c���(��09j�c�!�֙�]��y�ꨥ7�|���R��"�׋�����5�+!7sk�~y�)��LmG���5�CB�2'a5��q?�C����>�]�2r=��F'���i�猸��������p�w�YW�F��"���ʲMIm�#`xQRA��y��}=�K��������V������تv3���W�?��8�V�|� Ky+Y�X�Fu�p&���r� m+ݨ����,��HS���H�4��`t}d�v�t.v˚�Wī߁ݗ���4a_�/��x
�	�����g�9��"�5�6ǬN�ȿ(6�!؆��x�>Mzp�u��C�v��(�W ��������S�A���R1N��v�I;�����Ok�hB��j)!k<��%O�w/*�~��6eaY6��*Z�i9|5�Q�x<qBF��6A/�t�bS�y��q���tZD��÷J�p�ꭱi&���J�p`o�G��4h�פ��y3|�C"��'����^&��}��3�o���@Bg�P�+���}�P�^�?mrZTl+)�B�Q��b�x�g�H���d�O#���ʬw
e/�[V��j�'��$��c��S�N)0qR���<!f���prv ���̒t��\��|b��G�hz�� �s}�ߔ x��l�b[d{7L~6�G�>.�V���)Ҕ���N^s���|���	l��c�`��<� �:�} � �EN���|0VA/,+~�t�a2�t��d��h�m�ϲ��(�:Yw[m��֬+�)�q���%�M(|Q_XO�Xt�ޯ���O�\�Ԧ��1)��P�k���G��$�H��e����[Y��L�^g]4���=3�kt8���.�(�(_�7�71��x�1���|Q4y!D��h��ǧ���4*���X8��L�LP �ufN�[>�.	y?"��N�p�$�A�!���ڰ͙���
)%	����DZ���e�?9��J��ˇل��h��m�#�9�o�b�a���x�Pn9���*��S���~y连-F���[�(���/V05;
Sy�s�%���3�0���m)�>�a��\����e��)/W4�Q�/p�^�<S���*�E��4k;$�`� �����h��N�&%g�by[4l?(>b��Xy≪�¨�����;�vDd��ʾ�hP$�Q�^x#�ꪳ��T�(t�LOQ� 77��)���u,5�2�`��H�t����ސC�ih����H22�A�p�ۺ����A�Q����[��A7���H�����ZP��I�Ql��z�\bE����{ I�11c:�ETW1
��csE����M�Q�h�52D��Ɓ���q��n�H�g�ҝ��}K�X �;� q�]����̩��㪪�!�ݼ���dX*pi������9�u>^z1�n�� Xg�&����x���s;�r��\�w#� 5�9������fؗe[�g�I@a��������#���?���p��&(~H�$�����`K�sti-1yH�j�Hiw+:�u@��g����1�jj43����l�>�Ds����N.�F�h��&Q@�V$�I�~���~����6�.���P�_pI ������)��޲���
~�ٲm��Z��aDT�[����ۀ��6
r�\_?հ��%:�J�X��v�k^�y�%B����iu��9 �Tr�ù�h�;-gr�$���嫸�G?R�`RE����XmJ��?�+��_'ok��t�0ш�K���ڎ���#m��.�}_�O!��'��2�}.$�2
#Q��_�o4J�mL�	̛te.eE����E��U��.h@ET����*j<x�g
̿M��Y��<h�\?��5����r^h�&ƆA=p�T�t�����}��'��;��m�U=��PK���t��4W����g��M��ؾ��$�ꆭ?j�f�T�A��[�����v������.�*!��'Kʝ#%�������s�5=���L`�2(����Gk&�A�'$��X��q1Mx��8�z|bpu�]��a�Y=;�]���,�<����<���h+�O�e�Y���P��{�-Ip�.|�i`��}>��|zO��z�"�hEE\��0�� ��0�K�Uz�=.W	�z��n��q���c�Yv�#W���}��*9z]�^E�	���	�iЉ?fن�L�h�����k3y�^l�L�Gj��?�>r����d��J3���J��@�V�4�å�8�qU��S���/e�3���M_p�27�3;�����@1{�(~��A����X��~At�$(�l0dѯDk��D|,��eF}�Nz_̿ң�Z������fiJ%�<9	����p윏&"d;��*���5�g�\��$J�n�ih�f�#m�G��S���K�3�^`���^�N/��e �M`�3�j��|(K90�5��e���)����,!B4����2ݷ��MO�:����|����O�ᐠ������$Xf��T7�Z�dQ�ݜ�L�|�O�9���nQ5r��MJU����$p�a��FF��	KP.�H�&[�yh�\��٦���`�]@j��� /���5����B
��0Qb5n���V|OB`�q����}v�U��2S��I��3��La�7��R0Iu��
��C�$����O��d�o�
��@-��'
:;� H�����#�$� �wE�S�W�O�߄.(���b��=6AP����_�t��4�oݹ�� �1��?Wx���	ְOHRIOL�F�rH���ߵ�$A��6I��f�gG��Z��`��P����2�rÍ�-�7o��e-މ��:`3�ȁ�4)�\���3��2��?MORE
���dw~�tl)� ;��܁g��&�?D3������.��Z�̈���=�ʆ�-+d2�M�<0�CpJ�?C=���M��rA�����ʤ�����	�,"�#�'X� ��X�m���߹Gb-��S����*�qW�FߗF����Z��$bğED�m���f�hhW�ms2���0��QoR[)Ѷ#�w}*�D6�D������Rg�������\9�׼tѽL�m�^(��44S	��B��T&�m�\�&�Kn@L��8?�݃����P���IAc��uI��t��&LU��a��8�/'>��8p���=�k\`KN�DJ3)��n/G��h���5�����G�g�?Q�6���]�-�����=@$�J�L���.>ط3�0�b��V��H������;�mYf[�ϐF�D
-�"�L�p��I?ͦ�H��W��ea�е���7�?V��0�����
�pb���z��E�>'�����Y���g(ܟ�r�ain0aO�b�x�S����Z���E�On
&�v4l�<KF���oN��${P-Y��E"�TN��܁�__���$�$}��H&D�p���(�H/��.�J˾��>��©���B�Cf���w�cEK%j+Ő�L�P��U����%�X(®�k�M��#?Q�6:6wss�~�v,wҮk��S$����w����dL���"|Rۛ0Jw"k��E��"���R���)���{��kz���@W��U�rB���Q&1CĲ@8��:�Z�^l�p�a��'$h��&@U��<�v�Q��Fg5�k�#���P��q�hG��"���Fa��4D�����m?t`���;�o���K�.;[ ����U<`���V�$t!�a��09	��K��b���X���'|�Y�����o�Q�-�)�����.x�w�&k�VOp�S�:�5��L%w�(b��dw��Z���Y2�����4x�ȝt3�쳞�8wjRǺP��=�񒐲�RNk���SN�Z�2?�0�>�]���͉|��j�k&B�Ox�S�bh�Ei�Qɭ�3��Q��X��s��Q�Y��d�M���iL�n�V�UT�TbөB#��n6ٔ�
���ã�yӟ"�U ����R�c�;h������:���E�t��@j"�l7� ��G�g��7'_�1�"	�f��/�O��ը u�j��1�p��LY���q2�5��K�܌����O��3�X:�M����%���ȧ\X���j}e�K?n=�1~�Qb&�un�;����͏�-y�0��?H%���-�ڂR�!�ށ��~�2U^���w�M
����t�ʞ�2����0-�@-��l`a��!����'>�x�ݠ9
c�̨z��G]I�"�=p�kg�b�*�#-��g���]�{5��.#Κ�5Ӱ��u��U�.��!���d6p����Q��݊T�S,�M�G��[��Y��
��Kq,�'�O�|�R��`�����9��IG���	�Ė"}�������i5�����>j��p��;9���x�������.���f	�Y^=Ҿ���.gW�9���|�]]˼�|]w���AE�������XTbh�����:٧����5@�߰q,��g���D��Q�G�8?�Nq�����`���9��Y�'�@Z��k�ʺb��L��-�o-+�/�N�YT�d��)ʹ����&_�6�OK&��؟ۀ�<e/s��uG{��]��,�Es�P��sd����*�r��fٰ�5{ ��\��Q�f�u|}�s�4�c�x�°�oC�&\j�t���X��}�OdaF;6Ꮀ>m2�sAP	N���W�%Wj'AcW7�5qY�j��V��@5F� ��⋨���]A!�8Ҫ)�Q�}x
�W+��8&f��G8�
Ʊ#s�N [ٻH�|��=�=�(Pk��n�v�D�.o�Ҿ�Y�7�G�K�>��[��Z���܍|���Q�qУW
�jS�ɪ�CU`.��c�:z�\�Y&r�nD��Uޕ���_�MN����(Wȅ��tഹJ�1�V(I�2�Pz��>Q}�1-��^�<�?tz���H�>TI~��c�Z�?"��G�Ӹ6�����}�_�7F`Au
���5"-�@��$�is6^�U�q�ͪ�7�p�K������{���䦾��O��Th�{�}��}�
1֥�=V�ZazHf�F����(�ǝ��R�-6m�f�U#v����rt*+����.ڬ�Y��(��{����S���%���q܌%5q�E�&���l�,.м�Jf�MPU蠹錋[���T�X�'"�3;w<�����Ғ��ZR6e�R�
�n��n��M!K�:.�N�K>�;dx3�x�[�[ńtE�5�[�2?�����lA�8�D	d+�,Sn����xk"��-�p���.ԓN���49�[����Pp��l���p<;��rీ!����Ǹf�@ïA �O�����[9��T$bw*�'�A��OYY2Q�#�����)�o��yӛ�*���ӱ�,��� WB���ȩgx������,W� ${�R�g��Ayz#��'N������u�˟%����ZX� �:Q��Ԑ�Q]��/9׭��`�S�+�|�s���g�.b/�J &�({���-?Ne� ��я�X�7.�ƠC w������pI���k}Ц���.��M��3����[6#Z����B~�#�c\�׭�&g�|.s�E/7�zj�u�P���@��7�h�K���H����|�����m�Hm�薚8��n�T��&���f� ��Y&�"��̛��<�9��b�$h�gP���o��s�.ӕz��6Q�h�����/��l�z���8x�i(��ʊϏ�;�@�g�`35���-I[0�� 	��=N =QH�=$����TA��G4����h���؀A����~��|Z~;�"���ܦp)P{|S�L�* ��&I��ɢSW+�4�)f!�)Z�9Ra��mM'�=�9˒?��h���1���vЀ�����q�������G��_a�]��m��0�����g���<m���u�]9֖���NA��:|�$x�і}��m��.� "�A3|�b�	l�{�⓺��@%���O�
�BXor�6<���� q���"��%����	��7+�Ŕ�+�R<��nL[�c�Q~�*f�1@���\$#-bvK6C�,;��2���h\ 3��&Q$�F���ѻ�9��0T�,�`8є!U6?��
ZMy��#L�Mȏr4X��,v�.g�c�Bh�Vv�����=)��P<�$*�%#-�-¼���DNÐ�O��w���Կ]��Ԓ#x�	�Ϝൔ��by�I8�PJ��]A�o�q {�G#���o����|EJ(B����U�;��S��e�R
��<�?�
�6oNկ��>WlϏ<;�á���	���yoh��(�l����q�*O�>�_��~��	�pz���3R	����Cɍ���#^��D_H�*mTwm�Y�I@�\o��]�B^��`� EG�-[�\Ta{jM�#�[	���Fp���$���A�#�!�_�����NA�?���	�Ao˦���&T�W�|-~��w����?�C��ؙp��a2_k��c ��@�A��\t�ՃȨ�u�9My���Z�FKY@#���ۊ���G�C�1^��7Nf�+Ś<08H�\ �C�9g��g�4m�
��,�k� ��a}��c5e3ˡ��K��Txv{v���`��p: �Ϫ�K��Q��ʢr��
F�vb��Ν��-U�z�i	,�2dt�ǈ�?����ʍЉdz:�&~�.7vx~�B���<�*��N�񱸹�Z� �E��Kg��<�!/d&��:����kuk�_��I��@�=h��K���b_&e�P��P��.r�z|���H+�s�!�P��|�">�q�
�̑�����3�j�?!i���f������[�X;Ό�ƅB_�Zj�<a"S���4��-c�X�鹦UeT�VA2*պF<*�]�񒾎�C!�F}q�f��b�О��d�{g���0Yf���1�s�������'f���>6�J,��� q�7��#�X��O4VX4�C�q�������:P�A��.�%:B�v��������;x�X�Rz\�V'�6
E�������o�o]�%)w�
�H�(�������)g��J��P"#�ͩ�ϛ�5ܺ\i�le��}������FcSB6��D���k�l'v������9=��
�?So��E�1޿o��h/�&�&�P��r>jT(7��2�
k͖����^��W��ܸ(㩴n�F��;mK�/D���?�R<��"y gu�c���-Y�@p��Ա�uN�.1H5��z ĝ��h�R�Ǻ�^~J�>D:}'`��x���@�7�t��a��S���>���!���@#�E/�d�}3��e�T�"04�H;���ۆx�Θ���؁����Ɩ�5�m��.�8�*G��%(�)rE��7x��))�?/�3ɑ6ǡ4�ѣ��2J� �˻�6u�d�M)�+}L��`��t�njO���-�lQ77O���e1�x�R����H�Z�����;JUx��n9�eo�b��D�x��U��:�->�bsp�ƿ
�ߪ�,���LI[C-�8=" .a�=:�?i�sv�6��ve���'Q��G��F�����1�pO��kG��	���[����3�&F��<,�r�6����,J�͑	U����A�kj�0	A	5Aܔ;��Oؚ��^�G���M�`�P�i�j{h�>}��s�l����c?��^�E �*���eO:E�8�&ߞ2�I!lw�����H0�E�*�h[<o�6� *m�Uq��
�=�}d�8l�;�Rz��&;_�Z���Z*o4�H+7w��L��h;��cTV&�f�y��N��@�B7e��ǳ�w�pmq�W�,|����^�!�Q�V�g�S�S��0�?�� �đ����U\i�XE�Pk��7�ß�V͎�P�������1�D�+��f���������RAwgW�����V�|O҉ZSg�������c� ���֫��p��C,A�v!�1=����53����sA�[h�<2�DiR�ӧ[$F4�������f����m<��Š-����P�rXô%�Q�q�D��:z�`�<jz��3C�@C@'��2ƙ^���sg�VwơC"�M��R,�9#�Q�TM��1����Dl��]\Q%�np��w�.��sU�Q��!J]y�O\���hzFAǒ�7'��m�I���S�^#>���<���x��W�yUE�f`Ѥ2`���oZ��a�i���pU���
gX�`�>�n�Nr��%V����`3�3�%�9��`���;�M���$�h)Y������������*J��nOq�Y>��.tw��4RJ͑ #�v��՗���6�ച�HD�nl.4��� a}�
�QF�h�~��I�S`x��O\�2anؠs,��ߙ� ��{�3p`����}�o�=)5~���Ԃ> Ӟ:�Lх#o(M�D}݌����x���C���M��׿��9\�Ӷ�"�57��皈�}�cT-
#&�;�U��p��A?v��G�T9!��gZ�e��o(��������8��f��)I#�������d��"���c�����9�hP2]Q�Оe�ɖ�\� x��f��˨L��Ȣ��� 0�9\;����x�b�&�=��b�����5燵 �L�J��a�o��D,PJ��A��o�o#�ٔb|�"j�Y��z���[ڡn��Y�G`�M�ޛe�6����cM�:ho+�jhV琘����%�V���q��J�zY�A�|�!|�s3̔�/��5}�{�y�2�;&m�{:@eɥ�}��(�M���=��08؇�WJ�+������B�G��5�cD��=j7��������,��K��,$�0�-�ޙ5��T�h�W��^��
'j��&��2�4�&�l�4�����;'�>p��5+�4$��	��l%���|���?�1�t@q:�o����=~ɾ�.�Xu�Z,��E�/�8���Ӝ«��6#'ꨕ�&'q�AA��hl5M�M���b��(�"^x�o�WٳvW�6�#�&q���Z^6P»�y䋋�ef"�xrN��F�ԣ3�@��� ���y$���mKi�`~�ޯ�So������: ´I���f-�
P��C@�#o�Sv+���+�j�Y�dg8g:,)w0�|�s�j�P�H�
g���J���CHwR���k��mT�D �~�fK�D"%�쉜d�l��@ޖ�S���!�ɠ�|�D����_*���aS+��m���}��t�7�a��pN���N������"0��ypp_�o��5��ܛ��RXM��꜖�6�k���r9�[�
��H��:��АfVt.�����R��,�%c�-b����z�K�� ��z�lG�5H: zw��%µ���Y�S�e�XN��
I{��	�@��048Dj/�iP�e5'��F�ߙRa���>��+�%4�ݎ��#b�<��:DO;əX�xb�S��Pr�ʗK�|<�\�R� ������^pCk�Q��Cѻl���|c/���/�~���ϩs{��2E�WE`�<S�P2�%�Tna!%0i�a83�j�����#�|�'�pt�uQ3>��"�1��b��R$䚆J�R5r� �b{�G-�}����U������ ���D��c4�.�<�F�q�U�n�x`�&��S�&��sBH��Z䴋�Ŷt�۳X�ތ�~���=�KAR� �,���n2f�AG+3<�5)�1�=~YB��4ͥ+��`��xO�m]	�sQ�& �9�FvZ�6���gL�P3�-�g�~�	}�]��?�Ό#�ECNZ5�= �@�*��u�e[�ņ��(uze^�G轫��Hn��s� 1|������A�TX��	Z��ynG��.�:�я�������ӎ��?P�,l�GhYHl�c?Xw_�s���Ͼ]S�7p��	$��=�� �����mA�?��i��R��yOT]3���(8U5�Ql]��<b���#-���Z0ul��K|K������� o�Z�W'���I)�{�IHD�T&�u+�_�A;T}P��сU-��e������2�Q0�`�e�Bs�e�{�n�[�
=��kF�DZ=���C�(�������9���6	���_��NP��^Iџpz�3�iuF6�LO���8�6��p�|�.���%�>ʻ���c� ��[�>����� �K20'�ɯ �DFwu��d}��6O^<Ԯ|C��h߅m����@9���DA���_�V���|��E��aߘP �����.� ��2�.C�fz[�(ۜ�������o<`��P4�j��7@V���>\O��Ĥk
N���W�=��l�N���� �Y��E�8H=�s*&W/cϡ|p}���S���<�eiG79=�~?�'���\�ƿJMu��|��J� ��&��
f�-����tQ�"�,���Y��K��H����6��	��Qz�� {�����#Նۯ�~6��=���ݰ`�i�1��˼Om_�F�
��r�wZ��=��D �t8p"2}�Q��g:��QW��k��h�9xy�@M��]�"� ��q��u��Y�Ė��}�I#�SȦx�:'��!�xǬ��vc����n��a�U�}N�J�}e���J��a���tϡ��H_X�|����K<�Bt(AG�֘F͊��Ex�a�]:��f�M�ΰMd�d�0��q���?�b�����^�#A[�-�[�zGi�,�͇�񳠬li�M��`����`�ñ��q(�^}��XL@��h��eF�M��y^*���}�%u�G����ϚZF�CK&�qL�.js)o��o��_�IM��]��]!Ib(�~�2��{�\c"v�_P7+�p�>��y�sSa�z�����^[� �T����Ƨ�yNoE�t���	��V)̀��Q,��Ϳ�`�w#p�y9�C�u'����W���o���fcr��	���1�:��M�5�))�ʉR餛�Q�`�ޠs�B�t*@��+2��+�V�yNʙQ5خ�����(�s-���g�b�|��`�/	�g��4_��͆i�g#bJLB��[�Z�xB謹�<�"s��#0\#���#4���&i`��?�%����m`]f))�َi��H�U�!"0a�r��R�x�i�1���ZQ7����Y3�L�F�Q������w���"9��0V[��>ޠ��o�s�<�EF;}bΰ��=CH];A���7[d�6��PG=��;.�J��P' 2�G�`�S�Zs�ǿ�~��Vr{�v<lw`�����*O^�˺�f�)�~�����s&O`�H5p���ui�$d���Zæ�Aj������=�?��Hb���^���������ʽq�T�u��)w+��᎘�=�e�%�Ĩ�U 芦1㸿�?!�	Eze�i�$츦�-�a4�?e��&���u�G=/�(SNb�����BO;]�+6_R�==+;���]ꇢ�`���i~N�'��t��e��<S�2y�QۖH�M�r��ȥRy�otD��z7�� ���G�Q���m(R95���8�l����{~~1�ԫY�>{������f"�iR�7�=�����M�=�`Bn�%[�A^`���VbmG(�H���I2űd��.����wΡ��;�1����Ƴ�ȡ�p[Ňt+1Si�b~%�B��$�ݻg+�ϸ1(���G���\�
�Q���]bQ(�O�v8�Yk�M����������)��}k_N��y�������]k�f�=���yoZ���9ćj�mk櫃5,�l�vH�	�O�d�En7''/��ev�iv`*��{��U7]���s=���nZ�*e�n����v��^v1G{{h����4���<�ȶ��5�iIF��%;P(���SANY �4\����Ľ���l,�Mh��OӢo��~��Rh��y������܁F����	��Oƛ��xf�=�1����R;�D-��#�C�
�mȿ���:կa%�Z��>c(�1���W�������2+� �@P`��M�������atg����L�Յ��c��~�CTa'��9̂@�,�O�B>@���̷!u����=oj�|��s���s���ܥ{��}�z".��^m7�Y�=��p�G� ���Q�!��J�8��`��tN���]3m���L���(1q�G��HJEQ�6Gq�y�Rt������w\���=���̊�g�o����wh���Ƹ�����	�\�#a"�$�<���h�5oJ��Ww1�x��m���'�G{�}�hx^�� �; �\0?�:�ߣ��]��SL@mD�'�����Dr߲$��iO���J'��L�В
�ŏ��M�&øl�KwH�1��/����2��(ى���B ���\b�K��>��8ޥ�������Ђw��L�\����x��
t` Ma���u̒B+��3D�Wł`.�BX�����|6c[�R+�v�`۪��)�<ZnRC�cP��B꫙u!ܰ��um�C�V�&�gT�X��wϓ������׸�~�UՃ%mM�ӧ�q�.k,iyc���5���Oۦ��$���q����.gO�HŤ3\O���11��ӧ��"~�+�eQ��:�ͻu��H��/H�ژb�ö2���Cb�T�9J"�g�2�j������m9_a�*�B��)� uh�o�Ő��-j}�⦶1n�vz�MG��ЪO%l;v�_t�����Sz���-y3��XTu'���&A',K�����U'�*��8"�^���#�7S��������)J�h�K�C��]��ǳ�e�P�}H���;�!Ut�Is�I�F�7D�Hc�Q����'�ѻ�f�?�Ds�,���d�����G����2T6C���t���|�YV:5`�4�i$��qu�}�;l1��1�~5�0"R'r�a�rVC'dl{�(���5�ՙGE��F�;��9g�Ħ�;0k���:� �+��y�v�%�3	����ɼf52	��O!6�t�Xn2<��+a���F�	*7cZk���Q.J.��j\d�/z�Ia�c��L/�3
"��� �_�qӲ^��
p��b'Ҳ����r�S�`Կ���BQu�\�K%�ħiK^Q?O�Y�K0�GQ�f�E}ݗ`[bo��/�	��6�eBbt���h��Jd���`]��H�W�吉�E�w���Y��)7�m���I���!u�������5�y_
`�ox*8������8-H�����A$r#�KQ�o�(�U�,��Y:@?�������Dw>��C��$�o��	{"[��C9Ӊ/x��R�}
�7̾���Z��?�$�G0Xns�N�P�ˀ)�O�E���N����Eqx(�hδ@�,T%?���K�o�oA)�L�t�T*����V�| ��jE[�`. ˔��mN��̦:�ԟ���)��b��w��[\��0��^j�փ�Gk��V{�������Je�3�h���1��7};ncF�ݏ;�����1e�*�GqkP����ퟒ���h�0���q�	�ߠ�qR!.��m���ً%#��>�n�k� |h#n���%3[�N�s�lE��R�홎��+��앪X��.eZw�K[�A�� \��u���E���h�8IU��#~��Pa��"�/��9�*�ܴ��(Yh	4b���:�RN��x� o��T���J�hx~�-��ł�f\vi�T���D{ 1vV��E�VD�rEx%�6�*�Vzp0�
�O�0��_nh��BS���JJZ�.B����8`%�'��o�;�c/Y)D�MrhWA�W���܌l�0�>���9��G��u89�3�A*�i��)jZχ�=�'���7�!��1J���FI̎>1/�z5�}I8�+���6
\�
�;V ֭ڮk7�l���ݽ�8W�~h���7�H��"1��b�}?�G>$��(?��pBo]�0����1�ɿ��Ss�V�Q�����#�0�YL�g�Wۿ�Z�= ̙FS��#�Q�����W|� �w�~�*��5(��ĳ�W`�o�R8"����s���1�s�9��?ۥs<�i	����gJ3��I�Ǜ��.�[���p�?-�b1C!3���1
@-�5TW��|��4t�H�(�W�������_����M"*�g��.PR���I$�ge�g+�v�E�n�-C���8�O BS-޶g�^�A�;M��$���4�	���3��%f�(���Ӻ�C�f�������U x�
,%�>J�K֔w�%DMoA(��W4��IoCu��? Qإ�Š&6�eן�R.c�Mr#,�d�_pf~P88jԹ� �6/�Q6���I@$�Rlo�6��f!�%j{l�R֠��)H�I�Q�����=�9a�&���B�Jy �}KIO�'�)���L`�W���2�{�U���n�*
���9�T��"{E%�Q���@P��.t��Τ��g���*H��[��;��GM�V��H����Uِ�L
z����$@9Sl�ӐX��8���4<�{���[=����n���Ov9���l�:^��2Nu�C����s��/
�=r+�^��S\M�����҅"7��0v��Q�I[Gk�~X}|_��b7H
����ڲ��D�V	lb���me��iG�hIp[��>���!Di���w��ϢٝX2��0x�Q��)����O�b����&+���F�1P����4��ǧIlI�?
�KN�KE5�MD@t���6\5���,K���v���qEN�N"��N��G_�����ͻs-@�@=��-�D٦E���D媿�z'C�u.箟#~��(��_۾\ �u��{�ͯ�q���q2dЀ�q ���+��No�MMߏ�bn�(�(;g9�ǣ��� IA#5�����W�قk��	��@+�����R)�S�iW>�{|4�2�&�Su!��d:Z�<@���-?2����V�0=~�[~�/؆���e�s�0|������P��G�'R��4��!��D4���h^�<�V�O&Py��E/t�+6���y��P�ZxP<L�d��T5�s�wl�cͭ��U��ġfo3�$��f�o����_���&V��z�]��u���y�U-Ab5��c�M�Ҡ�El�C��ԙ��G�mPI�v�(� O=�WJҁ���l����Z�K��eGx-�܈$�j�T���ԙ���0����屘 Y�i�
��)�
�U��/>@����_��>���.P.f4_+A���{6 ���r��u�|YL��ל��I��l���-�p�n���ԉ1��=��r�9��*e5n�K
��碁m��̽P8
��]L�q��*�I^7Br�Q��7�Oi�(2��]ª"�
���RiǋU�˿�h�	�
>��njo|Z�ԉ��2�ڃ"p8#�y�Ȓ��Fd֊J�s�-9H�})f(pv&q�e�Y
����w�-\L*g��G��y�R�V���>�8��,\/	.�k���2�&78�@]Eo�-gC)'I-�>�UGw�z�F�\��[�G�J:�v�d
b#��Z-�!�����������lR�.8�k�&Z�x�̨������Uׁ�b����α���s�V�j�.4*PplU�h�e?���H���L�,c6�F����-� �d;�	#/�3��r��x���RT����дũ
_��Je�C9��@�I9	*K��U_dl�+�i�i�J^�"�	ŵ{����I{�Q@{7< k�yl)U�(���H=��wb�e?���D��s�vG����'_6s�e~!H��D�n�d�z��
���6@�g~Sr|��pu��$)���R�m�Z��g�\Xy3��=o;U�����i�<*��{`�?�9��a��Pޛ�;5��{��w���*S՟��n�BT��kH��OϚBh�]�{[�~1�A�a:GK �e�/��j�"�\$�O��Rk�S�.�θŶ�HS��8D^��f�yS�:�P4l���M�5����p8W�B���>�h�5�Z^� ���߷�ŧ(\�K�t�Ȧq�k}��K�LӞL<�I��~��B����]�Q��\�|�����fN�q�v*RЈ͏ؓ�����>hn�N&�_L�����=oԮ��]jm���߇Oӫ�l���zW����.�d��#��CG;�(k"P�E���¨?*�$j�,��q�g�����<(CX���x`�z�?��q�	�$s�.&�2m|-~���>��mӱ���uC��Kw��A��¨� W��/���Z���%�����L.؝��>�s����Ѷ?	l%k�f!��H�d����,��a�۬u]�E%�J�m�ڙ��x�"�m.��D�i�\i���,���t��$���9:�^[mCc�4A���u��̺!�_b��(�6��� I<�����QI9�[lp(�R�&����$lj�YP_[D�����E�'���Sn�@|q�1qT�"�T� �$P�nS1ͽ�h��}����m�x!�i؆4���߄/�J\N:~>X�Ԁxl�v��d���*D��8�"�����7�K邶�P.zŢ�����0ú���p���+Be:�CQ:m��i��u�	���0J�8��g�.kSu�X�-&W�3|^h��x`6�߹�tS��ߓ��7bcv޻��:�1/=y�tA�����S��kh��������򉱾wx�#E��?>}gŀzm���ڲ�������#�F���3X�=y�+w㷦�~���w�t�4�ES�	��?Ϣ&�'/N�f��i ���B��q�vv���W��:f�?��}��~ݽ2|�^�l�G�n�/�z���`;����^T���^g;������
�N�7�X����Oq�->����e<��>��!�|.1��Q2��}�6��h0�dR�ʴT}fc����Z���#�=pa�^�8vt@�G0�4��`)��� �6C�n,M�0#��ڥ��UOu��S��Zo�DY�]+?���P���=�J�Ԁ��U�h��V�g�(^�e����2a.�	�j�j��¬�m�P�G��S��Y��|����	F��x�0�7VnԚ��aS���;�H���u���2���	��V�BO|�QT����)�z���̈����zz����
Q�E��f��-�c�H���^&�O�caU��G�.=FJ�l��uV��i"��"�aN����z�=�x�}X�7�1��Rk�e!̥�P�l>�:!���њ-���5V��D@B i�I�QF�͎�SUE̘,�;�Uvb��-^����p\)q����{��G|+4a ��و�ԍ�v�K�8&8��X�O4�\�4�kH�`�Wn���&�&9�	
��M�!�琙��̒H�M5���q�F=zr2@݆�����d����}�8Z�X��%�+&�x�fQ+p*JI97�Q�����I�e�PR�V{4����fUo�o���!���Bt^�}L�O�����ђo=	����'�z�`cHFmdde�����``OS��׈�ԩ���0��Ct��Іj��&�����Ee*j��l�s�v�__X��M͟��`�4�2�rv{mr�B9Y�J_�c�i?�� ~9���f1���tqUd�j@�緹�|��*=i�iB�Ek���֏Sq�� �贈Gd�ɩ܂W.v�q���?�Wy�!��'�E�6k>y��+�s��y�e��Ē��0{���m�^�qg6�yg�Y�JI/а���&��2l7A��堨�����"�RC?��8��ϻ�����im!�Da>�p���?"�f�%}b�(ۻ{&�#('��=�IާbϾF��6�4������4�����qQ}l��\b�a'�#GO�,�q�ca���H>༲e&+8 � �j1!��R"Ɯw����%�v�U�z�e�ǣxJo���*����Qs��dV�rH9FƩ��Ar]�0�n���|}s|&�d�#F8�0x}/���Cc(��/fDt����w�2v�s�?З��е�BD��O�=�\�O��k�"	���)7EN�Z �@�BM ��y���v�q�m�N崹���E4<��!�������(ǋ �@<�{�������� �1ܞzhn����!"�Y�-<�ŕ��m&{Z���]�4�ϻ�b~��,11e\2j�Clʽ;�j�&�����j�Ss>�����=�'��s�U�E'��'������Dt��H_r���E}�^���������x��?U�����6��҅�W�����*B &fG���EeH�#~�Py� iH������y�y�L�j��N�4��"���.�\�G��뻀��#���h�7{5��v8Q0E�˪��p�Z*GƔ�;f�]wU�I15i���1_����uJ�r��\
��)����|x|v,!x�}IhJ���w��%��O�ȝh��>o��A�������+Ԅx�L��t�4g��"B���X���Z�qT�C}7!����� �3�l����n*'_%�a{P_��-B��b1��*كT
"r$�W��^���^�Q�;���h�MYU��F�t7N����p7J��Gq�{�ւ ^*��,�X�,��6�Yj�/l��R�3SĬkGāPo�M��iۆ�s��0[���@�ġ����?U뾵��H�]�e�YUވ�S�&��:� [H/�|� �h� ���O,"�.7g!�(fT�
`Ĵy�)�y�7���RyIv�}%���u{m�\ߝ�-�.3�#=k8�<�xV�&R';Y⾞Iv{�cVRg�V�k�)�|�dQ��m��j%�+D�+X�r�"�O�.�9�9�M�g<����M7�d_y�7'�Qٷ�p�u�7�G�[��뛷Y2Ȓ�}L��<3����{�b�D�F%��\�/:�/�M)gSI�)�-=���}��s����	��fJ�6�dr�Ѳ6���-��}����Q���)iZi�`ĳ�$	/Yݷ}��;^�_?��\^}۠��Z���c����a��}��I��ɚ�	����@�^���C���Bt�/Q����J��B����C$9�b1b���4��!}�������]��E��?��W�j&��E*�ҥ9�T<.��@�#
��ʡ� �qZ�XM �$������?N�͵5��.��;���5��"��S<NA\�'����1�&��5�
:���ps�"��4F��ۨp�H)M�ֻJާP�K���i��:��y�[�f���,�T�>b.��4	J�g�s!�8�ׯ��J��߄���V���������L�sT�9�ס���R����}o&�lz󫓽��+o{�h❕�
��Q'�x��e(ϭ���$�!��3ŏ&��M�b0���*\l�W[�L�g��
�6�����!g^�Ȅ�NS�ui����^O��#/�?S��y�/߼�p�^!�+ft�ק�3C��H�#��S�H%�3"�D��2��[f��1'���3� �ב	2[��V���]�ջJ�S�B��Ȋ�'���q�)%��TP=��J������1wK��ۡM	D5Q��EV� ��w�b=���Z�C�x
��t�����\��Ȯ㗆rS?es�#m�ĕ&�����h���hŪ+��f~�� �/�V���ӂ�Q�hyv*|�P��9Maw�v8���b4�h�Mv����+"�3�Qor3n�Ϛy���5�=9)j|�Q�������A���.�V)eL�AA�G �#�tؾ�{��.hތۋv��&r&�ʼ�n{��;,m��,\���
��'85��G>$hq�$�
< 
��5�k��<+���49�:�?q���$3.莾X��WƄ;�9u��~2I��|����as��\���8{1�'��zQ2;d�=�|�7	�w�wD)ն�룗K���A-2Ӽ>��v6r�Y��/
���`�r{�2F�P{P�ͥf��[4!k���:x|3G�48&1%Q^ѱ�@�ީ�2�T�����Y���@�0�KM(��NfP �F�~���߭��@��[ 8�OO�O쯃���1(Ig��Eަ����T�]��������s/�z��|4�\�t�?�H��&ئ��9���W	R�-.�+�jLJ�1��ɩ��n���mo��Y|�f���i��=/��6����M���I�f$)�׋ʕ :$��P��������EF;�x`�;l+GRJ�_ʹF��%�d�H�\A���6�TL��f-@Xh���X����0��T*�V��^�ņ�}ʔ��*��L������P�&�x"fQ�]�M�lO-]����B�Ƚ�µʿEޣ��~&OWރxa���v�
�������*䛼x�(T'���L-e����d�e������O{m��$�{W�*8�oIй��'F)�hY�'�$mri�|8o�8���kn�%�y�V�'��B��"���#WY���JP��K
��=M8?�\0T="eb�}1���gth7c;)�洏��X�҄g;+�:ר�FCP�V+l�x\Ӡ�p�A�S^:��T�m���y/v��6��f�C��u��
�Jt�zc%?�3Bb�2^�a��wnٚ�
9AI��1�Z��������D$c�&v7��ӽ�A�oˣ��7���4�v@T��K\�+���3�5)��'�ںE+t��u�
_�"�}d�崌�F|ï?G�tC�D�Q���U'� �t�����ƾH@� !i�����<o�3���|S�ğc���o�5~���0-���J5�A�ґ�Ueo*/b`�<�_��N�,srX���	9�Pw����e�9��{GFQ�|FM$G��)x"�k�1�	!v�ɘ��o��V��"i�g!�T�ܳ��V�a�	�H�4:����z@�n������.)�g�w%<��{�wƶ�1�O+?�C=>	n�Z��s��YM�%�c��G����&|�l���L�K��8��v*�����$7r���]���X1�賝z}fj���ίz皁�c3�p�{.�sj'g��Ҁ`��23i���D'���I2mE��D<��JC���3k�-~p�J�&��=5�
յu|{H��H��O�3�ذ&����08����D��F�	f�1��5��O��S�͋T�P��vt���7zȐa�e!��ʦ�aS��q�W������ϻ��VG����T�na����P��8A�[��S�t����%�(t�l5CL6�/ �=�1d9	����n�j
S��T}l�W���b���w�]� �q$�N�$lzgC��R��^Cc�9�a��$�36���z��c��P�-U5c���zi�cPo�
]W�5�zw��C�c�q ����h�MO:܅:�z��ғ������FU������Au;)��@��I�l��^�׌�x�Y�P�C��?�w`"n=iQ�1�x�������U��0���%�0|����=��;0�}��֙hX�^2�7��[�
c�Pb��Ֆ�N���po�jH?�-�~������7�==�re�njE$=Q�@�{:z=��#�;Y�Z/w��%�wyT�G�(�/�pi�;�#�>����L�ӗO�����@G�)���9�����nF�nn����ed���e�8��Əu1�_r��Cr���c�Ǧ+��y;�VW�����Յ�9�ȿ���{b^e����K�{��5q��f�5ɬ7��?�,�V��r4ʸ���^~>r�p��0���c�&F�9����LY��Q|!�$�r�B�Ў ߏ�2���|u:��
 �k�9Ѓ04't�	f)�]�@��azY�"B�$�i��.�x��
�T ',B0���/g_-X����z/Y���t�2�sR�(M+AxΚ1PVm%��k��(S�,t�p
Ϣ,�-���F��"�XN����_oO��3wq ���-�=�z�6�t*�s�d1� ��tHֶ�\hB��(����v2y�T���d➜!�D�YU�3�c��V{~*��V�������`H]�!�ix�<�$��s��ێ #zb��]��������q�h?����'N�`�I%*Cv*O�uT�M/��>M'���Я�f�@[{���h�^�~~�p$|�ݥD'�d�;�|���m5Uqw� r]I ��MS ���R��jgw[%]���[UJ�#�}u����-;Q(T���1�x��m�Q��=T\���H�st����R�)��&�ؿ�O�"��fd���m�*	�9��*���vHܬ1���;�~}B�B��p4;�6F�[�ٵG���pV�_*���;�K�9t���oa���g��]ruY��3�Y�^����Uݯk2�yǅg��F7J����ѥ�x�����w�aH��9�k�v	W"EV���m��(�pNΪ3�W:�i��/BҌ_��c��Ap�_��յA>y;��L�*w���o
��@	�H�ms:�z���X�>��A[��$������/�#�V�q�������2h�����"Q|��%kcA�&m�׍�g|'X�ϊٖ�d�������<b��5׬����|�e���̮U5��{�'tW&�y������#��)_��[�֮M�Sy7�C'����:�Ӕ�z	��2�:���=b�]t8�G������Z	�g�y�ē���6f���bL��B���gs`�r�oa�
�^��HᢢI��7$.Ͽ��E�a�����-��K�4��ߤ{�E )�t�ixbZ�"��@P|w�������[�p���igpR�޼����-�j�M��9�?����uy��?���]e�
{�ٍj.�6�u~��d�O�蒚% N�.��̧���OMHf���9]wF��A��M����`�ǹ���A�r-��0ү�e�=��0Y3��E��p݌.xf�g�'�Z�FȺ�<F���XE����v�]��	ǲՅ~�����?�Btg+�:�Z��,|w|'Ӿ��n�~T��>$�t�,�՚��d���9;�<)�*!nU�ߧ�#Q�J�=a��1��88�ç���f� ���VR��va]F�#qˆ���Y2ȉ�F_��=�k���q��y?E~x.U=&T?gWGq
c%}nʦ�c����{��8�YI���c�Bà-�~�CV>����gvE1YD����s0���F�Ф�G�^[�(y|h�'Q�����B�4O/cWs#_�S;�)���]�z�	���"B��7�MVp�/��uY���Q)X���a��'[T��'�7����GX%�8Y�靈���n�Jf���
M�Z<����F1DSjp��@$�U���ݲ��l�<�8�r)���G�0$�\2ڎ�tǙ	�M��,�)����Z���Bޞ� ��M#�u���B2;�����'<Y?�����̢�;�w�V1-���R�����L�����(��E��m�j�-Z��5z:y����@��(kܥ�Wpӹ��2��9��.��Z�雌�k:�$㓟	L�گ�}����X+��숱�B��h�̄��g��:>kB�l�}$伾z|���b0�! ʛ����Ս��5.�U�E:P͂�jG�2��l�޾} ���DE`7i��m yð��VZK��2RN7��M��p G8��OTB):<̱�|��	��D^:78�yKrvm���
<�rD/ �V˿���B��\�p-��Ȯ���e.X� ҙ�*P��mX���n��g��_�6.>+ ŧͳ��̐_M�4bj���@v�L�s���K�E�Ŝ��� ,'.�I|o�	Wf%��:Ε|RE�:���-��-	��KU7k,��bK?hyx-p������Ė�"���[�yi�@y�U0 �U2�,us{c��}��HTL�&�%�;�
��γv\�4;ɒ@2SWOn�*y�VrQ�v��/U8tB2�<h}G}�Le o���������uw�g��%}]���ҐNX#?{:�1�`���∎K.�_���Z���krH��1R���|tQBՉ�+��TU#�Փc6��)����I������ŉ�N��;ؘ�����aDc��R�j���<x.PXƘcf\4���dK��z���,U@�3�p�T��O�[L����@����Y�.�:�Ϗc �`NN�@��-*��ceϛb�k�r�ϋ"�s���>0 �>�S�f��2�SR�Ba���L���-[Z��a%-Fi��D�P*�w6�c1���'7j��Wע��7���#����âqo�Ҥ��h���g�i�sݲ^��w�r����aR*&�
���w5#���d��k$'Y`����2�d�9�ShS~���zIܮ����Dz�)�\���R��`��ڎ$��Pq$ڿ����y�c�(oq���L�v�� ػͧ�(����
�6�\�	Jl�U��"t�G�톕x}� ږ���m�C(��'�:�n��	B�)���qM@��$ ��)��\���30�G^K�� �޸TE�>����-�tĲ�'���n-�&�J\�5.i�&�J�	Ʌ�M7�1�B�g�fm����`��R�D�	�{t.��‴�©}-�a�)d9+���ą|�:�kv ��ܽ�������m���5aub�UW�xC'������*m7Z��_�� I(+7�d=��e`䟞oU�{Y��g�j���֬�{��-nwC�ۚ�|P��u�*���GsG����J?X]	r�ؑ>E�/���@�i`�d�azi��U�HFED����f���4r�7"��7�BQ����w����QD>>�u7��}2��&�L8��L������;M�E�Bi�k����NF�n�(��-@ ��vc!I;u���j�a�OVP� '��0\�p���uČD���U�C��n�'��3�P4;~ʱ�㤪�l!��A�C3����:�G��M"�����[��(�J`(TFS`%z����b��ߎɫ0I�7zG�dPdjˈCٚ`�	L�&��C��Ur��oRK)=T2�B����]�a��o�|1]i�z��)gi�K�i^q�X��K��|j� D�W�4�5͑?��e��L�seI���#G�O�3 |(��<�>f�?��_5����ȸ���tw">�#���.�9�vYz�Jdj��YJp�9���p�j�:BV��ۿ=�Y�-��BCb%�Y�j��sҕ��{-*;��/��GVO�r�����ūf�6P��5� ��z�=
FJ��u���LTTGϟ�Y#�a��F̕����5���_Z����ڧgX�Д�W��aY{G_C)bA�宜t��bh��LyX�~����z!"��]�|�f�`�m����y�n�Ax,���1`�<h*��F0ݰ[rP�Ҫ��������5k��Ǻ�o�d�D_�g�%d�佟1����,��\��h��'K�<��s~e�8�c�e �u�#�[�|�4i�W.;q��&���R��UYL�r]��$"�;&��(Y�mD���q2 G濿�6������˒!����g�h���ZC�`�TD�y�ȼ���3��^,�h���&�4�D�l|U�X=ԧ|�X�l�������m �mv'ǩ �),b��sv����W#zHY�X6�o� y8^�K���`�}ux�{�F�rRD�*�O�<vOtx���_�|�7ke�w�a�ig�rt���\O].7�$�u5��Q�	��Nz��G��5"������oT�2���#`�z�i��H�gG��IWL0��ߡ��'~nO�%�|��x�-K�/���A��gyPL�'�;B����ro�]���#�<=mMˮG U|`M;�ȌK�F����2��6��k@A����������E��������t���Տ�=!����#&�^ud� �c���+��]�Aa��䊲�ز�2�5�g�yU��
"%=�r�E��&b�5Z�}z�`�|	-tov��-Ah�1��L�SG?��t'-LͰӗ�(}��¢����Tٸy \^�[<qC�<o�Q~�5,�##��L�'U׸���3+ L��9^����KK�$�x�ϟ잞Z�y 2Mo���i�Dҏ��̾���q��Cw�n.|C���{�i�|咷�%P�M�=ʔXf1P�u����s��Pî���P(<��_}`˱{n�l�,� �1��k�g�Rp^��x$��:�d;v�;�/�(*a	�2-�# 8��R/�y(�/ܛ�[�X�E�/��Kt#ͻ���f���D*T�w=KR�L�lZ����!���m5#�z�'�4�-�~[�x�U���d��[��5À���~ Aie=E�6�I�k�m"$��\p)�f֒�d�j��@�"Y["2(�3t�щ�����CQfTg��ꏋZ��M��F�J͒� LfT��.��xl���g4�
,��F���x�4�`ǟ�ѽV�1��GM�,���Xd8D��Y��)l�Ƅ�Tͬ�$^��Nj*5��:�}ҞY摶���5s;"0Xc�	g�R�b���8�el<i;��Μ��)�j9t;Ky�>�?@W�d��Y���ҧ�U��������on��;[�\y8�w�]�+d��Z#FX ����C� 4�@߼����҇wdd4ǫ_\R�$Ժ������O#ލ,���=��Z�K
`���Q�o����#PB�Oy�p�o~=��ы������~?�����%�"��W�R�[��M�O/+���}+��hy(�^���[Krx#�W���n>�^��1�O�㪵����j!Ir���H�����Ч�����
w��7�ޕrc���b�4���O���~B߬��sh'���E&4\�=�W��H�݆nZ���IF^1��?�W�������L�/��7�y>�V��Z|R��`���]�>��Lɭ���j
���n�ScM�����	c�__��$u�U�k
�[qi�9���"�[� H�5�x5�ptɆQ�GSX�d��K?��])?���44A�UW��p�K���G��l!]�������`��$�|����*H�""�^%sB���h�����K��Y�R�P\�s��*�u��s_
kR��<T|%�hTh�aˑ>(�7)�I��*(��m��T�̰ҟ�ct"���c�׫2IZJ�A��!��/���p��{�sy����ʿ����� &��V�F�[7�	���[�'ח�Q�x�ʂ'���X�)��C��_.-Z��h��,����������ݢ�6����4�d���v�RF��Df����w7�d�9�-�s�����C��?���Hw�L�P߁���,�"����9[�Y`��_<O�������,%���@c�*�D�?��gVqob�6�Z|���N���xd~a3i%�'�@0�d1$�wR�^�Sy�q2sr�j�%i-x�v��IV�K"1�]�ʦ�����D'p����R1o��l���i턧�5M���x���?�9�>��E3�N��,��\'Y���⮻
���+Ф�8�~;|_��}��3�L�Zr_V�h�'�����]bA::�+���t0�Yv�u�����i
��+���4_d�����)G*op�|s:8��?�H���٨\�����8���"�&H�6�^`_n`�psX�����ގ���K�ʦy;an$o�)���縫F�aĿ��2�����(MR�hPɗ�H�1���f�&��|ݩ6���,Yt��?gn�r��*�`���<� ��R:L�j~n'1�vX� #F0�_���=�3d������ደ/y�襕yԲA
�8����ױFk?��_����s�����/l���O��
fP���D�6�/���G��� ��5��D�(C�/�U�*!����Ԉ�r�g�r���[���;��ݮH�t�F�[��3�_N�����3�:��� �ɠ���B[��~'�2�&[BPa��n
��R+�������;�q��J9���e��
��d���S�Ux��N]N���k:��T�6�-'Zz�v�0 �͸j45[]��)'HE�I��2������p�h�D��.�l�����CA�GE�=����+�"��.G���-�l���\(����&&���^�1���E#����Rur�����hx���L�e=�ڼ�s���ߙd�����NrKq�V�|���U���S�]�\B�p[�|W ��c���	�K�"	,�*'��V��܊ ��'���@OćI����j<��/���ڛ9��-�H?���iҕl� � �<��+����:��L�lo���A��5�_|d��z����v�����*--���j��&�Ԛ[��S�]�V>��p��>�39^)��Y�W�����{F�����F�:�v�A����q��_N�Ԯ�[@Յ>[t	SOu1�.(]�bO���P���f�q:�:րg2G�W{������z�����3�E��k�`�I���(����|~S���jv�^�	�,
Y������v�>.�h"j�X���6䝩B��`���􊝵<T�Z� ��1�C�^�o��K,�S�r���o��PaW��+]�{��.�~�����������h�V�l|q�"j������k��p���j���D�Ic<�6��y��V���i�]9$���m���")�A.6��)��alN��b"��J�Ј��Dn"���s�����@"{�h>) Kfś�b7����K�ĒV���D�G�	���>ߥ��@� �y��"�� r]G���,1�a���5/O_|�G�ޚ���}���p��~^��zZ4�:��6��X�)c��dF��'�d]���q�g��+<|rSQ��~�#�zկ�X�W��?�N:�y5���a�*݁i@2r�1�܄�(z���Y!F~�y��q�����L	�IM䠨hGI� z#��ƪ�|�!0ߚ�aB��+���yr�P����� �u��X��7UZ��]q�y�0�����x����!�B�XRUu�8��E�t��-�e�}���(�FHd�G����_�m�R�ad���g��!Z����瑯(*ς��N�t)<��W04!}��'[9/�X�7V�����7̦-#����I-�Eq��
�i2�j	y"`H��@ x�|'��%9Hx�J��Mf���%���@.3ģ���k�<}]���PBD4A,�سݱ)q�9�kžMBRK�U� �QO/�-��M+L�u8J\q�������_�/���}�ሎ�S���,�O=���z`���>������̃<~��a�\Q>AA�"y����h�QSz�1�>�)ފa;=�hS�j�W��'������\��o�TD0�H��>0qX�	�*��U�MK_�������v� �����Č�S;ݑe��
��1@J�Vc��������D��`���|��{9m�&�NW��Be7����������$?�v��P9���;�;����oI�.	َ{a�<Uh�<�vi�R)�E�UMVc-��fv����^sA���4{e�'P�-���j+4����ϰ��T?�ݱ>n�F�LN9[$�g�1b�z�����s"��8U�k ZM-1"���V��2b�N��R�s4qx��N�`
��rMV�k���O��S�f�pJg0mi��k�&�*�9�
)��Sa��? �����~Uk.��@��x+c���Q�9E��x�?~`F´�5M���	܅�����tO_4���u�G�>��2�RxH� k��^������"0�C�E�?��YK8�������p�m���C��v� :�=��?Ơ�a@}�>�Qzһ�v���*�:����Q��Q�ҧ2D0F7#�^�r������wi��GI>O*�YC@���Ev��G�O%��Z�;狲�Y��:!����d��i��~jۘ�}\@��J���Y�?c�}�h�4������‒�X�q���I�c���;��{] F�:���m�SH�R��Q�<���ٔ��)���ͳ$�=Ƨ��ѫe<�C.�@y^�X�f��ҭvSͩuB���x��rv����e#��Y��SPAk�Xd��C�g���!�t�0�M^<�\s�E����oʌ��Q��9J^<�_�m�9m���e�2T�9�X�{�8ҝ����rת�ô����\`͉�'������U���F 3xC�ﳦ���&)I���>���OW��v���Q�Ez�ؠ�do�?x���z�.bXM�w������x�`z�|��^�9 ��=V��.*��n����1V�=�l�z������P��7�Ÿ�F�n�y�3�S8;z|��<.�V35��b;��#,<��Ӵ*k��V��J�e�شS��� L�4L����>�+t ��ԡ�v&�6�N�fʚ� \�#k\���l����`ȤU�Z@N�^BN�cM+�����\�o1xf�����J�<[�`�z��s����w��\?2�zZ��m�������)&�=���Ts�ÍS���3�"��?Q��UTh�K|ߑW���1n��{�i�F\k^qA��������W.r������̵�:�W�!C�EH�2�s׊��:��'p���$�n�\��_��ח����K�`�^'	�	�;�v`�(V��O-�Pv1¨�qZ\۸��",�	��nC���}�sbz��*��������69�GO����4��iR�?t7v�͑�ZVɃ\�I��3!~�1^�a������<7�*�m
Ę�x����h8�;�-u�]�����/�#?��z'��,<a� �R�$.g0Em�� G�ܽ?0�� ��'�0ѭ�R�(5>�JՐ��yJG����n
���uJ-!�:�{��>s�>�U�7ȗ��5��,K�4��r��H��/+����n�JB4F�L�z[
���� s�4��U X�DDF�X����C0���!����B�o쬁��?��իzz�	ܭnƢ'�f�S�r�c~(�N?`'��}�]'=������~S�x��i��"ʲM9��p��Xy�W������4����K����a�%<������|�5��4H10������8P�����F���b�����s��?Z�n�+�cs�\պ����54?c(��n�I1�}|�X��5�(��5�NU��e�����e��ᒄ���Ӹֹ��Z ���\�$b�6WK�-�G5�k ��z:��t�X��nv�|#P�'t���:ܨ���vp*W���_��E:j��L�0�\�)�F���D�S���d>e���SW�Ԍ����0������<��f�i�`92�K�1�xB�s]os�5Oٶ��̍�n�[���j���J$��iO�(���uv"�������Ҽ8h5s�*2�`=A��1�i�< �F��N#n�[Z�!�|g߾1�i��t��~�bW��_~��Dl����η2���ͮguO1��Pv,�X�i�܉�d�b��s���t'y#b۠5�k
���P�G���p��q���f�.ny ���A�~h�2*��}��!��'|����4k�4z_^�C��*�~�b���7����UU����lEW%:Fr_*%-��ӿ�G��>6.U�]O���r�{ǔy�d�,k��
c�y4?*�uA�����W,��jp,���E����j0N<'�e��si1�;TW�/�N����)j:ܹW�-��C��/(S��L�X��OvK9�ʹ����~B3���P������zu�, �_�?���[4��UR��ϱ�:'}?�ŷ捛�c��^6<H{���|��oj���s'L���|���ɺ	�nV4��0H�X�\Pn��������X'��A{z�5ײ_��\ ��5��q�C��?A�
�m�m�*�@2kWջ�q�,���Y�D�8�(<���FaL��I��w,eN��u�tX��G-O��C͙ɇ��V���=�Ja �I����<����\�X�6�	�s��Un��(��ѡ!�}�q��&r����!V�7�i�$,(�$"&�h��[PQ �c��E5U�ڞ�!ʒ�L���vԙ�u�� )5�+PvThor����a�w_%;zz{�]^�'��Ԡ��Ym��Z����jliC���^{HyZ"�,��C�'��X�\�fȧE�?�dp�����I���X^�q�d���J.Q�&�7\HeS�AE�V�JoAb°i�m��MS��zg�>���t�2�Y<	c��q�f�<��}��#��:�HH��4ҡ!tU��a�v>W�����9H�j3k�N���F����'|�#�㒧z�$:��}�%Ld��,���(w�w�K~[� �n��wŜ�gD��"c�����]��:wG��Bڳ�os�R����&.�7?.c���-��&��"��{{�_E�4-�M|џ�i�>����������\��6!��0"�1��ވ�@�~;��9���P	ˉ,1ۇ�����=��+���/4'��@g��X��Q�_Wi�-�� C�{�F�L���f�b�Tpq���.�g�m�+��|�1�0Y����<���\�>���=���Sс��'���:o5A��ª�x��?�'o���],c���Ye�)�)��>l��� �$O/h�!��"��KHܥ �6�5��$D�nO}a���3(<�({��W����nW��]�Juॱe�pe�=nd!��wل���҈
f�+9{[^�"ve%�o��ə�\�&�d/��8�_��x��r��R@���P̡j~�Q��G��ʌ1�Z:���N�B�?���tu2.7�ˣo�S~�OGk�	�?��b����QӰ���N�)Q.��v н�;�Z����L���%+�"�&�*)n���|� �����4�E�$i\�!&^@<�����zIۘN��K$�|�q5HP#�����5t����f,���^ϜP�?�Kͨ�WX3����<A�����8�%�mkӳKs��ܝ<kGq\���w.�E��y�*[a�l��4'~\z�g�m:�g���W��	�{�9�n���p�ֶ�B�f����}h���h��V�&E��ǵ�aN'J=�86�/c�oa��\���fq2��,絻ߺ���?�� ��`,�V ���ِ@],��F�k�g�8׹8Uڥ`c����2c��� �3�c	��b�S�3'=H9�^�ߎ��d;B6ܰTš y_�u���a�x!l�(|�BU"��X�ڎ� K��p`\���șV(x"�����I����y���Cd��!������W������~b/:��)��XҿUg���nwJN�cm��q3;��F6j��I9k4~)g��!w엜0���f�%Ă�w��]�"ye����F�++�D�'��x/V���%�<�T��j�jz�(`�F�A������^���*�0��F�p����	x�꯴���#�*��
Y_�	.�8V��*���l�A�d4�c�=p�o{@N�:L�M9i��a�uc����ܓ�@��T)�]��9�0Mい;��������D�!
f�W���4 �=���$�����(�k������)q�70���%��?d�=�2m8i��Ug�lyA���kpA�u��t�$�$PQ����Z��_ �����&�����q�r��H�"�\���蛹K2�q�1g���1L���\wwg��a�'�'=����`���s�>@��l����v��z�ll6R(KQ�NK6�f���
�?Z���^Q�eDY1�/h� `e���1奰Z�$̇����8_Y��{J,sO����\ �A ����S���Ǽ����½���w+M�Ñ����y�͘�@��uB,�e~�ۮ�`qKޚ��{�;KB5o�)uM�W�
�ؼ�f$F��0&�$�gm-�D�^o�ն���G�V�ԟ���g��[D O�\��*<P��%}���oN(3��g���Kl6���21kq�~�p���*��gO��j�gBފ�u`X�>������;���r{O�-$� 6�Ƀ�O��9E94��nW���M�딌^`�ǻ�TE�l}�6��L�{T�2��R��j��
.�NDwh_��K���T��|*m�o�g:�j�H�=r�*���ܫK�u�h%�N¾�7��.�Sg�\�z�x ��B[j�\��x鈛�،�/t���֒eM����Ky�S��{'����&����{2���~� ���$DL=8SO$UM!��p�,��۬h������q�Ƌ�Gg�x#j��C���c�"�uA96u��%i�b��o�0��dޟ��A�=�L'�6E�Y�� ���#�`/U��A��ol^}�e)tӄ�/=/nK	�(l��D��t��=��h����NZG�٭̱��qb˳L	u �����L�!������Ɗ{���qm�`��ڧCP��c��a�*iV��h�y�4- b��c�O��O�B[yi?iF�j�k�ʙ�����.�E9TJ�Fܟ�e���	IΔ���̊��:�aVJ�7�E^L��6�4�ٮ�DPl$TvBMslg�<g���'s!a>����o�c�S�l"���,b곛�b?x-V޵�c��z�㥠l�rJ�D�ψ��t ��xmXpQp���-�2��ۤ�u���i�mc|l c7�ӂ�[�b�i��)7���3�$����T��D�?�k*5�xt��[�;#h��y�S$0n���	��ޡ����#oP*�¦>�@�֎7=��1����^��U�N�1N�K��-���Y�����+�PZ
��A�9f��7���#,DP�a
K�{�� �R��oV+���u�6�����A�L���U�ZA�s�L���sS��R�ɽ��M˶��i��.&Q��\�E{�v��ԭ�3yC�&RIQɊ���h��g�
���T�7��qmwKE��R�\������kP28���b��
K�����n�T�Q"�kw'J�ЈЎ����1��q�3�}T��h�	�*�<�^��ht[TM��tO��$I6S� ꭉ�`��8�|qe��߹�REفǐʞ]J��k<����U}��9Ί+$�H��I���9;Q���gͥILV�U����e[��?!��$���C��A�%�ܮТ����zE�Ӑ,��d��ú�gJ���9P�ՙ�D�IV���ZE�t	�+��kH���gu�Yu��8�#�go��"�c�'�d G�*Xl&М$�	��-=�������"�z��I���~������4�~��5����=+�ix��a�Xo9��C|�x�@����,��8ŉ�9y�%%��:��{;.�a j+�@Lo@�lL����|�����A�^Y��Q�AޱBj�z��1�I��t�PU��;M�MG�ɹ��xp����R<�V�e��j�I�P���(�ў��%W���6C��WV_��a��΋g;�{Q���#o49��A$�W$� Ϫ�׹�#�?����n����?��K��MG�$��.6�K�����Z��m����\����
��hĥ�G�&�!���3}y?*Tb)��5͏���&WIͩ%�({���[�r�Ro�W�ˤѧ�ypd'�L_M�/\�)�W!g����:<���>�IhB���,u �Ov2P!8���q��F�
��UZ����dX��<t���g -��I"!ƞ��\���	R���3��P�DbD�E��a�f�i�Z%�R�F�>sӳN��"������c��rz��T��5���AV֯���ζ3���������.��!�p�p"�yZ�x�$�1/��@n_ѢZ쳳P;���k	�W@ S�'5�Z�=m����6�iE�3�r� ��� |~@S�2|�T�#o�#����g.*M�:�"씫>�(�"NE��PHݞ~
�B��K:&���6	��ԚNo�<�)��{8D80��G���c��(��t se܌���LOg���v,9�d��I�^�|5R�m�����6��}6����2��5zܪs>�]��2���N�ϲ��5p~��0T7mߔ������T����lh����-��	����?�9��R5<f=��~�Ke���p�� tc�%q�Ƃ��gPX���˱~����t�]~��j��6f��q�H��q���x��������yjx�ᢝ� �;�好��SBrfGa��s<#Kk�O�.���0KU3�]w�t��:=B�u5�~�m�LW�D:Fy'���nN2#�4�Y%ߐ�c���nQV�Hj����(]X�P����^�����^�F4�¯���ہ�!�:ګ��#�
�u2+D��g��7�]�J�^���<Ay�d K�]{�}A08/f�b��Hb��Y�1�$ЩF ��Y���H]u��l�]��S�� �V�Y�b�[R�����`��ܫ�o�3u.����Fj0 S7�w��c[H ��Q���^�i�|�ą�#��V�z���o-%S�AA�__|PWکj��K@��z����.H*���I�#��l�Z��~	
��c�!�/� �9*�v�n��0����ޚ�N�T��$ J�&���&�c�-�(\;��@���ѾͣѠȗe7�<���5R,��R�O�s��2M�_���e�QE^M�h2�V��Tpi�sdH��-�������¬p�������8�M�T�Ƿ9X^��>�r�z�Y�w-]���g%|mD� ��;��)��1W���g9"Ä\�PK�惇$�?�Y�����O�Vm�k�����:e�o�[�|�Ԅ��hHdM���@�
��?iN[�����4�Z|�ƴ���V��a؍ƯH~G�b��ɔo���S�j�xK%ub;�n�W�Dq�U>^�i�qG�� �Ŧ�
�Ow4���D����聶0q�)C�ռVFY��|$���8�LJU:h/+���!7G_ZC*�*�&�����2ع��}�����0��J��xFS�Fa��/*���#hQ4 �y�d��l��T�GB7����T�[jY����=q�����2D'�M��������$�>��Ǟ2�,&Ȏ��]$�Ke`��qD��� ^�4���m��	�\��p��a�%���)�'0`n݉=c�'�zR��E��Ǻa0�I, ϰ� 04�K�����
-χ� �����2�=��i"f�P��zr�M�d�wOh[^�@G�d�li����K�6�L"e
@/�u�ͼ�;�_Y����NP��5���2C�R��X��W�xˢ�ݴ;�cα�x:��!iDC���#g�ӌlU�$��D� `.P���pW��>_H��鼓S���LCT�r�19p��P?gJ��p"y��]ً:i���R���K���(�C��[iuFK����Eh;L0�k_n����_�r�i���# �b�=zvz����S�u?ߥ�r�����ā�e<<9W{W>P(Y��!째�l�a���ګ������TҠ1��7��I�c�u�+�dJ����j}����*��S`��|�����е�J�t�?�0�+<U�3�+����}洖Q��m���g
[��!l�0��ny3�̈��gܰ����ۚ?^ӒTϊ��Xf2��vQ��2��q�b�q,�+������T�SF��^�G�>�v��p�Q��W�zL��&ʓy6;0�H_9�/7�j��	�p r�ώ}�B���A���s�iߡ6�p��h!�򴺈�j�ƍ�.��^l�Њ�s:(Q$ �Q���L��٭���&��C2vT>X�W1��ؙɒ���yD
Ρ%��(��Sm�D8�~|���}�B�4�I�}��U�U�
��4]���][zX~��b�V�pε)b�%�4�H��l��PK����]�A�@Pë��?P
��P���H�7��C��%]:��ٖd��{X6�,(�,����i�"��_�x�c���)�r{���E�S��_d�e�Efg�fN�B[%C���̨;;����G�{��_� �;q��%���ᱍ����X�m~O/ u6�u�c��WE����j�׳,�ɲ}���Xh�����g�|��W#�:��{?�'�֤Ȟ�ܔ�Z�A�x|J�������_��x	�?Uz,��Jv�VA=qa�U���ܒ)��E��ezE)���M6hIx�|��O.�4�VݼM#׳%��`jB�:��|�7nǇܨ�q���A��j�ʁ7n�0@�� m&�,�Š0{��l���׷�(]퇉����pȼ3���Z-i�-r�=\���\#���E(���L���A��G?�h�m}��Ȝ�A������2m���z��+X���Ѫ�4��It1���[�,����`�1��f��uP��K[xa�ʀ�uO�lB����ED�R6v��э�r��eaw�����wUcר=.�edP�mu`;��^���I$�$�"B�ž�G�l8��oWG�>"(��,�����VJ>U$Pp�ih9�{I��qMe�ڜ��Q	!���WOG�,�c��WM�q)���,�
��Y�9�*���Y�9��ɄOkl/2:��_�xd����`
ͥM�%^�܊ݻ�٫_h1�^Lڽ�X�I:�@8a�720 ��6�ȶt�^�υL�x�Nl�ٮ�o�-ä́����v9ڳ��W�!��k�TA��-oi"�鲳��v����9���8�T������!L�>�|T<|5�_*O{��o?O6�&��#�MІD�y���Y�x�@\��B=��%YA[�r8�N�pD��kR�W�JO{�T�r[-�B����'֛���e���dB�*�<�Q#_�F9��D��R�e�>RX�	ί$&�<$���pA��t���;J�Jc���sZCiN���<�SP�k� �}�Q�D'�raD�~�3�ӞG�W}$�p4���LD|ܸ��]��zN���[ۘ�#g�X��I��5`=Nz/�B5<�M�@���-��4��޴��"!')��ѨZ*l���h�ݜ�4HX$�$D��Λ���w�z�${f�n�d���&N?& �٭�ó�jx��A��*���OQH:w8�Y?�J�l�=�-^!|-��PއQ.�Li���i�M�r���=x^�Ǫ�����Հ�i���Ȃv�����)TdP�[�WD���um�9�ak����&L��
��*�}���}�)i���*˷�x�}����
�y�$���B�bʰp�a��O ���9]�2Qz�4�q&�<E�0�<ncT �v��B�/|�뵻����+�]�1#�[	���s?��r�~]F��4q����c��:8��-;w�^��\,��Xb9:kd��w{.���s2W�G��q�/�k\��o�*��h����y��Q�?���Ḙ�)�Fiͼ�PK��)u-M�"�7"4�>�<�J��]�Q��IR|�Pr���c�b0�� � 
L�GY:¯Ć+ا>pa�iAb��S�T%�5���!3jL>茬���wҎ ��t���\�8���[�[iu%��b�%��.Q�_�K�u�ϥ��I���|�py�������~SJ(��5z�p���)K+�#zߩ�M��"���=�H@v)�G^��6F~E�t�A��Iǽ��J®Gkj���܈I�լ,�c��7��,�t�2+M/86��SŖ�YP����pb�� �����]���&���p�^^���:�g�|g���������Hˇ���4��$,����f3�#�D#�|DA�ʔ��:P*a�y;#flV��=c���b�2��9ϢdT����1���/�{����h/�%"u�b�}�u��4?i`��1!7�!oS���^}X��i�[E`( c G��#���mSA��Ѩx(h�2� d�&*ߒH�����N�{����jF#���"�A��9����H~���S.�b�(>����Mw��Apl�P����n�1R-}�L�Sд^�#��é�1�,��˧S*/OV��~� �)��	M��ȍکř�}e�g~��ۼ?3�и�xE��A��	F��re�󘨷�ʅ�]����eC�o���)��,���}�𵛨�r�Wˆm�-��;�@l"�xKO��Q����G�ha7�E��v�_ԫ��o����P���q������32&�4����e�qir�I�OK+S'��,g��Rg(:iY�%Y�:���Ϟ1������/�����֘ր��C���L�A��tz���j����Z����δ�晇P)����1nTR�u<��i�Q�.��M� ����R�l�v/k�Rƪk;=�ʨi���
�,h�ccy���p��ci�/|���}�G[Qx���V��Cd�>���Pgg��75��c[�e��԰q�2g�P���8�pKD�0M�"��®�,�0���
#I����,<�GμsO� �&D�_���c��2�a!���n�H��t���A�?�?�@��2O&���߰׾���±�Z�QN��<qb��U?3T�?�	S��v���o�u��K�4��֏6m� �>�0�ڝ!����jL]}��R)��K ����/M�]߻*����YѶ{�\$�n�7(E�%��=@s:����ݠ9�=� (��y1FPb5��>{iC��\��>�bk"�y�7Ĺ�$�`jF~��:��@� I�����Zw�{l���d����nSu���Z����(�~�` c���/]��ke��8h0���E�U�5�jm,����c+D�:�5��%b��Xڽ�$kڭU�푘-�:P\W0�&�1�5�פf=(�*�����:� I}��j����kxsKF��׻$��c�'�H�N���D;���K-�5��z�+FI��yXqˉ�:���Ln�j��F���@b{����[���6�n-��� ��}g2��iO��uޒ틶�N�Β�H�����F��R��8�|i}l��+��8=v��|�F���b&���]�VnL]M�M6D���xZ �Sx�8w���AGFJ�8�P�����aj�F���p)��dј1O˷�-:���j������TÊ��`����z��M� s�cMdD��#��o�ဍ���;Ɉr�y�k�0Ӯ?l�p�lUVJ���L��c=���Пy�#Zu�yӺ�ƭh���y*�U���M1���+�U�NV3��k����-�.�:S�������돭��|�q���$��À�&&fN�Р��P�P�Ѫ_�Dnn�E�/:-+B9�xw���8?�9��,�ܮ���<�QT��q��C�<=��ɈB��n�E�̩O~p�[^=ľ�O6NoW�O�xk�"m���;�W�y�YO˭c����O��a��.ém�?Ӎ�?]̄�O�zq�e� B������3a���j>YI��uQCrG6q[��un��sai插����9���J�#�ܔ���v��N�i۪d��]�j�f9\̣����A���4$;<2�R�׹�t�]D�!����0}�G�0�iA!��i�1V��|^�c�������̅�U�v���k�yF�D�H�r��5���S�G-�������A�������OE�&�C�ˬA�$@ߙ��6�����K�mM_�Y,�r09��fg�x�hV�+��t����I��2R|d�69��D���W��7�4��%loH��"u}�#��d�v��#��M�1�DY��wc=���d�j�"��.�K��n�_�+w�Y1��Φ�R��g˙��n��o1=��I3��<J%��&Ę�f3*�cC_��z����ڊ�:os�1��"��Y��vZ�o���ʸ����,�&�����F ��p�H#��#+�G}��v�r��L��$�\�-'��-n6YK�n�@&֐���$6v�s�o�8vp�O�n�l�Cq����?��Q��XQ���5⽞�I�0�����)7B��9���q/D�Z�č�<�E�F�2jl���d
�-
F{ w?X]K	1|�h�%�+;{�N�+i���mo�@�2�j��"���=ƍ��iB{�lsK�5�I��
�ݕaE��T��-H�����y�擪E`Cz�}ˬx,�3*�ʠ�����?(8����
B�!Ƀ���_�拄�q�R��l8ǂѧȾ�2�vt���#�/���4��a���/�:�AK"�O" v���\hn��	A*7�bݳ��+�ܞ��&<ҷoQ����C��m-,��΢��֝~��Cn#�:.���k��W(j�"3���7|4BR��p��ܺ��`�$%v%�?
��2Z~7˸j� �*d�L���(-H�����ׅ�q궿,Z�@.Whe�m�������ޕ���U�9���#���r���[����5��L ���\��=7�#��0��Ac,v�UU�9��~�' ��lDg��� z�;��:b|L37�S�m�b��=��V��6��k��J�a�mg�|��M7���/fҞ�� Q_P��S��\\W�����XX�;�P��}��?*��;D]��=�W|I�O�)��S�"��O���M�\�MW8��Fz`�߈Ib�`/S������'��M�.��8���Ŧ�4%TWq��$0�&�!���H��I��F��@�� c���լ�fb�w3� �Ɋ62?S�c/7?� �A�Gx�#L�-�j<B�4y�O�f��𨡉|�.M�p"���殐:56kKU�zK�Bu�@���oK�68hDV�JJ�
x�7��7�M����f��lW*�F#a��yN�ڤ&#�~��L�L��_�/���e;�a�j7�;D�~� ܐ���nO��]�.h���=ʢ7�I�
=�9z�&p������%"� ���wk�����!>������ᭂ����'b�]b=�o�r<�0:2�j�s��ۇ||�k�IьDNwE/��}fO)�J��F=�a"JTCUt�i���8ρ�CT�[G�a�d�$c�""�L��|S�Yx됴Ya�M]�1ߧ�7.φ��z��7���'D@��؎��I�{�����"�.�D�3�p&ay��Bx��j�Lx�E3P��C-OI6�X� �O�gb�r*b�z���#KQ;s)u�g�-��eBp�Fd�����|T����8cpO� 3�|X	���`gӞ�n�?VO�&�Xf������sq�5�j!�z
����CS��7������K���8�m9
����Q���V��ح:|ռ�K�����I� �#�q����� 	4՚v܌,?b��v����!JfF�w?�0	,\P\\��)?^J�E^L���=b��>(1_���"�V��~�������r����I���Zh�.m���. �Di_3�6����e1�Ş�
��M�Me��a����v��!�~�(*�1��=_�W �'b����zDZ�+�t	�pג^;0ghL�����qTcou���D����U��"��~?W7ɸ��{�;�?^u�-�xO�A�F���5w��[����1�%��k�ױ?Y�Gu��  �c��(��'@�w��C#���D�>��x�� kI��ʢ�>������u����Ӌ�x �Wj\W�
Ϣ���-��#��f$b�w�7��~���0�f�մ���Cb�}[���j��q�W]r%���2�x3��Е5V��$�e�KF7�XyL��i���[:jg`� ��n��tÜ�K�0�o���5���(a�9n,y!pٛ��U�-~�����h(N���jǖ�L"#W&��b�&�iu�'�Z�x>Q-�ڛ�f�TuCB�*�)�h�E]8i��bMq�F�]s��������T��g�d�����W�rW�)�@b��_�`u��}$����>�'���=�78'6]�x��� ٌV�-�O��Ԙ��}��M��S�S�DT;T �I�z��~��$�b
��e�`"�} Z��&A�\�ʿ�R?�y�w$F������� .�]΁P�?|�0Dd�Q�T�fUD�F<��i_V�!���j�
:�����W����00prV����#0�>�vO�(��GcN�}q-Uۋ��k��O�UFY� 1㣄�i��6ЦtܸQ��Cy�̊4��Ę{���3�ѵ���ϋ6Ȉ�mD�?���-�GS�c���m�p<	������U�3m���"���n���!rbvGh��8�����g����r�J��ks;���B�ob����f�*R��qQ�2�~��1�*��R��e��x�?�K`8o�`��0�QFx��R&-�z�62���!?d��b�� ����%��$��F}8��!����D��]`�KIzݝO�a	�h���ĕ����M��; �1��܇��E =����%X�&Np#z1�j����R+_�c�k��oK�v���ё3<_�	��#S[(�3I@#u�Gxme�NܟJv�4%b_�(�90@m5ǥQo9Xg����׸<����rq$-aK��	�̿"\A���=L8��a*����|�(Q	��0k�(n��M�զ:�\��D��O�D�<t�F:v
KwU,��s�A�#��B ���ʎԉ���t
��,;ڸbBF!���(�Tf��&;��}�'i���6��W*��5�S	��
�L���2]�_l��Ð7ao�fi��K� ���K�_�j���@Q���+U\43}�@#yS�r�,�^�b�w�,�5i�	C0Җ���iG��58p��[#O��co@/y�'zR��i�����M�S�R���Kr�NT�|��,�����l��?w�c.��A�C��?�ҎN�m�;x�Z�/�F��U��r#yX����0�����G��1� �#~� �3-a�b���;����l��pg��*�=���}��oé=��*�y�"��Yo/���J0�b`��B�3<�t�J0?�W(XxŮ�\��@�������	��$��5X� ��G�[sӳ�k��σ���J7��o��վ�k�=��1���":̧�	] �<�_p����ݞ�P N-�x�x�r�Q�Tjl5��-<�08ӄ.r��	c�N��C`%���Qw�����ȭ�c/J:8^]?��X��h�� �)V[�CdM���#i'RS�a�6���R����?	��� 	O�7�ϊ� _�>L�)j�ReὃqB\Z���n��p�GS���%��*f/`!�}�g���h*�� ?ӏU�%�5�@�z���E��ݻ��R2��E�}��D=���������M����P�.�*��L-y2k�]����7z���Dh̊�J�\�����f��0��>�ыS!3S��a��Np�*�l:>��n�"�����C2�}������4��G������At{��6R����y�c������K��\��	
�ژ��~	�1�l�B�`���5���>�]=�=�wU�؂=����nx.�������T�V������@2�H-�x�`t��=�|��������V�p�؏�7T�E���N�$�t?�	SoT�R�n�&��9��UL��3�����
Ab� &��;g����A�����S��D�K�Y�.��� ���Y��rC�7�=���ѤNL�J""�"��M�9��m	Ո'�C�|����ߠ=5�un��`܊	�*8�w��qkA�U���	,&J��Y �H��C�&q��PAng�@��RU�����q�٥6Æ���/�P������Ž~,o��� �R��tt����F��0�S�Ч)���E�"M��m�Ɔ�����Ű�~HG�Β�捿��]���4�>j�����Ok�� RQ���c�f�����ʘpZ��@���3t�?t@K����<J�C@E@눔���tN���$F�w�L/0d�H��x�Tҳu�(7X�9�w&8[x�d����\�H[�JiQ3��ǰmK�eQ$�b�=�-��-6�z�qK��a�|���FeG9�;��T-ZP1���rR��9��9'�tZ)y),q���_�z3��Y���z+v�ޥ�D��ohUF�n~�y�ಊ4d��ƹ�(G�<BZ�����Y�#L&���g6t�:űz�~Ij��qtk�W	�#���.H������K���D6���,���c�;0�dx��Ō6��(h�وq�ԈH���P�>T%ф��f4־a�uka0\YU�^X6�Z�0zoJ���9Au���όU�OYR$���-�&n)'�ad��x?��`o��t�ET���҂&�FA�U��>���{~7�M��9� �N,Ch��5{����:UP��s��q��"� ��[ɴ����
S2ܵ!8�n}�F�k�����o�A~��xBE�� �%"�u	@����z�E�[F�c�/�Bv�u;S���͠;���kd��}�!�ན��&ۗ2I=: *��ӏ�(�ɇpUds��,B�����H!��	��5Fd���qp�~�4X�[���d��MBciy�c�^{6R�䴒�D��J2�$�&���B���{q����ŧ��Rc��y]{�\��E�}���$g|k_(8���N��f��Ѡ.�A�,c�Q�f��B$�dS@L�5�S��/�ôhP�a�W���o)����-������Vp��a�tE�Y�}V��f("�ETW����$�OQ�^{W��h���z��`��?Z�r�
��l=����������b�W�z��'�?t�N_�����H��R�:`�;���2�:�X��Z���^w�k���:��C��뤝�b���|�?�E&"%�D�e�EN�e$�����M��>}%s-�tB����@3�PS��"��[q�Z����VWq��J��[��|�-��-_,ۺ���]�\��ɴ�p��W,�}L��JQORضU��bI�n����]�0���|v^��?�yq�‛��e	���pu��:f�6���(��:��wцhH���I�~��˺I�=�������S��V�A���Usn�������-zf�\��_���0�F[b[Ӯ��S��u�<le[w��� �mz=j�)�Ңka1hh`��(�M�%����Є����(��XZ l�2��἖x��g��#S=c����fkSN3ۍ��:� ����]K��55C}?���+��X_��--�-�ŵ1.SPX诗�_�mx���*J�Q!�r���[�Y���*oqc&�`d4V5T3�x�:A�DQ���G�����Ӈ�`1#��=�%�G�"�Q�h�M�p4V����|�
�BR�dF�nÒɽ%t��<�D@8��9�t�ĺ�!�T5�o��i��Q5km��
Mƒ� g�؛=3���H]���9��?H�����b�LK��i>p�&βi���>TQ����ތ2�u��	ژ<�&�`�kH�a�pqƿ�7���.#ϔyO/����U��R�<j������fQ-T>%xC��	 �9�ia�z�_KĊ�b�D�Χs���{ZfI�`.TWԼfܽG����Z�G�x7���Vx#�W�|Q!��v���i�BN����g��#^����!�~q��ݱ>�
�EVѧ�<RIL�� �SsaJ�J�"��LN�����Jf0�Y���yi�AXI���R���t��h��N��Z���ܖ܌ߡ��a'�l��2�x���B9Z���Z{�v��v"D�2�%�Q�	��\t��a�3䢫rPKӱ�H��P�I�:���27��M��m'���>d	�8-=F���:�еvQS�R�T���ߴ�k���ΈPfcl%�5j`�ͼ����y�(Q���~�t4rlP���s\^�)(�h}�^�.P�T���AI�����Ǽ��І�X�W8`Q��m�����{�3�� v���������vw��{�)�GErܮ�P�TGאʇrkטj'~V;3��&Z��1~�De�p�q�_��C�%�4p1��G^=/Xb���",f�z��s�dG�z`�����
�Ps�z�~�d�/ ���'�+�pX1qK�,}r��3�>��^�2ćjW�����b^����H%��0uy�� oй4,&�����֔*�	Po
@}�"�����Mkom�*gY!�տ�Ǝ� Ǝ�C��A 4��Dk��>�*	5�" ���c�*?��S ��F�	����� �/��30��k�g�d�躟�iƧT�(�H�u8��;f}��HJ�X4��]GV��l:}��d&yBS���6 ����������{F��? �xʡ�:�[j�w���ƈ.k�&�^����p75����ӳ�DR�;P��:�`�|� #%��:A1�A�U�������A'0vo�/�p��	��"F�Q�+|B�g��m��V;��zH��>�GE�������F�N뾫9�r!^��hu�Ł@����cIc��4�.���Otͱh�(pj��B.M�B�6�3�����e��	�lI�����V4�q8��hS}�!t�-��J�"��99�>��hC���D~�r}�ҩ6�D�,�)9e/�|�����G �M);��L-~0�y�¸.��&�5>Q�3)�>"���qL����������zM�Pv䱻�o�x��*����E�3���� ^�IѦL�.	U&
�E��78��xƀ�	��ޥ��Hcėg�B޶ש႐�}���d�b���(ϖ�{W�vؾ��!~�Y�����6E~@����΀���&^�Ǳ.
CX�]dLt����S|/�v���	މ��|��H��H�EU=���-�N�S�{���-��-��(����Ț_�dP����@��L�%Ӣ#�p�C�E�c�����l}׵����@�#ig9���{L��敉�e�*	�×Eȸ0L�ùH���v����E��e�.qm��P� ��R�ʗ���UR�'"�X�qr!����VB�G����)H\W�V�l�|ƌ���dR����ǫ��iv��!����#�q0���}�|��b�5(i��óp z'(��/���k��j;	0�j�˧Ɓ�{%S.'�t�-�{,R��|6x��?W�ALOrCjT���n���ϩ�y7��+-9�X-�,^v�_�`�t%%�FF������B_K1�z�4���{���C0z�6,�}<ؙ��w/��j2)խ��G$�T�=��X�0	ꚏ�ʤ�[���&]6�\�Un'�:��X���ͳ̻�!�Sd�P�7&�7>���j����Э��=��7s@MN�5�MޢC��hDf��KP�1���g�9��S��S�a���2�c �7`�a��Б�ԁhRS^w�1��	��[��Nұ�������h����9�CO��,��y�7 !�"���Ui��$:(95[�/	2��B3KA�d�V�!����N�ϲ�G��� ��aL۬�����"�h�oƑ��?�ɿ54O��ƌ�78��"2K�Y�cް9�
&��� q��4����S�E�zetM̓�Dr�/�k	��l�2�"�?�u�k�lu���Ǌ��\' ڀ&� �۞]h��G��js5��J�碳r�JY�ۅ���!��n��b}S�B�j�\ٳ�����36,��'C���#�E�E���3j��YfZ�./�ӗЋ+<�^2�d�͒�#��޽V,ћl1��E�U�d"�`=K �-�?�E�Y���D�W�'.����Ѕ��9/Q=3�4I�R�0�l��
�O��N��@!Gf5����v_-#�"�7�M�5�x�z�_(P�]�^�
(j:��k�hqg�;�ፇ����RQi��[��5n�I��,m�J�zn���D�/�Z������G(�+4u�իSL@%3�5W��X�a.fV�a�v�cb������w ��1:Ə��+���r1�����iq��������Ǹ~�I�K�<����}�0|Ҕ����ɣ��Ydnj]��}�b]њ�^|�4��Af�#���昇�R~z�;# ���uE����	9e(�	�f�$�L��-[j��YRTJ�����������(m������b���I�l�!�D���v��n����$ȳ���7�+&�5# ��dy�����9gVl��
L������;�I���=�����{D���U�QT4��2������y�#K����=������?��eb���V����)h���+��;L�!<�>_  ~*K�	�ޔY;��C{A���_����N�!�)(��n�կ[S0{�dYX&q���h~U��7�lO���B�͋��e���F�㪗���S �W)������m���R��	k���9��-*��`!�[�1S��i�(z� B��L�����<Aj��X�[A▼�z�P-}�p�0��g�ᅫ�]�[�Rʖ�;V�0����Nk���Li@%�?dY��� <R$ʼ�BőΏ�֮J�Śr��E�I�Ό�(b�q�(B��3%����Wb��`^>M\�b��FY# o����Ye�[l����0���f�	U�jϷa��S6h�|S�e����ժ�N%�#i�;*��,�X�R����(�NPiU�hA���7G���>7^C�}�6츹��V�(�折Q��2���;Ĳ�I#����9�	�5E��43��(T���D��c��\=V���G���ۤ�>���fU<�V�$��w��uh2gz�xzH0����b�)ٜR�#G�&�Ũ\2�]��"��]�w��c�SiW�����~B`�Ix�EwfZt2p�\9=k�G�y<���p��7oc/��##��W�1�D��A~6W��9h�lz7�Ld�¦�^�谐�>P�y��$ #�v�����Hϲ�ƕ<5Z�n�G����Z��+W�0���8����b/j�%����-��'�%���ݝȕ��u^��}�5���j�^���P��XM�DmZ��ђ�8tr+���~���A�{@�}��`��
����=�g�G y�}VR�l���O��{�yǹ��J�f�}���P�/��	���Y��#0�AU��L����&�d�uq���"ܧ�����"Z1�S:����s��a=�ø�:��đ��,޼=16�3m��+��Ҿ�����F%.����#��=���ʮ��`��s���Ni1�v�$��t`f�W�hF�9L1�^o���א��A����S�,�=)�Ź�y�.�A���GB�;��&i�ͺ9&�ѕyDҋ�2�����c^��e��	�)�Yߧܳg�I��=��B'ԡ�0�$�c�G��!�R^���+�V9S��.q���{�0��121�3�X��`XxE�a0fi?�g��%��gE�$e���&�¯��u�lp%늵�8�h��'���m�)��^�����̃�Ȋ�vK�9�t�d��/�z�� f�@�#flA�J��!�M���I��,��>��>�'����<�]�a������1��`���U^r-��+�VMIL���(d21�e�}�5ζ	���MY�8Dhp���u/�Ƙ.�w�l(,=�]��[B.�B�Qd'E^�����G����s����%8������9��4�G�9+����ߊz1F�cw�{�'��R�%����j�bۅ��{�	�3����uǰ�n�>����A�b������~oD'���p��� ҥ�߂A���s�H"������2j�>����Wc�T�:~�F�̸r^2�Gc����j�+c��UĿ�]���4��1����Ğ��E�,7N\o�뼠�^����v�[��!	���h�������C˂8A,�r<�����j,QUz��`KWVy�z�����`���h�I�DG��'��߀��8r�׆<�t�	ͳ���%O�j�m��/e\�V�>Nh-�L� ��m6 ��Bc����4�{�]��8����J{�����q����A��"�E���m"ӵo�UT �Ds��O�q�L�,xq�⩄���ka�1'_i��5|g��f��g-Tݿ�����e}I���x*�c��i� #�k���@S�P�A��@����l#��������� �Q_���
�ݦ�{Y�[c���s0H'#�=c)q0#���r����T�(�?�b7�g��'!<�s��7+�">�����{_��l2�u	3P>��rS���GR��Ǿ�wA82
��pg���h�~�А�q�7U�~�_��x�q?���j�+�Q��1] [!�}������՟�'^�lnQ+BH�s��L�[zq�p���xzդʭ�v���	O��=�(��~G�c�2���T/u�V�)a�*טj|�#�VN���;@����-T��Ȼb�>�^ ��渄�ܘ�[�gҎZ8/#KnA��Z�|W�?��@/M>�}Ȳ�?���LW�+<��$�3�IJ]I�W�!n$;~�\������	T��3�Z�9���h@6�͛(�户-������߹sƆ����M�y��ta��תl�6�Y�l?�10kN�K4���9���3�Sy��d~��zz��ю(*p�{E�V3/�,��h�<8gr��=۞@pAJJg��[��{����}D]$i�v�'��"
�~���40ݫ�Xw��!�t�UW�Jr-�K�~{-�o]# E�M������-���)#���m%�j|��R#9ck�|���I�{x���O!O���2�4R��-%�=�����A�2����� =G~�~���vA����0�F+}�p���U��UWmc�}�{m;�N�#�4�mЀ/=�cʧ4{��_�M☪�.�ܘ{�)�� ][�-��&`��CI`wz�;@�=S�j�����Z4BK���6 2R��Z�����r>ș�ɖ#�>�z�E�jt8�?�TV~��>v<������I������@V�a�$JY�Y�|9PC��Zڞ@�L��P���
[=簄�]�V�7�^�R��X��{ٝgm�k0k�Ѫ��ĕ ���4;Sk��:o;B,��?�����+1�)z?���C�� &gl��%�gn�ZxHu�N�Ƹ��2�@V��];ͬd2>d�x�`�k�//��y��C~�y_��ty��Q�i�3[�_�+I�tC; �o �noޜ��6&���h���N��9l�R�D�����0z���qW��b��}yP���Ow������Ç�A2�![�����2���wkx=F&1}{*�ϒ�iΨ
�EW<x�x�G�fT5LY�L�����M����X�e�>�kz1Y8�)/��'$��4,Jίf-+{wt����QFm�	��SZ=C�'+���T��z��#" ӗ�?��(�a��w��8�ykR�+d^B�+rJ����
*!�4d��Yb�hjP'��(7����ڄ�F0.+½#�mH�����MkBy��Nc_FFzR�*U�R�7��v�1k�m&[��56�����.Y�[zi6��|��i��� +�j^S�mօ�%wʹ����(`%i��q�+�*��ůL9��������I�[�!�>�~�<� ���W�ia{����.�,@'7\?��'�.C��������3��#�6����~0�/�I��U�[]�y���DЃ�ߌ�~?i��}ҽ�l�W`�� �ߴP|Q�?�jŬ�S���M�-�+��)�p:<&���%�Md�M�7؄1�2�4:�v�g�w���Go�U�Ċ]S�/2{��� p�X�O��bn�w0uQ�L��fZ�,���N�\#�(�6L<RG�E
~�x�+�r���n�����3��#k28�L�%\C� �b�|=Ǝ��V=���C�SR��<�LS~� C_��X��}����˙��áU�����%=�E7os޲��"�V?�������o����s�zq�/���tP�6�eW�D�1�װ��a���� �NI[��̶��ɢ�X�����ED3$-����o�3�L�t����h���i��-'*�&��~�^˰��m믃W
�5�C��*����#�=�r��9�p��9bX���!��7�}��h�Ǥ}��|�Emmr9�f	eJ��s
��\k���k	��þ� )E�,�1Y�{��[m���A|�4��y�;�^���y�O�U������Y��W��0�d�#�(�
7���w�����T�}�#7N4D�8܏�
SvFfk�h���A�<��V��Bs"ř�ü�� %(�+���mK�(�+(&ahH0�Ev��� re��n�ŖI���Rz�ݙ��w%�Z�c4�������Ǐ�՞9��DX�u�W.�ta���KSY���u�?�(�����3�-ۼ���ՋЀǞ��d��
i�_�2af����m�G?$>�O4�D�@d�qP�f��.`�|����
��.?�KG{am=�R}�)�W��?�$&�6NFA�؄���Z���*Òf[�w��k�r_��?��p��_"�,�zz�Q�%>~�0�T���G���\,373�}yÊ:����-��5����~,����3C"S*<��e]n�H5�����AЏ;�t|*r��TU�b�P~��?����0
i��ۮ���a�A��z�u����os��� �_�`\��Sr������Gݓ��Ct�IR�sٖࣂE%�{�?�,�9tx������x���.ϰI,��^�S����
�N
+��'
7ح�r5>i�E	�>�\>g�찙�͓��ǿ	�ĕ9ίFL��Tyk4ގ���OC�T�m^� ��%z���ÃƇ�ӡ|�$�~��w�"�"�/�%���;˻z&Ģ��y���oz�!i0D4�HA��;Oݹ�G��YRYS���s0
+.�@ܟܴ4��G�.�����m�Έ�k�9��� ���n�M�vG�ː-롴MF㜊����[��.чvE&�����d	�l�^Q!	~�b�&<Jd1SҒ��*��͞ˀ�h��N�>&~�OӼ+7ܟO���(T���'
9`��t&�A�������c��KNI%�����F�y�F�+�M	|�Ghr�Qa�C(���п���S�LX�r>��A@�腀�F�r�i ���8i �z�����$.��xMD{�eː���Y��]$�B��e��Gf6�:=�]KPdO��l�G=�PA�����a ��5uo�UJd} ��.�D2�_%˕ɘly{n��!�Az���\C3U��1����6j���]#a&��Ȑ*H�ɶ��J^վ�Q*P���(ÆxD����w�� }�4���Y|$t���`!�Gd��"��KjA�+��&^7J�|�d�G�^���B��HMe�X�[�����CM(%6�梷CZL3,{��u����%]�q�k��gU��o[����[M�Sa][w���P�r$�7GW@ !���T�_X��x��Q2�5��5D�l����ѫU�e��x
u��e���I�p�%�osn?؞�\eK����+P���p/�P���D'��/J��!�-�ǓU�l$c���u�ՅTaw�	�JXD��M��cS,�5��<x���:<�=��&&���麪�i����j�J�a��8�;y��?�	���<��Ƌ�y�&>)?�#�\CLb=e/�����tݟl2�2�|� ݳ����xh���WC�L'6Dn�3G�A�ؖYh��]� �VS�����G�~u����4��sz�A��MUm�z2̰�rDߠ\u�/�s��[\#��2�SM$��+�cx�RH��6�X��D�o�-��{��T;3N'��C(�/"�[�ۜ����j0��m
 I���u7t�P�8�����j�@�l��>����$Ͽ)�@?F�X��w5�����3�Q���	�aD�N)���)�Y���8q@���s�� "�DQ�abeuf��) ��[�7���U>z��a̂�;ٌP@~�2�����\j,(y�;�/� �63�?ב��9m�����+R�"o���	mb��-E]1��G���k�u����n>j�x��7��0x��*/�h� ���#�9�)����3��� +�q
td&j�v9�*�@Q�l���#ɶ|�uM����f��l�@�O�<�9.��O�� JHt��eqQ��[4^%ݝ�!�޻�|d��)����߲^@)t@��T��eF�Ұg��n%���{Tm_��6�KR���懦S,!a)���}eQ@~J�WwB�J�E%�Tp`��K� ��R�&2�tH8��dF��ښ}��:X��C��l����v�k�E��P�����A� �	]�ߎ=l��W��,���3L#-��uh�ʘ��#JR�e�o~}"d��p�9��s�(7�@[ǝ�����9}nxa�.���%4
�f��,Z����d#	�t`��s�o�hWvU$H���Ķ7��07����\`<�?����m��袷�9���]zb��>���Fj��?�����;|�㬋!'�9pcNRgK���3��<�8['���n���L�#��g
���6�fR�(�$������R�f�'%���P���z�)2���Z&@��k���(��<��$'�V�Ȥ�?˟��?z����Q��}\W�ߊ�a�o@PGu��P�9�R����S
̦���@���]��ֱ��]:=���msx�9�,�հ%%K2�V^�-S�ܩ��:��6�Saφ̩E����r C����w'���x�A��:~�V�肆˻ai-�zJ;��]pP�3e@[�XR�f:�'��x��1	�4`����g���S���c�$ 7���HM7�����$��!�>&4n�R��zփ�'?[�2���X���?kIҚIPؿ��=�h̹�cC��Q����g�ߕ�_�,1`x��	j���p���������p��O�vl�.0�����H ���-�ŀ.'�}��k�N�H�����d�#�Kh��s�\����d�����mNE�T$�}�aqD�F��$�%�������'e<d����u�e�|��UW���2� �Qىޣ������������x4X>�x%]f��|pnN�^���\��o�(R�������^���������N�� T�b*,�Vn�2@������?kh���r��+m��S�����84$�r��0V�%�CV�H.x �ɾ�ç�L3wS���>aC�@�a�s8œ+�¬��~�;��Z�S�-%�|�b������E瞱@�gT�b{<D݅�S!���\Qj�v��C=�U�Z�+	h�Ry��;��:|��@9.�3��xAt��D.�'Qx���;8}%t�;���}*9d�H����w`�O�\f����Xq��Ӈ�V�K���As�,�� f&�������n`������E�Z�W5:*�����_���ǎ���`��$��� ��7:s�%�s���k���9���/1�������[�ڈ?��LZ�1F��*�<R�����&�m��h�J3RBL�@n�.�Xj��������A+�>��r��;��o�m�/6A�eo<���{4�u�j�$�I�Jvzsj�/Q�ժ
�s�Ӑ����=M��|�+��]���D��q�!����Я�7��ƫ[�MeuҪh��t����M��K��[�^��e�}=\7��4�c�G�5��� <Wg`�x	4M���B�����d�J[	4�Xj;�5��P��&:v�M�7=5���PE��I��`�ADҗA]�
��;P8��T���/�G���
�H�&���Z�+�b��� ���dqɞ�)��:G�՟sfQ>��O���0vD�ԝ�.�R�>w���P�E{��c����T�x���jf��eE�9:����E�Wl�"�]�rq����Ց�~2��8��ks[$0Eq�=�7�m��p�U��$��ɼh��҂�D��t<[�ynXl����Rs���F�ށ��ù�۩�~!��{�	gmb�ܨ�{��NPC[�%Df�o��gx3��C6�[jwG�8$�% ��m�}+��շ�KF��&mE;�á�dW!8�12���7�9����?WZ��8�-3wVO�[NZ��,��;S��u�^��)����-��ߵDGN̵��vW�L��\���*���.[�)�A"��x�4P:�# i�h�(u�z���% ?uRv��}2&a�p|��d>T��;�̳��to��o��J��F�3���a���!ˋ<�)�����sGR.�,|����N�6�й�J6^x��=��N4����'!���g��l�|�<��Z���w��A%\OށU��̀!��\&L/�b�Pbښ�"�R31�#�t�B&@8���.�����,.��)4-8;�Sh��v�͢#B=�*��ntt	�p�U+~t{+a����܉�Wv��n#M������ϩ��·�%.?��ժZ�~"��-�%Q�U���쫅ҳ��$��b0�������}�_�����s��g�׀�������|���{��Ĵ;��v�v�=�,%�ŉ�r6;Btp�H��左�=�l��,����p��\��K�9 ���?��D͂�S�×�CT�G(>�K���I�K�<)�����0͚�ح�x�[����AW�r꛻�r��i�4�mջC�ʸk/H�U�W��^e�)��{�R�&�H�z��6����9P�IY� r����U��m�G��g	l��@��Ik�݁�z��P;���3|y ���O�00�3���tJ��ٝiV28�ԉ��'%N<Ձ��xx*��0�0�*O<l�u�����i)e��0����VMF�v�a��Vx�- G���-Z���9�,�?i^7����>�XW�,����O��~���k��v������Յ�96픁�L��xy�l��#�p�c��&P�،g1��Cz�d��o�GK�U�� ^]8τT��l����C���5ΕJVm�Jb1Fr�E֘����c//��ę��/��(:m���x:���o�,�c�p�/���%F��C^?�!~h�o9�8k��������:Un���֑���E|P�q!lv�cvgSQ ��2� �,��=n1��I(�)�Q�I�_�9��^C����W�*����{���F1����\�P��*v!�{]@&\=�,ps9�I:yn5�Ӯ�gi��_�g?�%��Uq@ֈ��sL�D��+NLT"�=���L��ǻ<�|�3�o�뱷�� ��6i	g[h*���n�?��cJlF0@H-V���x�֎��M���*l �F�'&R�+F�rv�k��Ng?�78��D����m�q�ZK(q1���O�+��,<]ڷ�pF�i�[v�qh��M���5��aRc���U�$�*q,�~�g�^M�Dڬ��_x$Y _h� �HV�A%l��a�4��P�8�0���6�s�"3�PZw(�:�����F!
��$j^9��	�1�XY-�������MC�:��f%����|hl�.�~d�� Ot�\&[v��
�k�wkN���v��k4%�n�@H4����~~���oer��{��8����B<���'�P����SJ����c[WAl)%�#*3�1��+���>=F!7(X
�L��V��R�zm���8��l�� +���C
�
�Nyf}	�n�m{T���O>F(<b���u���T���%�q�K�`��v^���*(4!��?��L���_�b��>�D�'`-�K�J��=������4�T]��/�{��w��D
<3��Vkn�u�6�t/K�J>�h=����鼃 � ;��\���$�u+J��s#��w�{�����=����7P��������o(�Sa4�0P���9X��VRKa[ ��+7oݼ���b�jc�p�Q����0�!�^��C�N9&���Y8CQe ���b������x�������Y�K���������_X��T��b�C
7�i"�UD������RF�us�P�1a�&<��m�6�n�U�%=R�1��T�.͚�$�pT�����X������UfJd�����0���O��O����۞�dYǞ�7Llu��SOT�C;B�x���u��C�)��3
u�{7#	� ���PQ%&"�	'�:�%�]�N���tB�y�,�N"錱Qcb�A��34��]3c ;�Z(��٠���R2�KW�lx�q%X94�K����4X���.�}�Q��!jd��uI�oJ�腊*��F����S��0�\gͲ�y.�p{ȿ���.�D?k�Ϋ�����k�OS��F�C�4�^�)�$��5Y�{�7��Xt�����>�o���JFi��S��ͼ�o�Ҭ
|�|����9.�/������<b�:���_Q����7�w�=ߝ�L��A�(\y9�,�Mcum[��  =�u�:���eF�)Me4G鲕Jb0�}��T�� ;�	��p`V�wo��ԩ��3-��8�Ji�l
{�c8�2��;5���i��j�Q=b�-�r6�Q�C^��3ρ���	g"z~��#�"�������@���@������؟��T�td"�������p���b�Nu�'(ڞm(��8�R���&�`��q���4�iŽ��w�L%�ť��e��y�Mp���P�\һ-�<i��'��'�X�A�HpJ��?�׽�H�IF��`�o&�Rf��s�[!��9�Gm:��DJԂ2���ﻶN]BH���?ϼэ������苙qI�IrTy�,[���t�,�	�r�=5�<�k*�s?�<��R��������Pcu�q����McOTOdL�KS$��H�U����Y�O�����_���&<K\�+�6�eu��4��}"�#M�P�]\5��� �)Z��	^0���%��9
�X)��10J��h����6���^6�Mz��}5Z+�t^m���K\x��σ �z�׃a>�47gU)LJx�Ǚ�E\��dR�����S�x���� �p����"�g��G��F,?�q��t��|�\,�c����}!Z:��3�� ��Ĵs���!��É��k���1c;� #�?֜X�}y�
���86�!��4����F����)�@���ߐ�h[t>��Z{�|qVI'��e�g�bL!ۚ�[��)z�$"�o��N^T"'�q0�D�����>���e���>S#v��=h����=eI�L0e��`�0�f�b���>^bH�T=5M��e��˸$>�1@������n��+ ��T�33'I(1q��eM׮�m�uU���f%��*����T��J_�j�7,|[�7S����e~\��S�%��Ui��e�o/�Ǉ��ɘ��A�Pf�p�ֲ볹8ؤr��+Mo�ңUJm���{:`�'���,�&�N��:����鲟����{5D�!a�yٌ�"��P���%	��G�{�����T�'j"���g�7���6,n�:����b����b8�6z�u�k�(u���,�NE��
gC�g��{�r5"Qa�eM���b����΀�;z=Л��Z� 19����|1��jE!�������k�~]� �a`Q�&&N�)�ߪf��&B[h�泒�R���7���ܱ^�*${SW�E�~�d��9ק��K��P>�Q�H��{k{�-B��Sn*���.���Ⳛ�?{��"�&�p���9�.^ؒ D�8SV�jõE�V�&.���i9�W��1��)�}�&�8YZ���xL�%gb�5�~|�)�2�>�P#�vT9�_�������
gg�A6<(��gի�C�4�4��;��g��Ig0�ݿB��_� =.N�X6Л+��pۛ�w�����om�,`�l��o��* �������p���F� n��B>�i�>����|�ز
���p�hʋ>nDq��M��l�aP��GY�8�3(C���#Gۀ�H�[������Q���iM}n_�0�Ip�k�]uP�����s� 0<�K��TZ�����l+�(�?��8���\' �fY�u� kZ�F�86�3�A�3n�0��N?5�}([L��s@gNO���J��e�:0Ü[��$B"��VX�Y�X����.:��Y��"�.!�����tg/� l���d���������d��y��Nۈ2N�%L��e�{-?���o��7��X�V����B|��)��.���C�U]��^4�%���g'S��Fy�BwC`��B 2"��\��}ɒn�W�N�� �I��	��N��O���⓲剎U���Cxf�f�|�>�6Ợhl)�o�&��tNi��DN�^wh�6
��A%����8\��8������A�4!:4בP2���BźcT	E�ԢI�[�/�&�'� |�]�(���|s�fW�0����z���������36<֎�c}�<���j�}�^�+����{�]����/~��ev j��4f�4�`%0�0�/��U���L��M �K-��*�~%�N^f�������W��@����1^�"4,�W�	��BX�L ���o�O��x�"��F�����o����e��k&wZ��B�ʖ�2�`i~��X��/CjZ���RD5�Y*��Rc-i	�4�.����Y�(O��$�j��2�ң�
:���|�6�HWPJ#��r��If�^ۢ~�Ǟ��$�3lY�_Z_*XK�>(S0����-��9!��U_�?�2y�Wy=m��d��^���g� c��Z�!�
8� �lN�Ȁ�n���u�0��Yh�y�r�7رP�� ��#�ˣ��m?�nh�p�ø����~���- L�W>]z�5���Gv)Ԣ1��e"dh���yR�;ܢ�BV�E��3�H´?�j�J��s+�2�v~OCZ�*����Xٹ�-��O�5�D��6�$I����k"$r��c����Pz+U�NF7�Z}ͤ&Uc�͜Ƒ;s�J_Hfj�Ơ6�=(�0"$ndezPI��B8�Q���?�ϙ��1i�7�l� Yk5oJ5�'��7���l.իzxʞ�*51c#���@�߂_�g_h�v�bߜ���O�ts燭��2�v!$阳��p	4��蓯��S��s�������֜dͬe$,