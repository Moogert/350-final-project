��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���D��ܨ::��{:�6�4�'���4u@��E�o<#��|��h%w��П�M�:�������6��W����~�H-_B�s+{�LnR���{��q��ʝO���
	Eݴ�5�]-l z�2�zK�Ԟ��� �U��F�Ig��{���;�5��`JJ5;6�M2���Mn��-�+󯂀C��U�
��R%�����oxTO��نw�dI_�� oF]_#��o�o��Bߋ�֬�a�.���H}>w�?���~��i�m�]�����p��s@�⋓k�T<�M����^�L��-����r�V�ހ`4�	XWS���GjZh5��V(�Ǽ��mm�`���3���ު�P��1�36�L��>|̢h���	�àmK��]���	�
M�|�9�d�c�N-��A��5����TʀY(ņ �g摽�����>�I��mnꇊ���ʙ5�uu��IۄQ�׋�VR �˙� -��L�2~{�����:���J3(���S�[a��IHƬE��s�dԗ	B��@��_���ja�+����~��@^D�7��wQơ�a�q�����<�n����������rV�S�X�ۿ��@K�5�����g�RscE�U���6�'Y��l�d�H9Ֆ_-(Sh2�b�T��X�!�EA����E�}i���ƴ~c,5~r������Ĳ��?`�xx��cY��@��1��v��A@eAooz����A��o#V
�g|�C�ު)V�	qxǞr�܄��7px.E��c	\�f�X�^ B�s�m�g㹿3e9?��q���Y�%��)��ɀ�@(Y]x��Uճ܋"5��*��R'Hl
w����$�K�N^93��3���s3UcՌ��k�G����3	� ^D��Ў�:o��4���
"��	خD�|�@Δ��b5��Ԍ��oޟ�#��� mf9��ߊ�iO�U�=��A��?���1K��;} ����]��S ������ tM���T*Zm1ި���n�Ǻ%��-yc�����"��n	x�@Y��0KD�%�]�K@W�(c��oCķ%� ܆�s��J>�~�}ԕqH�ޅ�) 8�v�1se��ms'C֩�^�(�Q�"<�ox��s��JB�\��ߜO�����uX������9��r�F�u(��L�B�'hU{���%��Fi#pl`BkǞ����m]����`��h�V��~X����#y'ǘ�*��|_��Wk۬d��Ţ*�TC2?�s�ɱjF)�=��!���9� 卒�@��=6A�MA�3�i�&Eq�#��S`Һ<�_t�~{gȦo>�\  W\H��aF�X488ح%<���"p�������3��"���5Z���lԝ����Dn�}F��0����ib��;��݊�퐕ҢF^��ޏP���5?�Ě�Ƽ���I?�=c��ʒ�|z�K�R 6�b��w��zu�~65D��7O_f��U�*��O3����ʡ�zpi�����u�@�Z��­{X�6`X��TS���
�[���+#�u)��R���A)�2�C�M�$���R`�5���U@�&?��Y�����Z㲯��,���	��� _T�ܞ����m& �9AL�_9��)X���вB��@�:�8VAEX6��P$u�z/���?�1��kG�����bԏt��m��pX�E�Z�%����y#a�vb0�ѝA���f���vm���0��zɑ�j��3���j[u��TV˦ם9��h�a�@��&�t7��%<�q�%2��u����{ѹ�^�7�J���ٗ���J�gU���N�*kE�N���G��f��s�O.��P6�B~E��%Ky���aՐ��)��_xF3\%��>J�7�A ���-B���ˌf�_!U[���#����'P/|���U�X'�������ְp��!�涱T��*C�
x��xN���v�����]r����.l>�l����h�-麌|LOD����o}��5=��I�-RR;9h{ºYu�`���
,p��5��"�|5Ad;�Ұ���o�c�,�=���ʹIB�D쁣����0�<�f2�F�H�Y݌��n�]�C
QW��9%Y��
�
/�9nh\ò�_��wn�?j�n\_��T�[������A�C.�B_�����>��\'�rx��3>
��$��LS�B;f$^H�>����-�=VS��~��0��rQ/t&$�L��BOk���_G��L��U��#���$�}F^:����7T_荧^f(�p"��-~g�pb�����~�ҍ�L�)�Ձ6�?��̟MQ��Y�>��8&k2�e��fJng9��ۨ�՘@��Ǒ*u��:�eq�Vٚz5������J�
��P�K��$� ��v�^X�-R�3_�)|�&�LpD����65�Kmg�&�~q2�n�ti�,u>U��:���'���~w�БN

HC�އ��>����T0� X����՘ކ:���#�K!4��������y�mg Z��x�D)O�f�>��D�Rs�)��2Zl�
e��W�� �F�>��~>�8��"<�E�/�a$Y#��l���9�0��CaF�O��F��G.����G�؇[�Q"�����bR�m�@e�Hm�]5����N-�Yq7��X���I(�\���ˡ�H��_y1�]/���pG�h+����@&2��_>�6��a~��B����R�Z1�����)�9=�{9	'g�"h3Z���ު�a�ː�0�*�C��u��)0����q��5�&�ʉ��]�p%����HCEW�䏡�b<R��pԠ ��M�e�+u�3�Xe?F�n].#����n��O4��P��4��犛,0�K��H�!e�H��M���#s�lM��w�'8l�|0�P�V�r�宽�j�����[ñ��|���H�;�rtB�k��	��AP�^����w��sZH �x��r[�s�����Vrm�s(KCc,G��ٖ4N}X)���e}�4�o�i'1��- UK��7(�:E��g֕o�)L��7$3�2wf ,�l����*0*d�Jhъ���S�]�h.�>�he9@��}x{
K�`���n�o}�7�@�ǿ-v���x
�-�gF� ���q�F�O˰�J�B;
����JW��o0�d�D�gS!��_3�w{7|�@~�������z�Hx�3���8^����@��I]M�똝z���K�9:K�&���-&kD|����`FX@�&�iT��2����jٹڤ�y&�?�
�Ƃ��Eĵ0���+0�������$gOD��f�s+9R��������#�>Kα2�������$��SC�򗔒x)؈'����с�S��t.K��-�������6�(.S��eQ��Bejbv�ѵ�9+,���p[��E��.���tߙ�R��|x���U�[�P��م�`�Ι�Tn��Z⬒X�ʃus�=sѝ�IU�P�z�@�Λ�Y��3R/x��<��ϥu���.?X}���X�rМ�\Îѳc�$�9@i~u&cM��?�J�)�<LO��B��@t\ற㼒�8�V詘T0y�ÌD(�-&Q����[_��͢�5n#'D�z�<t5���*�G*��F�:	A�d�Rȕ3r�M���O��i�řchf�o!��櫘]�ڛy�@+����cw�|Yƈ�V�gw��9����ajR����^{�!����F�����)
q��J>�p��s� �NqPӧ$h���\�O��%��B��Ԓ�f�j�7(��3 �3\�+{�]X<*[rB6c�'�^T��U7�9A�j�
�&ە��̐��Kw�-���v/0ǾG��n�����O�6g�N/�}�/\��ϰ���㺫��sN����(#V�]����G�i���مuT����,�t�E���?��v�!ջ��XpS��@Zup{8&T�����_���:V����:^jAX.Ϥ�r�4���'ᚋ(s	�D��p��Z)��M:8�B�����PEu)
�i�=_E�B�j�#mGƷ����>��&�Vn<��� �xf���8?'��ٵ�E���Q��Ic�س��Q�yK"O��-��~o�i�O��Dv<���2��	�Y�}ٍ����(��X�^�<� x�G+�U��Z�-z�RL?<��`c�G2җ��׹ug7go{	��>���Q֚
$��Pe@����XZ�I�Gͺ�7_6�~�
�#�4��}�P�vU�آm��\��!��<ߪM�Q'h�|�~�X4t�@��/9�m$�(�4�uю�\����.;�7��v��1:�>�&�3���E�A��%(�R��]%�ga���o!�E*�}�v�>��w����w[hS�z�ӗ�C Q�o�V��&�ƈ9��)"�>���o�;Er"�Q��rcN0p8:��M��^�sR�"o�� �>#zI�[\'w}�/��7���;����)BVh'@	�֍�n�po>R]�؆^�ē���kx\u>�1l*I5xO��ŋ\�ti���YF���F ���@|&M���S$~.�=E��-&��N�rq���U�8-�aU��H��v/���S�xH ���e��_�'��[��U[����������ÿ�CLz�=�1Y������K���-�&�,����/eK��=z�X���~�����|��x�S��.�Г{n`��-�KX�T��<���|���JdgT�O�_�)Żm$e����8���^��txR�_�y}K���} ����SS<z���)��v�� ��zؗ۠����h�Ne5)$f"�K�Wϛ�˕�v4H�1��6�����[4��l�3�����8�o��<,	���[�Cͼ����Kq7���̇q�}��6�ul#'�a����s���w�N�a�?]�}P��%����\f;����e-��x;�{�y�)o!��G���X �-VG����Z��vp��=����o�i�n��ݢ݌i����_���'����lmf��?�Cot��0�s7'bw�m�)�0���Q�}$���Odi~� _�A7�泣b�.�����#	�ȲP]gͮ��sr��a&�9F��g�.��/
S�/饀���ٌ[�작�=��6^��~�qP��9��b���(������N�:���ӆ ��tP֠�(�CA�-�ˮ��PJ�̎h.9�|��(�2�0q�{�C_ĆߏuwfyGֆo]�LX�$�Z�OK3r����m_㧩j�a��79�^f~����º=� Fƽ\�����e2���k��04�dD��O��e���i�@�u�ܯ�>�����¿�y�sz+��R@Z��yI���h���824�{����GW4���/jg��*��_��G��^N�^_�=g�d�ֿ���)[���Ui��4�׎��:c:��[|1�	��ۿ<���!��O��J'v�q�Ӓ�3�;�{z)�>q�r�2������%�h��)�E��]b��G�Lo�]j�`_S���%&� D�%*l>��]�٫��a��� �Oh�~g��q�֊+#`�mJ��G�Fܹ�k�m��@������^� �)Cp�G����ad[#u>[��~��m>&��GQ+#��|Trr�m�,��]�m�+Qn���[J��P�b`D�
<�U����qn��*VU՛���u؆���7Ŷ岨Y�����7t��YG��&)����p��{w�a
d��G����vo��Nwc�:�t�♓ۦ��gvD̊��`�l&��ZD�{[��#o�G_$��\���{G��J6��'��� ��x	��ъm^��I (�p�y�
*9�|؉��Z8�^� cJ����61Vkn���*��EEJAm	�o�3 Cd^4��խ��1�:W�sH�ܕ�7�����p����`>ǂG:�󅺃�2��2/�2���N��_n�X��-�u�5� �V���n�� ���<G>u�%�Ѫ��'��J(��=	�MK~��2A�rU��>�:l�gCE+_�
]�;�?d}DJ�ț�ߢfc��շ^K�tUU�u����'�}����2PR �n�8`��ŉ���z�際��`.�Rw�Z?3񆏅7��5���G�鎺�ߝG�ظI;g�ڀ�)�L*�z0J�+�QF��h��+���r80?v�=��v^���@�9�T��1{5+���
����?��7��y) ��ƯJ�Mp���j|͛���u�T��YYXX����$��%�[��ݖX��X�+$~V���F�o��_w��� *A#����THt�0���	�w�Ϩ�K�uu	��{�ţ��ː�fq����Rk\���O)=�^0V~�J��%�{�Na���*Ԣ�c&'K��Zo0y�!��58�i_G��%{XȂ8�_6O����d�'[ȀW-t��XS�a���b(H5�����w���,�R��q�2x	��%ȇ�\��m��K����-\{�(�t���^J�r����ᇥM��0��0JX��0��Tv��ٰ@��˱]���jLv��q�4���Zl3ɩ�|ܻ�2��]�2Sb6g����W�nu�(���C*��(�w ��~v�h�X.�q��4�ST��<kFy?[�Z�$[�F�K/g!&�w_ٻO�&@��֛6ˢz�D�j(H��[�8Nu"D� ���p�>����KnA���!ւ�J��7kW�9�qt�C&Z?gD΃6�e/�`f�~�V����N��O�T���ӱ��j�X�]�[���I���
�7�2��[~r�L@��Na��;LF�L����ۯ����Bv;3.] ���d�E9hy$t�ޖh�@it%^�!F�C��`�ǵ���J�fKܖ�܇�
�<��>�nNێZ�����l1�9ͷ+���� 3!�Pn��B+�lMx9�D��埑�Rq+�f�~�R�A�R�i,���Zά�n�:{U.��|�&�Y��CZ�B�]�bPt��Ԛ �P"�gO��[���$oq���Df��ƍ)��>	\���!'����\����LsoO�m1Jzv�����,���	�L6��R�T6���,�����;���C����c����cd���W�P����Pe~��Ci�q���ܒ�9hd�vM�3sp"54#��w鯸	f��t3��6fCN�j�"
6�s�`у��o�-�q���b-Q��)飼��%A+���n��&�)E;�唂%���C+!�c:��Ҋ��y�}��{�����֖i��U�ޥ�'�KϺ��LVi�i��:�ޕU}�C90�[T��I�8�(��Wtmqz�q�<~T'7آ���xh��2����ZźS�"���b7�?����a5�c����p� ��.XH��"��x��V�-Z���(�w��ƍIx����g�B7�ӛb��,�0��M�q���je�'���t�+q����,PM�|��k^(�)	bM,K	M��i��xbk6
`���Z��qk�>t{?�agC!\n1�X����i��m�O����~�Ov�i�ǐ�����ߴmf�R���3ޤ?:{/&M��u��s�3�(	���7�y����0Q��[�Z�t�IHCt]�_���0"_�_���� �2wf-���2�vc��B���N��g���N�&���U������-��!=��Q%j��$+Z��Q��2�t;�y! ���4��w9I��$��.�H�7~��r���g��=Bp،�Ә��k�(��~I�jݪ�B�/�ͯO�u���e������͜�"qZ���aY�*u�K���*rwL0��^�m:�H�����7�ݽn���<�y\H ��J���"h��r_�b��
"�«&7i�ё���ee�k����Q�Kr� 4���MT|�7��iwpg�"�����dyG�X_WD��2[Q�m��_�H_f�a��.��r$��ڋHƊ�}{�^��A��l�*�݆}�['�:Piǝ����>I�\��T^��l�~�(\E�m>�����&��V��Ɨy��Pu-�+�muf�B�ٻnm��`����8����L��n1$�-7�4o�M���c>�>g�g�Gf?,u��՟DY���Q$b\����!���v�̣�t��?O����I�MmC����x}�(��&"�_��>����F��0V�j�]N�|��j�����Z-�~����S<(�_���#����<-	��s�W*��rH�ZJ9<jSA�Im�x��f�N�Y��
�/��[E��ibWP����=�V�br�\�N,*_��G	\��Ո�ž�����ҍC�����N���4���}�Dϻį�Xq7>:F�+�hpP���#�$�m���;V�}�Ze+g��JuT�V���i�f4ݛ��?�ne_6�t!/�/��M2����I��7M���c�ډy�/dI����2`��yN<��l+m�7<xԈv�g����ޡ�y�� "ԥ��#&?B6�6�;��A�u����!��S��� >CwL�d__��j.?��w�W��lC	GB8�Y<�4�ie�oBw����r���~(A���%�{�ެ3�`6 (W�[��LpN��EDx���+�������<��aԭ���s���<{օ��!e
~2O���:Q��D��V1A��'�H�SD�u'��^۵�q)<��G�=R�50��׉����c�b��P��0^�QDٌ:+Bts0p�w�`g;}�3%��]��ǃ�D8��-���m5yd{H �� �~����;I'aDP��N
Fy�&���f�A����N�s�ήX��x	>��c�ą6R�R�����I�Hp��z�D������ ]NB���uA���͋gv}>hJQ��[�(Z�+���g %�9�pU���ENk�2=*$��5G�76�9i����������K0Z�g'Z&F���u�3�HF���_� Q���c��'�;��br�v�e3g�� �y�c����422���2SW�+��eJp~�.sR�5��8��,(v\�����sm�*��q��q:\���c�hh�ZŠ�v���y���Y����T�D��Bi��ӨA����O���(��IS5������I����%u�/Yk�R���Y7�x�CPf8��7�9Y�zJ�($�2{��FZ؁ƌ{t�\���I����54��v���ވ�it�~H]�o=��I!3Ao�a	���~	[�)v����Y��f4&�N��غW>+T\,ra9�i��,�u?��C�yIg��W����q&�H��7-KS�4�[ӿ� \CXJY"�>E>A$���q���L������M$���"��]�Ik�gĐ��i̗t�nB��+�3�C������k��"pXFni��)�
�f5��I�&��*Y��Tc���H��Oժ�inV��6��DdW�������q���@ǚg�g\v%��a����n�XUYV�Կ������q����V%���.ȑ܎�m;� f�?N,'ec��ߢd�sN����Ķ�Ү�6��O8��?� ��f�(�`8�Z��i:m�=f�<N�ɿ�L}Wvl�Pؒ��	� �m���l0*�z��18ŋ.7Wj��7b��l��Ca&�P��[r�����{#����`D��.
�m����n4�N�]J�U7�ck L���D[]�#\�����щH_����|0Ar�/�G��J)H������G��:��6I)`-�!O�eG��[�������a8L�c��	�~��&����-+�Ⱦ����8����*�Ze�o�<�φ�v{����i�i�w�y�m��
fE�d����/Z�b��7B�$.���D�BXԦ��"w�=.��D|
�G�׳��N^����Si��.1X�l�b�#��̆�� �!��Ք�$�܆��:�P<]�lN�ؤغ��8�8�x!��Ev41�����b]��t�\�m���'Đ�	��O�BŽMb�»�~�s�hX�h'������K��g���fRFG�C��kxs�l0�H#N���y�3�D��*����`%@qw�X(����	���t@�D����s ���}ձ� �B�@�(�rx�In��i[J������$��O�k��#���2�*_WB�&ܠI��tvX|d2PT�����LDe|ʍ�/�&�Y�{�W�.
4�����Zǡ}�w�������]��N=�p��˧�4͵����tFx�M�Ě�}67�d]�k� ��d"e)Wj��,�n~;nu�M�c:����C!�^)U��k\W�G }A����9[sOg��y��x���oZ�IkM�T{On93��펠�Bl6������C$�*��(X�~��h��0w��	H�{@�Á+���8_L/nÙ뺷�5.-&����䢮�'�Oԙ��TPQI�g�3�����1�����XZ�P�Xў弑Ec�u��g-s�6�%�Ȟl�b˨AAK�������𘶄�0>�Qk�ҹ�{�����&�Y�7�	MEދ�(��&���CFzS�o;�|X��x##H�eE��T\������|�?�\�x�7�pFL@���c4��3c�!e�n��&i㔏�%�	��(G�;o���B�/M�T�4�T�@��-:ܪ���w �Ȇ���Tl��u�/
��0*)��S�Sp�O5w�����g
{
1�T��+���2��iv��x�G��7��(DM�/���4�g8���Z_��k�JO� \y4�g��X�C�O�iZ/�����s�\P�`���B�ҥ�IEs���CฎǞ-P�(Dj��'��ՙ^o9��PM��#k�r�0��=l>���/��;�UQ���I���
.�p'6��U|�g�1�Z� �[\HS��*��?�������2��o;C�](�t?��4:sjMA�Si�]�Mg'���x�6j�^-���1L���M�h�=���F��Y��2fi� �)��|)��2��J�C�Y��Uأ��������3'��^���t�A9���M�!���A�l�;�mFr���9�#��ہd�����匈�t�M�<��X�*S \�,Θ�<�YS��جK�±p$���`�ⵗ��o��]�^��I�L��KeMz��_���K�o�'vzZDFPOֽ�7���僗i���9d+�g�"��Dy�_7Rﳪ��?eץ���O�!�3��kJv�]��bçE�F�ڰe���`������m���75�TUUe(�d�0(�o0bT��n�i�a�ƎǽT�p��W�C%M��F�j��~�g���ڴ=U{���[��9{��-R��?;k-��^�-��c������'�/C� �q�r�~�e��q_в�~�6���O�"+��(�e�=2�H��O*�G�̃�"}�`D�ۼ~��АT��[5����Gx��3�!Yb,��g���9>�v�m��T�jI����Fzf�.��6o��y����=
���B\�����b��<(��Y9�7�9g�j.{�e�*���3����A@�lJ����=59['����pr���b�}l��xk�oF���k�2�)[6��u��eġ< N�i��������kA�8�;�/� f���\�Y�"�,N-D>���9�sC�5�t!SI��	�J@_����Ϳ�E��`	z�?)'�:[ĤQ9Y�!U�=�KM7i�<�2(dLhy	�M�~ <t�]����$׳28���r��:�qO�@�/�?� h8�ȃuEj�CP��e��KZO���H��>�KE�zT����=�Vm��c�Djcaꀴ�uq���Jw�s"1�<