��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g������*���Li�ĉ�3���R�\��0}��N��i�b�QO3s��N��㐝p�W ��Kl]���BI숹�(�a$����=ZA��Z��<e�TrRd���t�o#��K7�QX3��O���� eT�2j�Ŝ�5�| ҭ��\���I$��Ng��^�i�cۣ
,�P\��B:�CN� z���� ��hc��GB	:b�[�5Rf���il��.Q��</4X <�Z*�Zv[Sr�w�P�����˘��C��\&�η��zR��bA�AE�Y�w��\�7¿ȣ���p�A
 I�!�C�^�@��r�>����Hr<Դ�K���ﵘ�Q��h��Z.���${��A{�1��+`����P$2�W2h�ɖ�K�z3kFu~�?��!o��)�t�����-��Y!��!hr"h|b�����̦�ɠ�v��arLu`�y��4x���y�h-��]��`}�\]caլs'c+R)p[n��m�۟�������y��,-�H"|���1����v�#]������P5Š��3�h�M�$9��yW^���1�Q�!΢�KxF�,�+�z�� �V�^z�k.�E�O���0���Ⱦ("����5�,���]��<o�^�f��P3��$�Fɷ	�GGH*��Ѝt��Y7xD���L]9Z����YOp���.�bJ�O-�5A�Z������:�8�� E?�]�Ă�D���FO�t���5��`l!t��ۻ����[
>�|����:�i-zX��{w�$?M�e:uc�*���帗���
w�����"�琿���[�z1�m!�D�g���1d��%k
/�wy!;S�6:=�����e������� g�'�h��f�r�@��M�y��L�կ�;�%a�nw49��WIy���ͱ��E��	w��t��ɀ}ҁ�zNI��.�p��sA#Ӄ���{8p��	��\�J��cE���d�:s��b5�o��F�"19b4��s�n�5`J~.��aQ�	H�᚟�������9���������G �1W�(j/0"12X#�p�$���i,��_������� �?w�]�B�7V̠�"�Hb|Q�\}:�3bS$Y�5�A����V��3�%���N�Z��'t�S��̈́��@�QX��c�YON�.���#��l�iĻ��n��:M�SɮeM`I�r蒫�,�ާ;S�B�xO>�I���`�S��RXS�^��*�_RU(���
�cAVd�gT������!�]ԎNcs[������P��&���+��q>D�R�ε�J���Js6���6��v�(�B�=Etܞ�f�a�K���H7݂|�<�w��Gy�vN�X�{~�Ŏ��{0��Sp�2Zַ�FI���{�[�ØԨ7Ƞ�3��kQ(�٥Z�4��*���w�� ��U�9��3q+4b�._��}���^�^�(3QH��v�#0�Q�xE�"E�,�`�'�6-��$>H�����Z^ʝ�9�MR��AZ[���z�f�sgk9���+��Q0L��k�i�5Ɨ+�'gn�7*\�=RapH���c�鴙
�T�y�����x"�G�f�3pt3A*k�7������i�6,�b�	T���E�n�W��P�E� ��#�s>�� � ��,��x��l�#?_=� �H��Ԅ�Ț�����Ȭ�p1��݆�Y�,	9�v�g{�b��}�E1'����aE�f���Rp�;4��]�����	O]�o6���Wf��2q�[�b"Y���U��(��㢜����`���#׆C�gy�r�����޸�qk�y��Ų3lxq�s�L����]���� ���Jcяʑ�<�M+�TP����N����_�iA;�:	G���n�����%w\D���j�(٣�`�(��! !<oYrz���ajV�ey��SD5^U̿��y2�;P�?J�>����
�z�e�4)~yU�q��j��8�UȐ�g�ZR83v:��sK֝ �}��3�SN���~��ܽql2��C��r��3-�#���� K-_,M)���*����*G$d:iEd��V��U�=z�@�l΋�t�(7��]�Py�$�憶c��{Kڵ��Åty�`����f��z�s�Y4�;��o��&&���W��-��2��u�K}Z��v��@+1��#̏_�s�?57:�N�N	�cahb����G�T=�����Dd#���V��%�52��z���Ȉ�����I��w[ޢ��7�y$!B�Y3�4!Y�I�!�l��$OHO�É�̇G�.q:��*E,ȵ�\ml�ȯ��>E-M_�EΊ���o�x/�H1�
�pLB�C��0��A�J�w~�2�s<g)�L�5���]�J�V�z�~F�F�Dv�c���Wuq��F*��0T��Լ����{[��l�L5A@9C��P����.�|@�����Ps}�PO[��r��C�&E�#t,M�'�a���+���>�%�R}m[�j�}�T�So��F� ��Y��K��.��6���CJ
/�3�O�h1�H���xp:\{~{,r8K�\��w2J/��3�� �<!�]�If�$ļ��H������hg�\�Z-3�h��n Y�i�rn�q�h�k�aܪ-k
?���J�����q1���@��	d�K`hȯ�p"'�%�ԗ��( {Z7Xnd��.�9 �X��fPY-��9r���f�[I8l�O�	F1� ��Z�����O�hA[���0�/6t�����H(��t���lԱ�����!�S4b����k���'Rm�p�Pb����N`eF���IjޭS
�o�(Ib��/�Ć�Vnԡ�}��B�V�j<��P[y�k��X���K�uff���D�}�9&<��w,�e���� |�v�O�\���������/_]�b�̄{�{.�4F%a�(��sȋ�*��E��b����[i��0��0@�\������s��"t�1X�k�Ə�a�����d���N�SF�?��2������J�z�P���jf ؇k;���@٨�Ʉ|��AL�_D#���#�o�ܕ.�g,7uѩ �3LQ��K\T��v���9&�ͫ�qţ����3�G�S!F���	� ¢2b�-�U�O$�n���G	��Co�W�|���{���w�̅���Ь���9n�6M�ē��?ؔh��[�O�T�F.	M'ʭF�$x#�b�f��엻��-#��>��{L7��� �,�ͪ^1��5��fo�@�<�d�m��ɴ���U?]V�$�B�@d[����h�������N?��E��}���0��X�jurĤ�Å�:9I��=�o��;�z!7�ЁџM/��Cި��9�o�e�\}aZ2��f5y�*�b���G��Uبg���`��x�$�35ƭ���V������WZ)z*{�D�5��$)��ʻXrk���x��Cw��źu�vؽ�Қ��j�L���j���i@��#�c��_[i⛂�i�k��]�6�����ێ�܍΀��5�gg<�U��/a�ɸ��y��=a]n�c
2~�V�؃.<!s����w��Qez��g]���w��C���*Эg	�
qb �y���	uQ5�Z�y��8! )�i¦�x_��f]�EF��n���Y(j���6�ϪX�kEkmx�0�ړ�?F�f���~/�@���(�*�c<e��rD�Õ�KxI@\�t��Ld�>�6�8�9���{�Y)Y�xO�pv[�����W���Z|_��X�?̸w�������e9�> ���ށ8��0�s��)�=D)x�HԻpK��d`Ҁo�yH`v��
x��I��<4������E����'�t�^�F�g�@OWu�OS��/$�М�x�NB����6����_�P��d!��� �|�+=s�R�*���N�^w<�o֑0Q����k�ey�������!��	��s�g�R�=�ô�Z& �D�e�.�2$ �{ ����2����n"�@����*l&A�b��3�_�{i.u˼s99���'LU�K_B8�������	8p
�G��a#� h0�'��d��E��=��zi�}WuW�-�J��!�1�b�{�f�>��4!��(�&��T��["ž����!��uSP!�Ã�5I��݇���*d�׆������D�L񀊿�@k��R�к0{�]iP��Da%{]�Y;�c�?I<�q.}�Ŀ��h�[U=C\������c�����G{I9�&E�dC6�KG�&�f���/�.:�e��ѝ�x}�u)Nk�V������b�'����&��K�S���Myۨ��\�	������=�����;��=*^w#u��8��'TS�$�����Gd��A�+����=��F{GW7Ch$�{@1������Ckf�6�=v����VB)����A���{��|���� 7(m�1�%G6��[\�.��Zv�6�v��:�&�:4$�������!m�3�m�|~@�����0(fH�����Ȱ|��mq2H����O�W��-��\a,�i�H���%��0�>��V�v�vl�pF����"��S�'QS��ϧP�s,�V�?��t���I���Ǳ)0i����u�Lƌ�SY�����p�9B�kT�=��$��y�f���
TꈵR����r.=��j��	eKG��`��q�Sj�h���$^�b$b�:�!���8�d����$4o�9.�P�"�@g�c��j�7F�$y�E-(�37G��{�B��Қ�p�5�F�F�+���}��~������D�
����"�}&Cc�-���U���^��t��j|u5��f`~'$Of����O��l,"�R��CƖ���
Z�(?�����h��u����|mpt�O��f�s<ؾ�B!�4'��c v�+_�Q�u��m?�/L�ϳ��Ē�޴��#�o#����j� .\���#T�����=b���A#�Dщc��G�3sؙV����w*�B����C���dhA)� |[jH9ݝ'���-V-����)�^��;o�5��X��IB���/���RR:����B8��קpwۀ(L��<m��o�Xe�'	���8�^�s`��>l���s�S?�2�-+��x���/�*��#G���s���Ė��W���h�H���<��K���5[�J���x" ��-$���3dD�P��{�ryVl�+D�"~}u����r�6�;:v�N�@AhYaی9��_M�|Ws��9�����K����Q���Rda�O�E���Z���\��`�8.a=y��h�Q�5sn��UD�{DQ��������}6����8�{V-�g���@��d�R#��qV��L�Z���T���Y��n��^l�E�%W�I8ɗ>8�e�@�H�ͯ�K��8No2�Yz���!� ���΄ݲ��е^�����]Hߢԩk��y2�3� �[�y�vN謺�,Ӱ���gf �
⁝G�?�
��֗�u��xCU��<Xr�fr������qA���7��&�񤙮��#�2����%��n��,�X��K�%��0�m�b�Ҳ��|F�V
��qT+�cBP��]�O����@)i��;�x8z4��C�k��#��f��ۅɻ�1��f��cW'Y�#[���F�F��'���()�����֪ؐ�!��;@��.�D�PT�N��&��7ٔ��8��R�N߂B�r��;�$5�����(��]�����r��&Fɗ�BӬ�]_�a�e^���J�o�����>༓}�X8+����cH\��͔@�azW����m�Q*���*)�M<���c�xn^(J�5G<nJ�f���2����&�z�8I��|�{�4�M�\�+H�O�r���Fr�h�L9�`�{ۛ�\M�|k3�>Z�ȱʓ�ISLF���V�ᆅ�� =��E�h��|˩0AjnAŭ�=��AĔ�)&���T�d�V�\ϓ�(.��"T�}���D�
?��H���<��9{��G�Ő·i��,�;� ��eRy7ͷ��f��l���ݘ�s�#ڧ=�땘�Ӵ/q������:^ӓB�O��49�T^�;�;��w�^�RV�W`Ǽǣ>^�h))˅����%�!Wx�8nYS�<�`��E7$�Ȗ`p����|�<m0�I]��F��Wc�]v��>5Kw��R٤�� �ӈ�!J]���Gf������&UN�
�vL�{y匟���I��}�w;��]�{�꫻N��G�hĹ4Y��#�we��e��P}�	�|��}��Ύ����
=Z�y2@9~��;�B &����4�z<�Է�C~r�FLV&˿�)�o��8��ou�4e�-�dfD\S�ˁՐB ������af���Z[#Ǘ9��W��SR��f���B���lh� �)P6�T1��"�P��Q$�:��F=SS�}4��.�@���^|���OWn&y�ߍT�c�L�\W��x���m� �){��.��g�T���=��c�elr���?�So0M�񨏳�?L��s'��U]���2�oУ�MZܗ��y0Þ'p��]��6�4�
0/[S�cZ�Y�|�ql��!���`t/�;�\+X73����mؼ�{0'�`���>�S���l�����琰�m��j��}��!�q6#��Șg{Rc -Y'��0/3b���y��ʎ)�
�8�Z�N
%͓tݘ(����|G�c�:&¢���5��wji�&CM"pw|ٗd�bWɚ�Op$ؔ�VlV�TkQ��O��Q�����z��x�5��˗�$��Ү�D�rAԮ����/?8�e�7.'��K�:+`�\�)�٧�3ὕR Sb��ҹ@yD8�C�8ƲP1Ħ��w00ؤ�{�՟|(��?z-�|�/���>K�]tj_KA�q*���H'(����}^��p�:}����K�?h��w,td͕��~�D�b�3�d��:�ђ�:Y��r�@o�#0z�K���UƜ#=�������N-O:�û�0Xl1\7))����--�{7�~����p��k��^L���#O� [��a�d����P��?�-΢[	��"�P����p�����* (�OD)k��~�)�I��U2��X��k���<���*��BWHQ:(�0dm�p1�پу�DtРNf�U��ۅ�p���o�|�#m��̦�)<��v�6W��~���~FE�e���v<K�F�oUa�mF����>]\?$��0�W	J6����/��X�N1ē��{4.�@JX�A� PȈ�n��L�4�J����䷜�H��"]D��	�TZ���n[�j�\B�*ZE��ɻC,�O2�~�!�ל{P�A�7*,��Cc��y`6A3@���5DN�2f�u1
z<$���C�|���[C�'G5�����|$�p0V;���}'<E������-<gdC�����5NT�ƌ��h����H�J�Ln�k�;5pqϡ�XBv���^.w��V͖`�G@��~Aj�*;p'		�l����l�?�m�:���6P�NT����#Awi�ͮR>�g�|�9�}�ar���eEDr�4�w��0��|kd�t�����4%��V�4��Td����������G��d��؋E0#y��Cd�x|���yN���ݳ��`��P@��7g]�Y
#0/M���z���
� U|���^��@�b}F���D+w UT��ovlc3B)�'V�!Q�1�ʍ^}�����k�NhOQB����ނ3�6{ȳH�g�u��p�A�ϖ�\�ip�M�V%�<�������z�[Z5W�C��xe�%*v@�4,h��L�~�.����6"�CW������ڇ��0�V�6t�S�Jl5`_)WI���y�i�a�[/�)ٺ�u��j[�6̎�YW�3�IO�]�sn���ڧ��nT)� A�	ES��b�\$�Ј(�E�dك�@�0J��+��$�8�O�v�݄��_p+|ͪt��i綺?�|�#��v�'�d��r����(&a���G֤bQ��7㘟�ʆ��-5'�
n�������.!�~;V��\ ���u+q9��O8&�e�@��y�8�bR}�NP�4���D���j�f(>}X�q>�r�y���T�L�ҵ.�'������OQ;o��!��b���P�?��Ͳym?�e���4��`�]����L�*Dc��0�Ϋh�.�8���dt���x2�$�H�����k|�02u����c������nZ�����n�j�R�?�pc�$�w)�s��4��e��1��*+�]ђ���훚���T`��{<�.��q�T�_�Z�����������L��N�6k��UfW4D�^��x2�~tO�ؙx���#o�Q.����f(Ͷ$��\����9�
�k>R�ߟ�3���R�U|�4��9�� Z7��09�x�[�E^Ҧ��h�A�U��iB_@:���~����t´�NG26��_���C�&�SR����Uq�������f�I9���m�_��a����r�A˶�����Dޛ����5�5�c6�rfI1gD�w�v��!G���n��e�+�f�:M����&��|9ST�����p'�ǫ#=*�.ްJ���#$*1[4A�b:.������R9�Cc|�0���6��TLO�W�K��Z��-��uJ(�zD7���Y���g�[��+_$$l�^5V��RO�]Y~��+��.��R^�U��H�_�&�ӫ&�,#��j��D�Ij���V�V�V7A��u��"-��X�m�1cD'"��,��E��lC�#(;�j���m?�k��z�1G��^�5^'Vʤ��K{f�"m{-|�T�u�1��/��//��'�� ��+�3�	P�RU7�{oTL��������B�H�~�K]�n1� �Q���i
�	��'dkiйź��pӇ��{B2_�ۿ�����	��4��׹*������e]�~�֧%n��8Ȧ����"l-��h�85�����Y��8Ƴr�v�������SB:}��1��RT��(>?�P�`j	��+w���=z�6�]O���_����3Պ�#WR�+�C��/?=��:�4��"ͷ�em�4cHP�E0���[Z�w�`Q��\������'44CF����U%���P�M�k.cH��+��f���g�QfZ)���FT(�䵨����xG0�S$���>~�Pq�Tl�5�r�����T}_�qx��w�s��G��O�����ɖ�ځϗ�;���
б.�mM�>)��oo��'8w�[z�k�SWq���v����~]��KD�8#tH�E�'�����h���Dᦖ��D6'��q�8���5~�J;Q���������]8r�Bż[�����*`/8X�Ztcm|>:*�L�>�9���+���i�r��i���NL�*ۤ1�j2��a��l!�)/�;�g�doJ��Ko��U>���VH�[�O�ԝ���5ia#�vCT}���i<��`c�&M���Xa��WӸ�l7���z��&�_Қ}п�Xg��ӹKmxt1���)�E� r]�;0�Ǧ�oI�ʞ�q0�u�J%U�h��� ��3��^݌���pcD��	w!g��>�~�W���Q�P9�8�W)&�sۓ�
�P?��"��ǅ����z�A�w;۔��������(�x��zl����g~x`��E���1��9���4����k(�yD���ӈ�<����U�3 yz� �f��������Q��R����Q�~��m ^��D�nhX�A���(�%�W�C4B����.R؈���!Gs�Ǉ�|����櫠�i�;H?�9�i���?i�mz�
_U��	��T+����H�B#.��� fT-O�x�d�':$�؜/L�y;�����mPp^J��#-��H�Q,�?�Y��P�=T;�=����.6��|8�����i��?����ϳO�p��K�y#����� m�)�ЮO�<�q�N�q���\/Ԑe=N~}�֐o;�ܓ�5]��ݘ�?q�i��-�T"��
��+'�!�A���~C����
�QIK�D�>1�wH����o�t��S*�oT}�P���ő@¸  $P�j�F�VE-D��7
X�<t�ݣ���5q�W�:��/�Zua��V�U|� ����/��6��4D����+�d`�Bi���`�8�����`g�MrN,b2����B}�3����;�鍝��_O��~?�N?�|o�����Lv�vH����}b�;8&�	`0�ɣzp��mFX�}����B��lMP��'E����o��N�'��5dl�sI��%�o���ǝA0�~���|�D�IM���~R�;��%q�����8�{�������
��4�<���=��n���^��۱E7�?���N��ː������y�i�>�A0�7�ޞ\��M`��wr�� P�\�8�$�V��|�}��C��У%��`���M�{i�j	���G  ��U�Ds�<gFdB�\��|$��>Xie8��<X�d-5��Q�FZ`���r�����k�G���:�y3Sk�,MG@\�4�������Fb+���<݇5�����d����XO���P��s[\'I������o��������y���{S>�b"P��/[o��!i��1�&��b;��tv�Fűz=Br����#I�!uZNȰ�@�ȯ��I���f%�'��@b	y�S�A��K��W�Te�R6�j��U#�����_a��"|J�&�!L����-gц�I�y���K���L�S:*`!9/p(���!����E�~�婥��Cބ�[��р0x{ю�ࢱWh�n9t�����=��p	u:{��r����ﻴS�g/������nE�,"���f��*��K�	 :���p�#����o�p�QܩgQ(ފ��S��8Ҋ�賽an�<	S2{c+ �J�*>M��]��~:���������̼-�����n���v��Z��J򈘻���U�����dn*"�)]YʻI-W|�����0�lz�fbGZ(6�O�	���L����(`��t���V36����D��d�5�������htt`�1��i�APxI�j�vP�Z��@$�w��{��0�b�h0�uF{�:����:q�Zc6Y�r�T$���s����q|Z�xvp_j�y׮����r,&;�2���^7RH|v{�Zŏ^����	�QgGG��ڃEw�W��aPw���g���v�"���N��ȦBO:������ӳ����M�^��ψ"��b,�_@��Jw8�����U�b����Ő[	�G,�w`�]���5ɪG�^�!��oa<� H�8���Ǖ�K�:.l5��n�i]
��`�6Ҫ�
�~�����V������WR����ϱ���3�����J�`Dc��'x>�f��"-[��.B1!sY��TG���[<��y�`��`<)��#*6�Խ	E�0�}�t��);%�H��V�FqצS�o�W�؄�����Q~�"�!���3Wm�d�w� r	�,Mkԋ�w�Mɿyr:&����vf��fLr���)����M�������A%M7!Yq�l����TB�S_�91�CWL{�#*Dh^5�M-�+XW�G��J��E|-Seש�$�����r2t��L�	~�gh%N��\A�����Ѥ<,�;j��i7M�;h�z��%rY}A��ۃ4ɗ3�zY�U�@���cw�M�%��Po
�2M�}U쓮y�#�Ce�vr�N�N� "H�U�S"��<�(��S���� �݅Ѐ� ��lѲ�c����I��x�~��U��s�F��Q4�K��-l�9!l����Ȱ�0+��IO<>�|��ɎO���,*H�g���C���B���>��5KEr�YGa"� r�#i�	�:r�1hC�Ȓ�H����a�ώ��В�MtU�K��ǙU��ݝ�;�w���ƖVpi����^2��m�^�ҵӒ��$7a�"H����ҹ�
d�IңssVXA�����p�7��y�K�<R�J��Y�<�m�o���^�G�q
�;+}����<⦦䭼L	�I�wu����������o9����|G���o�!�����o����G=��9D�] ���^��Գ��U�?��ޮM�a�Ħ����%�m�py�!���W�?�Xs���\��i�L]�|�ы����җ�2�!�2ip����/�e�6�Ɂ���a���������\0xY-���V�t�#Ns�J)0��:�Z�g&r-f��@
B@�.����7�^����_�z�e=�)�iq;���Qy.W�.}�^������G#�\�����Ƙ����4f�)N��|�� ����g�����\W���%o�,Ob�Zn�#,�Q �Ѫ�Y.w�L�3�t�C�en3���ڸg�v�$I�l���iD��2�7���p���,�ᐃ<�aOS�� ��|����ÙS�}a��2��K�d�L����8,�~8{�mgV/�*t�:(L�v�㲬Nɿ�\S�?���)�C���o�a�%�a�Hq|G;�ֈ��&Dkc�÷��-�l,O^�j��
��	��-�H�h�x<q�?���h9�OJ��ײ��V���u�!��<ѝx#��"�{ ��]x)"����Y�Uɡ�S\�(�0M���������5,i2�88}7,�u��{�3d0�A��|i8L���^�/%��u)�k	�yR{f3��;Z�+G"�9��gRY��8th��[��"��G\vm�@?#����vnp}\��#5�8��A�:��xL{�%�c�VE��Q�pߡh�ޅ�bWM��J����	�+���:��k�Z��q�ȳ6���=��}]�4�M�7�Ô�x-Ru^��L�dp�/A�%�:�`�O�`-�gyb�ӎ0UǪ���b�Q�Cx����������gPD��@'zD�S[2b���2�B
oc�LS�a�_��z#�x�`�x&:�}5���� 2�)��1���Z�w� ��=\2�#� جqĽ/��K[H����Ԋk�D�Z(z�mj��x��OZ&'�~�%�W��".�r�8�_4����� �W�{ X��X�[G-��@�xy�b��1�w�&P����/�m��K|�Y�����%�fq��c.�ԅ��;ϛ�����F����aj�~7S�/�܉iK\�����%��>+2���y����Y8&�{Xg��w���m����a������KO������q�s�g�~������s`��#�~2��+lq��u��J�L��sJQNy����e����ۥ�!��g��zE�E݁��NV�J��I�������Δ��6�0�&	;	�V�ѱy���"�Z��\m��q�l���$?���٪��,��:�;����a�"ǣU��_3��O]�#5zBE�����|��g ����P�����EEl0�?�	<_(��Z���Ԅv����8���JSe<v��ۤ L�kӽ� �3=�Q�9Bۖ���� x&��8�@������<C����3~#��鉨P�E�ie�����]6�5Y�]p��Q\�!ճ��>�VZ8�^	vl��i���2ܽꅅiپyl�l4`��"ptƋ�ό(�-��F�|"���I�ݹjR0#����V=j�Z:4����$\I�萱޷d<�`��p_�'t`g���/�yO�����nMA0[n	�/�Z�Q�.�B�����i�).Q����͑ �`3i z7V4�r����T#-l� f.-ը�2�qc�&�����93/�UGNJ�mA����rM;���y�+�3��� �$9�����Bu�+�$$Lۍkh?`�5�4�*�Jx>(Q���s�`�o�]޵�՗S	���/CE�S�&��:*���76�W3"D�%���{/� �6�!{ۢ�L�l�y!��u�o1s�S��`�|La@���u˰ĘM���`ѕ<i.Q���{]��"C��*5�pe	��X�I�䧀�,U�������#����q:OҌ����M�Y�}��jP��B��UA�-H�Q\���󆹰�k�f �j�}�[V������ϓ��L�w �f���,Mrợo6�0_0�d*���X�αjx���J�cW!����l�!��,�S�0<<�	��|�k�Y$�!�UiG� ��-X�(��;UB&2�"V\�bS	p����A)=2�ֳ��$a�,�^5M><_h$wY����g��ǣ�Or��,��}�(G�-�c(��C7�4��\V�O�D�ƒ!���5~)A�Q��y���J+��o���A&��
|ɹa]��mk,�ZQt3"&��(c����7���*aI���w��F�����9W����P���ͺ'v6����~oik�%����@�h�I�tyѬR�ރ�fLG�M���d��}�8�d ��ĹJ�y(ƿ��f@=C*������=�M�CCU�_
;Q�C=^$g�r�W�� YkW)$���J��nc:��A|��۶�ťS��<�yB�ܼ�çzfz�v��)��cF��)5������Uԟ!А
53�jh�l�8��C���ax~��g�������tTJl�>��g�r(SB�ѤVK�:+L��R��+��l4AP�U�h4i�|���Ʊ�#DvO���S���� ��-�j1��9l�gܫ}�������^S{�K��9�)ڞ�fUq�����9�Ѓ���?���k��n����)Xn��ŗ�3��4=�V3��6��)7�3�]=�Q�|�*2��!F
�N���_�<KC�]=��2|�r�%�,��Җ&���2
���Eo�<�l�?��C&��#�d����7�*�/Y����6@c�%?	W�Rš1����_��l
_
�K�N�����U(�W�������������x�>�R�5�#�T��e�I�#��oڇ���՟�V>NA2��~�U��c ��Mk��y�?�/ ��nx�Z����^)��{����)�+Pv91/@���8�\��p� '"����x@{��ǣ�$:���N�˶�4>�m���	-��@�����實��a]F0��Ž���@���� ��k.Z璙����v�����	d�?�8���(^Ӽ������f�Ʃ>uD��A���r_)��݊q�̧E�H���A��@����(k�e�u;�ka���R)m�����ЪȪP��gt�?W��9��N��<=2}( ��w��G�d��J������M���˳:�T,�p��a�6TC�(���7��${�7"H����L�mnC��A�p��;�t����xP3�T��r�������[���n\��v�5�����n��ʖ��1���`wگjrω�%�}��ƻ��)rp7���%Fi����_�=z�]��(�&:D�BG�|��"���Nl�`5�R�+X�ss�!�x���p�w�$xF��#_�KA�7��ك�!����^��-p4��f��)w�B�AQ�'��v�j�3Z�����8sλ� ��Q����ج�8�Zf1
�!���7OU�Gx.���Nj����O��k��ph��57f{`(�Z�WШ���ƚ��{�m��C�׶���J#- ��)�v��#v��|r�ek�Q2�O�s��/������ƺ>(C��|W�@��������rU"��Vy�6��?�d"��њC	�6����|g��:*�B;�Uf1�fA7��%k�T��3��D`N��a#�8(L;�P-�XId0M��=�X,�d:j�R���vm��U�<���P7ID�.�F085+(M�7 ^�g�ekO[���dg���T"��0:jz���hU�����8z9�wƇ���' ��D9z@P��P���݆�S��y/%��KT������K"y�F�	�C��e����m��f�+�mr���¸77r����D['A�H���K���O=x:\�|�n�W��pU�;q��*�e 
XXo��hx����ڔu6��kҲW1NY��/ZޘZ�0���+�/�^�w�e*v����T5�2u4��<���d~:C�$T�b���g9�ne`��Dd'hԮd{��4X�`�����Q�z" 0�~��F���J��*C����5=����ɇq�Z��	5�
����a��r�u3qv$������R�g�� \�,<D~��@�-��L���V�mw��3����X��.az�?9��Ap9)E<���J�����R�Zd��'��Y����`��oZ�c>��O�"7���6�0D�7
�(owX�aD����%aX�W��.H>G���"U�(��W��q��"W���ϐ���N�jy����Qpaw!��g´Cc��e��Hb6��9�7O'SEX���I;NS�xb���w��(`���Hew� �S�W*�Gl"ڏ!ޕ�b/X�%�����Y���9��3��M��u�i�A��Ϲd@�}h�J��(l?I{�8�O'P�~c���l���VA�w�#�e��?�os~�����Zd/����ʉV�*��R7Ppz��إ��%j��x��,��P��`%�ucUj��8��"��U�K��0�$�!�����oB���>p��<�M�$=���W�j���儅2��i��-B�ܷo����C�Zf[�.4�Su�voFJ~�;_bQ���,�ϻ@(1�����cg�����}��&'wҗ^����d|Sv䞬Y��hQ/`l��\J�Ȝ��V@��Y]W�_��?�A䚘�[�xO���H�tq�5)�[��lS��GY�$o��p:;�N�%�۩�*��k�e��l����9D�ߡ1����t5r�� HG�����l�R>��s��9�׊�Ž1�����?'����t��S!�g#���ȳ��*<.=�[�1���=~�gqd7����1fD��[��4�O�kW�P`91�i�$��p�g~nv��=�?x�>��ޥ*�_G�]��63�1'����	�B�o�-i�gM���ڡ�Wv���g�3�8*����H�mÙ��/}t�*/1e̾R����ZY��
h-6�,��@>< D�fIw�R�fK�5�Wo.z緸��L��ДKR��oԘ��:����S*�j#³V��O�ަ�o�27�w^΋�Aԗ��g��k�0�i�p�J��#	g�� 9D�e6κ»&��^��ę.ϲ8�z�bݒ��J��6|b�K�k+���
搪ñS�㧩�=`
A��Ы�D�
���A3��H��ϸ�N	�]���S?���MW�+�丽Z��F �� �@{2� Wh[��q���������Ѕ /
��%� �r8Z_�f4}}�� �R����&�}���s�Z���jNu]:��
5St��v!K�}���H�͢�6���&s_\?�,�X�Vt�_+|��~���z�� ��9�G�4@*��H]��a��ɌÆ��s=���LBk�I�'���)�ؿ�\+d�Qܡ�-) 
�o���5C�x��$X�Z}c/Ҽ��DG�2��JPޟ�+%賂��+	4����W�P�J2���9VR��Ƿd|���۩�e����(H��Ԫ��TJ7�|M6����/H�,�_�1�C@�NA�ů�i�/bk�� ��y�A2���c��4L^�x���=%�YQ�0���[%K`���f�pX�S�kaPQ�z`�sxBh�ZXz	�-�?F�#x�޴J�hT����(K
S�eҙ,?|q�Ɩ�n#�Db�ߒV��ͬe�`�s,�f���<�P�Z)�2;%���<~-��ĭ�[�3�:������l�����^TE����얪?j�a�������'��0�.J�<��.o���."cc�?hNٌ1�m�1�����b?2T�!����s�2���� E�����`�Qo���R|w�5�͔z��)����\S(����4�(�Z15���=L��!~�UzGzI��>� �ܢ�˷j����x�������a�T�i����[���4�P�:�Hf�%�j�d��Km�Pl�h�W���U�|;��һF5f��$�齲���d"�0���ˑ<]I�l�{�R/0��Y�}ep�OH�a�Mf=+'�=$����0��@����G8�K����@�ڵ*k��Zcw��)��-waSY�r���<Yu��� ��X>�$�Q�0A�&m� o3���|����fa>g�ϻ�>Ps\*�l#	Tyy)ӣ�!���I���赓����G�	��#�8����Y��869F�,�c�O�����p�[A�QP�d�u�� ��b��аi`3��@i�ɥ%�[��[�`�����@��+il���"�ya�Q�@� :��-�1����N��{h�e���=�17�9�1v���*`R���)ևE���I���iMp��V@{9�0�ӯ�E�d�O)} ���L��2��)�o���b!��c�n�w�q���Lv������xȾC4��#��b�����j�a�����D�b�uH��sD��B��C��������Y�*8!Q�>B�=%������	�����e}L�����3�#���g�>L���U�V$�w���Agj[��x]|�L-@�Y��gQ^.���~��I#[�;�����}D#���;F����,v� r ��p�O�O[H�db��8' ݠ��f&����/[0��l�3c������@v�j�������f���W�#%Ѻ����!�k�k�k���*)�����
q��=@�D�����?Z���L �c�,��o�9yG[)�|�+{74=�ox��DT��R�le�ov���2#=G�~,��/� E��A-(58�4�M��K_�r��[�(��!���K���Ǟl*���>~f�Pr���IM{�YO���ΏQ̗=V2i�贁�.���1{����}]���8{�s�d�`�_qA�1�C���������[�S��-�Wl�d|)!&�y~��RT¯]�\t��R���˾���;�`n��b��f�Y�ޮ9�؃tb�eՏ��¦ر���y�C#� l(@�K�5�f�d��E�S����K�0��o���ع1� (o�*�.��bGʂ��� Д�1q����3�$�a�������G��~N�!�~.f��,R
vH=�����@�N� �g���p'ԻÂ�i��a�������	˰Fd�<��@͜�w����n^�K�Z�᷹I�͟6�`ėџjP��@�o&�[jAn�5�,��Hm�3xP,&�W+��rZ��P�p���'�G(����Eg�Y~t�ul�-�޵�Z_7A(t����,�����u��y�� ��%���|����sl�Ե43S=>�+׻op��ؾM�]��27]L�R��!�g�	ο2#��Q���_NI?O�GPu���o�)�^p����&l<�f_i���2K�~	�C�D��"�Či� �kJ�W]~p�O��dj2G�Z-06���ҏ�P�Ө��璑���A�(��\�H���e�_�+�iUk>Қn�?��).�!da�8����fslD1d_�a�,Ӏ'���[*�{����)8�!oE�ߵt��Ktz�UB��-�3Y�9b��Ta��=,������(>0uA��aH�u��AK:� ISѳ��H�2?�������g�?r���?Y���<*Y��z�d��F
��R Y����
�S���M��GCv㚓~/ ���V��*��xb�L��J(qE�6�>k�7��^[>>nST�Xj��i��}<�'�0���LA���ǈ���QC{vI{���d�3��aČ�X��ƚ]"Wy�%9�QptdV��ړ멽ީ=����t�)I�������e��nG�4�%ci,GQ%�#Tf�+�̱�R �\�32l�-A���'�����寁�A��Gm��O^��V݂,(0s�����>�(���9���SOYɴ2������z�)c*���z~9�T�s��9G���L/�ʋ{,�W�[�^�Ǵ��~��W���!A����V�y,�|9t�����m2U���|�����sL_56+p����r'^)����c�nkx�[�|F5��?�@ʚEM�k(�7%���<�W�M>5��� ����A$۷�O8�ʫ��t��?��Q9��
�H�"K��^�P0�F��"���24ç�]n�-�w��=�_��ֱ�e	,�ƪ�<ho
!2�1���bYǐ���Lئ�� �u�¶�Dd�uH���D�j�v�H4��b
�#4e\�$�NK>_�O�A��	S[�G���F�z]]-ca�}*p�7����B���`l)��	��DV�������v�uS�~Ӌ]`�b��Q΄l��k2�o�W�M�μt8I�!��덅��#��2���F��P�������B�y�jR�-82A�F��4ɳh7)f�܎��>�p��0m��`��X|�l�.^-i����b�-�H��F�Az��8���jJ@ND�J]:�j힥}l[�H�?���ˉ�.Kw9|Z½�Β�%CL�Y����fM��VC�������E���f�V-r"+�z��v�w��3��_GI+Q��Ԁ[7k�!�xKO�h��[�tE�Be B�}Qu]<�Hy�jo�=�(�7I��y폗y�D΁��
��k�o��1����M�Z��$4 ��aW'��'�{b+���7k(�*�␙��UU�Ajb���!��aJd�I�(�V��놀��T�'��s��i��G�W�{v�������g�m�ss{�9�--C������QcD&a,���ߏ�>�קq�;L9��A�x󵾮�&�kStǏ��c���]j����/�--2����\�_� ��)��F�������߅=o�q#�@8|wI�Ѹ��7[Zďn��+��n����)u%C�H�
@�-l��7�	�'P 
"[���7�[lLO���Y~�'��n�u��σ�����[#�0��]��75�^}���uECQt:� �	��i��`2)�ch�	$`m�l��2�� �� 7���^�s�j�1�fՠ���N�t�|f$%'e�>�����`�mf�Qn!J����j�A�+�$!�'(��T[��n�#� ^K��\ÕQ��M/+�i6:%��|�zE��#|$:����%�T� ke*yз��	���A��CQ��H�W�kf�75�f�
9Ek�L>D�)3�ϱb�\����&���~gA�hB���W6]����C��$��Xj��)ht�p/�=�m��I�D�G����Bq�#��a�s��e&�,�1�;, mo��1��ݨ�l��*xIR�K	N��t"N �^%K^("<E��6JSU/�ZW1U��$xQ�L���F��c���`���}���J�W�����U�W�s'K�.Jth���{Fme|z����k���NW�<��/D2�z��	0}�'�ۘ�;��c	y ?gy�/Q���	�B��-�پ���WG�+�ۢ���?���C�a�����>�D+�}84�*����#ӄ�*����"bw	"ؠB8��.�J���Z���?��"�9= v��z���5�4!	L"�����o&�8mA����^*��Yr�!��Ë�HQ����A˃~��^Ȱm�ÌE�80=���~~���n��{k��ϙ�.�6*�1��R�66�Hֹ��f*'X�g��ˠ�c�L��*O�WV6ba<UV��saXGޮ(��>����܁e�b/��ǂ����$�;��y�]�hZ0ƨ�w�|k���`��7��RZ �Q�W��o?	?��?x�a;4���]���ϛ�L�y7qU^��
v�c��J��Q.��@sD����bJǠ���g�f����U�e<1���U���쵞R��=���\��$�+}�A��@l̠������9'������r]��X��ɂ�7��4}�e���2	Bv�*D�v�7��}-Úji�����d������y��(�0šEW[�tV�ϊl�4��֭A&m�܇��\]V�5:��е�n��=f�i%s������N��c���.ȧ�qDZ�,ǲ�L ��Qc��.���;[���2���7��nSL[��bm#�cm\�w��Q�W)�1A��%�x���ۀd�o���a�Y��d������5�� E��W~����Uui�� ��������n�KS��b� ���k� aZ��.��9�FEƜ)��Ѵ�=;�o^�y��{O6k��l
2�hyE�)�O�8�'�h�ǜ��!�#y�%��!�A�5hnx�[���PO���ߪw��y��>��>�Uy�\��i�Ъ������gG������x���<�#��$#7��G�<SȲ�݋92�U/���	��Ɓ��$Z �Pƺo������L�l��ac�}�\.iQp�Y)�R��:^����u��ւ+-"1�ges�3؊�?����8\7U�˚�_�`s�g�|{q�
d��S�K�i�7F���u��K�}��RWI�r�ȩ��Q����K,�1Ą�;\�xfk5&`�s�y#/�;5T<s8L�X2�5h"�p��ҚĿ.!%%]���i+��p�n��A�������N��918G'NK��j�!J��Ω����ɒ��o�,�����)�c��������s�`�������OfB�˿��̩��Mq�`֝]�D�V�tT �o�#�Vr�_TK!`�*!֒�#%+�H�)�L����'|*��O�� &��.H�+�ӰA���!�O-�1wm��7Z�7�@�&����k�%oq8�I�ՎOܼ����q�G�
��A��������.�k21���ccڏVY����h�Z��t�����F��*��RL����BJ��ьꍚ���@��*����d�Ȁ����_��}]dne�(J˻�/��bmR+��\�ʂ� �L�[�<��L�i�a�ؓz�N�=��{��I�LB���U,I��p'�G�ʑ!OQ�F���]Lŝ �|7V2����.����ً�������t�E�5���U�Dv�	$ywnϺ���c!���Cj}#O�kp�����j�1[#&�Պ7pA]z"�6\�\s�-������"p��<(���R��nrM���_��X�誙Aw�_�������	��j��TWӎJ���M,�OG�c���I�4���#kuF{
�E��"w#Y��x� ΄��.�s�����'?�s���"����%Y��ci���-��b��툁�6�+O/K�XB�맾��F�x/Er����)�Gp�H���xH�թ�ʣ�r
ՐJ$��)�E��ge�/���8��@���rú��T [�����Y�z�r&\�2AU�k�<��S����`/jJ��C����H1�cmY�
(�5aH�;V���O_��Q��:�H�q �[��[I��WM��%�D�~��l93�ph�#�_�k��p���6�t;� N�&�K������B����X[�X�tD����DjIm�)�a�K0�K�k���zL1��h�Q�X��v>���䜌U�ǫ"a{��rBǻ��K���J� �}�♗2��!k�i�K�z\�9�5(V����Nm5�m�ŵH
��N�:j�x���޼�A>��MWN��Օ��cw(��ؕzޘ5���T�J�{N2�F�j�G�_�`���	�i�O�����X��|l��OwZK:���	�D�r���_q�j�^����-�;��Nb1�:eoA�\Z����OC���^�Ҽ��{tlHY)Ev��h���2���zA��c]�g�0�D��>>������b��xQ.	��C��F���j�v�&y�����"Wnv3?h.���K3ؤ��������{�k��CU@=�I��Ժ�ڗ0�avn���:ޕ
 heݯ+N�����[�[0o�fu�K��eq���V��<�r����G�����G#��)��%9s�Z�p<���;*]~��EI���m �����QibJ) j�ѫkE�=+��`�?��8���1p��o
#��w��ΨZ�zk)x�H����D��j	ҩ5�]���� p��޽ayxA�Lw�qp�u�X�J3'��T�uf��h�X����F
�-M��j��t�MÜ_��UO���k+N4$x�oGzP'�??��3o���N��c��V��mA<���e���}逺[n��q�q����j��\�t�!�Pi�������꛷����ۍ;���p"��<$}oΝ��:���^�Q����?�l����s�U���P�WJ�U�D�x���y�tV}��ϥ[�1����ǣ��U>�iH0�IS:�Ą�%S����Ӣ���qgQx�㗞v+a;�(��&tJ���9�c�k �o��~���Y�a�+�<�Z�Xq����_Y��xe}1���=�ߖ�џ�{<S(��#��{�,���al������,�{r�M*�9c�G�,���'�!��������C���c�;��A\������G�������Ă��	@�Gp�tX[H�H���s���8���g�@��=�#r��Q�"y�U5��ӷ����IgXd�v@��N�Ώ:���J�Z�����E���<���z`�5�c��	�pwc���Q��ݯ���T[��l����9�8W#,�2�+v�f)���� -�4��wd"w�J��;\	ꊎ?Os8�.��J_�_Ym��a%�31�&Dbh���V*�T>1F���U	�s�~��:����[�*�%Đ�h�^��z�3�jѺ|�Wj��@�#/�.n�Uk��Fi�%�N��!���~�8~g��,*G�ڿH�S��~W���1/�Q蝷���� <�X7Թ��u��u�\᪕lBX�&z$��9^��P�b��I��ه!�g�$|�7���-�v�`�{���2-����1`��M���V୆	L�6+�{HRų*H?y<�!�O��ɢpm��Jȯs��ꋚ�xX/�ȼ��3�uΌ���R�ゕnAl.�`z�dn����~��n�!+$�&��؟^1�,ug�3�����/�}����r�|��É�<�Qa��;m�U~/'q���;�R�-'u����e�А��Z��嶻,�L�m�������`���bN�fs��w� �*XBR>H���b������	��} Y��%4���Mk�Cf���:���w'b,���]�c<n%�b�J����@����?4 �����#�]��P������ŭ-ŒmG�ؐ���S�ä�=�b(��T�l�]�%�D��tR��@�@}~����&'���oEVڧ��^=S �M,;G_��h�M��*\~�~݂-�7���b���>�Ο��w�,��%L��b�i���(�m=7�Z0xl��S��=H�/_��Q�,��FL�bG�ͤ&0m~�� �{�������fmh�T���2 ߩ�-_�y��&�L�g���k/i�kv��k���+��-�&��
�9��h�&�hr�~��i�]w��j���+��}O���+��v$Z�D��u���B=˅yD��dD�zc�O�]��~��,!l�҅f�y.���P�q/0��+J8L	.�w�e�p>��a*A&�m�N���1���z�kz�>RB�p����[���[�i`l�8��5)��ߦ�e�~���;�)��YГ��١-ev�78���������3��'�����#_`�� P��d���� ,%�D��h��;�xJ����ӏ�6�wa�C(����=�{'���M[_����0�.x�繟��9��F3u�;\�^)I��=�: W��ob��g��f�Ί翗̓�I��v��3=B��7p���,���L��z�60(�#���+R�e~�4 �#�?�ҽN���_�4T��F��� �~K��Xn� ����ԝ�����GH���Y�P��~�<�[A�T)�B��v�O[���Hq���1�,�E��ό;c��r#�ʅ�x�S��/��j�;yV���1@}*�����%�]lN�'�Sg<�:g�(���d��Ts���ư׎�G��x�}_��V�au��>�7�vKb@K�;p���뫶p��!2�zDB>ɯL�X�s�d-~R��$��
Dc��=ڻ����;�F|qX��<�n7(�]�ĵ��$�dN�aX-�^yx��������S�>�8V2�񋪈���Z��$�9׻�{g�Ħ��%x`���T��V��np�y��3��:y	"/�w8��3�&pZ4��I��\��al�M���,���Ϩg�Ϫ���Vga|(J�g���.l��{���fn/�e|�����Z�1��5/8Ӻq��g*ڿ?�Q�6����r#�o���x����p�W,\z��`�?�J,`<f��;�.�u:�ry �����wB�C�����!o[8d2�<��cqʝԮ���/C`I>�����aߵ4���P0�۱�3����k���b'+K�(���E�ϥ�d`��u�U���xT/ ��M�������@$�4��]'/A�r8�Ӳ�G~�\b��no�Es���|>�8�!4K�R�H��JI�#�69^:^����w<sA>�^X���Bm�.Dm�C��!�-TO�\�h���i1k{�`�EFu�}��E�Ll� �s�f�u��d �;�5�c���rM�zi�&�9ѕ�N��p��8CL�D%P����=&�p<kZbd�ػ�vV�G�S�=�]��2LY��L���k����0x�5�΅H�d��R��B��~60	m����K�L�ہ�ϣ���M����� g�ijn��X��8�(����+��JQ��	\$֬=���b���ԊZ�ˑ��C9	[Lq�ߡԩ�p-��,Z5���sDՋ=�9�CT����$�����L�s�2�lgE��U2$,��uk}���3��a}��Z�Bt����'J�Iuƻ��:(o�t4Z��:B��ř�	�8#*��)m
&9�^	����Ѐ���Hj�l���B5� .�Ā�� #Q�uoU &��S��K�Z$�hD�(��ߦyqzwk�1p�T�&�x[y��wG��)=���Հl��&C�뭢�t�������,�3Ϸ�����cBI�ӛ:�P��q[�nT��c�N�9{p-w�V�Q$3��1#�$�����OB������'jmvL�h�B��?��Z<�RO�?���%�Q6r[��%�o�M��&g�d�l�̙)��y�K?����-�׌#��]|��{�38�+Hދs���Q\$��XV[����.���2�T��i��[��ߥ���#�=N����_�o�KIY�D�J�����!���G����G}��΁�s�=kc'��]Z��@�+��J�`-��"�&��1��UUyu"��..�@\fs���M�Z�5�Re��;�)F��Y�1k��O2�����ζ�W�zL�ށ� XO�������J����3���Rr��'\g�r��]U�T���cAW��O2��ڏ�k
�Џ|�d���ߖ彿U��4]ŗ��K�;F7��},%Z��a��8v>��=�D�B�}E.MyM��b
\��~i��w@ԁeRG`�F�2/��yh�U�Q��?� l�Ɵ��/4������B��w�����]cC�� D`F?f��_LǬ_�L���,p���=W�Yo�:����;+9r.7���e�qhϕ�(�ws}:;k���k�\ԂӴj�^��r�F�<j���Q��S���OOz|E���8N%f���O[��ng�;҆��`{��zn��pBmR���a� �.������{�l���s�%��H�Zp��s���倜��d�eH�h�����U:T���I���Ώr���j�����5�ڡ.`w�g�����y�F��@Q`�a�.=��W߶ݲ4z��,JO+�T�*0!b�I��ē⠊�6���w�^�q��T>�ڇ�f=�K��E���j�� �+ޕ�a%=z��dS��wn�CJ����*��9�.�[��㚋�#�Px'�`t\�{+���%|�5 #��X`{��˅�L1�O�81�~MX��g$��2�-]��|�[C���"��	[p�Y�D�_@�+����ru���(M�o�8�٦<a����/2P��p�v��E=��"A���2OSEtI�Q4���q=<��#g�^g�X`��������o�_�l|�U�t��@L%�T��b^ZÏO�(�+.��6��-a���g��.�!富脉E�G���� +���}�v�O��0��[�O���,#�uƋxS<��KS'����	�Q�\�/�}�-��^/o�S8�![���O�8����@Vh�F_s45<��;�X�r��]n3g+`B�{��X���UL���1��C�˩8jF�@���|hʧ���iL�R	m*�R��f|UR���Y����Ť�Lu�*Rڄ�Dd�f�N�|�x�|�h1�"�}��֦�Wc�O��q�wD�!p����+!�, }���
W��[����i{y�"F���:�h���R� ,{�"TAܸRS���k�
t̡ꛤ^.)���A:l�X�eҊ�jj�с�ck����S0�n:@�b5���w�������&6p���z�{H�#b����dd5Qddv�A#=|J���!o�&U���2�c�6��WK[�̨��jf�x�/I�7�#��w���`�i���w�h��(����e�1(������1=���p��N�[����0��>"I��l@
�!��1̾[��r�{��i�{n��w۝n�������zVI"eC��xd�7� ��6��{�qf���Z�6�Ak��Zxm��zk��B�h���#�6���{xQ�V=�K>�@����;�^#��*���̂i��<^�l���o!q�\��Ҋ�i�VS�4��ośY�b+; T'����rXG�'�Wg�����Vx�Q��Mb���e��
g}��٣�'�t��xp�2�Dz`��k0^w��'�L>�v?0c�S8�J��w� ER����2� ��J��ͻi(�}�\G��C��#} �>�?�}Ku�ޠ�d�q+0t{�=�1S�'U%������9L�&�n����h>Z_灰����8A��!'�'�v*�9����,uE/'��.�B�"j^7ǜC��k�H'�5�^f<������5k�=���J�E�;"�����@eaV��X���wߒ�t�_�al"�Q�&V�c@r�Fǡ[�,-����S.�̜�@e]��h�jx)"�5W'Ho9Xy�	�)��BM-��i�W1����c�37�����C������T�PZ�?�KL���x4�Z�E%�u^�����s��h�$ÝF��c(�O#.�	���(9�M�1l�o����m`!��|q�����R�)H����]��x���F�E�E�Y�\�-l$�����Ͽ��Y^�!1�sɏϙ�]��T��`��tH�H�8B&�l�	z��Н D�D�Y�\В�@�Ӏ�o5	K�y��w�hg=�/XTZU`w���c�so�N�x�%^�s��#b�Yu�˼<"a2+�S��$U��$ㄸZ޽@e7��x�\���y+���;[zΫ`�3PFwļ��D��G{�3�??�^E��uL��YZ�����Rh�h[�X��)�T�Hf��F}J�G�;LW$Q���tLݥi���S��<AV���h8/u��dldΰ#�BIʉ�4�H|
�dR�,j�ʟ� uK�y�����m��p��,�Yk9�@�A2<�g_��CR�>48�C� &�JWId7��@.O���!@c^��-[�V= 3��fC���U��ј�@| Q�ڕ�y��|r�<�"2�j���a9��$s�z�ԓ�V1�k���r|�Qn@�p҂���	�� �o�vi��j�ӂ9R�U��`�����zz��	
��s�a�A6s�Μ�=�������(a^�X֢�JM@.Ǧ�K�!�Iy��
������ �s|ٯ�
�b����])Dlu=�;P-cq�T�Q5q�J6oXK��%�o���` i,f>��5L�&��X��_'�i{_����8s< ø�
�t�e#���$��C�L���\���S'��P�0��#����!Ι+[���7.
�C�.����@��o$�آn�&ڀ�S�{��k�v2QVis����{��N�SU3˞�a�Y9bڛ�p��j���}�n�$'��=�1(P��J���!��8�6f[��(O�Xw���B�{u�h���|���.�䧡���2#�>YA�H7��,����A��t�R�o���z�+C��/�)��H�{g4�p_�ՙU�L���}{'�eg����.�h7��\x	d7��#�3��c@�J@�b��p5%~|V.x�7�0�.��<t��M�A��Im���I�Q�_W�bw��L�w*��̤0#W7e�;Apm��}�.�M���ֶ����E�oR�4bn��j����
�ܝ�Ŧ{1�
�	Q6S-��+�Λؾ�K"-� c��̩��Á1�Zl�E�$��u�s�6	��b��Q�Ů�ݍ�Z�X����;];����p|`5��6�ED��Xp=���7�$�^mG+�b��o�r/����~�"����~��n�.5ݒ�x"B�Ǆ"$�G��q��/�i!a���rnT�M��m�[A�A�-Vk�N�.z��*��V?E�����(`w�~U�V\���+՛6�������c橗/7��cĳzWqF�
�]�B0b�I�Y�j��1��YՐ��"�JG�o�����N�{ƪ����Ƨ�5��AhStq7���*�n��c?�dg�q����!��i1(�t�(���e7Սo�8x�9��Cq�($�[�`��8[z��;OFTwC�����J&���!��9{�.��CV͢��|X�|8�Pb�4��!n`��
��Xg��!h� �le�U.�| �3sh�R������Pq�Pm,ҿ�����/�.WD� �H����y��j���eP9/�)�h�2]b%w��ߺ�r�;��S��@:�K��,N:c�Z�%����h�e-9@�W5�Q~+�7�w��"�z�t��2�%q��%�:����d�%�ID�_LE��S2������&7�/�Y����c�JY� c6xv�{��|�����WSUB��ȍ���G��<�&�V�c
ٞ'�lP��e:��c�̪Ĕ���#��=|��S��A�R��풛�9B�	�v���9z�{��`` �BB��FS��,5L�.�۾S��m�ދpW*:�cY-â�kÑt�b��C�oy�Y�e�f�5�q��H�������2����;eB�[H��]������
S@�y�Z��o��R矨jTf�����H�_��X��L2E�Tg�ڟ�&`���"�~f%M��S��@'�^�L��P^
�X{�S��(�e�J�&����xX�7=�/C
��9��E 4���p����&`��!mq���UKnC�i�j��������r#2�Z��[K���l��5�b�`4<������z`�%\ۯo�b���t�����WbeG���I-�MKeU��ƹ��n4��T֠ͼ&XÌ%�A 9�#ļ\�����R/Qp�a}3���'$r>E���^fs�(+E��a]� -T��gj��,�51�j\v��P��z���/���X���p��(#����.��˓Tq�g� T��9/Y��՝;�L�R!�Nr� �f���<4���@���'���"P��D�[31�K#J2V��Gַ�X[���a�q�7P~:r�TftN~�|�J�{��a���  ���W&�'�_����9>�}�%R��i��U�3O�?�q�L�����5�Xk	�P+���}�6�)�t����9WוX�:��Jn�����7vV��2 �?�����LA�`n��'��ɕ&��[Lg1Q���` "�z=�w�ڴ �d����{.u�#$��)l����>��=zb�ռ�,QxUf����	Ee�� ��g��A��<�	�t����
�Q�^��+���M%U��:p�=X���X{��4U������@�){[I�x��Ά�K����;k�2�`%�-*=Z����M׃���ͷ����v��P!�����,�$,���~��=�p� &6|��_��b�Ue�r1H�8��㮐C'�0����BK=I�V=rU��!�y��	^փ�9�]*� �l�d&�p�=�	�YrUt���n�[cx�q�F�lrG_BP�E����� wˁAoh�J0���%��KʭpV�B��G��=�,T��t(�zv41l�#�u)�j�w$Rt�~����zZ��U�y���p���Ϸ��u��c�J���B��jx�4�t�"��k	�Y�'˛���.��=����TVj1��3r"��T_Uw'Ǯ*<��k������^ �*+tX2k�x��`r�yZ#^L��@,�� �[�|p=�j�u�hK| �FS�۴-��7Ox6������cL��a|b�e��;��KD&&�)/�SY(�,�C��)�Yא%JH=�}�iU�9!�|c{���V�>܊8�f��\�ĭ��!���h0kڡ�a(#9��
 ������+o.["�B��m!н6��}���֭ޏ���Ԉ�?9|��U�����o�����oj�U��j*#���*@X�'R��Q�ߺ�j/�e%W���K��i�eE��p����㢺�F\�K�@S���_D��7�6Y&3�F��q���E�%k�����)oI��B�),��Lg�_��n�VP��"_��Z2싘I�Y$�E�'�g�c��i�ǃǎΡZm��=?'[:��]gډ:j Hu˔�2�-�+*]��ץ����۴
zڗ�����Pv�g� ��r4ՊR�B�G�OƎRّ�e��qk���ü8��t[��՛��&�޳gu��	"�+ٴ�j�ܠ�݉;��׳��چTV��Zz���qL���	� ��?�OF�fEś��]Mr�}ر;�w<����D�̐�[#$C��,~Pz�x�]���	��[f�&���a���S����$�8��A�V/��K�-: V� ��ʟ�.�sI��#���׭NO��u��L�G��:��$�J�=.�ʸ��[����1�`x/eO��.fA"&��fE�.��ݫ����d�� &�#R*�n�V^P���J���~�}�):�z�W3��.�A3ĩ@�X�>�9�GR8\J�,*�{������.�r�v4�`N�S����d{'�:��DĹ�6$�f�E"{+��+����D�{����g�]�6��d�T�W�O��KҲHK����F]��A���/�?��fH������eA�T�Ir�V]\wJ�Z�%X���%P<B��b�@֢tY[�<�o7���<��ol[3��ȏ���Y��)���T�^��F���N����W�^�n��Nx2�X�g�3�VpԔ'��Ǩ�����i���fIa��c�$c��W��\)y�CӍ���E�H��[�ij�mG���X�w���3�\!��!���d{���:�{[A�Af�b����_��i�$��4
	�dR�Wfݍ�M�/�.�q x/m��u�!�u�X�D�M�<��r���4�Av��o���)1yX3��s	�w1c�z@E�7	T��SB@M�c	m%�=6���עS���Ox��31�
^9����؆����%�tryp%�ہ!�y큀q%�dIӵW�����.(A���%}���x�9)�X. H ���7�n�B)�"��<0Y/���/!e	�]쁜W��%X�p�.w/�z�)/��.$�SPi�p�����&���h�^��%�Ð�zC��L����F�۽-�	�޾�=�~oݦ���a��y�1!�кy�w�����q��S�-��8�퇽������_1T^Қ�ظP&ɵ��:�2�)����~���� y8�s���i_P�z~�����qQ��R�Kh��a�
���t�Y�vu��[~,��k��TV��}&b�-��|�+��]��bƛ�9��T�L�첻�$9SД�p8ɾ�}&�3��/�$	x�HQ�o7���W����
� �%��N��X��G�u����u�����NY���{K��[���В�^��H���/�3Y���ns��ȁ[]LTϧ��uX���}T�<��S�4��c��Ğ�V�E�܎b�h=�����0�H߉�^�Ա�RҾIA�&(��r�B�|-��;yo?$%��T������ ��?���	��������J�<�� j�4ꥷC2Uu����Dـ�G�4=��7gS��Czֹ��	یZ�g�܁�����`a�v
NAr�So3����Qы�dţ�p[��(H2ȩ*ң�/
4 ga�/�@d��94�`����Oy�M>k��	C��˔(^�'��Զ��R����%V�py���w
���x9K�����^8b��ZD��i���((�Zڙa�A�cR�D0ȣM�G�YZ2�,>��R^��VS�]~�H�Y���g,5������K�*�&23jF��d���
4���r�i�����:`�&\U|��D��Ø�y��7�j�۠���-� C������K3�|�����ꏎ�du��:���9�q?�C�MH�߲MA�\�\����A�u����
��|z1lѾ�~N�p�<܈�֚��M_���#�L�Ԛ�/cK�#,�s#v��g�����(BE�J�W�1�w6�������w*��D��>K2G�^�d�zࣧN�Fk#jw"b���8PϾb@���� �D0t�r0���2����-rK=zi��V.�-<��έ�.CC�x�0�a_r8�l�4N#��e�ǯ$�i�+���,UR ��&��r�<��GH͕=���{d^0�`���#o��"�2���<�N+�laN:f�k�B~�Dk��N�˔�W�|��p�����9���0������6�KK�􌌷tC�V �,�23M9 yI_\%Q�T2�V~��J˙-�W���A��M�ϗ�h*,��������!S�v\͙�xM�<�*����n>-!k�_ �CV*Yh�U'r��z�k�^�Io"����F>cJ�;�G�=�I��J��5p�Q�?}φbZ�0Jr��*�}� C���b�9�����)�<-�b�s�u�k��#6/n ��:�$�g��ׇ����c�վ��]��߁��ZR�=m��ղv��=��6��n�����-��� X�?�u����� 	�>1+��l�K*����iw���3SDO��ҵ��[��A�x�i�/!Kn����Lm*�S����S�xfN�Tɠz��EZS8��1H>�y�y�-�i	��3f �2f���о�������ʲ���8���%+�@�[�AC9/uG~i��.aҲr]����<��O�Rwh�����4���L�u���dY��S�t�0�֧A�wO���E�&�c	L�.À=�qNM�(ؓ�A��t�$jS��\k�{���/{P�������Mdr&�@
��Z`$������C�W��Wp���E,�PU������l��k��_�B���ķ%��y��vƯ�?r�#�e�%��yNF�{���qoǤ�j���+�d�G�8�K���Ii���.m�Jx]����� �U��P�Bh�9�*�Z�7�c~-l恦�k��GQ�P{�Wn"7�Mű ��O�3G5��骅��y����Ѫ34ܯ��j'�O���%$ ����Pi��3ڠQ�k&M>����6bܷ<M��;���.h.���j�Q��wN�uqT��#B�c�L2��qp�I�Y>C��U����QI>;����S|������ߌ�E\5?��sƇ�7g.)ÚmN����B� )��:p�<m}����~mA��`ȓfu��u*�m�S��N���z�]3�`RUu�}
S�_,�Q�Y���ݹM�e�e��� O,SI;�8�{��~��� 
��ht�괋
u���q�e-����N�~��G�@IG�a�xZa@�2�b^X�����+��k�/;��!���y0\��L|�α�:��=�QO����et�S�+a�$|�ƨ�T�ߘ [i��o��A�m0W��(��	�DdlJÔeMV�3Tl��I���8�C�
�Fճ�
!���h�@��#=&�0'A����`�4'\�˄n�U�W����ԁ����:1�ڼ:����~�vJ�E��i�(J��pa�4U�[�R� FMIX���C��K��p��}��G��Į>��2U	)^A
�-g�C��f=�Ԓ[Km������J��s�" +k����-
K|�:��V���+jͣ��Z_�}7�#�>��(�������MV��^�P%a5�C'�:3x�x���ufSR�eMJ�gij��(��A_��>#,\>-Z��>
�?N��?V��8%��~+JB��O���8$�9���;��}�m����B�ݾ����1�ܙ���憥�԰eS������mm��7�,�c�a"�ImT���'F�V/�ƌ7�-�;��z��m���P�c�9A!�jb��8�G�:	�I����b�wf�ՁɩM�E�y�~8JR.����k���Zy�x��Iz1A��~s��"�����l�(fvV՜�V�t�� �~?����zE~��+T6M^���v݌�W��X`Q�@�)�W��\a�(y�%�t��9� 4��O�0;1ʴz�-��m�vϞF_̜R���U�J*����J]}b�R�����ĔN��*@uUvo�:��zT�&]{d�l畋VmdM�f�>E{k�d�
�z�\^IEC0dg�s1�!���L�H�i�w�n�b�`�����J���U��@����	Aj;F� �T��tmGr�o��_Ce\��rN��BOz�a]��oe�@���1��_@R �&s|����~Y��k�[%C�Ը�e��X|Q/����D6j�7�/|W�As3�F��8��+g� ۘ�$�Z�g� I�%���T�;0�f̵���o�x$%'4�-��=�Ʒs��Ƽ8m���~[�mt2[�Ѝ�� \)-Q�7��P}G��'�p�7��b���f�����y�:�d�Qܮ%��^鑺F�x��^D��X'�J�HA1ëy+�EЍ&~�>�X�O�G���)��B�u�<�U���`2ۻ!
At(q�u�-e�5�O��@�G�c�y��b�9�����O8����}�Q�=�SH��ê̋Oؿ(�A�|��r^7�H�
������߻2����췣���VD>N��(sf���욖l��}�� Q �t���}L;�-�'�t0E��.g*R���ʧ�L!����O@���3�Fr[�tC���3|�O�}@����v�H�@���@�yk�C�W�aH��?]#���:���Yv�Ë�K)'H�Q�����a�*[�"ݟ�������y�[%Wed�eR]k��%�_��k+,�^Jv�n�Nh<Kr�����g��>H�De�D�}
X$�㯦nK7,�X�����5�)�D�E������z#�d_�k\���!6c �@?���n���Ĥ�5/�*����i��.�3��Mo�|�V��4��8���U���IX{�%�u^J%N��\��	',�M���,iG����ӽ��̵�0�9ݻ6�hۚ�%#a3��n݀T��x.N���(>a珎z"4@�4�~�a�-�>3jB�tB�xl��BЃ�/f)Z��&o��M���c�������۰G"�O[���.$�ѻďhu��3X�{" �r�}��m{�����)�L�]�T�r�:YB��f����2\�?�����&XV���<+J����%0��l�%HTG'�=��R�y`���+���K�M����v'i)�9k(�A����.�]�kz��	'"{�1�%>&޴�M(����x�Y�ra�*gM&�a+�/����⍐&2!,�wʚIɻu�������΃�2������ꖘ��L�*������Ӛ��.�lD��D{�c���s#E����k�P�G�߈�N)�k�QW����=YHt4DF�ɥޟ l;��_�{�>q��AC �N��ClO���~k�6p�3����j�&uOD2CL�S m�NM�Vu�����_��	���T�ՆP��B
�Q�t�����_�b��?r�(���m�ѳ�<���B~V�4!%-%�RZ1GI4'Q�٣	AX���</i8����_`�\�D0���pL�y����9�Ř�? 	R���Zf��2����e��8���nT��9�J��L7�>���
��5�2���;����\��3	E�g�ҫ���ׇ�v�]װ\&�!�@��#G�zTҢ�_=z��)�-�|۸��׋u_.l*��8t��A~cD�����â`�EA^��$��q K�5o�8�5����]�[�
%++ү8%]��l�0�����X����3��a��.��}1#��R��F�M9`/j+�-��o���H^]��@Vl����%���b4m��ԅKg�S�X��A�X����=E��c�.�՟�C�|{[~}c�G���P���zb�@���m&�f��@�]^!��A��D\�pO�&�Ǧu���CЮ|i<k\t����,�ӳ<H��u-Ȧk
��e���W�5<��ž�;X;����� h/4�UtI�"�_X�dýP�o�V����\�F����YI2�9��1��X��_7�I������(�c�j��3��Z��Q��M���=E��zD�т�)j�����ۘ��z�����;Ey��f��t��ב�_v�_��`S�A*�8��`��7*�e6��M��ؚ��3	�g}W��:�&�:0|p�NM{/������V,`�E&�=,u�A��;�
��x6�r'p<���ţ��R�5�6�<��D�ߒ�ڕ�2G��t��c�w��Hfz�?�����k�K2��ڊ���Ww,�Spɜ�f&�<$�f��1Om�]�fM�l���@�mx<7���Q�Al����Z�Zt
u\������t&�G���6��k�ل�sf������4�E���Pi%dRJ��{T�O��+�ǶB�u8����������[��0h��P0�M�| ��I4�9� ;ӟԻ��,^��v����lE�!�Y��3�<3כ&����o4�o�Ԣ+W���s��f�#3�18��(���%�/�-�ӽ��ó���sY�ۢ�z!�H��B��mI���/�Ô�N�+$gGQ�I��|��9"����ڼ�!�=���)��м*F�pL���#���!�;�%7�4!^��|J&ݵJ�H�R9�~1�ĩ�
��
ۋ�����P}�GzYk�Ѣ�i0�Qc�2�aڹ�-б[�©}Gd���,�#���~���Ai�@��|�[�h@)4���Me,����ǩ���Y��Տ�k���J0S�kd��˥�CUb&�<4ʷ4�2�-`�-����M�hl�S�⋎���¯�'k�	y���󜬏C�*�ȅ�\ͨD���`E. ��H|Ӈ`��7�3�\e�.	� �xخ���Q��p%���=�(b�Em�H�C��-^�-"� `\����ÿL)�[��P�Ș�R-`���^n�~M��Q�|�k]�P��L54lN�N�g�˱(�zWr���8SL5���:�U���
_Atq�'u�:k��~g��P���4���^���t���Ǳ���Is=�n��O���;�~/�J��i�m�xQP/^��e�1W�z�*$8cb�M}j��K\���2��MR�)5��leYa3З���EqI��yԘ��,G�m�S���o�Ș�nF�w
14����oՅXT���wi�4s�?��*�w�i<J}�ua���;/4M_j�ݗ�-�VLs`Uɟ�x� ֍�T���̞��ҼCS ������Uk��n'�FY��t��
|*u��gJ��J7��[��Y�|�IpݏK�c#���yMU�I�0�zQ>o��k�8!y����  �Rq���ٛnN���]!R
OH	���;,ä�T��pCΛ�=��a:�ӵ�(�(.E����Ư5�tfF�ENLK��0�z&C9��L��Mx0k^VLGx���&��]�y��&5��Va�S�15E``���;N����&��� �x�0�1��aV�%xw�ս���#F��-��&�$�ѠMui}�-�JRoΰ*�G���uú�.�<�MD���]��=����,\u�`m!��L�{���K��?y�oA-q~�?e��(�m枘h��"<�A����ho���{���cs��B,�&�#���]-��|�ad�;ԘK뿪�b�Gų�ljl��{�݄H�� �rZ��ϗ`_�K�k�]���ɖ�B`��)���]��`�=�ߡ3�OI��/�� m�s�]���X3@��)���]�Js�BD�&���^d��D>�5VA����.��ZG�2h'u���w9��`���}�f��1�A"p�)�֘Jd�&_;��[���e�[k�[|�>�C�g�@~�0r��F]�V��"�6̆	tޝ�g�>�?9�cx�4�H��3t���B�����ѯV��XX�˼��劂�>$\�?�Xd��jd��67��m~,�Ds|�:�%�PI���E��/s���P�+� �œ�O|�_��Pt��I(����0��~E(N��x�N�n�hA��P~٧ਏM��,U�l�AD|�/���Hgtɘ��$�_n!h�XfOK�pᎊ�~,�[�=^ ݄K4�I$	��%��Kf�́<����(�w�.CB�_�A�>YS���(����Y�b	�w��7z���?�"6i��m꿢L��|M9C��!K�kǪ��>�<�CE�I"�w��M��-�8�ks��*�?��w��EXt�e�5��wQO� >�Xf�n󹙷X����4�Ȝ�7P��������4���3Y��x	`$e]:�&:y��^n���+u�Az�2����1i(o-sWG�E�бY�9���24��o�C��d�Q���$�NM޺�0�*r\f���oR�8S9I����ٹ��l��C0�[���h�{�*|Cm>N�r��"4�K��:������퉌VP��
�A����CB�c"@���v��0��'/���[f$SH;���w�b{��k�IuFh9@�X���? ����Þi	������-�&�k"���P����1n����,�B<�$��,�~�W�/���<��TnA2;g��/�Rm���w��5���W;z(]�*`�/P {�zDSpHT�gS��B�@R�䰎�f��|�hW��W�~wE(G�_�iV�߲�˥�t�.{=��Cԏ&O ͛�t�v�!�����o����JNہLOG�P������v\q�2���=Px��.�?�o�/�H8e�U�`d��k��@$��<�r�~)�������@5�D���*�`�(#��#�5i<�[���8���҄vt���hez�ءUw�c��ߒ�E�@R��[G�o�o-)�)d�`3V�<"z��ÿ���`2_�&�m��)j����jݾ�3�9�'YʍvFظ�V��zAv�t�y��߳X~�12�i �FòVFM���1��|ݖl�j �P�J�]\6��3a v-�5�I�����kaN����g��7]�����+yW�X6dyN�}^�KŊAD�/�%���2s��Y�>mF�Ajқ����㤓fg򦸳�v��2"_+�I�uwU�[Q}�SD��-��A2F�Z@��F�`�^ oû����N?l[EQ:۩ y��n�dO���rd,m�z������m�s�n�y	}�K��#���n�������T��愲�-V+��oX4�d�
��7���
��!��^&�.�D	.��n�R�l�J����7>���;���}i� m~��#����L�m��;�;����`����mz�&r�E|(ɢ�p�6�9�J*�I"N�OwC!V�{�j�6Be����׭'v.v4�jP7>�<��Kj]���ZfB���瓄��Z�8��XM ��Z�o Ь��x�;�ە��P�IF(��'J?��r�e�୷������iӏ����o����h��?_�a~}�E�>ot�l���15�q�eQ�{zЄ�����H�ZW��,�֍C�0����Gn��`�8�\�Ȁ�M����h��9�%��,faN�Ժ���{-���G,;vdyM�%-nQ�&��[h��Ey�%���JL��dd��PB��`����T�V,;��w�ֽ����bU�˼�*+3�$��	~�o�ipׄW��7�D��7�gE�����p��f�+A��m��z��'�Sg�Ԣ��h��i��<#�>޾d]v�[hY�CE�Ҹ����=��>&�s�cu��^��|�,@E�:ނU��s6�ӆSwɍL��Rr�Lϛ�*�M}�n��#h�:CJ��wǆS9螹,���u��p�x�xa��ב���<V>\yf	Hm�j���D����٪�i �|�X�z�i�now�$Rq� ���]���[�B-�0WB1>�����^���x5l��C�8x>�p!���*�	ź���(bCȕ�Y�拉f+!����<�f�X�Bb���lVI����!�٢6�O��@��Q)�6����x�Z�̭D��f��Pk
gk�}��m�Ә����ꠎU�
�?�ч���b������F�75$�P�b����|[���q��iR�����"��APa}��$8@����[����'A�m����ߍ�J��Y���n����0d(�+2���P+-�hz|�A!����an��/vz��D�%��{���:�@a�CŔ�6I(�o�~H2�L���Y,����rq%�R�P�s-DH��}�-��Y4�%]@���U�*���b0�:��=W���Pq���!��g�Nh����/v�~tU4h3Z�Z�� ��"n�;�w��i@K	VwSu��#s�Y�M������}*��痞ۘc���\��;��Hvc��� D�?�ʍ�G���;.�\��8TV#����<���*QLmi>�^�k_�i�h����Q�R��tS��y���*n�{�[��)ZGP�C��Y,��.��p/*�ހ8�DA�40�,D(�`�NX|���Y�L��HLB�����X�ñj�\O���	�_�Ll��^����Z:vCn�8����|/BmDSV�[�05����8����[�Z��`:�	Ob;a��>�z�,�p�O� Sh->���w��H��ט�K�fJBx���NGS?$�2�(=h0��n����1^�0�ԭ���"������\�$�)�{M���K_|b�i���fW�bE�O^{9�GZ<~:w�#)r���*�nv��o��8�T1>;ey\���1vHx{5���n�U`����c'��/����1�*�dkb ��6g�ب�0�ԷQ2rx��4�o����
9eE��x�0�@�V���l�h|�u���2N�Uk�I_n�)�B|���#����4���e6��'c�E~ȏ��(-׉�
?�^^H��(�H_lc�SO���H疡+�7u�#V@�EB�� �j8�ԫ#���kr���qy�󛯌�Q`�7kgo�����Ns������3�/��׎��k��2/�2>��%�T��A�]p]�@7���
K7b���ٱ�e"�]rj�I�9�G���T��)�7<� -�5��^�<t���"	]�Y�}!�+O���K��H3��n�h���CJ3�Є��Y�`]xN��}�*�3�Ba���
ƣZ{Y�G��5A^���0�[��w����ↃU`��.�A�5����kծ��P��p�}�%�e-�o�R�.����!'Da���85���|� B<i���a� 鎥W�"'��|)�}9��FtoՅ��Z�9xY+�D^aѮF��#�����$5"x���Ȕ��\9jz-���r�Z��z[ky�&���'�0=�D�r~�xI�F�yk�珛��܀^��W����b��k���2�w�YM/����������?(6�t`�%�k-����H��R6g�H�B>Ϡ����@�ۉ�^4sD*�%J''�-�*3�K�k5٭��̎�(���2*��s.��ћ>}l{��}J:6�R���#T��\�6&;�5q2�耀�ؤ�4��F=CL�ʾ��d=s����*Жg�m�Q�4	�KcT\�O�Y>�^�K͉�Ό�q�����͐%n�pa�HpЋjFx���Z�_���N�ް�`�oE��"+Ap!+#�����g2��;�EoN��+��lb�����{��̥3(�� }��A��b��Ê�&��8�Qː��sh�Sz�3h��Եem���|����Z��I��*�v�U4�(?``�Ft�c��0�㉳�R��q�or���>�
�rᖯ���J$��$�T���-�xF

�����������_���
E��eLE�YP>݊�RȎH�x�F172!�.*-p�$Hʍ?�K�8������*sN�9�v����$�HEK����d_�^�t�c�3���d{�0W���jA�zSRX�أ��ɍ�Z��z5�n�����VjS@���Uɯ���1e�0-V!���/��ߘ`B| �x1��R]�?�@@�>��f����)a�,7&L��2=}�l�T�|*x��j�����b�\|��6	n��l��_ڲV��K����,�X�
o��x�������;�`�=�[v�"HJ�şR�ķ��W�bw�v|{/l��4}:�B��R���\�qS�ի�X�Nb��	�~��:������*��� H*[�Z`<${K-ʲ���I�V�RD�[���k��}�/���g��]�j�f��MDXӨd��x%5t�m!�`r��+��.�"�U���_�<CM�h�5�g�W�6.𠥄��7��h��m0�=z� ᰟu�6a:Z� �>�e������5EVZS�'����#H����%�Z�U.F��H��v�4�����v	[�}N�����F'3�}��;B��~���Ƅ���ǣ��*ý(�T�������9w�R�I��Z]*��d<�^[�^�,Z{�UM�z��ט�!if�Lp�s�'�nuϊC6���8+`k�?���`/&Ԕˎ{U<|V�}�H����
$Ug�[Y��_��3w#��m��`?1�V��qX��U$O��{����dp=Gd3��)�ji�mr�ҷ���	z��ͭ�>�{�["��cx�~�C���h��Vd9�~m,�8�	������0͔��W0�r2���:�XpB�]o��e#�A�찼3�=�ɷȃP3���������/ ����+g7W���� ��Q���)� 吶��=#�e�q�]��q���ճ�&k��W��a�"WDǑ1ޮ'ێ��n���Ɣ�5���dÛ�G*H���ޱ�6�);n"MQjCI��Au`O�]�؋e�WiNp��j�6�K��]ث'۹����e8�qc����j��&�*/��:*´�z �}�ەc�c��_@�Q��kq���R�c��O�"HV���Hh�P�Bhb��GU=EO���(:5�)��Z��/����w�j�):D1\)c%A�I`eڅ��Zʷ��v��g3�׻]��hF�m��Eݲ�:���A�.��Jn�ڪ���F��>*D�[r��T
p���<���[E����p�N����b�n�ˣ�\|�g:����˷��J�o贒�v���P�~����=�)��]w������Im(#�qt�)�x��nFw����\�-k���@@<O��c���U?L."���C���ce>e��5��{cɟX������h}��� ,$���E~�@�W�;�vI�]�0N��g������&z�A�X�Za�tf�R���jX��4��o/�����n�W�%�}�\WG�x��-�� <,����G�b��j(�ҹ74��C��Hh����W�O�Іed�� ���+\rY?�w�@L��(��o*����y�ե� S�JI�x�Պ�{ȶ�|i�>|�,X�x�9)W�!?`+]�u���dT�{$)�?��#�cb-�0��}�GZ����e�ޢ�|>
�A�w��A]�-~��YR�r5$H	��ҙ��$����s���䈠$:�3��Q1�-X�4J�d�G,q�T������0J淽���+[��q;���B[Q�+K����e��9E�A�]6"�J6��v$O�`]�L����B��q�#�%�\��h���[1��/`�%�>�*S5y�j��yv]qʨ]�m��Kj$�D���u�Į����AXT_�<�t[҈���$[���0U �M��gg�1�7���������nJEJ����H��F�yC3�
�rV�0G��h�N���j����w���zyp����v@&�Dw��P��G*��ؖ����jv�k8K�q#`Ne&j/�ٸ��5&���>W�����Ky9rV�SA��ISG�F��R�'r)��A+�\����g�\lD �P4��%5���J���=��Է�|�޳��e��c.M�֯uFp]QJ�,%X�tնwC��W�'>��=�� ?J���Ե�S�}���+����9��>��Ν���f��z�m�N&jUL�/<AAt�	&�������H�C@��߱��5�_�����24kCb�#��A�ֵ���i5qm=��í�r\����f�>M�����$�T)�$d������[�̚��+!�A�(g�B�J�at��K����-�imj�	�h�Cミ�kA�e�����Yڒ�J�����Rf"��	Z�#��f��کX���f��~'ܧvDP�\���ޯ-� ��0�b��������
7��z���	9���)�[B̦��IG%�W��ʿ1����tݸ/������Y! �>x�~>���]S�
����ic�3%0�B�:ke�^Zu��z�:���M�����n���(��Z�� ��P���i��p�5� ��@�T���F��:�2@C�~*�jā�)�@.���b� ߀��! ��s��_[��`"\
V�PM�*H�u?���]i��O��UryMi�D�o'W�,7�P��9R���}5�F����,����s�o��1��N��G39WV�^F�M�ۿcPQDKY��ʕ�)��Ս�GŰ�����H��,6��0�~�,2ߝkBG��/�%r�
�D��@!�|�.p����� �=����۴�(|�I�����l�B��:��dwǔU~���I-��*~QL
���V�`�=\�J\����Nð%�]�9T@�l��b��i��K�|�u3�1Z�훀ٯ�Ee)�]X_�cC��N�|H�{�7]���D�%��`��Y�J��QC3X�+��{��;��K��C�?~�<��S"r6t�C�,"	�V§���e� /z���jһX-�����!��=��LoV�#�I��=Ȱ��$�*Ժ,D�Xn��E�\��;7�MsS��vJ�ۆW�a�Y���-����=�'����![d�e�v���mu��\O���-�W��s����n�&�f��(TЉ�G��ƛ����>b����|�#�w���W,sfn�BT������kF4���Y��r.HQϖ�s@tI�Ws�uoΕ�����c��e��{��F��5;�qUY,jJ��|�Y�R+�J�K~_������3��y=�O��������� ��F+���+�o�N�@�}��K��٭������y���`���P�k��H��!"��f[�D}�Gjf�X��ι ��ٿb����xT{$�P���� :��}�
 y���A֦��A����i��7\��+�XM����۠c��7�.M��3�&�Զ%^�n^��{��*�-:?�ann�A�y���W�