-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
F9V0QxEkK7cw3xJgIe0Ax6SCaojDP6E8PRh64hb7ZHbKlXYUGKEFVXazYkutXO4OqeKGxbgbafmh
vaRleF0Dga51E+ZSEtb12ulKRCYBtntBQ906zTAZQuzYJEIXj8+vwWp0dpZyZO0FGFYXA19JlTJa
Hv+XS6t5hlmg3TeM1Wyp4l6IJSLJBqC+xUs8u/UrOBiREqqNP/3qlEuQGhd+pS3JpEE1+2iB0bCc
+YQ39J4Mm4l0n9Qy7D9lOR3ZS1X+tGeIX3w2BAeVt0O4fAmMMD+lO0g/CYXpPcIajJhyBMD6W/Ne
1zd1PK6wl30WgXcO+pWJfeMYcvpLJOaYbAw0HA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
PmWAyS/VJKD58A9DbioZ4NbwOYYjL0CdSfycEJIKAlgwa671rKuwRFsSBpul7GGwYzFNcwvSboks
BKl8duNgRYI+oa+o+qGEXWNTH5793miqgdiG2Z0Y6oqEGsGE88DJnRjrUfQCDvCPe03DlseFTjFA
NrEIVojFmnc7Mu5hW0fcwWFq8rt0w0IW4G1fDK4T11z1gbN+D8EcM29gW54863xbq8SDpzU6EBsa
lNSwA6uuEttNHQqLxdKwMdDZeWaSE0Mdvr+4XqzvTN7FwWmqTeWRvkFrOm35S9Dh7648jAZP/1m+
yEMf3C/GHd0hwh1UC6hHlIq7EVOEcPnH+DnLFsSjZdWPLTvJftSbhg9NoJNyKf2sctiEdxYzQL2r
v6Mw10g/1wKNxaTSFBrt7tfVLTTKJtfS8cahm+7CUHoYLpI5xrpASn3/VzFXQblhMbksWaFHiWYL
QR40RaOH/zZi5kgDDea1f9GowoIe3jO5v+FKlRjXPs3TCEwIEmazWAPG686ISBRWjFdVqyoiVrgI
mb7F4aWHHXqp4EZzEg1gQBb73UZgVctQrFjX/TA3DdsHmiR9WtVxrc/NZOGN1zWaUD7lfI0gvgsW
q7uCnO8wyEUVyTGos2Y2NkJy8Prz8ckq/k8ifhXPNBOQIniz4FhDhjK88IjGa0Gxu4UBmR/saK7c
oKxEjjr5NJiiKyITDY6bJaaRdUwyre1VcIOd9kR+72aXdBPv5lspOiha24QiDxi4S6kKIWq5fOra
2mwq2dz9aUJIBVDhWErbPiG2UVyOzSOVPnjx0YcQOEYqLJpVqsm8UD8mT8RbxwRcvCbcoP8TaOf1
/AVHpr7gbChgamPOiD/1h+1S+bFtvn3EE+OHf2t7z64RP3LrIBpwUuj3QZ06GDc8Oy6IRXJ0+4oj
0AZbVErKesE5VSLRjPqAGXiKP7/qzYkQGfNwdyGfgqGtg7huyacKyi6k6ARrwA5d8MQHbvecWepJ
RWXWAw4Vd0+eGdsYkZ3oIKWGcoXu2cxEl2w2S6BGknEaIk30QCHX1jJDP6S0TJU11U4LIyfAG55J
rUZeiTw5NsllmrMtwTTouKv4FX+ihQbJzjF0RDfkpvYcyh0sLlVFPDiY1EZfZTeYfGWsVb9K66XT
zzjhYnSiwmpTgLiV7ShXCx8+Zu8PD++ISArw8gK1GH+DN2K0kpSOIkTt/SCqcE+t6Ml9v/Iqv2Iw
BiVoiMFTBADhaaRQlGh13pJbllehqhc5gaw5Hqw7kNgWUeoCma4CR0TwLxbt/EnMFJXKNyMvnl3Y
nhry3mB5BdOapXKIpUGwYo+AfZAHSu3gCcqLoAvD9vGWZj6fqOWPPAmBQOTrgYB5JSY9IjMq8tYF
8UhC+iKLhldPTqppJ7r/iCUsM6cPzbt2LbmIoW4zod4xlZHPWl5WDVw0qj1sv59td+KwVNrrONaR
e6dnoX4X0yR8H3X8FxxiwJae1vAojRvJRTZaMPotgXEMTHTtxrf+eNfA8GHw4Vf7cWGRG66rdCEQ
i0j6n5jqMbc5ja/+pfjQr14GJI4oHfQxfkobjLjU67HYTkNUhhBhj2Z01U6/mlWS8A7CHCxuoSDw
95Csau76DowachUtQtn6EcoceEGt3N0xtJjvb4M5+aBYwaE5OJ/HmAzHDLk7MtGVxZ3OI6nY1dS4
aXLJveT2TbWjn51UxR8/eU6+4JeFWxcfDffmivwZQXgqpsZ/bAHvliGrFlg/dxXF6AKRnMI6vcky
cw/u8theJRuhdDgjjtpZQFtEeJnasw2K0zRDUALckZXAFnZy8LiPpe+kG+2IHG+1pXTJfSET0y89
N2vC3+lH6gzvpqqv1GzNQM8xdbe29smm9EfgHFbGyU3nrIu0UyzQgUW8lih5+V9TbiL6FINH/JmP
ZxgtsEROUoLg4uGKbagUtHt8bHFN67lajasJBC0jnqcAOK5rTYJduCwvm6b7p6fDCVIw6Zn4S6pU
oOm8FDG4LvYDXZoSjceUtJ9drWMeShIHeksHgLevBuxfP7TIJDL3abAfu9L+jRl1jog3ysRXtjR8
scaCTEQjNnili4HWZRpQ3kD8Axd37uLAJSFJkNPEzAjp4R55m9C3xgCCnRrxq7FFtHA1jFiSpaD4
jVVfehxH0nWlwPWiNKpKIEulraik6oOLywJpzH+PBeVUqCxkeIlufzzWP5lAgV0QuFun2rkGQGLq
/bVka5HCFjlR7kx35s+TOWgoS6oASmk4zLKrdWKk6l1zOKehkDtoHEN+AQPHzU3WDcD0IxIZGGlE
d7Bl5ahc0VtWLtbQ7NBVTtQU3EuIjfcrSejBoy28oeOX3YxRv1LGjF6PRhSSwhHxKB9u1ZdfkWJ/
wCCfrny9smoVnoGHjYhMwM037jVH87UL4yKKRUxYnHJjpw/AFELFZ2QOVxqtGru9i3GIZzvUTCA5
f2l6J3MXxJF3+toZRwSVUxifamGXw6WfacxnTO2ysQItc2j3bW3c13kKxfUQ1EqbbVV9Vf3sTPR6
Adjnn2RqzmDReHCo3U0UQm0NOZO1QmJacYROQLRaBksS8P9ftWiN2GpA4+0fKgzOZe6Ps6FZKeY1
Cb7wxup5NRcszwhvtoy9HLOPYlqIJcW/1TgXDchDjTEmbcCPQf/5UlCC3hiIRYR9HelqzEaAFd3G
USjsqDLGvFe2ppoSv2QsSBtyUYFT5QDHfENmLuLLCXILkGTwOwoTozVwAIqGsxWGiheK71eI0c9h
BsM37SEJikEYhUWCLzRRaH+HThxIcSdiPsjD5ajPXhzItXigYZHZu0vE6aPFol6l8hUVoporrq67
+/XJGBxOYvFJlk0p7YfAxTbOQbr5wpATRnnuqol+y5ecnAwjpQFD0mVZ0TVqavd+nHoA7ygmc0GL
k7MG/k7fUOUFUgxIxeZ5JlaWBU6vgRu5hKhk8jyrNDIG70iJBc468AiesPeSUc/ST8aYNsLyedz1
JMvx3ZLohaJlrlzIzC4v5IHuPeNfCLVJucFf3iTzoWWi9FWOZyKYfvO6Rcrm18xGrhhnir6kNcy6
uAMgzO+dtcO+j+A12IbdJyXMrt34fPtNeR04LJl043XeISMkN8pFDLIpGqv9Tz3yMD6JQlxCo8XU
LalAUPeUlF12V3GTnkpRj0dPuWfy5rkcLGAj0JjwfoCsotlBQPiy/Rej+427jz+SqQU50ljNH4eM
505Si90HSk4in5e9uEn3i/a9Un81zfmmba1CFrCZugwShz4ikH1HK0Z/YQS4TVIAhqVXPS5ZKGXo
XQHME28LYPVrn3t+qmfkTL2tnHBX4ZnrEDWwJGU4549fLajsNg1YiINy5nmZN2Jl4v4S2st1wWXz
X5Rz5gyT01KMqiAeNJNItbL0CBhFrxIeBW33fvaX3diHEHtM05GvFTE9iphypW86LKe5jb9jxja3
fzx9fw3+Y7aKehAQPX5PU2phW7lcDT0wgB5EAOgBMbmMnVyfvFF/181uDZL5PRombYAndL1h9CDc
Zw5QHnQUi4Mzszg2zu4cZ52iSnJRRDfnfzfALCxm9blOM6s5XLBeI+5husA82Ae8yM5vreLLctrO
AVJ2UbVpdXhclneFqFjqq8Qm8rhmDtinCohkLGG/w2JAnyDYqw2HLh69pKlL2CQyd/SEHdfk/lmM
9FkLi2ExumAFDS+T8LXIpvkOHuKnurLgGPUGsHpENEpaLVAca2BczK+FIRaapX6F+/EL9pXduMBe
F7dqcralfPHlObpBJoEKJq1NA+S5BGoJKhERqFrlg8N1HwiE7K0KtJpDd2MgMD3mdUECherG3gbj
iovJEDFTA06PlKIQNFJGS9LL94m5agrK1gdl+juRcRNs1rww4k+eTN1rbnxgQOsrwQy9jDkw6WpP
L1kaYFgj5awFC3d6ftuJJr8DYffSmPnQj6a3tipXYl9YTg24CKkq7ObiWRR9ugrz1cLsPNPSKjbs
qlO+MDvIGOEav/l3WcB598nqF54nlpRtqwlQDXZ+IsOtXHm3jAvkz8xmgRRJr0zKTSorh48mzLvu
RYMBwmnvxT4ZtODMn9nqpVzHHtcn4PI09/Rsy5rLF/sWBOeqvArTWPKu1WecWHxi2HV0GWK90NKu
h003Y1s0luJK4Ef9EDLKPXelH6MhF4s9oGbh74kxeQ02kEjf0Im+rpGBN/xjeSbp58GRDggLSS6Y
iBVsDk/r/jQVlsJyaTEa9P3XK9iUYFIfCP7H3fs7T693NoVUHuJ3Ce8m/dPWC35UvR8cBnrp6kiL
C8Eez+AwaVLQjelEo3eY3AQb6U/83XpIo0cALAS6HJ1Qb+N8P6gQe2PHgYHQbsPHgampjadfVqko
bsI1pXfFZC26xI/fvUqgWhLKlzBcYweaVCfdgmGTBs/rklCXmmxhbJOF+TlRLy8iwnzTe/2HEJaX
x5s9Lmcd+ZF5k/ZyEhNL+HuYaTIRLQ3KWcJjRJIOCm4/+piubA6Ev4pLVe7Q26XOP/N9GfVEz+Ge
ohHpXSPyhdR+dJT9OfzYGmFv/UPjOBcekoJ37AuiSWhwdmjWuqSpVnibzXusavMbxM/Gs4DN9dKX
z/JhHJ3wQO8IPhkI1n76zsLGmDQC6VRM40gKYjAJla/fjGUEfQD+VE2+DIAu8267Zpgr7rH7Ax7H
cDMjX6CMilMArcChHBGuUaE8iQUSUwy5g+FZLyb3KjX/32VBCirDjIgHvz21rOw2e2EDayXo4BNX
mbjlAHiZthR4wOMAGy2B7asol9GrnEOikm0P3vq40ZrDMCbe2gKejrCKgreF3RpSYRPEyvx4/Tmp
achfJmL9OnK1DBpMAxWTYiHIkEOlPP7I8ly02Zb4HYQzOPkudDnzEEfZnQ/5VHvCUfrxT56gBYV7
BDdMY8idQ++6Md4dhsZPw6HDTaGr1TmSIIlE534RGpusCR1qW9rZndgPxQ8WQ+IDwlkLBxAiFUBY
CltZlIv9N+4oz7fsa7mnatSXy9gxPqNiEB0/lcXAlFLS6SBbK5vdH8LAf7ZzzqODu/dJXqcLWmZE
Dwysxrr9qsCBJuyuTK9LElxuEzJZzJb76J8PUxQfsR+t27HxdNuA0eZ9RXpWssbLDRLyfJPad6Fn
d+da0PZd8Hk31bQ/qdD4zb0PHCqOVJ01G54cUYqnAdEVeHTExHGKrLzSq/BcQ6o85coUCJf0q9+U
GaiC+0CIHCC+SiO81UAao4tpDwI18xAxmpOd4mzWDT4uf0dcUvDept4cXNOsFHSL9GvKDVVZVbYF
J3CCSPeMWhsSstsWBqbmGz8+wwvN+xDoaKhX78x00oSQaVE9I69Spq0X3ipfA9VekBoVWPaOwisc
6ehR6kPhr+w8cMaCrgO6q2pqXZYUCIGkf7rQOmSkM0bydM1FLPe1+zmfZPZ1Ucw6NHQhRXq7gI8q
Ml2fOzXDfu6kIIIRmEu+0sK5mXrHPz9HOauy27IpSxwjXQmxuwTV+6fL2eSH2KnTc6dzS0AxtBEy
9MtHfkylL6pGnwvBIsLfY6H75I8UtBLeoCO6lZIEja5aU1JLXpJdQL5TJw/DkEA5Z6ZzS7mCNLsW
wjmnOW2hMzzKO9vKNAesFnf92iao2RSIwAA2EgoXrvzOTjrX2PesFXjxCBsmwSZgB35s3TQ1L/yO
I9Wj3o3jY8//bE6mhbAQkT0MaFRHeN1wI79X9bQh4TDHyBfO2IkDPchVINL2+xF22lZkWJ4+k3VL
ARtZlYLF8q+GNgWVSihKrgl6GtpySiGmzKePXVTbFFju7VGJfL1ARp4kBkZnAutE8L5bhXnBQPc0
LlO3h6Dm1iMwsW5efPHAFhhmzG4PhKm11Bk7t8o5RcnRwMyS5S3m7suPSg0ulVXTj1gk05C59jFC
Q55MNThkrDoedfLnapqKyG9hecpHeipj4SGNmRm/QNlvoatEAHchBObZgFAW/ju33kXWvDLSHZly
Yfgpsackw5qRZjYRYxJ9BvxZbvG7txK/xi4sqWbVw38bcMy5B1fHvTUgPI0JxmOJvpjM/YdfwkKG
PZ2KU2qjXgQDPN8mUW+S3Fos1pKr9AiCKMXQpaZlxqHmv1q5d+Gkx0bGOGVLEYd5pz2xLtZXLQx2
d1TZfhNwlr04u70nf2AsFS7lfdSb2mtztwmUKecVr6Vrw1Kl82Tqj2zGjZcHwMxRTdq6WG4BI988
K6RbkpP5o0c/Vqu/52Ybj1wN1uoMpVxr5R2j+W4HELdS+Vd64/q2L9uOgb2saan/lS+t5W+3WEch
QAYbs3VaeQh2u8W/ViXOdBdZDwlh6/zJF80a4hvWjkBG9FM4XdJ70OqMLrsaH1SrtBYaOP1c7f7Z
CYSoAwkRVBTEj1yt0z0hNSGOM35URsyttBF6GSrNp01+EpkJxUzQGOm69+a9XG43QZo3vk/ehkJF
gm4bEA+5c9nsgZ5j2vHT5yrOsr94z6kDzNTJcmG8PfB3k9ALxc8q8xSfz7LNuTd6smxHOsoRf+7y
c2ETVx5EtmKPzgrigMDzBxxcusjCEmm25yyTXn7obyU5kv3d/n28eTFUs3ryvqxM2nhQfT2i7/jR
eahLwF2dLrt3rZfVFdgasfSRqyPnLur69aomu10euTOyQwDQmM3udnk/BM/HXgydgRCI7AK0WR1c
2qnAmlF5GNlI2VtYi//SXiVEQKy/MgzootHDBY2q4am4jj0yGJhUkxkpyvwWUXJGCA4aDkm44yXG
5yv6Xps3Bu9BxYh+3RR/80s3afcwQAYwM3pHlUtWzgaYf4nDJsVzfsNvpvwzm607fqtd0Wi5jtc/
6P2HgHfEKPA1rG08to+SSH2lGCVY2qLYdBE3sRA16qHGv0z1cut9paVjgjDK6gGl3rUJPSK1sUDJ
5uhSiEhT40F8qnZuCAbU6Ukcp6zdreCW2slHiTcgECbiqKSoPoUoAKWrm1RW9u99te9MLEW0C3jK
FkitZiQPuMMBZXh8hSstxKU5OqhYd4KluFEKdw1dEqOdycUGt4dBq5bzlZt8asJTJMiehdSoviBJ
W/sc0kR9uXo1C6cGAG4oT/peUkBo8dW5n4L/esybxbHQtEbWP9n+BWHd/cQFEuRRQokGg1eQDapu
AHQItKgRaXikfezfu1QnXx1XRJADno2gO0LL9maLp+a7veCL5hY5n6KF1VJXL3A+49/Tz3U+bO5q
e/6fU4jp5nfZ+s9S00Y4Zz/siEqa5sQNeoeGRLkbVQsM/NaQLQ5j0HcSOttG3e/iWRSJ5wDA33WZ
Fv0dXAFLCj82MLJJ57N9Dm6Na5sd7JlS/5358Fr5OXXQWKSSdD9CeyVb4YYAw8tr96tM4pd9my/M
+p+J/nsAfDQISrM2fY981qN/YBsK/hcf5xylJAMdQ2R4t9QDlA3VtUo4W7w3pqSxctIqipk6/Qy/
lrZVwAQU5MrVk6tEMkkILMCOMP2SEywp3IhuFykIfOz9NA8mLi3BLKpsFPUQbCooFv/IqHtUclv+
eAN0B8nKzLWYZUliL8CxNUFSNWjpOh7P2YJx1TaBWb6OybRgKTMOtYY8cxlgYfzkt/ZVfMvzl72c
uCBdl3VyPUMeE3Wggp7Vllvl7GEey2Uf4drJAIhiMSWQfMKi99qNxCB9uKWqyH3GizThN9cP7zbe
tKQ2cg9hrmOcf2jWBldltX4kLCOfY1yOi5rSceV2BBNa3wPgTT53YMlpvhsVQbfvycdjMGFunARK
nWOna9DvhbkU/bSxgqTIG2KIVc4RaBKOuvApi4WnNtMYdqnqnLh93bmDT2SpB/GTJxmd8MBB/Zrz
2zPWHED6KPnMIbFOxVhPnxrQf2DMhdVDr1fE3bdHcbltg1HOH0JwnO8iUMIy0Cu+YIHDPPlh1b+c
Mhm4PYlQJaLlXHsgyTl/GuQBRgVyOzEUPn+xtz7j2q3FRurSEM+uWBg42oLgRVfgS2s5emuhQDvA
FBsuEacJxz6ePe0ewmid/AnWxkmTTpy1ZqXFAnQ6hlExplpcRIBb9g6lApGPm1CoXC5kWQLKBnAh
+Wp+6duxOGwcZ1fzDEwpINTpialKF5DOm01z7LnXORnf7yrI/TVgW4axmflYYJlvu0TV3SL4Bhwc
QU1BXy9ikI3eapcfdrfyejj41kEgd9vsE/EazW5DdCC8spRBhywU0hmrYGJVDTcI2AuikQnWejXa
TVFMMQLPH23wKktmazNCb7iaO2yXkl8ztrOPcLOhNugKe4DwuZVBfdemS13OghGKWVwlX2CBBjfu
jeUQxbIcw32coNQ52bGSh9hsN8S0rTyfguPSJU0Edquy8Owtkpm76z5Zvkhb1ZwySQeww0vB832K
0oMmBBwFaxztnaF+VQToATtjyC8PFGbbSmj5rR02V1eH/Wk8ctyADG02QzdFMFKKIBORW21bm0eT
//LctDrCKPIwO1HvJDioAfJCXScYcODL49G/+FX403TQi8MZLP0V6o+HgMH6X5wt4XE341u3qbPT
HA5L981w8027ZVuBI+betNhSwBxZytgJr1442v4Uz+4JnmRNXBlcCg1K+vtqmsYFAflb8tlh58cu
m2MHcKktaXr9no5GriIeY7Q/2c0NbZMyOP74j8aKwqw1ho2uWo3hv+5b/TMOmVq1s2nstF9TcyJu
iF9CYqrT8RQ8qasAxgI/2c38tZtaHavYdtG6O8k5kXnYUA/jR1+YFehGLv+Q8YlLYPxSP1htuRbZ
RRX2Jl2fFm8DWZdsrADyx8jKU1qB/P+vT4tAkvsL9h06ZcJlxb/WabGOvZoezBdLVAjS11UJJ0lh
C8uHAS19BCBAXuWW/Y7913XHXGKXXOpIFPARC/NAMeNj6qbv4Ohw/vWREmcGTBi9UITigEtIT+Yy
ioHbFIY2DiBRHyKJG51c5/bPzDuOXWjXe0o3p0e3efZvyrhhGTXagzMtRb26cKXmf8uxR94wc4Vx
mh2jukQEbcLI0Oah4mw//q4tsjntIdvA5bqUXKNsh4t0hJnxew3CVedqqyG008xh/zRsGftT7sn3
nPJm1GwhIHZ73i47HWxJfxXHIflEpsBtN0rIa/ryhfxjboO7pCXO8SvPF5oLHOHLPuwIaglmqxTF
6jX4t+e347yBg2xkQnpu2vbVGQn/nr9JqbE+ozhOIT1Yw5A5gpyG0QGgVCgArmmXKwomBd3iI7vM
ksq9/xjOKcqSFZ6Cx5PdBCHqd+Und7/P3bkhJA16bsMasDEzowEwPBP98PQmbR8lAWzO3bnFVGdZ
UUp6AH7RoB/J+lzgEVf4+6VMNgarNVC04W8btNNNsVzsGtZCv65uaOactuQJeBHm1NhTTqTFUtjD
ZFMwcAlhaaOTc31iY6xGdk7qQZsY15ooVhA/MBmMXUfnCwPXTN0nuOaY3SS1VAnuVEfdX0FeODeD
1wZG+fTiOy7I2czYc5SrYezm3yOD2aLmWoLBaqNiIJqoMCeB5OJRLKDGXLSetuqGZXX65qOax7KC
yc11gHAT7/Naegoi2F3aIF16a1T8lIwhYPWDCEqcfHCMABvjCkittVn1+EOF2oYwA3tm05hqCsOX
8d3bmfaJjQTH0zLN7lB6fEkM7k9S2heHYqBltxnRckMgC4x2HTWgfMkosAN1zknnWldme+PcZWOH
c0IJEevda1vJPXMVKE9H/9dj0ZGGuM39ojtVGi0vWt8tjgJRVLAgbTs3DathXbal9tKukEi+rGpo
lMNBcF7p3XffOXrmv0seml7qZE7SAv+5pxR/7nf66bv4/9PbPeylSQK3C0LxC792aDKknVJny06F
pHYngL89JctlRnecsco+kVJduDJdvvAXc4QGveeYCcNES7XVXIsYCvBMVJvThXF1Gh2knFrEbPwB
pLGcrmXCGSyecU2Alt8wr7lMPSH8/UNPRTpkL6jEYnahPB1SUQe0x72Yw0rH8ICqKuBO0FfwZ8QR
zqBR4sxOfZqNAR38XGxF7lLQp3X1iNObO5oBR8IUEgEy4i061j3Os9CdrCe4AeHD+Ghn0qekqTyk
HFghMfJwdPyQ18xZjSS/1T4tC62FrztE3hQOpCiWH9Mpn/nN73aqTQBYzeY77bne2AbkCp/LaT4e
2UVlBCD2CHlOmIfykupfZZinjMnVdO/3lSiPZWrpr+sUxpkmXWU0r1jlYsSEO0hMSlKWX3Wt27lM
HFUbNtdYmnWEADGIjuyVbyELDEZkUZ2YEnOG0bzU9+S8AJBUhL+Cgbay137ywSYjruguu2Pyq+gl
5+FtQmJlPDeugACO8/t+595o9BY6OsERinLkr51yeDf+umxSRi7ziqd0NITWNCcBQkStdA0W41IT
LFoB3iaZaJUyGhKUEssDjqVdQDiI9t2e4FjT/5OCT76wPeDfrXWuPTEIYUf0wW7yI8p03K5fTE3M
OtZ/0dDNIWxuofnX0jFwx5QTHb+fpcn65IsjIRptReJhggSTh1bU2Buvqsvzz4wSPo3frrY218d+
VW3wxff/ktlgptG+Wk1QWT85BLzPUDr5nY2K4C2Huq/ScXLpZEaA2NlDI8V/mXhCA5hBpaiCRf+A
wG0z1WXEgKFnF/AlhY8xRJi3uqRa3fbR3/Kf4g2hQ5ZrnJBdMICe9D7coSn6AAs0IkMNT6/oOxt4
vwqdzBaDg/kl0H7l/vgcDqBrvetUMCVfLnjii6z/QXvCGZtLduiutlSJzWmBTAyjB29xGtzrXAC6
Gd+vVy9fRI9VSb8tTz2mkVHR8XNzMV5g090QfjkFdXIM4PA1l8RNkfaxMDJAJgYYyU6+5g9N/XdB
rk6tkwowYxwNiKFXQ53f6OmeberLjns5xgUBd5jIWOcaMqd3ShvXZobZGprqDS9vWomx4v0gF4QI
jiHCBppFqYeSGN4tzQQ5cvbTOqoadNIZ5NWs5/raN4FYA857ACI0p0aiS0MIcwOkweelx0MUIVtf
G86rhGFMyDuRN9yf0R9PjoMvey7FGcsrmniyU0sPtjO99Zkhx7lQ820jbejAEcVF71JWZY8FZWy0
oRhjZmsFQSSlJ0wFAnflCOLICpRu3Zfu6pE/Q3rn+Cr5xU8XV9L7x7feh8D27+0LqTZocaFlTmBF
8bqlR2MwXt75mkslNT4+SUjKF3B1X0t4/vjsZGm1v1oKbsifCjDUNmM/rVkb8JFaUhot58SoFU/x
EoUZWBZNvKqiMNpfmRaTf/nHLgkNR8OezZ+UBSNLjyCObNQD8hndp8IRTnG3NPbKKVX/dJItjNsI
VyYrz//U12Smhvi8/ZGp5TC37C+TXyNiy38xnIqRHRj2Q24HsDNYqMqsexVolk37AA3Swo1ffx5G
1kawkzevUIcm3foNU/oHoeyirUP9JOj5/tMGEBnc36HMQDpRZUeTQH1VCIgnV/DoAGOGlKBNJkFQ
+uKrCzAlJt01VtYPRezDexGJVvATMtMpZ+62cl54NNoykxvpq+cGTNRZtYzUKYN+YwgZ7mKWitrf
/rRyvuw0TnkkO80qlwklf67GIhLSJrIWYLam90NBTyC0Uc5qGv0n00c6YHeng7fLJjkfIqpA33g5
mXV8sz+Clhpf4GkHtJka7QrpKB8tXOfQcz2r+Un0aD9IzOEv8Dwh9jfUCqtrovlsn7ebV98x24PX
JD3IQP6SW8OpGU8Vj17YrgTBzURMaJ3L2Qq7uw/AhMSdRDQ2SIo9VP8IKQ45G8rw54TMY0rkBkmi
fbTYUOEKwXTULmayTMAZMRWgNyt9po5Dmtsx16hpR+D0MXCzji8QZzZ8PB7FVQ5gC7ozGozZj38y
F2C9ulxflJZZUEJnosbxr/61zgy166jtP/SEk2FcmHqGcL69uh4bpmX5d2vd41dGtej+TVnMicdo
yQpl9aEzuSNKlZHwbQ==
`protect end_protected
