-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o0MJ8bFRHduQRC9vNu7tv7YQlbehVKM9zHWQtH3zqQC6V2nWfi7I6evT405970NZ9A6HMVa82lsa
mxhoYi489jO6kzOnqOqYQd2RjBQJ2SthMk4ZXqjmzDKlDChCfeL1MMhsRZyHGYGWcyy81sT8os0P
BcgZThZeJDZPrNo6hylzadnrjlTrrimgGvgS6w2orNumE4/192OJLFph7Jc2AwsFaSi8MyKbnnA5
0jwOV9NFPjH3MrGuV7feiivpseYnBIRLSG/Wp3Auk/qSgH2vfAluFXUhSmINiEhqSXheX37zme1O
pHUT8NBINZ8X7G4cIO/VVmYJljqh8d29cB3CGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
/FygmR/Or2AG4YqupyvNxTQhBJp/ykJ/kQEREC+w2BsKoI0AsZBLuSSgOx+8aPIEev3lYdXrtn2o
++IM66qNN/vskIdlIzUn0UFNqD9D+r/NkBEf34gorEF7EXsNm63ikogk9Zf7XD8Z4tTeF4MJQ6Be
Rlq1fKM1uidgctRNw2M0rOVQmITrAykQVIdfkGDCQwN90SuDLZ+Qo8ufFz9c9xZCNWiAIVvh+KBW
b/jkOU4Dr2RxdYpfNIN61ueuBq5x+czQWJYqLQZrPgKQptKMIvznrrZ/3I+kLYtYEAXv0eYuDt5m
kUiD7a7F0A+tvoeM6iN6LxwqlXjwW1xD7QLCoVILwkDv7D7EmUVO9VyEBfctmYfYCjAAdutyACV1
dwcqqCQgCluuCOpCITF8m/7jq2EVjyXbNpMAgTgU1Kn0lfck5kaFrkNtaAXrCgHt9bQddjX1K3fJ
67P5mz72Wr96u60jiIWqOEmG1q71RaDQVK6dnXuza0XLcWJexTu1mTlBxpZlssDKVupuQ38TEJOl
ceJHi+rvq9zpHrQjxBMo2wrg5fqS4gFfjUbIEQNH8yU4izsC52uSRLTDDtVWlXi3oh+6z82aGLT4
XtYeK58L04P/NUfdnIiANjlH7SxpR/mF/qArvirTdHaZuuJO5ZDSHJdLPfcyTpoRVkITHF/n+dmG
IIqk/QQYvJUAIsoUiXCSt8tPdjSQ5c42cfyRufEs/jnWDm04nRoG9hXS6ew1adANpO7Pfy5bBgMH
hunzw7TtUu07x7xjPSRBOtTnhM5oKRnOR/qbkrAQA1to9LBfKoIKsODkOENsanriN62gRGp0QS//
URDSWd7LwGXQuCdD6JCRbflR6Xh3jIg3xKt2CpARKJ37hRjqpX57rp0x0Ru+zlYoUa5ZoS2Dz31m
UAaB5re8ty50RWO3C7jJiYTFamFZyytANf7krMkLdTj7Wy6gUygviFdQ0Iw7dZ46beNFzozlevb4
imKTluxcRv//JowHFVpaSUbjiS0BVALlBCM9ZTeQlBbIp0TjJGIGVYnduhMnqxn0/rzVmhOE4I/5
YCescew3echXpMPtdrTWa0DFaLv3sV4Zk1hGc+0DYJWQy9GZjvPRFt6mgN/8KuHFVUbv3ap0LzbC
/6CrfQK+ie9iUwcimkJMVW7r11rvEnWX7mTLrk60OEE4tAZCUyc6fUQ6pj1yQSh52ehKG7KAH1VT
xV37tHH42MYvWi1RXhYEajgGj/uf5bO7oXtqK8vWBue8Ms6s5+BAhh+/GuliKfqmMfr0MVMkdEfz
rZFiEoTLhPkAfddoiu+foAD2k4qL/aWE0NUIsClkPXbboP+E0WpSVesBxbqDCNQGoTGlanLUJEi4
i7AQ2dVMfvZNBFctm9Y2WLcDMrBrFHuLstd09Yw0qigKBgJR9cNPfAZKh2IDRe/20vXCa7MmJUiE
VEejJVUtdRIUUYroEO6Y5b9sOk+lzE+WAmWBySzXybX5db9T1qWyd5KLNfetw8gyKIcrHfnQZ4Bp
YA26Yh6cEnLAbaePUh19wLCg0DozzmucENsK9v7C2Jar0GC/Es96XslvnlgKnIZN12zTdMivjp7I
CHJrrVbLWajX/tjTTvDAfBZnJnSV3pOgFwwfo3dJ8Rb7vTyBN1llHa0y0y6KklNQ6qZJEGa9QKIw
EOW3qhzSuRJo40bQr+J9Wc09HR8yQmP22cUCQSo/HFYpfVGdAIZFktI8H9jdosZGvKXSgxYP9V7G
lIFmvEV39CsZxiNGffiGfTQxfCk3I8GF2V5zAulwB62ZujJ9zNo34mwN52KPxqy5dPI5NhKcyPCS
qQI05o3hJ+jKnwyjCZ89h5XaVWqRrjpXjr0W1NbOSva/3U55TUj0XOs+43kcwu6XX1XOt12laJfn
JgnSDz+1invirNc4kbojACUvgJJJE/i2DnTgnT+hc7hKWmBRqPLuzeVRXM3HsVdixtwjSF7gULdV
HpZz19NRDnW0ykkkpoDxInaHcHE5TEdb9ZnRyWs9YeTxwqN8q2OrHcSthoMQkJnQIxtkkF/MoZ5+
wCvIKYhMzAIbXBiooMirNvFt/KTTBtmQzBoxX5v3k15P3gqTbpUg1xEutebYlzNY+4HsybP4RKwa
iOgahuS5x37tRQplBMpBZCzKwVLU29LsTEypu0DRZmmJu/JeFvCEZ9SZQL19/qJzLCl4hnyguK1a
32VqtyhZD9WbCdnL1yb98jzdc8nWV6SSyrPUI0x8gADy866ZMlEOoIpGaivqjpv+cc21hiNmSBEg
dQ9xQ98CBMbnVWho0yaDybT/ldX33C7YvmPsO595yWO6mv8GwFZdIpTajioWPSV/MAte6ZOTE845
9sNcwgVtrFqxevJEB6hYERxKijQ/nuXstA2OdM8ff2cSr8ovmqjfbMav1/q1sP9I7HQKS/0CXwJg
pBBfslmRultJfv2dHBsU2tq7k6BckTYYL/Kf3QV/kLUl7q1hYk4FUChzQczVuhviOmF8hVOAL4QB
UKWr6FhiGoYXdiZ2hLLTFyK/tsi8tUp2VvGZBXsxZ33/DSC+6AmFXMkBkoZIkolWM2slV8QMrf7P
RXIR+/ymKLoo2R39XyLeguLy9YJdPdUcW2+45SMlunR2fHxi56P6/7E+x7dA8GxUQbBuYvuLWX/0
s7BVfTey8/6HJcO4/7FNaTowVBBnowjomjd9i1sGtjAP4wpaVjYzFANyV7pnkh51d4QCr/BJUuoP
QiitJSrreSDEt6OY0GDGFIEXQUDsrLSJFcLOiTAdlyipghaHI6BgZve3xb1MKxbT6NShg+vJjnFl
bgsY3MIVP/oeJFDZy3hbTw+wn1hYMbp1OyZig+kmjlNNJBDVZdJoqx1HqV2V3sYMMDL7AMDWLw1Q
6co80+O/Ezw5U49Md+oQveGuHbZmjhlscrtnDVMeU2ISB4cMKhYDyIZfv/WhTvwznLg+km5yief6
6mgneJgGHqC1mgqO/4TyTDlDH1Ax3Z5tJXaXdXLTW233CUggLbtBtEw3foaBZYhET+hd3A5ONgoR
O8jpV06xCbHvtBc5RV7YhegNOXkndvVPv+0A/hcRmaQRHx/dte/hRxISRzZ4eDhKqf4yGzsvad3l
l1lL5BJDlTnRHyLwbyp4BF+NKk4Oz6W6i2sJCiOhEd+kHDQI9ZlHzYNLjJbtAoIuHZd3D6/5eKJc
6qlgqnEd7V2o2GwpmbaK+HxmKiVVCTsQ+6Wf9sw8fGtEUcyJHu8LxU45/PAC6oEZGKvaWAxpp7JF
R4IFzGAgW2S5TF6dyYrHPGd2tL8VZd2gKm9oFNxrpQ312zlkXjmej9/y0nEi+4187FmLFPoNTLmc
X54B4CkKvKBMgqWIPNhJS/SeKhJkUzeTvBIjf727IKnj1SNoEb6VdSSlKUCmywd0ElyRaDkLU1Aa
5A0gl68xkzDK+lE+3uwSf9AKpK/K60rLzGNtnSMmRKZ+HakHIMph8rMiSJpXTsSFQzuYF9jKuIIV
Z/k8H281LpvjWjpgzhw3BPUlgZzh1wMSTFj0/c1jM4ANhY61wvjbJe13LOP2kJUnIqOPGcOt0zM7
QHSgNih5WzZxyulUm/UnlPwO2dzNZafcUQF39vNMU78Q48+u6EZflWpo6yyOkF80ZJK5mJ3halkT
GYTh0LNv2ZpyiPRr/vQ/5er2H+Sa+Z7/Hl5yHwQn6VtXOiAgvelHOpNnHuqnQFFovK50N/LJ/lRv
k7r68F1PTqKMc/o1TCnD1ajotJwKSCXUKzd+ngC7IXzbRqYM11olaZRXPx0Y9uHddp8CQe0p+aNH
nXNHE8ih9rAYMeylm1SKdmtW4G5H94J52FdxDOwksYqm9Wa3eNUK9+5rLYX/d396SDr3gVAY3dKA
QwVurIuzTVLyflxNca39WK4pu3DtEL46OcFFjjZUvW7DuM+s0kpAzJfaTzdydfbQJnYxobuCvPQD
sYYoKhBwsE1JotZMUOLx+Q4GXsFSaJaNBv2qKUSiFOXR+s+i/tFdk3K185Vk1F+qxHC4A/e8V6Ps
032OcH8LSB1FUSdsjqJV2C7xIKuNIJNBRsrO9ljREm4+wxGESDvpM2M6rMbA833LRaj+WcM13Lb0
emko48sUxaXLny/e6DCbIGcS1ibIsIU2zmHFrEmcYM2yB3Uq5TjWhk9VwbMGSW1nfsVtSZbhAI+U
PMgPb2197GOA0+uPCz96GYod915jEW//mCFOaG2D7kdtmgmSs+QrNRjxeS+HooIy0CcGoBQAk4Nf
HKEAs2ZzEw6po+g7eNmlXfrwprymYIqK4Ogms3qLn717yFpbu9qIU+814RutUHjGbnVPT4ur2ATH
3WiH9vFaJJe/GUUwmiD2/4Z3Sm5K3sva1MoggFh4aBCH8+8sOXdpkaTJHDL7eJ/SGs4xMG2egtvK
n65+aRrtvk5wpGBMNWVae/GOakJwr8wyXFt0f8Bwe4FjJcW4G680xjscJhJzhkmw7BuN23UIRxFx
wEsJcUnauLsaR7G8FsQnnE0kyuzm0obD1NCPm87jUhSXUDgJMXp68v8a/gkXozJQyfIqIvIHEfxT
yRVC6Msk2nzM1Ob0iHgBoP3EwPVgYufh7AYwJDlhZAnx0zbAhOA0vxYzvpsmJkZoquC4RuQcYenD
gZ2YxWzAa99ngA0UtvnnAjG9NfZ0VNAklkZGNK1ZXs1Oev7Vn8xqF97YPbVOmqOMRCrmj+AE9Qyk
m91KqwtkmHbAWvpSh8tPQ59HR8y6zFatjPXMpH5NaItDloDvBul6Zankj8YRArEMYmjLIWBDK+6O
R20rpKgkhSOGNemY4+xByYxUmv3n+FHF+xgcY210qE4jNGLPBZ8yweFGtnWHrHWiotE+cPle3JDu
g8NRKrEl1QkpG75qf4WDCdnzAamoUsgFwUrO9DQhwz/ele4VyQdtRKB4SeTOH3KYPxnxax/hCB7L
kiBaN2Hz5JqkHpN/ofJKcFIN8h7wqKMhCfVidLs+DhSwooJR6hJNWrrgXEytBHW7MnaBLDV4HE6L
TUok5txWJloKjL5zbjXBI+twrFAE6DGBDVjah7Dm4qcHgUAYbUuEdjmRNSst6jF+Kbrd6tCRf8IX
hhoIWAl5V+yD4DsQXgtAmtjRkf119RaRqYSju86kZZgju5ZkZCVhkRr+DUgyUC+JrtFMFP5zk7rK
m2XscRDqaDMSEYOID+eQi7gCb/OE8jka7XGpvC4i6F3jwjhPbTx1H9DQ6hOeP5cg+ENF7QItaj5e
KUAYezGkvA1MOV5sxfMb0gdSjkdHXDPndK/yYUTDtnSrtKdBi/HZi0y+55k4PurHGOMKTr+ZnUXY
xAG/KG3QHJWTbl1X6dphr/+Csc8XUESNapVFpdWL49OuUbpzp9VZ2sbfEjX4Za+y6nnw7YnGCFS4
Aj/szpGyy9kY7WKFcmDPyEaUCZpOcNFOIV1fHrOdu/ZTVhD5nMtE0dKqkmOxN6/OWcRJNZ6L9krX
bx1mCKW7BVUc9EeuUXjVKTM5oPZMVPdCBgNHKOO1QW6hMbNsUF1ELdOGMRW1PJ7xMbrjAykp5zMe
4mH+q8T/1DCwQtPP3qghtHNBesI2OthYnvG8FvGOEZiENLtd7TPqyh92bioGCmlVJmbs+q9r7QZQ
PuiKZ69bv324PbseRthZXLiAvlMFhg4ht3DNmUa5KMXoOlufbgnbyMtQd5VVw2i0YbTU6s+tX9xB
hz8STqpqj2CHgcueXCt+SAHWI/6ymMLIjZxN8sYKmXA5TU4mzBjw8Tb7fx6qAcImd7+xw14njq6e
9vE1qfkePk1KCNDpsi7ZoszjQGNdedo5LlKnzhhJqV7bxagkqdiR6GJxgFvvQAJcuTOlnOqkG/FN
2MjLQ4ka25+V+t7dPK15Y+0BfPivp4JY7to9gKnV+Rm9IRD6JtRt+BoRduXzKrEqWpGl+xyUQ1gG
R2qCMabPimAjkYtbzBRJ9IhTCN6Y6HXtHuYUyM92qHYKI/A1rCXvge27LppbE229BBMtKNiYOXyp
0lyp+eXvtfa3hpa8Zd+2kJUbXyjwQJ3VPqyC20sZFzFYZWCjcjSqQBr81gV9t+qwdwOKm23zzF2q
rRTqi6jz5PsAeufXg/VuCOTq7uh4YAsYlquL4cKlczyxW/pa34X8lt65PXYHZovByiwb82OuEshu
DMFskSaA2wvFSgig7YbG/xu0JA+FIxnK23DKc7WkvkbEqAvx9c5HMzCir/aJKT26/uLdNJV2H8eR
thZWtIAoOuv7mcYww/MtGdkqKxI5wHK7v1LZdhPQ02t5yQTiVVGBjcnmmiK967MJoeWpeaC9EWY+
uhFvICtyNGxrAb6EJTCiGAHVurXnTn0KIHhJbbnIT7VlaCS1k2fRHMmPGFM8xAISxXxKYMbeChQM
KIGet28jbT/5k9hn1Ib8Aq6RcmLSk7TmHzulpsRHjr8DAx+1Semogwdjm1XSge9toJt0O2cGa3E9
ObL7PYh6USkjeqs2sYpkim9kPXuFH/IN8W94x+nagvYLKlZZ1fTSMqhOjG3mxMKDpFFd/Ajjc5DT
JR23Gm+aK5EJVJsBCrXG08zofJ0oRNJ38AFKw/X0WX74f47MrxTbnsLeNGBUg6YP2n/PAd1zOlJq
T2TUc5kgk3Q+Ih6F7YZPNOPcuYObMpieC2Wbirdy/zadfvAHeaqy/swFUptc5sl6Xue06LIRhWx6
V6002ZtO5GXkNvHlkZYr13AbXcJB3hEiNsK8ZRKlxvyos8TbL/PsgCFMs4z/q9Rtc6on+kYfBbHx
yBi4kAcKIN9yrhDP3o0VG3xwngp6iQgkZ9JNL1/mH5wonX6L7D4n2eCLcFYlAOCM93yi8LzKhuY0
4jTbr/mwh86B0SDeVUH+lsdzJgtI7Zcp9fZModlzSKs6xTtjAhnghUa09xrZUYuL4AGwbl19AfGi
5RrOHxWBZTG/yeqX0ygDHnBuSAH9ZGOrtHldoi+Mwu2WDQM2ouiUpBqYupGPCXwjsOUw7+41MSbT
uUGxH3pe2IPFRVqAPxRLGF6O8WLshkeAxhApeXMdrhL86OEeCvnyzEwiwA5FKL/4CmrWWyIlIhfi
OMPNnD8o/aU/9qCW1o4JQOSeskZ2Ox8SaYEtatOhEwZ1lzkO3mBjzEF1ZEcaDkYnpErzHzmglSYS
AVsqvVgdINLb5JmS4e+L/frt/+DfJZY6VKPUJRq/umroBU2bZLUEUXIwdNa+LxqOAyozBQxPTIXr
z1KalxLLhFSc6HFL6SrXx0vlY+4IU9vZ2v6YL5t0EGZjji7AGryZAUqgXmZLz7j1CxhLfKJsucQX
GWp/zQRjtMBWeR8nqPCPv7WKOJLSvehfO8ONalRXbVAqXaNN9agJs6i6/XDuwRcRSRQpiE2bY5xn
0ezarFZxCOKrMr0LEN69NsyBUM3w4nVMuxQe7nSbygHvz2INPJUB6xjpwdk1TFnsaVAlnt/N+Fzw
81of1H4YOrn6UnlGZAEwJYHvm2jP2z8CzMbCU/b11aqjQwRg2LhncGl6HZ3eQ8ebq9Jydw+vQ0s6
5vtsIAEYN71bYaH/fcPsXjgBe9gukyaLBrr1SSPtb8RuVvOYOyWgiHCAniAZsy/6cznRH5hY93Kp
dJibBWSs75hCsGnWz0A3/sdJhy88eOcQoJ2lxsiSA13iAuRBPH5sTRyMvh4HgIAFneD7zeKIsSHg
dh9xkphOsPndoABkYCJfQqkXxmGAeB3qN02u5emguMNMg6JJcoekE+XkBQovT2ySYLVMO4KhqcZK
LEOwO3mJzO5sp1CcP4N9bSMhheguBpjYTGJ9y7JBUL3y+vdhLpRtvfPb8/D81kCh1QBH1CWSDOGy
TsX+Y7WFCaYzc5mKq8BhwzTOgtHM3loiCXCV8SyBzSVbmXNaJYVl0rWpavQV8IzA0Ee/yRqcumA3
qiTacKyonA4oj3eTs6hUtGRGg8eSMIP0iHl2ILR/f4qgO6Dg/pSJDo3YvNK1YsLj/nmGE7zF0Tl8
v7C4I94j4sLSF7BKmIT3cIPQIVAIV72YtAwY7/cUPU2ASv5pLq7uuQq2DqQYDm9di8tR1ZhpGI55
M7Jvf70lL1FjPP+ACKeimuTbU5Oal4Pu9D1yA243oYmAZv40vzYH0K/qyILLlX+5GC19D4b5JKNK
R/hPZPBUa6kYCrU5JYsyXCRklF9hIXinB0mSPMupG52pLhOzyu1Irv1jna9eOaEWHmwzDY/5jfkU
Mwn1+CgOPCU0GAfwxMmbDJgbMuehOsDIJq50C4jTjGMen0afun4S85iDvzkZ+4PryaM7v1wyHZF5
PeBD/uPnLiFy21rza5An6RdKerphrKfUwmbLTZh28VvesRTIfKCwE5AFuoqSexKBGdJIWFUPC+XZ
UTSI3Rj59TDo/IrtguDAh/LDP2Gix+5W7IGebO/fhwaRbzsWchwjsRm6+Mdxd0cpG9yBQWZjilcr
Z/bYEpiChYpc7bB0omarMVUnP18Y/BdEBtRRiFAxNdibg5i2tf6atb2ePB/c3AAF49beiNJq2uu5
JCa52sXl+UqnDGj5DgfylheK5iCX0KGodsIItJbY8QcImMOagHIuodk5tSUK4kpnIfpQw+u/UDw7
t9btQM6MqCEUen7Rn/0nQkI6rKvz/OJ3ryJHfJypa3uPY2lHWD7hob73mcucjhhYF3TSUX8oBM2U
fnMY1KXoCp3olkiQ+XndJscT/VPd0+URd9HqImka4KQ//qVK7ABJ5c6iHJm8zpKX0GrCNeiiJwGR
os2EzZUonL7o6x8h9nmesGw3+inu9aNjvRh0SCzohmGLcD8JW3nJSz+bk17PpcgESXpn8u4/N4FI
VgKTPgOyXQ5STxplFiLE4sQqmvZkHmZDRgJXnRiEFrVyvfiia/7kMNnhNGcTfUo+XoFsaqFZbdtE
eEEkY6MCru9EFHrs+MoK2mHeGCfNGbcs8KulVSXcajVOoFM3IwV5Dumc1WanBuFQwOObyOwi1Wms
Gv/PTcFU0UP/sgAbO1pfH88I5B+CL2nHXSnN6tq4fHhigc6/geCFwpkJo5wHIw2KvAlFBCmieBqv
vGIJteVbo8NvWIJ4GLKHtELvC4LQdvhoa/mFfS3N0n4Je5pFSvtfXzwhFXz5Azjjl3gWaOU/lUox
hd2TQx7FgCa5Y+8JOXB9mSMs4MqMok+RRKmT41PcrU9qGRPeyed83lwXmze/tasBuf4HHMqfMPvH
DnBBjiefZb/Vj16uf34ADeiBFujpEGSM5itxGfNmhV3HDE/CkV4nZwozdQqzbkU1de6lqADccxP/
GyYLHty2hmWt+x1+2eN4Dn9neVBMZ4IqZ9NV1cbuh/3riDSvXMRcrMkkaBUqq5/LenT6LhJxbven
h0y0ENC7+hhpywoGep3Dgy5Mzq8HQ4QMB7+sZbyhroWtLtDjisVETS/ftLR9/KoUoXuZ8qX4fX5R
GZo0A0kGu04Kw41NSgkSxFt/LTGWvlaYjzbFfY0FBDWLvLvYrAAI6jrcoZ5/NY7L36jwbHd/0srO
2kS8TELyzlBg/IwjyxV+DBXMFLhc0iSV21UkHeZ05Ys5xNxT/X/fJG8MBmKHpW10IjldtftnUNfF
N/c5IM53/3I6WAexR10h4DKwkKLCIOauEFtTmWpqQiBKjc2l0M1jeSatfjbBhl/MrLoWif+d9Pp5
VZ0HadeEyineLGwuYBSQokPIXKodFDgE+snU4PSGdcn5MKP92QC/V/zPeekvJYwGB0zkS0UwaUjH
hGHryzW1VFfo7k0mT3nUd4ssNlBjfVA95lpy26MAahWN7Wg5Sy2Qv9Aiqf0ujng4nWcP0goaY5Hd
d03zQiDk45tRdEFKuhDSdQQ5UL2T3xxWTfSpTI5ZOuM2ShwzJz+4FCXbazDkni/kxBK+XsMiCtek
d+z4Uqth8uTFDnomZUwmDCJ4mZiO4U+7ZTi/5lI+Zn6hBo1mheXiGrO1sUBZFbe0R+5/bZw3DY0+
EvZ5MkwV+fMW8ygzvSsvSMco7UizkhHyFjJIhiPrRxTR8ucXw+FVR0ABv0H3rKNaZ10p0+shbnfX
36rWz4vWZLu/QRj1PUP0pz231IOTrmam5YDlfW9rrLBDyD/iLOy+XTVOa07JwEqa9r2anlTqwNnv
knKe0c21sxEUgT241sVKgLOk2M/41kk5JfLzUMS58IjOEgIcGQSYWU1zpAMBfBY9wA4vhiBkFoFr
FcQqtuIktn1zIQs6XRFXfmYtX51zQNXbhyuRFD2XXv7y2tBcMMKfMMotNDntqpyW846+KGShYeWa
iI5cARgZIJFgVh6VC8qWaIiN0i4uJZJP7uA+xHnuT32izhAN7fTOOCw3w9AU1cSmp9hG2aJxNzTp
eFA+XglefPVturjSRj/kFBLNsSbPtlE+XnDhG4eLNou9O4m+oNc6BK12QgEEFLC9PEDEMaLaglvc
7/3FF03B+3HgDAr7Y1c5pnaZSvN4FbWBQ6WByAGtokvg8PhuKpgyiYrgNBjPWgMNnFUjjOrG11V1
XSCyqhdOy/pzzYIaQEiJyuIpd/bOBHUqfKlnO+yGekFOYGQvfGvmXQ/GeWT0enAbEN7o+Zf27rRe
YImTCzqAFpduLJvdh+QvxtX2341tZ2iz8S/pAp33U/zaVtBSYFjswuy9EP5JmS8W8oHYLIRzLb9P
DXcHRJxTK9fZSnB88jny0Ngp6AWQXoRIRHUvQeNOEM5mRJEo3X8wAjk2Jqy7P/DEdehsSqBeJhDl
3eC4IkJTKcuBgKcArRvGQRMTr+5B+NAX01qU+7oCVbA+hcP7JlvmyNb5ZCykyE3OGajDOB5+mz6R
2bCSTt2QgVyWSzivchXpIqp6aqlq8zlotRxvdfzFfWrv2dlMd3DEz+iUsru9W8ushcGymg88LiHE
5mYnBXENwrVTZqzF3ZffGI59k1Q2kEIYkW9JKLBtIB4iaFYdCneoW3CrRcmzoOTrup8/zpOIPWkY
nk4EuuX8TRVg7VWEra0141tojvr6RKVws3UoPbNvzXngBMNI8qna8InGxPy1CnPheaZ4xdkNxjtA
EQhPhlq+ICRkJwM9PkqaME4i+v7JdfGsrSrYyrodjcZK6rTYpx4Fc1EI90r0cIQ7WY1AkCkf3AF6
5udRNrS5VN3d5A17ccznFVTiiC09+QebKfltZdEW5G7wIvau2C4ycKWBZpt9aZ0NaKWSnBmoeXQh
fzMsHloV7Yv8jo4MmlyPVSIb7hE1RBNOW7xw8yEgjc2PZYXs0yDV3lxOl2T6X7LAPfiTy1DRdZL/
n8dEjwIh8s7pOzA33NehLgMwmvLf1CehIV3bhL1wUwQu2W/e4bj+4YABHlHoKwIu6Y7XrUiywyvk
B1DHSGnR7/4oZMoB5x2BuQxhm3hdDsUZxewVj40chBfySvfW2BWCLt5Q4MFTbAf0sW0oYoxzdmfl
SFYs+LFO8La02xt86aamfuqBoCYBk/uHK2ejzCmXqeYTrEHvmEFldX9X35EX/sE4yXD86TxbKRqY
SnN1Nxfm1no0SQjqFMMdcVi0hsdZrfPy6BfKqu3TWVjvg6RkERDc/0kxCEeIqhWz9mMnlgrPE8Jr
hMdaXTnED321QCo/PWNr4KNktrKj2nnz55zt5N8SfAo45d3TDx4OcTp3Vo9ZYUg+u7exK6a0k2iV
wGfrl+OjGyfuWGmrV7iWi/jzR/MB0NlFVXXa4Vwk6N6L04ZRzaZHL8Q5uVDh0HuTAqc7usWi1L5y
CBHXWh/yae/1C74w0lEVOMulTG61YAwU+2dAthH59AWSQRKf/NcC9QfVpOBVkfKKdE9Q8JqDWZWM
/3zoi9qqAmEuRtaTMwvqLl80PWrKtrP/LDOX2pYOm7Qp+E43/hWdb9BvgQ3f8VZoQFAAw1SEYmRD
nRaFcWnT83hpoU6Ys1PZH5ECXsimpcJ3ueYbJw4W1PyLWwpRvittD/C2MPdH2MsVU1AXIy8HVrj1
OcD6zUsbCZ9Wg5omEI4Ez6xrHeIU8N+HXjkIftqWoocFVkUxUK6WXGynU+4uxqquUUmBCQe3GGbf
SPsS2xGBbacjMhw1o1/Th+Fsc273qRAHRYtoYeB9p/ngt+M8OSrmFcMvh9YP4y4pYypwJ209V+kQ
Y7hiKVNyQPBaFGpz9cbA7drhIvIs4JGjQa0126SFKIL6ysZ8hWAXI5Mka+7xN+L/BzNTJ6YnS/SI
EhkoUexF5KnNZc05Ti9SdGWgAXSkZvfWj7wHoBdFZnaoNzZkgsC+jjdl1I5vJfXNmE0jNigYE48L
mYtsmNriPwb8N5ftKtdJvXUBzVFjGQJzoqmRAl5ApLdjcWXNwL1WYT6vUjV47MoXf1BMkJ/0kCB1
W+QuXcyvtjSEq1/kOInY6CeuF7NNUtRc6ztH6qGfSufZpJrfZLoc+2sHNq+cYKHY6TopHQY1EFyb
ciYF/xyuGTqJvTKctLR2qzIHYok5HWbO90GG/cQEbyk50YXwjDqxnjAVxNU5bZ0hEbZfz//lZWMm
kZGqn4EGWT8LGrBJPvQMeL/9eeOBYCuyUmAJYm7BLRoEIBVsKSSuBA/A42Noj8PmLeGWJ1adMBWL
aY4hKWIdrxwYfXTu8FWXxwUQhg==
`protect end_protected
