-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
L805OZ68oywL9JVXLeLfIN6E4N1LmqjGhlhABn3l/p1Uzx4n5jhQpehYMxQ3PGZZsXxjjuIcQqC8
QNlHVIdZM5WLvO5qYch+Y/D1AHBybE2EeUzDm5bxai8aJLq5eTBCkCmEsjvCH1jBVYYuAXp33ykh
spawFzfF5u3LqCGl7Kq8KUSdA7cgovRx3KjahZH6xFw35g6j0pZw/v0suIuLr7+co5rAbdCwNvPo
MDk0g0lOjvIJl969FA/RgMFbkGCW6StQy9f1kvf/4I7cf95Wt/WYzJrIwno7yERjAVXeHZYQKTdr
1nJU6MkcsrYQ+Llwe4Cw2RISXdbuBgdWJEe6Eg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20560)
`protect data_block
DgoHMpnRnqpfWJXEAGl85dy8wQFyWDGzjOZE3CZJN280mu5tLbs0wzkVvuHmiLqxyffqZG1+KJKn
8qFJZNKRBKXPip7DqnqRqVc0uxO0iG05S52WRGj0i+R21VTxT1ozuet7vrzhEN6ZEWedSGl+8dHN
pOwvtepoxE5GIV8gFNkn6YAaZ8Hx5pNHBVhhhDOq5lXaz/5vq1pdUm7q49bRFsv7nDd+zulyEXrU
gFnUiAOng3wx/2jyEcxQgVtP2blcIKpQo0i+eko12dFs7+na9PKhp/KB1D1Oq007+ivR5/fbea1Y
oMv8NUSkNuXlHCIsSBWkb3cSiyuJvCabKH9fcCX0ZfM0qy/aFcuEqzV+BgeLotiphfSjhmdDKxWv
2dAD3C8Qn6XVV/kEVdjtLYnPA+cWD+8aZV0Huum+1GT3HXYE/h6bloxWxz5E8vkFRtxi9wNIKVZt
2Bq73vyzDk9wTohTnQJ1NbhGagyoEYnx66ZI3hcppnltTUmYEy7XE/x7nc7O0fFz2xBalkkkXiju
0XoA92kuIBwP+Dkp63phFBJPvMaqjsFew4MRs7jKkzuKUTESoBRqeUSh6uEsbrKSAxAoq3YKFD3M
R0vOPFPwUCfPSSaLvg5CFYC2spHDLLNq3pttp2fHVOAoAcLdppnCfoEkvn+rJiac0oqjBYNEM1T/
w+tyRPN+dH3N/EjwWe2caUpYls741TEHFvZLLgNEif5Y0x8+BKHcDd4aNHV5wesBCB3+49iICV4Y
uJGgrXlmmYxvEmkeSw+xXl3vmD8RnwKNi3vPXBsW6cIbYm7sDJIfPZ1hP552a0d+OVAly7MLUFOn
fLNsLQn9sTz86kaGwwPyvQjjuYTm71DQXjDUrX+/LHsGzVRazkmk5WvBGfjAsZ8ZGdvh2hk/5TiP
AGjY1TA/5PeFQiuvntC6t3aEfnZKSigGXuIeG/5nFKP0dTZFgpNWMhzMeyTQEybXGhZ6mOe9SNL+
n/kuRflNPXwZFZX2zYTMz9K0lUgX16x7jMV7j+LRBigB8JPsWcPI358sHMaq8JSg0qdu20SkskNv
BT9lLWd1yE7LniyeCKNVtYtiEp48o0mVI4lm1+gGY5hFulD4QcKD2oQXPYhMJJfhnBnRibQ82H1k
8k+7DwOqOwnOYVKJSJZGmpR27+xtw0YqAN6HDNdE88QlKPup64e+4R/qHtFYRnnTE/bf5J7DVKm6
lJv2E4302JxXEGArDvJ+ZY6XfmnpbJxYN19ZyYWkzCk/kwRYqthqr4TxlrtRkP3lzdwajA8+/oa3
zo1Bxttt/2hpDX5j7oizXNRaYMAcvgRZkQIR56DNgUeaS6Ugw2WeKByCSEdEbljXqV/xHEKUiTEl
sTqU+P1mjf2XAr7AU3pufCyIJgISGhot3qetviRIDMOAzfuVHa8oeSr583gnjPOr44OAs2b3Y951
3zsMHWkqmg6KG/4MEHkEYuzxARTvuUZ21Eup0ZjAg+l1R1TgAwD+dszeI81IsmrrOrPzVmKFVxDS
kBV9hgQawDSmio/oGjQwFnScnwvnFc5GE7DUUmTZIvhi2H2XdF0hpQs2dw+GKR8VadjnJFzfdVB1
LcL9UXEXb3GBvEzmRIozG4Ju2WvNrs7FaRiVDZxbdzEfOChts7BZV2Vin820IbzZqGBx9eIXYrlY
dPYK2hoZ3dMhPty89EAQ21p5dP9f0VzvkehPSV/rQkmjAW2ecdEXC5ebB5AfNiMnjL5MV4TT9IcT
U4nuSO7u0O2niH7S0zXE1SuDcujb6Dd1Jv8kKBB7unHJ1TRSyHP4njw6cIZDokERO5Cen+95mMTX
3krxRRbqMk81eDbk6ljWwozXFNxFvAwtAOHe8pg2b984mzFffHVKVAdKBMrc3a1fKz0L1dS/7zhd
xaTd806/ilMjb3U++k69x85ta5sF3Iul4kB8Im45Llbe2So9/szWcCYwrsYOa5waA7W9WVGlsQ7K
vvZrf4qySWpZ6fuNJCsbEbl+KQP/kYgyswRuH1yjnZ5G/u2LmhyxShJvffXZc4n1PVNYmrUEq3bM
F38sUlvO/barM4ur8E/nBRYlUd0Ya+ZPzMfjESOucKWIjESW7dgeZAkjo8MoWwaKL3zgumGFW1kQ
TxIcYhXfjuaZRb3npLf7Kq07EzAgT1POSqaZb8jE/fgvTtkiL16LCGtJSDrFkq6UH0EIRmtsOnrU
SoYSlaC5q7JySraF4zNlArDUvkBNLb4LaQzgQ0o205d7OqiFrYxrP7rJDxmY5SAulBqxdPXfj2+1
TQ5tSAduuLDUMe/Qv079euukAQYDMQIoZyVs8xQ+n8j7S2RG+/iy2fm4cpJyYzqyYb3uepxKhZHw
VMg122oKIsn24H56P0NaAtg9L3U+J4Gw4Va0yDxLblw/QXptfcgVMs0MufdU/mSwvnuVaOOnjpnw
ytl4CL0gTCz5da3BiDcVoKe5qdT3sabnqMbs+eOUhTs1Miwb+Ha50WoD0QUofVWcNa385m4w8RpS
fmxdRdrYHmSVNq5M2AA5lqeeuaUSGzEzBs1d9oRPtmdfF0d5QLfom4yOiMSKiDnO1fOHnFM9ChQ5
j2sdVlJiwhG4MPu4CSPJ2+9hVRjdAEaYHxKML9QF2JcgRQVXSgGWnkz2MMR0Q4EFuZeLIde3qlxV
ycU0mn7f9F5rritdgCxt1PJjW1c/YglFjkmj1PK5PSwocYzKDpBDmINYV40k/krKi36mzksCrIET
/yfZChq0k01FE3ayEgPIrm+DuHB3pvLFcixFg8EB5aTXdPsdMEgTuVXY0Dyt4stERKR0yB84PMKJ
mCQxjQ55fSMB91lAA9W+ykSuaBI0/CJb7/hfHvQCiySxjypv+tT+xAKCcJjXUobJQSfhS00xvMww
RINn0GX/fS/2KSD1KkpqUXkc0p+xXLNzPrjRsfW/brOupwopRGxLoFl7qn4eY9W3q/l7+MZEmYyc
q+Lj2Ikn2l76YzHirituUWDs6jPZgdl/cev0LWg5hbxZ0ggkY/wgzgYtoO35CUYJDnNzWeoH4gWc
lwo2vXP6gAKAA4yN2cPI9vtY8Z2XVwvC05O7HHyX8XJAfgwXckdxZqmMXxd+2oqj8eg9L2SO4qaP
rag+ETiuMG8g81o9J/iQ0wX1O0/zEX4zrYdnR/Hkg+bdYAVKQvojqVrVS83X+Bl5vbZDsrpon4Up
ac7OOY/tRQfJi1MqMLWpH8tCLKVT60KzPAW4xJJ94FsOzjPmpvBTqQ2SQaWlnW8HNCcXwmHfLoIS
7MTNHC1dM6LyC1ZakPnVdbuk5UG7dv+3g5G8VEGhSC/bgzhLFeUD/bgVD8lrgtgumnpTFCa82uSg
G1raZhPOO7uSCMA1XT5iPT6TYE46AE02cIvi64zPgbos8rtd+UiH2H8FSJbJ35vnCPBorXiuNd7f
UD0otABe/vHjBfk4mUg25fOhZdxNx8MrShzD2QPKQ36C62IArnDovcXmtJJrCwDRRCuTl3qnBLw8
mBV/eY1vDORPLSylc9LVc8rBl9RoKd5fHisThgCtRtqmagC8n63TH7tQZQ0KmdsSxb3ZUQILTJGJ
KZUNLPqT05h9/rOEj5HZOxZinE3G1Ff044sBK/525vJFVttlLoc8ey5DYWqXxxaVWn13wwVgdx+8
nkHFydihftVbGtv/yxAVQLAeQM2Bxl8XkbReuTinvam/lc7CCwsG9nwfE084pafM+NeIyCkhhN4+
yhV7CKEBCpTBnGXv1sZoiy3VJso7dufmLiyrMc73oGRDzWZihqWXnbIevCjg4CA1cn5UaKgtc+Bu
z5xdyMMCejK8mKr+OLtHQB8axU2zjL3ArgUjIhHJS9OKKA/RSWaO6SB+D3gqnava7CENTdw0w+Lu
AxCG23GRYPfyTqVIOMgQouxJ5fhBdCA4frmEbMenlet0xBEolLap0fDS9bDKotQbbHlTV2ygL7tz
JkqE9pz/w81NTuCfyUGXuB3t1l3e8aO08Y5RKfbtRxIT58cmYnvbB3Pcjurrvu/gTcvrlUrJDbz1
gTDbqV6460y3o4CSVIaYg7n3QA1botGNVYkvGbeESlMotPHsgcm2e1XXiogVQoVY8cWPtKjxU8/0
i88GNQEUawXL+kLC+zN8yjFIbeJPt4cLBjHa7UKbRWD5f7AgfEj8uTyrmqPUAX2LOTY1df0e3iZt
kUpNsc4qbopBE+hs20RFNFTiqs8DYf8qVMz2zOk8CKhc+Fyzsziu1bgI8HwIh0S4tMwxLQ1HJCiU
9+gGeaah4HSlru1i+5WPKuITfNTlEJhC2XpZgH3KetJmy2T0eb5AyX5PRMnsWvCcnm0gU4nHf0U9
vAEw1bqykquvL/+mxrw4OWIduaWsjnp7gLQaMtTcsUtBpxcj8CVmgW1+uAXDPSoMoBvE6+w3wYMM
0jHv6gNFag4PWorh1jXaF3324cLp/+KLxEna9G4th+/IFWP2dJO7tjuSmfUuKAqVjB0nwzASfSEL
EWBBVl2/jAqnuGSXQ49EMRC8nOwQMkVFUctKTMc9mZ2sdF7mdul8SyidnjwkBh8xWtEQw9NInLmc
PSQrvqfSftefulkkKtZ/96GwpCpxvtOaMWtr0hZ8eMZOQ1rC1hbvu+Tp01SZHRXu7mr9MKbc2bhN
haCfBe/Q5Lo1SKIcUGbOo//VUd5V6XG2opzxrNGv22sztniDUs0iDzVNfQ01h1WiJcJY4r/kai2k
jPv8iUfSNDg3q1ec0YDcY6+EdjTPu6cJYdDuFzzUuuH7ignsB0Gtduq8RsaPcmkJ971S+zzXrXUR
L6HelsLoolyOBag4gaX3j1An/Bw8oxMUonqqAZXIwssbD4rYT/xYj4vJMqp1+62CyOblPxRCjBkF
dGlLPsjlHYa51FcuNR35t3q7aIYa4ilCMQTcUgvhJEsWm8Myn/qr0oY1bceORJxwHGa+46JhXSCD
1AL58U7ILCaqKHLyfzvl7a5bHLMnotE6qa6JHjrzNlnN7N78mqtFtqNP0dVZALHdk8kBLbyv9V+k
A416C3MOvQNefDaDJKKx+/8Fkot9cLY53KAIm3dO73jKhdbYwpp+VQepqvbr3v0aHdxcRwYF06pL
ZbQ1PiSOaqpyvK+Y/GWYzUiTC7ZSnugkESkZFCYvjcWe05l3O23SCzZV7u1qLdiFsT9l+tNvBv9D
4w+cixUFVcfj78gYJrQat+10jwfro3U4Lv6+AsVyraivL27MbonnT7cZExU6gTfjntDQn0AhUBOz
vd3WN3okHmvFLhbPDH71h2GWz3TfTBciWihLiI5GjA9QFSvxXjj8478K+ClyAjhh9wZRz1xoW98r
tfbqHUa0FiytpcCo7MtfIW3KncLCWekJA/OVEZgLgPoVWhvOwEsUw3Kie/9NZj0yhK1wbSNIkEYm
6uimLG2H0BQOkxRfgITSinZPOxmMTRJ3BQijUQpdcoNpHAb4vPH2i5notTWiQPJUZgT/GW2qch3S
RtFXIH1zNj9bNAr179h1RVWzms8JHkzvlRltyMouGK71o1RnYQ9CZ2mzWEUbOJgrbaF0OgZHh7T6
Rw2ud1tQ9TDWUagM2/z5iafkrALTykC6qcua8IaYB0++CLdzzS8ILMr5FXbkOScyEBDfLoKwVWWk
n4eXKd8VN6MoQJDDzv/Y7Ua+nuv8twjRL+mAlaZ0YuZM9NRtx5iq7juiQBLNIBviY/ZnQOnb7ST7
Jia47dMsKZDhpPmuDcijYhKzPpVpODCVODPBz8vi84tN3I+CkaqUy1IHufzWhWUw5f4UP8okir9L
c26Q+e3NGcyAtS0R7t9YNTgjqAb3PpuEh2JkRPrxNMLNjlVMuVB96OzJkQvEbs8T8IDSD6kfIB7N
JWqazkpx1N/vETzT5DNU5KDa+pNNRVvL8Uw0gzD56u9IArwbqGjsu0KPYQEVGCu96nMlERSbicKO
jfbKTBjk2DbpO6p4Cb4qYr+ZtGNAPqY+WkD39do4ZCQdwzpy71GOF+fEj7h0vQTVwL+8XOf52LM9
0eZXJvZfQOO3basafgfNkp/yW5N6A9vgB21RmC1RRsoY8iHAGSChdfDQZHL17ngV0BPbIXOJ0JNx
MW1VJ8uWD6d95SsTjMKsbrTBULl5fbUrG0tUVMiYTX05EF6rpMoyudCU5+BHYgtDK/ZiIWh7/hEf
flqOrBy4/LK+LCF5KXriKn4weXlC0fspoKaFELOlhstu8KtGNbY0byV6HdP+vusN38VQs2eJk3Zy
2wGpDpVn+FoClo+Mluqsh8vFb02GxBKNrXuztLBGiLAh5E+FgPF/32VWk93Lv1AP+xAOvFYJj5x5
bWWsMUpA7P6Y42QtgOwVSsDu0RnBDBCeO3oJshEwN5nCG4fMvygCSIHyUeSC4jg3SoUQ9gCWCNeQ
hTGacaxlb4rxF9wu5sdBFJI2kDcL4Qmpv52btgDO4KiykHCEV8U5KG/kcxSlIL3EY8jo5Va/frLm
MisFF4vxt7TcIlz8W5+kQy/jGYOTNvFPoeGRlU0fP8lEnJVssy+zqtTpGbTBKC/WT9pe+y2c2gJT
XELDJVPzcXHIKja7kxioi28ORIsQ6vv4QYCENZnw59c2r/wmJ9BW/eZ41IiuICaX21kv4Wqt/9Hp
94XrJUE7RZCD55z/3mY0Xl2BFhn0BdqqemGNuYQsGd/ewMqU4YIuNwfhqSG8zujslT9VbMyZHUaq
FYIlO0O3K3tBrZw3amoGvJzGfhkH3qkDSB7UNhCvbZHk86f1CGtLtHtdUU9THseBJwQEFarmVp2j
NXK44RKjrXf20AQXbE6vlOhydL8eRPPgF09qvomayCO0/6v2oRvESTrC6gmuveSk9/ZCoNkyTbpg
Itq6VFNyXYgahKmK/ZiFqn7PfMYwE/ya8NvosUYEr8UxsbCQY7HVbqmtHFoClmYOCYE2Mylrjx+1
sm3Dq7YQIE5vQsVdskUIRtHhiqHvTJDpL3G9waBiX2IH+40BD/IgglJQmy241RpdiRP77IHliIvA
0zLXfj7+E1w54+WcR0gwNlhw0EVJxEXfhHm/7/76rnIWwyZXRJlE5xkNZEEX3GWLXmOr9CMY/fgx
MLE41sQEqSJ+0rJRaRBQFtFDJWrHvYE31GYbtSp6T3IEHxTGWSiXqlPnh2SPTAMWSI7OJw+SLcYL
YTvaveCZDq2bKun2/vcsybzQt+CDZOHO/wFyNg6Kj8X/+MqITWdJjNE93K+vOS/ae+Nm5vyxHIX1
7bE1XbiKaxSvNE4roIoKq4DkwPPFLRta8uwCcVi8cl3YYgnSq/n434SP9kE0ZRpvm0c16TpscWhR
0A5L5RM1KwvkcTVgeGS+rPs8mhskWvjc7q5b0zVQYAQYQ+/SM0lUmqH4K2BBf/WcOHrOEavGYq0e
aOOZyY6nPRDoW5eqwLfYV4tJmgQl0GBFPrYhMMcag8j61WfPuoNlRJEPXIWpZzeFHPPKru497Bol
TmVn89njrN7FoCHfe5bVn7FeNUCwnqu+qgboTGEG0iK8lyR2kcgrg3E+ku8RRWgYmkulYgqv+7wl
cO9rkcvJmEcENmXgXV+FcjTNtTurzXiT5jEHwPrVG6VuYJItebuJjhSOwf7Ink8UFfMr9SouJx3R
998oIMrHHYMVHUQUAL15pFJcSdlPeKvkMMFgvTisKwZWWIHjuBtQSYtKmEGIrktfbE7IZgYre3iX
gwkxxIRukVCOya2grYBfwe/14u1DMsff9XJl2Qj6KWQzU4di7ha09ET9ssYFO5KV59U6okdE9Agf
B0o9XDwnxpQcDUmBx1lrWh+0rjn2DjV21cvzIwHknLY67G6c9h5cSyi01ixwR0QhC6fEcMFdgsi+
+AdBf3pX2wfpi8W3/OQz6hI4WWChqxtTM9HYPk+QHZ+p8R3YzrOVKMje98gUvVaQnYinf1tPWRRl
J2WfGa2dFNkOQLyKG8IkutJ9BQNAJU7dywekcAS2mJDgXl8b8YiAGe6wGAFaKBWOr5Gcj3vGO5ci
ilCEyn8PJ9YLImlA2fFtbMhmG2bOYW473Pckep1/I/acKQ/LHFlLBvgpnZtKykKKrxaPV6hEK1Y3
zWQCwHdbiFgQwrWifMWizJMdzjWSMcKTMSczmS8z0etHxt7aC4JteTzCOF2Aat/VRU93JPOf8KXb
hvsGU8aD0HnS/FDBnUDFddEQVOrhyUNCTTdjUgME8kx6pKJ3LWq3Ue284DLdRX45LxIC1Hjgv1IX
K+kAwmhGaD5e5jrMFI/WkxGE9ndJ0ZoHliZ0zJLw2SH0BOuFDtFmtrYQ+n2V0Hjy7qxmBYA0wdx/
RX9Ji8/vfnHPIlLBWgTRlZB/BipbpWNq2i6Po9pJUiosgGjjAp1V2LGb5A6o2ZPFxOd5SHa3JZf/
SFzH6lviu7dB673uq+PF3B1xZ3H9L/ZVU3ncQBW7xOkKZD8ijVUl2s0d97/1YHhdY3ytJXRUhVg1
KDOcCg8Mpc8mkPp+acdiBj4PpVUz2k+dC3ilR6KSBmI780tGoFqWV1BaBtdtlne7YWlkb2198UEW
31+mMg5DDf2C0iDgyEfiPEwrl2IqSRIqhfVDrUzit/YFpDVaeyBNh05vTfdr8ih9Rge2NtKcXdGF
5v5Wc3TG75iUjngQhYljiahtXmQ4yn8Rj9r84KtvVdnzLxOXyPlZRUjsv7Fc1QYleLPLaJ+6Zfdb
/ilIdfjphtv7AnRIKumzOpfyDSN5R45/IwVVvk5o2MNplfnYS6w4HqC258Ag/VggrKCCylrTImG1
kSFxbfDSe50NQPDyS2txIqBqlT5LY59EZQne3sfzqwGvabAvUDStvwxqoB0EUG7B3q0LRxINBgp9
onqeBmf9df96B6mL/GwPpG9zqOTLZtqd7e0Panzi+waYge0qK1Ydz2NYNb5rD8DRDqwG75kvhi6f
TRh+Vp6yjhQ58icjk7HjppemYaEwTrszzOGeb9f/1n4QxZVpNAH20HY0j/MNNxUAUe3iuaAwmHEf
Oy1aTLdZNZ5zvBJWcQLeEIPPc7qk8nMi5jgFkF3UFys+Dr4attmYe1YZmgVcTrOm+zZhNppZ/UaA
9EvK/dbMmJqXDljIaIVR96ZelFCKs5kS4QwGWETR/YS0+7BZQp0Fcc2E1ugd5XsWv0a1LBQXryu9
pw5srynp7YwaZfGEn1TRp4CdYg+L22OpHZy6cKzZK0W1s5nXpvRM8XD/GoGdyU7hsE+RIq7dWt3m
o7OGV+hLMpNzUvRk7OMc7j8lmwog7Srln7vm9/QVjFMaEpwCzsfy6WSPiLtIL2uVRezowpjYYKnf
Dn4uQDWq0/vpNbv69/E4wixZ+jRrWbS39Ul3IL6iHndKzN16QRGx6zFdtDCzcTj8LuPS6Baoh72T
s1boQBj1qbfa/2OShqO3WBMxCaInYWrlZoKpM/AkdmA927YJn+NYX6v1edXh+TOUKBgb4QT84PV8
aZga2ir+RsbkYXX7ljN7W98M21/vuGSy/GBGla3VqzYyYobIVy240usZ1swGStWtSEy+CvpFw2Ac
ipThyrR80JfGmN7OtCNygHfnQkemxLzsVc8Hk+qwQVcNtIZ4k4E2w7raCErAxZuuyJ0YFqB369PY
kIvXivnjxIFPuC9FzRxyIhX/remDGpSKmruLzyeTEeaxHCqIQxJ0i7cc0IuHJn8MCedSWo5F7xvV
tXASYyHrVzoft1mUQxKl3nR8hHghQABxttwsL0UWOhH0Tf3XDC0dZ/A4fJBXfwLVx4j/0HnLHbdH
MVcLZqVFsQlIqi7SrMInwy0wUozTz4jpho5ZgFs9LFEoQt41FaS6UsNmzOKRC3827XlPzWvUYu5D
5EwwvBXCHRrEpmdDBglvWFb2lkg63uSe1c3J8Yj5Qi75ou3eX2VWnA7/3PZFC+Y/oVsh82azjewH
UCnTqauEeipCN9S7iSjM+zEMRFG+wIVCUWdfr/RRiPebuCx8/owEYCYCodOBiFOiplgzPEkm/hvj
gwo5g3jgwdX1INAnBM5DGq9JMhJ4yHWeji9piq8eQpRlH82LEvxanDVT/VllF+rtKdk1A0tbZ24+
LymK78hXCQ0nT3oS09/whj8D5+kfkKAuQr152uf/PbjgoaLU1web9/OmnPbI3OFpgNKZRp9zvZA+
9w8gEKMjlRSRhvEI7n0oMS6zQpM+rRCOWxR6jW3yLfgp/8Gy80EphlEafv1dbsT5nmdPFnCrPIKL
+JdrESotTSASpPDy4720CVUmDf6Ujhd/AYuQMK0bEP4po0hGPMN8lDBEyvwcYiJODWnGN7bcCcNG
jU/xBzV+U382CdDxSGNxkM8s27h4GcbqISVJRTllwOTbmcSoHxa30LnBw9J2G6Er8/Q/DoByHFRv
94XkhMVi5d75H8Qqu+lPi+VJkPWxRsFG7ko/ZLUqE1VbXBYdxajqy2ErwbO6+zVOejqRVRik8WOh
OKy+7ld4cbRmS4H9/zRLFZIvfQ5rGM1k+Et0QRvt54HdFSlw1lD3HvjMG/cPQ1YHL7bUSgd3aV0b
N0Ok9mePDKH7/Yab59NDzosFwlxtzuguV9kJ9//IFY93zUMlJNRaTq8aFtRoZdw3iP1drlZAhouU
V1ysaOxMlHUWOWw99mVMbkj1d+D2YmFQz/lz63L0YtuTolovHGOyKwnDBBOKKGvWKWzFBljVhgSi
B1nenjFYQbzMDUBXMm234JvbYt5+V1mSelgSVJS2xNk7M7b1DvmgXMWwqnNEOVKiJDsxIdbnT7Ux
NvNtOyAKjr7YvegcPFIlBd0C8i2YDGjJDJgUyR5+TGbxFbOjyRewm0kBojWBr/d5Ba0wjOSOXim3
/wN8kcDpwWJ2fn/sOn4UGtV4yNDjoqWb6YPANQXVozGL0S+j0UNDZ+5P1TVA2CRHO+bAyVsWjNdP
elhfLWt69DjHgx3fHweDZqUAK1JIW4tWYaMzg5iy/eiZ8pydI4eYyf+zX1VV2PmGYmGtKA411vvm
laCOEG47mojoRlSDDs2cQRC9I+WGuyaSrIT7V3XxOgN32xowW0901Y8pOFw166jXHM9yNkCzlgD0
txAy2dPdoBlU+Bmrn3/NQMhgciLORWKmY80D+Un0VwNj3IBoF6DLHC176D9uzcqafh7SQbYssPX/
Zl7MAIVeVPHrMRt07/bvo8YobUu2qw6D5yKa9Eqtvr5//3De09y1yL606x+PtKc6YbaBymfnjruo
1vexyiChZ1Ime4STYVxZsEPNkWvFk6x8eWMMqiuIk0IofcRpztl3lOhfiPNnZRHnbcI1LXCRlqyQ
hGtbpw748H8my+A740IkWFu+8ZsdOyF4EOggN++bySRAin85j0PUl2ZQqqJzDdbpHiWSMWIYKkBy
caUeDumASpODlh1S4rLRWSl95LpHotWBfFStslzguyaLjNRzME69dgHBh7jB4kWb1vorYaZrZQvO
8OidDOwrJNfL2x1wmGBD5unNAg0ui8spOUc5jJktXCHxOJ3CJrQNa7cu9o/yRBF10fT2dWFR20IA
JZhZ8q10ietx13NGUwY0Dle+X16nvYmq/i5APrBPM0GrNqpQS/5/mhDEooV5IbZt6uigRtnJDdvW
0XuUbcjFwtMqjVUbtFIyIuqeLGFzSOODsebUySLfJRwS4dZ2Jv4b661lJATkQaOIpGaesdEwr7mC
kASi32N4hpIJi4ICl5ANDA8K5hzmhD6ZN9CJBzayKK09dPBEKXS0r4vVmceKy9TaZrwfhoS3aTO4
f453MuQZlvgTP5jeLqU42OVZkDftmUXBa2tWSa+WyB9W+xhXz19zQ+gHcnz4UH62D2wuOwGVgNNA
iHNS8GxPEoODovaGgagSBKAjNMxSE+Ah1aaSlXG1pu39U8yr0QLWcT2BldxYQo5YNYnkd7O2cn8W
Kj/e4LQ3LMTLMDBw+24NCXb3l6kyUKCu/kZgDO658+vTmav3oZn8wu4dCbazJKte0QJrVJNFWr6J
A3Sv6yr+UqYvUj9G9c1Jkyi3noGZxYEJyq0AVQiC5cT5LXK/eczjmQ7kEI7bRHtvSJfj5B6derOQ
pKDhshQlg+S/ypcjI0lKCRp1o7mP/n/5fBftoDCbmTWdnyv94Bhgai4AMZV/devfv7/7wPsLPHhG
JyoF7HjEWZSXG+ogwy5sOyjogDKSCLzsuem7kdBCzbPQqvkFPaaA0H5EvzPnMnwrtGTBiqRu79wQ
U6yVePB0Co+J3L8PAiRRCyrBTs7bDvo9QhfGI7wVWR+MY+h/poO+ehe9vKk4oArvfJ8n2cLAF8rZ
/ffp8Ey8lEfTRsFzbLj69oSHM+VFFt62TaYyxJK2EqcChD/Lhl0PUGHOYdsNAqSvADmtpkf0fKDC
RDfPRWQVZRp22ZHW+fJWSxWyOnwZMvUNQn+zq/xgzyKQ9KbzWMI8WqVBcvvjnhxWDr3f5pSuWjge
a+LoU/cAx41v4IFr12g4izHWTQ10jdu7AFOQuH7I96MDKpN4MAWNPpLewwaxV0or4/2IyCbSDOcZ
Vcq8RjgW803RbYXzOGYwKvYpNXz2rIra+U9ByyFcyGY3GqiEstltBZgQ94A1+oem5EoXCvKlaF3H
oM7dNJUOooSwvqTYhC6DeVi37Q9qrBhRoQT8jFaYK5/BMfomLXIp+6ep8NPSfxwkVUGpl5kfvN6V
Y5RedCKrQASCXqF1FzD5DrpknR7z+wKOamq2W/+MM/X6rSf6KHPLDHi+egSrKA/0J+OarFH8u8fY
LA2xr0ZNFfx8UBscidxRNEdYmwbEy3hT+ozpwmL/TsE4VkdaS3PabiPmYnT70acRBVEtaICPTUAn
4/aE/lWA4NF70vxxVSw12LtIRRstx6+4PuuW8G2uqjcnxx9TrAcy85Ucyc9HMrAK2sWv6n2I9rln
ygaYwe/uSa3diZbdprTi+N9G9sIBwYiRWSMUhB/UywC4JNgS91p0beIMiP9Q1L67ihKVKBVWK9qy
BvP82P8dG+VrluzKuVeFEuj1qv2takRJ0BOEa/PL8qzJTCxhp007F0apWn8qOYW1KxPNhfA9XlnJ
nWtXZO6qcJn5nnf5raFA7dr+1yp5d3PUdVbjrts0EBgVz6vB3dvxjpHXuUnlByHOTJE6eepuegom
NNFrTrUzSFjGOD4gPjLjhKk3sc366OKer7Vhji2RjhmIjD8O2S87V3gll/RR+DU18J+yF7QkUHoj
C/jEOb8LY9BjQRhPqseodU7lHDHf5lUNPN//L3jTFpYnojP7l/eBnDoH77pGoI5OinGrufDWptF0
XOjphh25Czfm/7N7KY45RwJZWGdlje6gmXUc8CrqjNpLSAO5YsI6aVQfvWduZvAvLqBioO8ArzKo
pbvO3oePVWwEGATPWGLKXwqB7670Dl7xr5BYmRgPsX+OP/nnK4GzhmfyKzyGe7+AS1QTH0K6fzxW
uN3YWyUjPf/Hf8D5ZHM0As3r76Epy8qEZnvTnSp3um7KQ1P3hfkD35ftxQBLA/FRzsE1RQXHdxBC
hMtOxzZSa0xLZvNXal04FIMRorUdoTb/41O4VzivSgebbeW8uXLzTCXEWuTLjH20zWzVO8BmPj2y
OZilFIH+QTQBMwPOzML3+/w+9oszQAn0XllIWcfapiT4lZ25PdFrQN5QxBpsvCowxpYlQwuZiup7
pNMTM7CwDnfzxwwHtkYqsdh8zzh3XIA4qVVsEr6DM7OTePPslxyq4mZ82OHCgr3PwsEynpzRLfch
nmmPj3k92EPopdsY7SsLWFcCbwAKSBCyxFyVbgIjkoiEqbPN8Bj7rLcUFBN0Faf4/f/UGD/pKC7Z
DQq/n/S+3II+pqSY5LnuEFk2xX+6fajgQzp9CJyWVJ/igL9485g0MFrUiKqQftWS0sv2ralOFbmj
hU3ivkND2CMq0eRKyusipBJtxTHgnc2Xf1kpI//AcF6CLAO8q9hfdD2PwrjyBw49HkY2SPTRpzq3
YC5QkIQeGAtPnDZCPzqJndZ/oV42JL3NO1acTMoCntJ5DwDYm/OR3AHTAS2akk4G/AYt+qKrZSBm
5dNXUl7UNMpQp9XAFsv3lh0LkViZjbBIBtJt73gSRv5IwQdUCc7EfF9RLwYK4kqO4BUogcSEwC7h
RI+FTrcdvSPxBKsMzG8pXxdlhpXVjfRWC8EVt3DGv2yzneewhPKJfpgV20am2WBquv2A7oz7ZU2U
DEv1PFEFItSg1gmHeATCNuNEfu0ElLl/JgAxlZ/4+KzULvPHI/NshdDWPPPNZY0KTuCahfRiPRUa
r1H1HSfTGE4Yhw33sxIBXY5Ta6fQ09lrRIPFalB/XqfZsdRzjTilyAkBwTuNhv/LwXwL6RCOH6AD
kyb36ceVmNlu8JnheBzfVH7M/WjZvC97Bm7o6R/QiEf9WiEMQn11fzCq9V60GkqUUhp/0XpXHeGV
gRi4lfqACEb9FkBHwXaxLwRTESUcl1cXic5IG9FHX8Tqfslpq0/S3W6ri1IIHgx3lr2DKsryuwV/
rQ6aH0E3biE7+7uZHkR3pKhbFBowsWuNL6R0eVeJslGyrsxDGvDJH8buiMzeUA0QCVIJW33rxDyZ
L3GDO8k0MeekFWwy4Ru7ewSOPN9ueDcyMef+SXjgVn3bg+0tHNoOossmUXi4tZ6++gIiiMuRDtoW
eNoepKrIfdF5hAD0y5kiiMjy8LZyuk53pyHabV+Hi5Arc5HDWxitPoRCe2RDSaETYZ0g6p0gOtAG
CSgVfHdPQwarYxo2qnUYgHZ5XkBWHV9ZWvF8+kUmPAB7LyCOua0Gb71DsIzV0Y26dD+sml92WN2a
bZZiHoeIt6SI29SR4JeHvtpahvJ2UVpN0FiHKFQJ4AmglAIvyijTjKPiin6L3q3dL3yz0bvZXB5T
yB09Wgeu31kS0/3MRUkmNv9QhgxFXq9BJSwFPmaRWJUQeyxTlZG2P7SKN60qKxwy8SIW66QIQ4j5
jso8WZltLCLmrHOi5XV1AAyq4p8cG1gG2+q+unbNMMCz8BSD4Z3KKdqDAMkE9NUYXswkGDwM9gb9
7zABH9SpOrl0t+g/elqOltS4OudTKZD1mticGzrTK+9C+Qg7qlyn4donAxgODVAyikRuuZmJ+7HX
SLpU05Y6SCBaUeslqIc91AHfQL4kUCU4MGCAZfcc6WZ3Vm7i0dZt3PJejoRQkaNGQvAbA7FgYiTs
/gBBng6kGpfINO4fOV+0OaFyhad2/JHS5GD9w5fGOcnaPTUTX6Oggiwoe9jzqD6xHRKgmffzKiuP
Up55BG15RTbZXhrTQsWjh/EvgA8WgTozA2x2YUtaOf+k8w8uZVhiG5oYgHTnPRTPqEqdl+AscBIj
uLBAjiC5+R0WTSzXSEsj7kBue2jw5L0zCIHHkusy7vZH8abj+2leJrZorzNXpT1DhJa9TlwTONVc
BPrw0LZGiPE4wfL6nDo9ikllbNP43kB3dhLqcMIlydmm1y84UDbeUwGttPEqvc/uUp7LnqejhU7o
AkSu7szVnKtGD3AmEi8ddEE4LUOI276V6Pe/0GtaTAgeX3qPj/KxhTbfYdYkfWDEwhSLzWOk5zwy
8i6RNwg4R7cEHeGF+s6vqeuyk5OVZ30oKlvLggLtCxRC82P6eWfECcpVbu/S02L9h2CF5X/gMqrG
ZbultU6eZhzE/wZNrIvSAescm2K+GzQ2NlmXiy2vWdaA1CaW3GETXkinh5Xs2yctaTd9DwniHF4o
SdJcCKjHvYg/dcrNKBKzBNPr4UhnKTwJO71rFXFsG/Y5IGUT/Q+cCnBea2ndEkSml8veYjP2ORZD
ZQod4ER5fysV9VrzDSLhbOpfD2qPry1joBc1r6VtONtzsQ7nOAJxf3uOy612ASsx/sV4/ukvfqQy
5Le6Le8izgU9gziMDg8ya1PXVQJDw2r5xHLK9auowGb3o/IQi74p3ypzojeYM9uhkMZVjGZ0wnOK
ZewqE5gh0OQ2QilhPmBlhaG6U3641AA08bbXgeTdfr+UaAsL4PTptERjrTm+ahYmUOwmGW/6Feoe
KVxah2EeZRlZegPkppe84PmikgF9wsOtiXLQ/agdjUug2tqyFC9lorbncqioeqWzXbum4RZqRrtp
fMAIeezRfgmycqX+fLu39n1B6OBwHCGu1/1TMPRPL40SBSfeuenSTeXJHwUA7hvjd11SCKG4TT7C
M/O2BLJ6yj1cpplVddR5VMi3e5+qu/gVeTlMIYh7V4b6zkODg21Wok2d/QS3BaxolNd7k24tSzSS
RkgCcecnpssXHP1e46V6MaLloSIaDPRcMM3IZgUZHTEpqcPYJYDdc73Yey8IuAkGUw9VZTVJ+YN/
lVpJSEjogAHDwlgoV9qWIHOkPuoghQn7YpzJjwjtn+UsIBSyVn5tR1hhX/LuWWKvFaO9Rgn6D7TI
4xwwMqypshhB638OqsV5VclUxWHu2pKHSaNRVfEO9imBqdM5c2IxJwTXOjd/fmw8eWoDz0PyeAmY
NHIrcLOPX/RgabVkJcOjERUqAiqhb6ASkxPlCngRer2EehHUcffyzswQ4cNXfmX2zPx1N9P1A43e
DVLppZv/7wKsBIAtmgDzzMl/rNma1xB+jfcZEPQzW8p2P6USZm9VEhJwmV+1ZFqUzoBp9cr7wiSn
1IvMkxNhZoUwzrQ/jwpeRgaQWgQ970LDddiMQ81XkWduBV8nPktg/khy7vaHB0lnkmbT5zWXXpzI
RvVPtm82mAGXWstQ6i/GBX//IV0jBhB79569RCuHOPAdP6MFbBmAkdcSHeAki+qfb5JIXX+LU4Nh
a46LA/OSZPH580N/X6EzcnU95yqTiQisQpzNm3/eIMY1Fm6mMDJFTnfsB0apRud9Er//+Tr3/UXJ
C0VdUKopQKKRmWstAspWGcqKmIM0k/rreumfkU7purRG9zxodgwiMa4q8xjhh0AR/CjAts0XeDMM
o4KRE6FENSgwkYpuKUiUV2VAT/GP717mk5d06xQXWCZehu5qHRvA2jr8I0BRFilJiNfVcfrztCNR
+yFJc1FA7Q5V3HFDDXqNzY0qATrpvOrg9QvrGHnrHJeyCp1k1+KW2FcItHkUNsbR/3IzVTLh5Lj3
EWIoXgdsZMQ0lnozbAbCtiMeXQUn9DxGHEVcw0y9Y/X0O2RMa29Vhc1LzxVSMXR5nD7kfzcrzyQn
IeVD8dqmcZUqpSjQ9JUANFn5O/kdGQ3mlYo7+R0q0zEvfRm4vNdZ6gdoqxM/DMI4my5Rr8yNm0eE
Lfl3UcFTrY3i8Hia29Om5FgTCrRwQAlTBXYL5Oy82RcxfCq0IvYwtM3/L9h/IG8QYQ5uSLwMlKT0
SW6zUyeP1Tpd7XZskKtNr8X496fmf277Xaxc0m7Xio0TgNJdHvnOp6Et5Q1lP6CcAyi5X7+irOk2
xytjCwImeJlffg5juapkKKxx0SsHqcVcmf4Qvap7IqBOZSFmSNvmtcQYQ3ncurU5HXJFccPCKuEG
7FLnfCEtBBPjeNTbFdjWpPCZXY4SEQmDYBNSI3EG+vk7YxC3kORxEBu4EQDLdVA5umzq6uYoKs1J
/DdjPPbj861kmJgrsJqBYOBdAjSpq/FYzliDZOyXJA1TWcFPtJDttv01Aqc6X9FtTlnb8ftqPRL/
7CquiThPm8+UA8pOirl/gSBOcdtRBgbEXSGuK8DfDK5uIaEZSVGMBGhAf7KhyC1XEAQD4bqjue6e
AMxclpSV4vhGgONvNqcL84YSxbrKn31cmQ3pZq2UbqiFYbQIQ9ME9aElqU9D+HmffNOUodYZWEbg
4qfdG5fsV03UqQzQznaTUVkogVl4uc4/+VXr44/wYI5JPoxGXpAwhO4NXbwBX8Mq6bL4vBM6AmCp
dDy4VKknXNxP6bGtrWfYaqdZGeZBJ4vzVov2Q9FeqJlviUna6NVJP4UC9bqnhjJ12U5RDSITpizJ
rdogg+/HtmeyXw91NoUjh1Zo0Z4T6a2MpV9feh5BH5AnIjUOLlfK67b+W/ranW52q4Y/fGAkkC9R
XRvvs/Y55HQcr20WPDqBEFoeEOIOUnvsyKeGSbxpsjx5A0JCvq78UBvDgcbcnlGY+urHQ+E1STFp
AjlZwuwk34to/UpHW0sWvlPvBX8Y1mHaNBpXwPRJs834w0sZDrZGZ5piDPz3mRhn3OOTAFrP2lhd
Pl+gBW6dx8mfuR7yyNhpUBJJ3Dcsh9jmJjv/Zk5dNGVSKkcO0zrVF/GTGkrCTLn8Q7ih8w8mB8M0
LpDLUvG1XhPPVoKKZ2iIh6ij15qqsCd6n7mIHcOeplLul9XeeXRYwHkdqo6GviF/3T5hWQlqq9ml
xWXahPydv+OLJh5+h9fVXgmZz4D04uKEXMhuukwjNU5b078nRtBt2GuTrTESf5o6Oxxftpluz8jo
zxHZBt9OEyOvTXV+p3V4NjIVklUi11/zc4LsSET5p+Cr4L6TWKFKk0TYEDmBAALxpLj33a3b0Vrw
0JTEBSBUjs7wPxyWLt40DZNIQzjvJ8Ne3PuEqV3EEtmNGcD5AiGE9AoB0DcB3DP9pUdaCS5dLB2H
CHSDbACjpCvd2W1f1OG6bIdMmx9K2x2KiesVBX0I83ImqmBfh3JhS7m4TLTg7wwzYCpJZn/y7wKs
18J0Jz27jiIUxzaDKYwhHv3221VSgG+hMnsy22B826nq2TyPJB3VkfFNazxFCCsdIFvaiI3dRVfI
EneBdrdCF40sd/sROoRikNwGGgyPC7pPm1VsAv9IqlpMpYzFhvBduxyuKq+V1kyl7ejeOTn4Ns3I
vY5LDTh4ITzzVAp2STUOt1uL8HfjaDVw/fmu/RMjkt/L/FUyIlLKNF3ThFPyDu7P+gt3Eaf9Wb3A
balzqD8qkOATps/IA70nagM1lMhPbaPjYrT5T49Rs0qeEaGhY5TrXmndoNVVwpSRHMaCht0IA3J+
iSntNifkrLRQfLpl9JGatCXcdNoQ7xyVB88PXVhvwG5vQM6SX22ArI0njAaRlEfuILX0hJcOyDZe
m7dMcSiT5W650FzveVFVrWV+pSPsySVtNyIZAh3w3EEs6Vu3hHobA/3huiWuwlOuRVjJS0L6jBap
FDZNVVe5E8qJTgChv21zH1yo4UfBDWa2/UzmH3HAySlnK6SRpDV64t+4t132/754R4V251UGdLdU
md73GgjeWE1ToRvZgcxH1IHEh/biYnGHbw0iKIMLfV1E/2Y4vSMJOK26oqwx8GYggWNqUeX7j1OQ
72hyHo78dZEnYSpZNdiKqx7elpJZGqVSrfaHRdT3ne9b2C/akz1+/4vvdsWeBN+nV2oSInGdFD4c
W6lrsP7Q21ITbuz2mM6SUn4CTrnYKyfXTtsyxj8tBuFx/NzSfmghsnnrjkGX9YR46Zo2YTjWa85X
B1Hu5freXRCj6Z7vht+0w+KR3+AXLDveG+tiuuRgI55QjRQAspNk25jDgjTe3Gb/rlkI6AvH/641
dP5C0r8jTr6IwxZQKeKHleZVEXhfKJ15DgExrQjBm/WWdJgReNpmIWsYuIwIMlh3cJGA3K3mhe21
C91Ag/jBy25mt7A6kljKtaeZ08zAWrBMtULysMgvvHF7AIjQfHJep3bXYbZd+Ejn9db/Z6AKS1Mw
VLxcsv3a1s3oO5bCygWNRDdRegJpwMim8obXhDP5ZqVo8VQ8ePR+csOFly4Ef7J7jk7p996yWx/C
1fJZ2fi+ACxcZwvOQ5j1m5rfDR5rbkAry9ZLxMzsLWimmyQc523lNov3zfgqROlb5iD3DR2QOFmP
vouITp3apebTzrAahBtn1hTZAQqNcvvKo2uV3guJoU9hc1vuic+4e4pcWZVqzCLuBeDdVAD9twT3
W2chhQlUS+NBedlWdPsMqs4eofGfB54qRIdXVSovV2BCk6a9IeWzmYq0dJRM4dNCFChTIdXXnMe4
G53+tm9VTqmpadC/nRKkbWFcwSgW0dCRjYpW6+hxbMsHxIpXYywlIXIOhqkt+NRh5gfV3AinQP2E
KfE418ydabFgGAJmSbYpYI9ZWGTYb10EBBYBbEiUEBjE/H3597J1FcTCdU7eAdcsOEgI08o2kQbR
jMmxUmd4iFQak0JwDca6ILiDd+pzX44qlOOkuiNv6sQW4NygIC46XuBeC3vb16IxT6V16hSwpkrp
kXgx1/cAqkJtMkFR7dB+5CGTt/hi4mkJwvdNI/U6os//tMUo2DKMQvXd1CvE2yT25NmEDGPF0i9Y
CpmOPdkApOxCJE0w+gF53OAIPeDex+oE2oD5KhZdrcjmQ/PfyekMWfb0v5PnqeVT6yo+NDvpvatc
xMObxZ4akZ3lLbDUfnqkqEB/UGWfJYl2YIka4chrhk27RZmdc8a/xEqRIxemks8lOdOwlel3MqiG
FlC7/2f2hlwWPJQMSlXmSTRbPlayaJ6wMgvlLCuiQOqdvKPBeu+T1ePmirnJJRTzVbM9f0/vOG+D
+dx+KdA8pgIZZc17sv/QLgSjfTV6CRNz1mXXtzSaYUAffzbqN4cgW6XqiExqNwkXAy1bTPemic0Y
0qnTRODfBdZxWVqk9BZRKGvPnpnWYWRwiMgcoA42HCFipssn4hEphq73gjcKNtY0ixWMGdf+0iOE
c5q7tFLqUKYe17jYTiD7EnyhnlUOoxOb57FH6XxFhUA/pWH354jNxj+oRQsHDf5Lt5eXT4WcxP4X
2vTUdMjvvtX2ZsZsE5UAUvvda6gFhQZ2iyx6SiVEVi1TeRvsR/hSDCXIgFhdRKnoLd5ze8C47UrU
+JnROh7AO1RR2N8mduiUmS4Jaoc5OwU5jbNj0q6xf4e/N1D5uzt3S0Gz45scFuORcsd836Ccjmgi
tnflHh826oEkaTjxpMRavwkjHo7I9cx4MJsnPpIlQ9w2F8v40OIUcVPB7HTb5tC5oNpmYFr8DPQN
OldlSDdq6PfA5ueNZ2ljTNNVvIZK0TViMJRKr+xVi9qsXr1dLYQU1oL8cqttPvzlSBgDbLP9Q+UX
1SOixbYkHqnbRJRUfPRc+8lC/CR8BC3+Ksd9mkB0bAG2qG3zsORSZJE5NZI9WNXWyRJHkdJ2TVVi
DZu47FpArbuqqqFhAanIs7oo+rTfegAisiSMa28PLiM4wIFhfiB8ISN18OhF6E1Mgr4AHeLXHib8
CJgHwMnshp2Jo32vJP2ZcLq9nD8xOWKnf+ljzwiocFMxxAhgu46cME5LT77HAPfmVvUtNBfdkvlU
VrTwYIZW6xvHM2YFZR1cIgeX0ncdFqFV4wduUisa+Z4nvMMvAn1GOLm1GbEGDzgs3epyUW9k4hxQ
09DinSms6RG2MuE0Z9f1u80KsQq20+/vqjiWSNG8IVDFUBT7Uaxn0IyHyPrF+j7dwrbidyrfarCu
nhjPvsScQd72p9Ma8GkJiSaj3BGleBl5B0x2Um/FfDkwXG3n7k74ScL7IhhJwbpraczuDR5n0VUw
UGDYiv8rDDLsf5xJ/7vS3qNWBaGY2AVQYHVdPOzGNrcqseJKur+pY7PF6yRygN1e+cZDrGiKw56S
bGGSqBMLe55rooEHj6WbsZdf/mXBv2Q4X8BHXqYEZ4qcizSIOWvkphN8wIm80CXjwS1IwNYZC+Mi
q9s2rIxUsPTIytK+NNjceFyn2qbPp1ieOUieI/StqvJ7wuc0jLKbCGBTTBtn2JrnDltQQlSaDc48
tdsmSbAhvZhH6hOSp0n408X2YdRCu6CTyszbEXCtNSoRAJEnaLZnzqxjYgel/mNF9rvq1OQ1Tze6
gT7H96EBcyKYuq0Rh3Oh/jTiT7mIFG9AtS1V0BViEPN+x47IAPzWWehFrb8kvM8mTimR1afhkbEz
IkEmozKi5bNJ/NTDt3dcrgq7WA1Hf6SEBM2pA/+SemRWzF5DE30//LqlEk5MWPJ/ckA+wpNdIA1k
0fprjTllqL3Ny16LDmyHYZ3PRXw+2Dycu1n+HqEwXO75KcyYHTRTdYKRFnyyA2ROgQcCHLD1UmAj
hxL32iDxrg2kmDMrc+nG0BeL+KeN/Agi/B1KfCwNHhrW8gcPpUM2Hvh2PcXDd527Sf1U5RfTtZ/k
XjZjTmJv8mk824W2Z/HRKDkTyPrdw3mVuZiVhmWXVBE6vYJ+AMJrY9BbOKkCzoVOIPSwg9ksyrd1
vw95Ivmj5idbIhpvXCmnUwET4mRT1Iu8GXK7L+RPFKkS6DJUc20J8uwGb2neBlO9qj426+LLWaPG
M83yHW1RRiefTpOPYqJAP5qo8b0P4ygo+y1snndHuhdKTSxr92QKNss9nhtDBxSmUo9Ix6luIMui
yhntwdQshQSJCsl5kOf2dIvwSHZ/2THgNUhhkKvBX+DTURk3SX5hEipYCMpIBTtd+jwiYuqFd8iO
Bl3uUImQl/jJO22LXAhwMJLJbST7ytebK3SuDtTVPhrbgWkpv/mJPnRC1HntQ5Sj5wNvjJg6y26n
JFdxFOar6gWWCkas61Y6mpu85PPD67K1xXhPRLraSD0uVtUjD/L8R5J1BQh6c/aOUAm9SFgUPpuK
WqpQKmLp52nz1HlQ+ZySJFWI6FXWyFmEb82XFlbRRw8AsoLZeiPCf9Dy3zdd71BnXOhBe/xF8MQ7
MZ6DiaDU+l+BAcn0XG9cPs2NsVCkQ3gk81Qk9QEb/ppfcNcY3NujWCPpoGPGnMbq0dThTQ8JS7jG
wX1LLw/mOqiUVvxsUgUtqvStBhKPon40NsJcp4Gnwb8HaF1ED7/72p4BUO2dB9+TSG2dUOTstL+z
ixNy/pWII9kx1qnVcJXecGuN/Y34c6i/bRs+2yb/lFgJXXh6Pj5V3fT1zIKp9LcEgLp2jSo1BASF
GH7uo5QoT4PXwp0bscb4tMKjxHDnHAyurFGE52y2g1eIq2khFWCz+KwNem7is6GV0l0/q3Djgirm
k7EzHWKYxdBrqoZWUNk7NrjKV3y2SEkzoMVNsckt1FiT835xd1Ck1YbHBCI5naXOm0NsyvxIFV80
veC5oIrXBhw0/U2iSzaRRWJvxzWMecdCnskn9bj7P1TrstJVzqXGbz2UDgH0sSjQ9YZxkLU2siw6
JKVCC8gG5HylpRJnuKsLPNAWA5fL+KW3K+XF6MMYD9S+0n/GUNVzyOlznmizC0REydwD/q7UqIcl
ZxoZBYIhZwJZmdnRGqWDiwXlaLcIho71xNWWKM+TtaFIzFhR170AJ46VQNVdQnIHGvSM5fLLD6LY
KB4F4zLRCxGr09m5tXb+3fIm0i0KJhHQU9gaQJpFb+kkmF3HQclqe+nVtYtzzhgcyyRMHfK4oFxM
z8DpuREx0n7fGRy28v7U8aWXhmRzJ6IfmvKxlAVuneWo+DXBnRnLnd3gXs9io7k7ZikhFNeCJFue
/buqhOt90HL629r+oITwpxP8iv+pepzZgyomhDh8H4bdfMnK7eUXAgdNNLWMTQ1uD52ToUWbhR4A
XcM8WTy1l6TttC8slTmDfl/kAaJ6m+9tspZFkPwFGjMTndUK+IgZ5AUzK5Bo5e3hBucSj7wtovpr
UEBXCJzzbTJcjBYlOZSVu5VWKKDYwCiyLASGMGzp4C1EDFJZyoYFO05M43RLlYkJZWm4OGfcnc68
OT42vumikWf4G1pxcdiY6eQdvmK5PxvhpJEMNkMFMbjW20BjXrOeT72l9W/dQEVdwtu3gxOSl7nL
zTZL+nBn4EYcgZmFcXgGT1m6JM0VjmSmGt0jXDUnVmrmZZyHVpGH7MRos2kCikMCQkaAauDe4tcT
snDud05y9jxYMqe6KMvhu/DDnKsRqDqpnRXypO3o9udByKTBr9vdTsRoVR7RqBGjqQ0HD8fJ6V6h
tJx/gH+RGtv0S2gttYVqAAgQfPlAOzOPCx6k9p1kodh/K1GsQ8ZLnOIwwyCQQLKRNdDUy66c5tvs
bHt+UgJo6kar/LjZSqcxbrvAqK5zAxC7yKakT/9ubc9yphKFU6NJVD064oZy6WR3enKFl68jobUP
/iRpG44+7RDGGpgCJYMyoVnEagbHCNL4zsQKuJhznEtmfBiDYVMdW4MnN1tTOZAva7goEdw2KuqE
+MwB6Of052/5fP9GR2l4f8Lno4n3+0Eflb+pzWtlvctKINkBHNYiDvlqaRG6cEcDPJXy6x0pWLHf
NvtGR4ODuOEEyIXZS2vy5ca+OOgg2X6nIqvCkUxQNv3NwOPbHdAaeNxwEE11orOrvt1nNAg71gO0
gxtHQcR6Ue1Trwmp4SrVRiuDQktR+/IrIBrB/qMA8vlzUYUhm1e3ZzhMMfV0MYazeCEkNJuFnEOk
C6Newmfngzp2qHq7/9Vopl2Oi8qTAl+fZc37vcGybDesXl68S2olzFZuP0gcnHooxc6V5h3TKMx2
HHSnrqGor87622ph16rzz/wfbh3Y2W2q8fVLSFI3i42s2DJhj0XKP/TYkQbS0cYXTbq+UELIyuBW
rtGQUsahBgptrsjA5I3SynfmqiiTgZzyK2bst+uKKz8H3Aq8pqwzXoFnKJcNbW2P3M9PgrgVqEu2
ZECj47dTcYMt6Dj695cpJrF6n7jOxmFrlSU9KIloFOjGcOYQfmqHnIhUmNZgwfkAL3ALAgFEkxdZ
Gog7wvtx/fFJhcsO2y6wNkGClhjVykjDkTBb8G+aBm9HMYnZK6hFF5ePNAUkMkxiiXP/UN1uQKBU
D2Sq3AU8RkHB4zrPbsXoJYUaVI4GyB7zHZXGy+LlUXZaLj1cRnWrPdOpDav4HaE5n4bEoxyUje5h
3ToeWb+UtguL4Uhw+CtfE9Y1qAvv58iki1Jtn+M+70cLoCxb9JmdWqoJ0pss8hb/beP1v6kM4i+R
pchpE16ozwqCFQk6KASjze7x4cWv1X5RbrpyNCK26LhmxszD+C2bzsuAeg7+wm+YdOaLEqGLR+Us
vBy1iGpmwXjElUH2+FL+Y7ayWs62p5cKKXI6LKUcKcRgWNZCXtHLxW1nQcsZbubuS0E+bYif+Tfq
0UJtP3r4trs2OOTpMe73xKtaWMYR17DgJpGCIhrJTmE3MZghDL9qYuTDbIWXz+Vt9vEiTbclvZm8
QThbUfCVefEAWyNt0Dgulh+4zXWQSsU/HYy176y0oNdpMMOkiwQ6IJFSUQ3n3s1emhXoCrxKdUx2
RGDXTAf4m84GML88dYcCBn/wf2fBloPkdnU2JYzz6bYhEILsd62djvVAsgplkvmtsV94kNMkDkaA
SidtbsPD6CwYcrivXRyzSQUB/+67gO4ODuaacITfElkh+YQjaOJNg64RShGMGjAbUVBQHAO+88v2
YjIksK+jqvwMxvvVCf4GGEIs630XY+DIpc0l0rk7kmskI4gKOB3KaXA2intN7Txnpv+NG9xiw84y
VTeV0tGYNYcXckMSYlM7hh9p7/+2FdwewYtTKrhEZXKsPkddha+0WTH+/kCcihjBVk47f4qpNftY
csabpcPEr1BR839CTQ3wnEe74NQMEO2oy4dntrp/3OYNiiEi/xRFb2ysuoWwk16KIo4oTmWVSYBs
qU/Y2fKwMPiGdjunNNKx6PGAKB9nFJ1U1E2I9weZ8nog3LTR8zuk9DIvyJyAVg4TBq/kBnYmNx92
6N7qauXis9pTKKuKCQE2+I57AIUI3rQIDA12kxpvg8U9aj/VLCQruEJA3EZktLhUGqsq4cF+p55C
nhRT62AprU2Uv/SxHaPlkwl+DUwpQmVsFmZYWfwCkL3HzLFHVnaz2Bw5ufit/zFaE8pm7cDQkxKC
Hv2XU1htBJY1cQpVifXgvlYRfM8i3t/DbG5+rDYXXz1GM9tbt2ZLw4Xo20x9VkzxQIEvTwkGn2MT
avpUa99xDfC79BP+CPkNyj9bv/f2TIUoO+pR5GrQe0hHrxvlTxh7uoamUJ/TR/unf2wIprBK6tZJ
Jj+w/BPMnuk07Rx3/TOlytOvhLBJYSoog78yn2mMOV9jnwdjUC84poueOeGbpSpcXSaa03K86EPa
xK2OE/QEoNgL+bvt8ZfUBzEFTNa4XUpfxLlhE97saYYQGrIPc4RmPTogp63qR23mmcd+9i+h8AWq
NN8DvmrVZjbcj3TsWSRYe18pHQgs0xcvh8+vvAJRmM9Cna5fvACJZIEqsGltgEEfFqJiPH7Mz2Pv
FeEdaukmlAQQn7yYRXRKv2/yjtQVHGxMrJ/IHZd6LpAdnQLoLW7EQcY7sEzufZMROPz+9OFon9XF
x+dgblghLPL1qJOw+G1N922tpujUB+P/q1nLpGZ3yU3vLnd9UmhdhMmNtLaPdqUX+8NkWigEsuZl
kmdfbFS8Y60ZP/TEntKMaAz2yFuObRl5uKLh6beHcyYXc98+I/HS+j85d3RrjLklS5uAk1vftvqX
LprvdFJKap+o1rg58eJZ7AcGEJ67MZXL+HgSuixN+7+/9EA8hYrkjRTjsL+L9XtWMQnuUp3qcG/u
n/dxbYjY9S4B8BQpDufg4I6cqUFBJsnS2hM6QZfcfDHCRJX4lBRyoPHwVMWRl6wONwazNt2Gw2l5
+VbUGgoP24v0dWkbBWFFF0yrZFvybdW0KHezbf4ha9e/bW06bthB2TeUMSo2RonU5YEeYiDgs2bC
0wCWmjwAFx+IpLCUVRy/padA7Edk6ZnNV0wSJVbX9cqWBdi1zaegdMji5Qk/9p9NnvZn+NwsrpDB
AS+Y8FZtAuiVREmumx524rjloCLzYDXHkEWoD+O/Z7YSTGcY22gRXnBy9ltvH34miQAbCLJJu8b3
5RIIjE99ReN2o5gtGRXtShbaLwSl4fbM9gYRmeruMtIrW6QUYvrvsvRe4LHJ3YJFclRehr0ZPHJl
VGs6seb7EEqHJdKdyQJTUaBfe7a7Y41HXohCVuIQcV1IvVMc/DQwTZWKcrpbZARRA+vzDhjRvbxW
0gyEa4B1i4GY2FHyrVrr+LXwoCo45Ps1mCRLXUn087KsfR5R/hqWts+QOJHCP2o4WUmKZMqtadWb
diJ3lSmhLgJWsR4jI1HwbE9uxBkUMFH7qiL7ouvQLwYH/ZF0vbZYqEGd5Kb5rr5fvmDslLQcvQOW
eXolZkiopIG7bAyV1TZdmXuFwLkv2/JRqKjML/s6MEgz8uVk2Es8jW0i5+fJR2O1wm+Pb7zlAUAt
NzaAzYwKsQWMns0Wo+XzrNMFosd1WLJp/0HdepBbxb43dH4B9xRUvLFtc9BRoPobFb3qXCar/QJS
PQPXE4cwhtxdaLXsSRLX4LUE0tZqLu8vOv4BKlAu9yuEsZ8ggAT2vrX+ehs0Lt6qasNJidYanLbx
GU57Xlv603Ad/zteoy8uTIg4ziIXcywEOrh2nS07ri0q8wY2jeb6mTiy4U5cuLCeDekh9iGqcFOS
dM0dMwembS/vYFB2wD1jIvA+X2jrC/d8dAF4zmnLBmkFfnsPYbjXUGSMKHdeJa8M4JLBvNHzhPdm
xSD2GoKataqnaxqqqtw/w/XSnJbgsblaKQr576Df1xjE8EeZpuN5vaqe7hXRfutEvvVd5BnHvegc
F8oFN8W1g4ijm1n5sACtRnLIN+TJwjZyqLB7lYgtHtTTm566L7w93g==
`protect end_protected
