-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bUfFuBqmcIVLfjjn6FduMaLeaYX7px50Ii1C/RPl6VzNMIAJneTi1QvanZXLlFhe1Uz1DiqT348l
rAd74UHltsh7nffJwM4DOeXt1VOuWPEXia++Atr2TtTgcm0gUWlKYWPrSrZYYhMWDrG+cbDGthwx
eDfsARymRzQ+0DQoqd24LH9qSTvBX7Hgq7d35W1flwdsEzzCTJOuC616+kP5RY0OxZ23rHwdDSjD
qSFYRaxAjkJMncB1qpZ5ij+IanEuUfR6Wp8DBw/iKLsXweMqbZidaHS+ECUrttGMiNQJhTByJSkd
gT4sf6abN7g5c5suDEnhiIWTO8/vo+jY5haPTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
jrfN+ZJuYhODsQTq+5xQb8d+Bou1csvN5Kt8o2CklXzgtFXsJHi4O7F61OC0PJnQR8EWyQ9pHLcB
gxZNm5zCBUBDSrzr/Yyue75EtY5a9HKWJWbQWmnHTGsNUciAuMoaDocD493FH1flShqghMguakbF
JONTk/qcJhvK0agqQtBVPf54q50ldE+6ZfWQJ71aZvXeezXytNbTpEbDkl3tBvezza+6bEsvwIt9
4NVQwxngOncb9M5U3RiUib7nvF8AcW02BmeQdOEwspQQJPZpZfMES+gJit+b7mVWLwUP+G94RfvW
Bs2LoQPZbD9YXhtemj8lxMnjWkXXrJPaxFrI4mKBLVqTHm3a6mTZdNbebm+8iiia1fCJBsBwE8LZ
QiZ5zahL8XxrakKmRyQXseW0tWz1vNrvjkDzyXFAyRgnzxhMT/cwpxyEv0m5+DCIU33nYFKj0UcE
Cdn1imIDl91fniDzAh2Fu1XV+6g+JfDX9zKGQ68KUmtBvuQaIY68rEszxPT+jVcjVfYXVqdAe07h
g6n5YSGuNWNwMsmOrPz43C1tdab5LdThIVAVZer31m/rvMEhdd4bRqGYB/0D0G8eV7cvLGhNaOiv
3h6LGUbKZD0uJzaIR0rLKNFviE5d1HYYNy+li9x81GKXpAkXYW10fyEHMVCFi4xtL2nbwlSYeZUY
ZYwK5ULjujAfbwY3yrxy7uRHcyPNQ2dRxe7ooiBpazd7MCA/ZhNG+Y6tYiYu2fIjuLMjSgOsaTQY
tN92KqRrHwo1rA3oB7K2ev3zphwngPMtmF4kqGwz/et6jRmlqCUso9q9IRR+0N1/QY1wwV/XzlKV
Al31C7V4VIBL5JNmZPFFPPw2qQ/3Oq9l3Bi4B20zCN5uuWOkGF+tzz/n901sEe0ueOeHL6y6v/vM
3FufHVzil6d38fiK3+fJX+jRXSYVi7bhJEg2e1nQ/JSbnvo9fJvJMLiKarUzLaCypUNW3Cf1vMzH
VdKUwSzLi/zIIIVk7tGK2N64CjYvuHnG47r9OXgqfgVKj6ynUt6rMRBTO9rWnfuTt0eIi7MHOvqM
Oi5Gms34qYDRIn6tUeSCYwxyDH1wDWLeM6v/b0eadwlCNWlbwAoOYxOkoi0w+ZM03vipACWYI3Pi
pEUbTs75aiJMs9RLuI0e4FDGCWtQ1M9e0/7jeU8qpTj3Qk1DKzdGE2lcq0eOvBku0O78dI/WNYG8
/d/yTatg6NiXMkmedujzvtyitrhhPzcgGDAteu5l0DPR7aH5ledx0kCYDkmu4emxgedAwy7U5jJg
mHNSHC69sA8OoGbsd77onrJ4dr3QB7hlQVQ+1JaElANmFtqJdgceJ914wdqnldV0ym1Fk4arqPnE
lR6EAmS9gEZvgqLA6RYX8srvNYN8DA4JXuA7JH7x8AgIgvmOXSUcAfP6J45vUJMM6zH0fNINvd9O
KQUNxX2HOuHCuXfnLbCnTjRG+4k/ytBiyP63Ri1GBbgtP/mcEHzuNVV20MDU4jY6zz179+ZZaaYA
hTB3/HpXFBEoPXBIrEYrVX/kbULazz25p9CaZLZK8a/H5p3DyI6MC4UrxWAQLzAdVZ9PA8KeQE6g
mbrk9UZvHLOIAAZUP/gazg7EZPWp963kGVGBbbS+MUKl2rR9XlHyAZTWb2vqM3ZQOsD73uRsC26C
TskK4G8IBSASn1x/DCGxRKOocA7o20UPuheFq0oeFedeLflSAj3CArumdezBVEgsC7n0G2YM04F8
1VtLxS+FNeaK1A75DfdhbHvHfpM3YExD1c+d1ML/QuMa8SRH0tigQ8uLwGyDobAX5Ofv0Ti8pjL7
q15dhG6tW+iCYqBJLh1YbyUS9t9KCyfXNZsuCJxZyUU/Hg7DCombHKgHY/RrqekqNMFI9j7XL7ni
BnB97YEqfnuDk55TUsl2ZSpxqjrrMABV1QQ+0lg73PCfTDkMy9OFGC9/lmTaZJfaUAQlyENu5Udn
RBDxY0QFZjj9on9tmcqvE4p0xez+B1bwkAiAgZOsy3n1GCuv2ABOJHUug609V56kug37mKI/EIhf
9n+X82W547ufi3jkMzHXEHLZgcSZsevTKaaCkmZrE5WvjGE5Qc/g9agAWUnITRwfM/ImtZZVbtOB
ifTmWm+pX5iQe+pIx5bIQkALpyTi1+tsfLnRnyLRGzthuyKNnrIIEWAr1T3x173qQG+489OUbtP3
tQesdfh0TEbwJvMwqiUZsEQ2JOBOovJZNje5MnbTvfkGsyCfihqI2b0blefFOt83GjIYwmkSNagr
KF7b7cTTW8uOjvszAizJC4/DN2YH2R3IvNHBfFOVPfYwhZlMRBxfHIcUbMPhwugI/M1ZT5alWNlp
YIxt9uU04KvX/d90J4hH7DmdWvGqNjVtUVSseMGck4MvwQ13upKi+vZ3xw/btz1dHVx+WIdQAtOJ
tMj9fTchyx3jXbdXrMcnYeofeDewqRGRTO4xQ1i1JqknNPIBK4FfgLUEVSrfPcfa6//wMr/SG9mH
Lc5N0IgIMyNJVuDcswoo1MC5WOrZhRbnh70eZEnYIWue2vLzsfLheYkIIL27WNAnplgU6WEIEG9b
P1WnxN4pAEDPj4xErjwHC0ZCpQzlPBPCE1c+S0sP7KG3EIwuXkZusnPQPBYTzGGSQ0MXCrErXMH8
ib4HDtj2mcUd08pZx+n+Ofsk9IJG1dVo/LBNl3PQ23y9PmV+R5pBmclQmgYhj/OeWNLbVLqFSJ3f
iq030vwBQOShAFFdGwXoGjeQIY+zPf04ZY0PMv0ynrqXyytPTaA0HFWhicg8Lz/7D+9sbOuwCus7
6o1bKagNcUfJ8PbxRNSPXhsSIkfVTAQf4tGKVg6ZQuQAijMLsOK8iOpHdfoSDXRhom8hoif2vICa
35YKYWb7PabGeFlGHhozgOXT5dvfNSgFlHLA4bYLi0/0kycMdBcWOKW2nZfq9svUbPdKs9ciZpv1
L/zeMmkN98aWrO3IqDve+UEpABFd5dMvicE9eHH26UXnRJhEn0yKtYJT7o3GJ/0KazWoFB56AyIM
OnRqRIV+qjJ8hVZpSGi0h2Q6d32xjYs2bnmWV27HLj1/bMbkT8T1CYbNONzu8yIOhoEzm9hEiviF
3WJBQZqiMc5IXcd0PSRgPQzkCYTOOUgTDwyGplkWXdmhftycerkS47LvOJ38AOhv10rMGJ70qWa3
pzi/QzAPc9TAWXeIlf7tR+tCud3pZA63sMStEPjufuk1l4Fa14aYTi6M3CrZQs3uyqqh2W5RbAvi
ASzBOIsfRxfzVwes3mU2kKbjdvWJSI2A/B3hhs+r9y3O1AVNHoAGzxb37b82xuPpyp2r4yhAwD9q
kT/88tbXxRqskWBeVNyC1SpQLN7u6ZQrcPOexOnB2/tNjZ0czW1UmOHW1vkEOrjxa3+PaTTj5E+D
sdzia6Hv31sWm410U8C8ORJ/PF+6nc16opMx3fY47+13jCODGV1gMue89zK4HRoKX3EirBEfDGlb
zZgEq8K80Op/FE+MOvRnjd7lV4RDOSUh8Awl9Jbg3TUMdrpXrmwFkSn750KDe2tm0FvRUnl7YvZY
oG0O5m1U9S3iB8cOREXLwqxjOHhH0LkBCGnafxc09V0sa15euq0q7+/lYn3pK3i9n8OcWLfJy97M
rxqnz624DVk+WdHQELBFuD58yVXsOb+hN6TqgD9Fsn/8lNBSABmOZkvCsQl215/5HyGuMwi+L2l5
OhXy35ed3jjSXg3mQmE5keAg8bDbcmACrDYqXUI/3UdvbWo/o07lng2G7usPT3KiqNyRpMl8aQRn
dEkf1LcT3spsYETPEuQSoaGQxfWSRfKKGvq19DDj3j0R6AJO+5Wwg/w4jUOxp82Yv2VIF2rBMo+Y
lvyPBV7A1yNLuSjp1pn2SPI55hP5lxpnJiZGt3MRkZPjRCWXjDjPJr0wyMo2/2ueCVJ+HCPvTCn7
rSoiJyQl1tDhLZWLRzpRg17FRIqCUMAiGo3+gigBgEjrFWaoc8TBBX/rFH/xuFYgNe2YHEa2Nvoh
kjg7G6zyxBOZHa5uVFSu1gMdR5y5YMfYFz/PtXYQOquaI3yH0xieffOOuDDRVPleEGONFu4uTRa1
R2wGltWWJTtL84JkKs9vbqxpipuicE0ZdTVFzMEFBqZqqaM7wcErbuP5CeM5iiq5l6/OXNrAydJi
wq4CBhEa4a8SXFp1vXiyM7Mk6mfNfuDLTUNEy+Xu0NNtv18u7i8fCguSbVqQVAEbDUUT3YR3eTxI
BrZthLqcXrpU4npJ3akvAolF9a4wGBwmsMWLDEvl1AVb82CwuLHmw9LqR9aonnRMU6ov6l2vp/jd
lq7yyj6tLpdkCTAREyaAV+u6s+oVxHLF238SWPSmRSA+Vms+nQfm/JhhyFDa+dMdU7hi0qb1sbFo
/J9VcEnpIIE6EFVzsHGFX3mdFKrZ6aACPSPuGx8w8X8WcixfQkt9kvuDQz2nNhH+w5kg4+ZQGSIv
lhS2/TSt5I1nV1t2J4KTwQ/id3jMo3FJ5EP19u89GI16+KcbdDmQPKzOIw7bxZyPn/9LIuA4lilV
d5VHN3CSWoitOqEa6T6sWrTvF4lwXt/Qzdm0MaxzCdiAsPa8FlTY5W4Ed0drRqZvgfeNSCi98G+t
mrUDbyZVLWbZuBYXkHeL/VDlFmM3+YMujG9tEy0tUZIWfWkOUTr4QQBVVZeCNoUW+mBbf7wJaKDh
KOz3vVWk7IJT+4xAyOFe7kwKyk/vxc8BjMZvxNyeNfcPPNc79qJ8m8ltx3qwBdvYlztlWOeyBkZ3
opLEqwF8dyVRR5TbJglxM9EnjieXvCzXMdjzEGejvNnmiqeVM3izJVcqcFTN3B3C0Q2wpjnEmYm4
IpkfoKBV9OCUR8BX7Xy5a/a+ed1+hyaDj4FkPhQB2qZZM4/yCVwok2wIj1kYULOoPMzguGAqaMFm
vKtIRk9+MWNvqWYGgmXdgfLH2xm/CD0F4j1iVxxNEsi+lEkcasnnZ3yJG/5t2+POgvjZpXn5siK9
nLMS8V7GZRGzrc02v1RGj64yfQq/V/DYoVHwjFWjxP+Ct/BIVRG4vsAl+csVCpCRYb7fbbZl6uhq
3zWh8j2nHPvUe64zZ+EvWP0TdrXuFelEeHEI1eSV5TOeOOgMkuxO6Ew+zR0nsWonxwoiWWTnyEqN
VyRr+hX7qUNZz73AIZMiYgYA9kaJXvXakjORe4rai3h6LRWwsndAFqxnyKNVcbLmLd9kuIlCADFb
POxYtzP3dY1RVJ4RtDixLZEhGK/Cwfa2X19MlHDYJ5t+DE90gwknwK6ZTV9EJZupCati68MRvZkb
KMnKVAk/mHumaj0Gh5N7hqGM1oIWrcJD7OvTwxNPTGNK8vjZ5k2vQuUCj0VzOCIitgOvz3wJYsK+
duWK+/91FascDA8Ynzp/+jiZnK6FFoWtF/oyKmRBVvth3WLriGCC/tJJXjG/wZ5Mso8Iy71/JKdV
vrRH1QeoviXPokdcwzkio7XM3tF1RV0ZFghPYxUjq8wX/m5zCRWMR2u7B4VSsRnEYdah90g9YAbB
ARgRGE/4sBOVx+OzNaI5rNQXPjfGT4zwxa7M34MKY+y8KM+REIwn7kqHqaZPbf/kwoyi+QaJ4oxo
AK0gvNkvd01BAmGCT+Z8tz5akDJdNO7VczBZbxVVRaNJ74yvILP5rxINWUxWgsmoOvJldD6CTXxp
m4vWQEo3aXuBPS7Dv7ZwX6k0NEwxuwdXWlh+/A9d29hg642Oi8lRAg0DxhYMNYzQ4ylgEs5keX8J
En1yNtplmDnPdyAaDT09lfausu9j4kB9b3ojMs+jYrNzaWn2WoHPgMRezBq9cONM9VUwvg32vgap
SM/KBqcC7yBmCzOKVba2oni1akhcj7f3lO+TLxNQa2dbI8BceQgi4Lt0QE76rjdCvbrTGdaRqP7r
0b8jzXZdjbPUTkdiBTNP9WE8DK2bIxZnXr5koSAl4wrzIi+H3dapRlIt7N8g7Ki5D5hBlrki9Qrg
7/PhKGzZeyDmKB16ztZwZXjHCEIiQ6vAVTPQtVojC1l+g51q9T30XaoXmtVOX227cmooP3RWMPhh
lfFe3n029/uMYHP05pICfO4aIwBHs/biYohnhyNhoKVwjnsU9M1LWu9/N+FzMeAro5kn17U+ZrVz
EifTRt2JBzb3zN+6vIe7XbxgA+DmoZW8uvHkevaZLsHd058dwmbRDaEECkDtFHGKzdR5q3niQhkT
SuAijxn/+nv5fwOluDmFg6VkSLytUwWdG2HnGsCd+EPrxfwCz6l3rx9kXOLjsok2OBr/JqKxkAV4
LLV5HpmxlWWqIHHLEmWHBCnLrbjqrN/V7mrvLWCO5NVpLKbh1EcTbHqzLvb/PwscQ5uUYGgGOASd
YMK+k4hvVnKfvRSQv4VQoSPuyJoLt0l+pdzUUOVA8w8b5AzZ4pzmgMcpPDfggE+Ybg72zRYpgp74
hklqIbUejE4rc94wOSJYDF1GyC6bPX2E01wCMN/k3YYAWYxom4n8VjYA80YDali68kIZZf7Zd0yh
GqlDjR9rk13S23sDo4BG4/NaIlyT28YdDaYz/HQobyk9OGGyNOKRVkVmKxF+x+LsZRgky03AVieK
9E2ekD7iPODwRGXA02k74OJkpMK6bwclm0slynb0JG3BAEwhW/0rIUVrbGlO4ZIC4KBDNnADJuUL
MwHSvX1G5Gp8CQbP7uJ23kwMXZFq2N6c007UVgHpS0e/BJnJIjZWa5S3EhPUO45dssf7nXFyZP7E
1EUvdVF3f7ENHtYfKRz727Ud2pSNl5UXLY7Tb1nhOiuJwlqmphQbwfsqjmTshRqoljOKNm+cWQz/
NLfPCzVxGyT7YutF6hsrgOowdbODqf4YwUFm07vmw2x3N9AGGJNkF70wYdNt1OYPtwKG9grerawV
COB5kAzqx7SdWuSACTb2g3r9++00F7lELXi2Exgaxh8GPZtd5sK89dA72W4AEKE5u7wQE4o0Qa3A
aTp6Ttm92AkayYrcvyixLboiZvcP7e4DBcHFcT+MqGk0vNv0G4EHJNZ2Ac930CVl7W+A9CfSHnBu
06Y5koLTzkGNcNMB7L6MiXvbx454HsqwWPApkFufByFlMfc8VQcFHzaBi901ZfuXP+IHt/I1Jl9I
zbVkwPwYFa3IqtDl6yVNkePJ9N7cqgH87O4Ob4v9QKKf8v6Yo3gktyOfAizint45A+AQGsBsruGX
60gMnXLSOuOOjXumHRLGFP+o6oGPoieSPeIcYAsvcx00QeF3Rd4IX8DFE/Ltn0VVWraEM3B56HlP
gu3dqHKrYZFLf3qeN36Xl1A8EmWzeWPYkPJXuMAhMAu3GuKE2mERvpJ82XnHx+RT00uXLLrtKG9B
cKtUA+C3BO3Vd42MlDi2zVqbSjfU40jsTE2MQGwPd6l4q8SFKfrIRdILNQW6hJpbkC3XauuoEwUN
fAF+abLwrUK70I5a8GPQBquIx+SxmvN51KvFbRSXRZ8wzlSoNsXjtWsQuBXGGB4EH3XHm+1IiJU5
PbJk1PaaXVsnw5YQK/1flT9dACuTFXsGOjQehX2wCiDhrVo5QdV5/IWCvMBaJrb9GmYSMKxLJWC3
X9gRdG/+ZeZvy4m/oDIiyomZyig1phCT6c4XEEOdOMNL1Rni0+k8wkmhrsCoxSfAJhlywWa3Nh0y
PsqrDMi4/bmQDMpG4kclgNnRJVwT71dp0WVsZmxZcUVmNdArw7lT5YhVdZHKZXPrRKMO6rrjHwau
E02LznDqnpRPQ6nJvFJYSLr/Azo8c206yPbgVg42TIS26qpqVHTSU+DxDs6KhL/8ujYr2+u9lg93
LswdAZZ1NtBjDvfcmeibU6U6wzbqExdZ58Wjxq2gFiaBPr5IeG16L9ZmLfQR0tpge/14KArooii3
KS8VJc5jE15YM2aITZPg3PikWvSvGCaWBSluLn7C0wBxrpbqOy2QkctskzN6towk9eLKFebvbF6P
efeVjtcLa0+SKzPvHChxCIqnsgMFHx9w2Hck7IS8TolqvftnyqayMwnZpXwDw1sNtgiv2FKjk+35
469dcNpLOt08d/M732utBiKezthn+ZcCLrhQOl26kHPu47slS0gASmHzpsJI43hXHe+5yENoWAY8
skq+M3LI8+w3xuBfu6VasNBSvv8/xN7DC/ynb54gozjqCd6ycOP5YX0BPlOpjiUtVQNAc6VFSS5F
Qpi3GiwR5hC6En+eRzxmzomJTaPDryoPcRRybRCyFk1E5vTsmEBo+RscSN5rcpMoKtDikS/o3wmJ
+HGoJz7q/ga6k+DAJhUoDGvTvXT1t7axzQf7sw3ZehL6xDgxH3uwSQHcZJEHxP7tJ5R5qLP4SMlx
tejgc3YkpI4WbvWys702o8xMuqbLUUDm8HLJlzMsFEQYoDBCBw+LxU+OtdRxVn0afHrXkrgqAZcS
LZw7tho8579q++dixhqFdd+SEKuvsywSWwK3gelKIVNscCeU92E7PNe7jXCJ62ZiU7QT4lv5KHBQ
VXDp4tkiTTsl+PwG3/RPwamlnik3f8pG8nLubZrG/i+pEOFnP47QhkgBkh9h3ihFh6nkGe5Cqe29
MVZgRnuMn8BiNz9dmbZlbCRoMurx6RTwcengUoW44IIbjOBLpC0XjyQoDjHJ1hw51vB5SLsqJoio
vijWyp2uVYzop05lb0sjXzrLF01ixYHrYPthP3DHUi20eGhw4H0hBxYtjVRj+URDiur+wfOsJNW9
4nh1C/8KXD7lFqvFDQP7fZRHUucgDqz+0CrxlP62hSL0/CoF3DInb82Rd9w12D10De/P+/pLELO1
8o8z2szHH85IVGAL05LkuTYBfpXHodKb8Kphb2uXnFnaFh/y0Ly/eqTK1M/FveVhaj5enp2ogSvs
M06T1f/UjmNKlvkEJo9AiHb7cHtCRUvCYqtrzWq0QWSu4KnaL8HEz5yoJexROWinkUbgvy94Hedr
pHMbgFe1bulZlJL1aBLxNXGS8iz0HrrsyDBexBbe33trEPN+qShKLdhqMhI/DkreIX16RN5z7ZUO
ZLLhoZUS6AhXN3hx2Zhzhsj3Guta0J0TzNqAVs8Hk5H3R+hTMe01bzPByIUTux8HaTfLNKaFbnAy
s53q7qsghda9Qn7zbG8EdEzTNmdQtagCF6tUjgAa6+cdrMET5fxANe5Lemi71rPqYYzQX2NIy172
vz+cPoV98OWkVn20hdfqpmROFad4jgNynP5wX4ne67zDjZ/V+cb18PQQsh2QP+952fRlPEwExGZv
Y1L2tp8a+R7e87OXe2QdnjYCE1klWql70B62LeoJcSXooa6ZfDJnCk6Zc36dP5FWyaTu/4W25ppi
MM/kL83AllV3Vn9jQfocgm/5eoQ01mvV+6eX3q0BwTK8QUjtTWvON1SaLNSr3ZssWi6Q1uZ4yEEG
/RoLb3sqdkO2O8/Kr3IArLhGo8H9jksERQ6JC17uEJt5UyRdQKCt0IIGqfTJhzvT8daQ23uOsZq4
ccvRVKXB1UWIbwvs3fTPDFSLA+FKZJXlnSrB3U9qRN1MMCCs+eOONLbAoGFsDtzuqNKa6UN+EMJf
1/NZnfxeS3+xNJqurkfcHrZIsbUlLwReRyGYkNBU9+qnyieBYJ6faCWXLUyo9CPITjlgWZRsCFfo
Ka2CqYTKTmsQBKaxbsGiQPtgCZPgnBwp/nurlzah1J1QyyHCB7Cqbc9TwoiAiny5umF9tE9Ux55i
82n8QzXzwgJR6mfc3EascOS+etS6uhdq/grHx7qAGXPts2sp9+NODW5jmij5uBzUwK2YUA6EUn40
n//21dfJ88EEUAb9ZKYlAnFrXc08+RZrd+ESrP+kQtcjlq7E+aLw9pM+NmneIQAayrJG5XPak8v+
AFaVwcwY3j8WPPkgE1gnR3l5Ga6yiKDdE8n+wjyXolzLG5deq+n8qTfP5Mi1gDwl7N/NyZFm2ZbM
lQ1zjE+R9Vi8hrA5I0q2h5OBBDpHl6yznqfxMLgspiSkeM6ZvrvQzrLaegdVizuEShT2kntgan0n
gFPIjiZixSThjsCTFCDIZ5yKDh8XAMngYkFo9hbqzr4zQ0XL+fGFzAVh4uAAgl4wdclw425NMkTN
5ni0b6fLJr6/vaEisGYQxAyFRgbE5IPysFDvC9/8QhJR38EoUD73W07f7hGmfRwlmvIaZi3Exa4S
eTWC5ZPp5M5yiyCxu7KXytFEb0jChh+AADxdozpzZ2HKSYX4oHjiYs9nShRPUk7mDjrAkNuxPv8/
k9TFEphvf6fAuIbgFTm9it2Xg46y+Gz2LlzYo4UR/w3cBYMfjiaKc+U6QhLpIvfZV9d4p23pKGZW
2EGt2Lr7aCh/MpNKZisiDyj1kSKm4i7cSC7EltBn7sOGf0uFk2BhUhLudis/sz/ey0EX/RvCmxQk
MojlqgykZxG/D767iAoo+FlJiHxy3mzhwYIKp1gzUPcp0wfUjCGaITmxxrHDjLdfHIuU3tH4YYkL
AT2G+Pb4IicNc+tyKYSKw5bmQzAnqGQ1L5TrXTsQHXK8GPvnP8ehe8WfwnA3Zo1ud41tnaFoWvwV
WQwgXv5krHfi3H7W2FsCNWq4MpMzxdvRMh1ad5UW7CnxDuonWMhlvZ9jt7l3hal94rZ5CnaxY0tH
Pz5zXjGwSe9oyt1OzR5KiW8vllFCcxhGLSPGtdyVRW6O4TFX/oMfmkXR1DrLQMnRo1BczPaNjwN8
DCuxzYLF9gvhvJqBK1nedNyW1f3/oHxpRUv2GMVXxcgxc338HcVLaiCHXFdpk6Lc/0clrMNjv++o
bRJ9y7nrKAoBTkf410v8+hmyNabqJGP5WsKbZ40S1TWPqnUBsgNCNFWiF/Z648phck6o7iJm+FSP
MnbrcEK7oFHPWDjzbbzCwrtWGcVF/eTC8a5wECEYqh37aReAP+zB82tj/NO7IsAZ5XIVKdRPTMvC
L9HtGOA39A93aCZ0OFCcga4d78exGeGWvBf3L98iXShn6ji4OX0Ie8x2fmbb/UnOV594AKklcQV4
79mBjXeLYITbXwOAKvJu1rsz1AT33V5UWC8S313leZ4a8/28MDLibnWHzCS2Yl/rwzeGuLE00RIM
+L7zBEwzjIOSZoZSz8AFrTmKFot7ILd5dRCW4X5HO7rDsL4pF/FCBzEqVoy5ZlPe7cbq5yeHZ9ov
iYYaoi5IQ8HKBFo4LZWN7PHYwna1+7doxnCL71qFWsMX+twYMmgLcbI7PlipvCp8QbTAY1S34M1H
Gg3m1LsnyO85SxwraYSCvghRz2HlIrc3NjY1aPEVThaK0p/6N/DPr1L4traeUbQdi/BMzVf/0oZE
eghHnFI+dgu/6hV0OeqKA0HCE6icYhJVmJoW5uN/RN7FAuSA8oOBXGUn0PTXuZzdXoHtDsuiSDE1
YGjyGFYklbLzVZwoQ0CO6Zz3rl/nd1f/R7I+1O/npWYB4NwkzRLrEiyA4eRgdZWD7aCi/9zel5V1
nRE1FUZTxjMbKu9b4VEC8fceEEywKKvjgGMQHYl5exUkHEHBx09XRMmQzNKTdM1IbNt74/jeHbLy
dHeL5jwMJjmRpzbqPTjA/LFak98uCvgEVMueNwsL2t8+bqqZy6fyGiX4/oHqqacGGb9guEZg56jt
CmM8NQwlKSHap9x/m/w20IhA9iF3cwV8mPYIKVsdZGRKabkcGmUhE529ZlAr2ZuT1SxfW+MO5vLM
m4KpwRTvJbDgIql373zN2/MmaOu2gYtGbQfHibwo/r3dOZiy3qiAvl1yVBptQnrY+8aouKKoIZXj
sHjClbJHpsdAcppttn2Ywh6rgIw5PWg5NFbzPq7Jsn6zkOGzJG0UTT0/4Qgf+d5y2T4eyvOpmfaq
8dXIQ11Z6p0WX5pBQL/uS24Cumx4hlce+siucM046V7g1W99dxPz9gssLsZefPLe09qIxOX6BOa/
ADMn8yAhPNPw7SVxXjbGmTa4Fw1tvbCsHVsoGYBvYT3iWifppOO1gprDuJloM0oLQmzkpGWzU3cV
z4etx3RMx/I+KY/lcZpy5ofA+p00yVALB2VIF+ymrBi8uUQOCLE6QJ4y8mW6dkOLR4g8aNt4moUk
jP41ko553rsaIzQ6J771FxhoSFX7HomuUQDzKQzS4uG41wsSuOJKRXiI2wK3rg+vGqiv+FYHiRZC
7k672/5A6u9HjIZpu/zvHzv01Pu2TVqWW9ZLQF77YzKLIejTGMqjtEGbWg6kseLimxsVFpJkFDFq
D0GVoHFilcm4ozAbhFdbMuRPOohm05leSkssIhoYYIg3RAtYXjkddjdteppGjxJMsCW9hgyi2Gdr
GnOYpNFtfbnyOwvEj8T29SkjTuOKfeFqzrafwcIpXoqSvP+rBDd8NbS1RjG8UC1pFAuMI5AXZKYT
3c/JNs8jBmmyTGhV/OS2elrtY5QcQ3LObqDjYETfXrSY9MoBiZcwMjLnIwNmBxj5ujPiDMBQgrGm
c4FxO/uHsUheX8Ijw8rlCupA27vH0QEsL2FUuP+QNqv4nic0JPiVJwX9j2EsvODArH/7la8rzW4S
O80PMdq6isbiSQN2/NWcJ2yH7pHKynhnrs5vg0U8v47YHbfVz7+27ZMGaAtDruXkbeG4wQdzGGVa
WGA1eyf2kG8ts9/cgQCBZGVvJOJHu+w+bNcwqPac6GUH6aWkOmTegPTisCrDxf+Ctq5Ok+VQDtxf
i8Sxo8M8zN3shTnwxdyXuns7qrYLtDiMNuyN+tBsTfGQdt9xmNzvvxePk8eT9hK1hwCfZdEqqolP
D2Xbx3uMpGm5FWjVhM6rHQP4Xih1zlBOQ6jduX0HT7RgVtPI3YnA6zfHrvp7l/A1TUJ6NVdkZ5zt
AfhwxOsu1/pSzl/fB8xdaCqhKp7Fj/qCkDeAndfLANpH6XqqYypyaRedm545NIeF88GoMEq4a3e0
ka37DeTbThxwGJnivYsUYH1f3fJLqGGu43yMwr49lZROIsQya9rd7eeHburSWpPmM6DDFyMzWw5S
y8jt+pkFcTmcsqt09GaUzDOv8d74mY3xQhzl027iCB76NINWttSgY7dfbzM6KmXeiKy7lo61ZYRB
qUPRWKuEUV8AZUcP5ySbAxIzXhVe0AiQ1Ti+het18InLVGDlXHw7QxIe1/XwZEsQ9Q68TBhT3Hti
enn/Z6K5hSY+qMaiA0pBu0iNgXQ6HYRXl7sFOAg+hudoo3xeJQE7tCcNihC0KMYEJQRxYT9TouWt
wc5azUbNkvFlesYWtrsh58gewUNjdSDg0na8+k+/vnSq7SzZMH8L9mavHOcuMS0o6Ujdtb1k0MB1
x2QtLxGcwKj7sn5g+XM1xuJ9adCL23vcoeJsUtTeVQgIGlHr5Oa3VJ3e0nP+dV54OPa+11kBJZXU
E5sWrWgJtSUa9Hm1eavf2edkRw5WMvEXIWv8xWpjMwQz8HHQmOUcuj4rUcGUs533QdB3hOzKulP/
e3vab0rOMB6FyxDDH/qgdpVXq8U4VFdjeHaW2w+Gu6U6765kNzqgvnHYwS7OdLFkFZwvYv8T6cJs
Zcve2abuzXuG7BWUoZR3ql4Ln99l99ZSGuLKYeKhjYh4N6kbCkcqdrwayATbOexMjbZ2U3JsI39e
n5TyD+dW8fmp+tsgHrV9bh4UMH1GTCs+hysEyQY6fBOFB0tjvvCNr4pHY5XLggDT18xCSb3yyIgX
IyhU+ZKMoYmY9zG7qUKw4fnhoY94N7nNriI5m8+2iSyggqJovj12wCHqaKIyGCiBlm7WYSPTA1Se
Uw5hze0PTZSR27Kj1yimAUOIzGGigzcr9pDLxVWWTtJ8gFUI+sQ1t+dGpte++B+LNWXYyR2/CCjn
no9YpL0Lp6n56BQ4mjOIqNsyUkBUJgFpSEwxclLC9zuyglKWyU6LK1YIeSEzTlpWaJWJjGrGTMPv
089z1VQzkIPtCUDgf3YwKSqFbSt+omYc9ZJGJ3EgHzuFdMwS8KXjh46V15nRg5nOc6ciLIq0PY9C
4egoeSOWHP/hrSSjOrpS5d621mTgpdlipptYg2NkrGW6KtB7Qd+eht0xIhLAFlbHkXAK1ndq8mdh
BwwPtuuEutrb9/4oi+MwqgsYJ3wZoTq9xwGrBRbLtZ8Tqi+339i1ruyk+KGQqGbF0lFiMnfnv50c
Hu71nqsW63RBWi1hXs9B8C9N8XH2IY0OtGkHPef7C94ZEx7JSqMcy9OiXbxCeqNNmKOAiOjDTG6z
9VshyfVlksn5whzVjP++pvZc0zTz+yAvLPymK4ADs6aGYFsVTKqdsM+rKPLUkXvJhUUWEac/7G1Q
zp/7eyO5p8ZArDokij0WfsdZ4hCgxqexBb7JRZcU+gCdOfULEUJq0FrcTWgGupVlTbQ9U6QKp9lK
Rjnz/UBT0YNobdyqBerUpxjlF8uy2bdYk+Ur9Fr7Kgrh77POA62UvMec6BWfYcNoz2t1GaCpaVwP
RjhirD0IkjBmYz6IHWn8ojU++z3oINHLsvuXBCb7p99Y9LMypdJBIkInaFPFVkHdppv6CZ3nGyFy
z+zGLMAp/suNEwFk/UYbIP42NZL0FloufTjaoaAhv5w/gPvHmioUW214yXiRgCOCOaVc6WH38As3
56qWDTQOJ51vULQlAk84GBx0YOaXkYe4Ip2mUA2HBs0qM4Z1aHK/l8SCs4GZwu/lNSFlLgXLkgdX
2eVozq5/gY95rAPZEWyXLpykOqpG/ruAlYGDt30bMplk8rYAo8Vt9azBY2r2G5I8hcdRVx/wswUL
/w4QzMPkNNblXhP7kAj1789gn7naNPB288WqdrXNANOvh3DiuFvdTXQ7FK9FPM0IE+mYmxPHGLDh
+5w6HH1OhTLjb4yqVh0SWT/IB8phD8oMnNvSl9PA+GU5M3cRy97p6555pd+EAsnO8Fia5L5iqPWz
l94lLEKwy5dzU+PkBsLoCMnz4vr9tiror5NpcksOnNE9G/Urovmp033BT/ms4OccoCCqUFHnJbcy
ek05BIFyKj1l0hWeCnt54zmMoHu6IniW6YnDiDae9dzQYWS0lu7FjHGn2Tdlrktgxwi7vA3turn/
OxO0gzMR9Z019vzluLP/JbOqBSB+ZBTsbziYgW4oIzFwAHxriEc/g1PdXAdbGa6nucNxH+LaSwae
+UYFeZQZeIsXgwVQZxU2xyrcww8mvWCY39cwaH/p2ODaguTHO0rFlzpM0gKqQB/empMcth7pUwxu
CrVbnPDXbQ9IxxqB5ePFcLqnOhAsAhtTplmQajh/EoTkh1s1pEpJ4w1UVPWFx5xoBYNvCwHo5Ydd
eLPUYV00R0DDcOEgtGauAaNFTFvJ39jOzmI54tAcNEPBkutE4k8UkooSCzchrvm4Z1TbHa+3QCz9
8gYcD2W0jT+dLADO1CUhnAhqUE1VOb9OFKJGDHo93np6a+BwmXrzla96fZhpKmHaA/3uKWvj4qCV
siyneIDnil7OE+4cOfreMDC3I8njaoR9RNhKJxY7WVQNiqfuv6SKRFGKX2ymgYqWFd3Qhn7UM1T8
oc5xJJ9E8OhguevbKCNoGcBdo8tyUV5ebrRd5uB6NZQlzE/qDZE8Mypl3zNB2wVcI+pNB1/X+qmo
WariyI6jxCror4y/P1jibkmz2p+cv8PtHAOud2C4yQsHz2tZpy6dTcLWn7rG+0P5YAcHc5WufPy/
gfVSfeq0xTeQqfbmFgzPllVA6ttID+OYHg3NhG/ZWCG++RFHESfu8sMGjNPJbdkKLn23lynItxrG
Xjj/Om325qqcfAC2gXNMhpbBEtefltmCDHRz45Qo+SwgBU4K1Vf6iWZ68+cQXiN6PMjGLbIhh8kN
ym2iMmgaXfvITYPHqYglItz01NIQkhVNzE28gKFqQNDd/Ps5jr1hz/QiigLcWgCFIjzOtZgfgRXq
RclaIpzW2GU9W03tr9D/qad030M0Uf2u/KHlPwjPzgtfU91PiCTE7hKYbYtRnF2L3vOVaifrbPLj
eDvJdIzGEs7FsjgRIzjV0cwxANV5+FG37wxNCxgD+fdK4tkEyreeoUSjCmhnO0Jm2UlqsbTZSNlr
6OO4xHbF+RK8/arnd2KcPgVkZtYFtfXfjATw/rQe7fqQ+tJl+54nBYR41omXXj91GCYonOTO4MaA
G9UKuadm+EpWyaE1dWbPLa/iyDQvVF1VTBChpgy0mXcip+yeHqXML9wQqivOCN6naUPkALaQSWLJ
VjjLc390Ppq+NyfmWQc00Gp3DBhZjv4/QQ44eR7yhBISpIF2FS6mliJMc+KTK3KwtOVHqoGLJ0Zp
rfBEv9prrVTawrPTAxtdC6D5up3fi2mex2GL1BRv5kxXJlQp8MT5NBElkivLkiZPWUpDygn6KMHx
s7fqKPnWZVO+zYjA64G/bGCc/2ZcuLtTy+tET5qStjUuVfMFmSNXFGNuYG4CDXpShe2NMclduv0k
N/Q893Zx8HpDuIUnAVJSpNwBO4U3FO7vITHs46uOzMRnOwIrhFhBlqsfZPCNdAjNrtfKgQDValBP
ordAiUBOX3HdbGqMScTpYYaolf5i7IQrHM0x9UHskA==
`protect end_protected
