-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZG4xfU9PhjJrPzcXafsujp8Q+3i5Ke6WF05GDM/5Pc1rnY81IduQGq3ExkPLEpP+nuiTqJBxUkyz
l7/ZDFgxd60etJ2QmlkvzIoYOLo/9H/v6a89Od6tf1XeCb1+nPqIRnJ7lDdPKMS4VW74/FjXo8KF
vN05fsjlXUa9aGIGXT5noMDyxW13SyFVCNCQajZSNm50IezijhjONZ4Q4YE9zpFR3DBK32+9fFYE
VbGRw05NNJOXffHEEcymmnCt+3bs5BhkdRWVajyJ2YeZv9cOJZc5wCp5pg3CUrjehbk/xrSBIfTc
aCfewCv2V7RdwJyNAsgncaPYci0sKCnaZ5dgHA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4688)
`protect data_block
oY6jAqR42Yx0EkF/rhfoM/07Ja1K6qJQfa443CiZmQKCqlPKPXWI+EmlYgzFh4RExvmFzHICtYHX
21ahrWtfR1wx0f+JxMEaPGo6BIDXN931i1KuFq7za/inHka0GtNYGIl7kUlqN/YFSOT/gpZMsysG
3kB5kSmwJmbr6ySa8tzAonAsiz6N/NMRJGVnBDAM4KjYf/cI9aXiJZ2K6yAgmKQ36vhmBIX0ZY1R
bQnPFAf4LbcXGViHww+aLP00+wLNbcHCcOZ1yZji23GD5EHHafS5rGULKFIW5QSAaRm00dz6/+4c
Af+uQ5J7Z1bLvVZuWi1kiykSA6vQZmXfiP2WJzbT5d4QvaoDqgfIpEXIsEPis2CV366DFHoxtgGs
YB8zIlUxSO2dRfjHBHJpanTPn8ZwNZ1k3XxnVidseg/azFBX6fbkAamDGVY1MNArympu8AodX7tV
VjN/bktWTyvjiQYBCPge7qHltjSB91vG5WOvW6Ky4HjEwhJIF4T1U5wJMGgzCZGK0H5a7GnrxmLI
Fq5pUQV3gdkCKT05pXB1M0gNFl3tX7eQcpwMA3krqAsme1soybbYJABUrVdxN3t9ByKTF9CexAuZ
cXMz2vlxOt6VEI116QdO22SvUl/kVQq++nke2ueC0+230B2oiO614eYspi5xNDhf+zl+EvOvGApM
TGOahsg/9mDB8Tb3oCplpoLlZoI7yca6ZdSydYz2DnIwLLP6ypzYH0/HHyq5fKN2qcr1lxJ3DC5O
kohlmxn6Gfv1lps/bftqiDJfjgPOki2mlshRxl+Q/Lbx7NpCYeqMksi6vzFCsNF/+IFhXD+CnvER
1NqqoyiE6OCwzUCzIAneaGv8RF86NSLUDcfkvKTxrYmiKz6/MdtRo7J/s51h1PNqV98XuvQOHRTk
0/q6xKi/GwkGMQfC/2bUlfo7oTcwmcFEDBJ1nd4E0EjyEVHnkG8hCzugdcY2KyiCBdYxKpqAu4wl
19u4JOXjQtps2h/s+piYS/6zZgBxbKXc9XrekC9OjqB4FRpD+5EvUlPCUI/XaXAr9jlYBHPd39rJ
7P8GztY9XGNeFVL8mX6JnCwzyKpz1oczI9JlcB78L7uW/ZIEPTHWowcoTxoofjji/A8ZXf4ljHgI
iDRGTVQ3Xpd1CJYYMuMmvaR7xlI56EBlvQKPNN7BTsYDm1RxGUE0gYnZIRrQOPvCJRcn6cqsSB/J
rkkCmcsILME949pst3+IRBvaTcJ4u4jxpDrFnT4+V3lq6aWfaJtc/5sz5i/8ijiTMObVP+WCPicS
FDZNzvnrtf72lOjHAx87DqAKtuuhySAYeFTfVbFCQIGzLV/ZL/gqOwztMDIZ3+p+lu8s0td3aNzM
+LuA5/WCe6PvZ58g+TSIMNbwbfD/dOzt5uzkaMq9qpV/5sqcpQHZJrNM6Re2I9KrDilSpFUYWMf3
PgohEt95bf0HYWhJpl+6hiy3irUV9H1hS73gKGQVtoBd8qGFeyrxakShSPHwRQHiL6eWWABM55Nc
RorD2F4jMncvFjR6ptT1RrAI+tJcA/UFR5lT29ts+cyctmqF4NTn0jvqkk2w0P3kPCpGaNmunq9U
OkRpS49iki54+xJhqCE56zWgb5WAEXOjOUlRRixgBo3KV1TEKUuocNmBkgnJx4xIHN/uef7hiOEn
HLLYasXUZlqV0d12sIjJA5CQCRhQ35jBr5ZaVIUbEfB8LKUyxoCW4yRFhhKu0UJwgI7IMon2vWYf
TsmZJXMsaDoDC2Mgr2a3+0XpfELviEppOOW7YGKJ7b+A0IVR39IWHWars9d2Hfw3PleO+hd2g6u8
fkUv+JtAbOSCFDTZt42cLdtRJt45LfGy5ObLSR1s9jTCw43wpVjC0VYQ7yyUITpdDBjpXb6y9HMU
hN/MU9mzcEBWH/thCcj+r6obvSoIkz8nHL2Vkn6DD8PkNOwWvagEOKtzhAB+ms7dftQgPt3kHPsA
zlbOKikdGXDEWL1MZMxtzcb6xKSfTBRxwwHjc2PA+ZG0OYxZuvmSXuNXdSpNDDRKOLis+NmjOmPa
GR3PHF0G8PNFl4YYBulilXVsBJaHmRqO9BgHn6EOkoCk04spC8PI/K86u9rV/8WUhl5wWhpbOydL
5DP9R+kIyNJFnbFT/VycHncIyGqIblMAb/38Ao8KtQGAfgJzogkfNc06httmc/1CBHh09jqKeflv
BAF1CQ+Mm4hKlaDQ1x9xs2raOs7IJQro/gwCP+wpJ9b1MI9sA1KyK+irsJJVGZ1Vlwb20KnzV5Oo
2XGbm8dTgM4o6QZmIhs6k6bgHFjPLYfvEyLKYyo704GqDVtXyxVd9KHTlYtas2E007+bw/IL+AIb
Wiqgb2OWneI1A8H56XQpau9ALl96pPqZrHVOurrFsAOXBmwM6BVQEA9oIlihGyg72ZndOzALccSX
PZlqOR5qfYeLEgyI8FLdYRCfL482eY64A5+8gnnnpc2hs2GJ5sjJ1lsAYxehtv2tjz6JwkiDMMcx
Vx2qG8XJQfB4tUv3YAFhZAsxnkfS8n50OPprEzA13LxKNe8RXEVwgEtcjlWQwU7Pa5Ffgu/75bkI
4HXeknDzAWr1/Gpr6QiIvl0+ygTBr1ajzUkRsuEycAfnWNd1acCdCQV+oC/WNfkJN1pIbjK9dHOb
41Ce2+kGQogBhutkDqAcx+AnpXcDWQ4+RrdcRB1YRephhQxlJ0roHlGqk3YYaSviZoUMO6z+KvjM
SZvFoio/9dVr5Lar7I60vDv2v8kn1eV2hv76djINV+c6kxeTonp9/psopf54dRzGViI8G0Hrx5ct
CoGOjZFF5s+7tsubRG7YRtQHarCvs8ntCItCzr5OVtRsWqI5kxd/jfGUMZPH9biSWdnYRQ5JHPbl
mxBiof9euMAeDkwbd/DMgbc94HiowbGTszCLajX2Q44/gxTXPAWxgHxrfpzeTevep9eM2Uwlo4Av
QqTKFKcifmtGdHA3cKwRq2iGvrGVcCKIFuunWdROm2+BrfDyJUjRkI7otFs+3Kvzd7hyY7rpHh39
GWk9R16+R4beSc8HJCAbjzD9JUGkDaOsvBWlO3Jm6kujQTE4EyujZkQjVa0jsEbW0IuRNqvSbTDc
elKIyubhMtZNwDcpPtwTpGGCEV+vcksNGgICvZu6FzXlugqIW1zfVBXMvtRAJHL7OEQM2uaG03Re
+rxbYhuh/ngFttKr1LpXDLoFo91iXOGUmlANb5M+OudeHEMGKcBrx7oZocvNHtFUMqVoEz8sb3gF
C+qOPoXntizpcbp9WFKSNnJizWs2j6ht92PNJWaKOgTVjD2Dw9YDTyr+DFNwGVf+tr69tK5uedbX
BsmdSGUBRBp26TLsnG3KEXPDLTnzafKAc2n3e8Lvc1vGlEOCohjQ8SOm3fhB9s5IWgE2N73zonxz
iFUIEjDDPiDOksNjIKvwp3mu/yC8RnmtUyD8FgcX0zNOMP9NqolEA5gGWtcKYsB+wBVQPEURz/Og
4Ed68iCUu0hxzYkD7gkqWnVEE67ZZVCXWe0J/nuMAFhotmvizY1ZrK1E7wJNhgaabwKpK/wLTk84
ncgmgcGgP5UE8S3DLdJKXh8YQFFfulu3W1vyi/G1xD5SJeXTmKvIk65S3T47nlUpFysv1jmzMhDu
bCecQcd0ucqT2IjrxqAZrv4gK7ndZKYg3gabW8rcaqFb3/HAGcZJGJJ/MD1dZnAVPQemwI8G5S01
zViXyFJQJwQJMphk1D+IArT1SaLmK8gnOtE6HtNE+i8EFsJJuAvI7WknTyf83HRnaiVQttN+pAUt
p310q86RZ9lfOuIhLDd6Rkv2UrDRFzobL394LGBvG49AWc3U6hrYYPT+kkkbnr1FL8D+obGi2+Bc
VulE8sKzC8aTQBg7aAFMNIMCNhtAYIkTFeYVxA/g/p0uB7gJTMQjWzzSyHeXoPI2GukyFrVLgKL9
S4wtdQHrBALkLtL07I59rIQbZtG656STNqbsaHrZcZ48a1inGKYjQ6bfL7M9/DdSoeM895TGtwY1
i3I/5DeGcVQIjUu++yJrCFNp5XgtgpeF4z9gQ6X2jjPDO2zR6nIEWwZ0gMxsIvnFkBfF6QGXH7Le
LblEog363G4BspCCVLiDnvrciivIhMk+ZGoTaNgWqpcRNLM4Ejf49pQ4J9SZi939AWL0Y9wItS3G
LGfBR2Q9ZGVpcJtDctEnlDDGBTbuOdxKIFQOU8CXUos48AP2Nmmx4BNjIx+cGHRXIUa44y1ttXc1
JKqoZE67aVmzt14TaQB81In44+A6cXzbUfJyp3dfaQsn/noHYN7sxacavNSQV8H+HPJeiTDHJdwL
wtkSogHMAXWLUxG6VcF5apeTO2WDlQT5aD6ZB/a5smv3BkWoCD53lL5ebrLTGz52yeHnPzU/UZ7t
fR1zHXSs5XA6YCWcPy913d+hUaV5a0ahR6M3L89XqfwDwrYh2HEE/n8KjChC/Dc1mDYikVrW8xSU
8KbfnJl83ok6cqtyvRlok6LG3kSuPlOGJ6Z9QfIz6wNxJaVES14S8oQLaLzc3gpcs1su997QZOfi
BKuwDCZbDARa6MmAlHdWmfPx+nBLWoKOUDnAx4y4h9dgYemTPjkZ6dGzkzHPJTtp3eNs1Ro2QesN
whgOYqhUuw39BetA07Zyagm1tyRP18v2g92rvcb0r5kz584kjFgTWEk2nAdvxm4Ao7FN9bzis7aa
uLzA2gGi3O5QALWIpD+tLQU6s+7aFyFwyn7K3l3aM7e93G2LL657PqqedFyNJ1hzcRwJNM2TQlpo
tZzcMiOAH5nrQLiP3Jh1vKPcvrGa5a2qSEuTI5P9rUhrV6hJylUxmV3amhsKge3QZpLD6MHHUkE/
xam2mPrbn+mIOIWyFz0cXcN+HjICevjGD1uOS9qJs9lcU3/ZOOY32TrWY0SysntXMeTMN8rL/4uY
JTQ8I8FTY92HN8QSSQAjCdktSouZqArA1cKcRLiYSmpmRE3PzNmzWzfqX4zsmYQTcwFEboejbr/2
oNX3FWg0r3iGXbOiBm8eXokeCjY602b0VC3ZzcCZTnBkisKnC3nht0TC52zxzp4p2lJJgJqo7ZuX
z0GMH+HillGol8qUi/tR9vJvlE5icIY0nXNQfljdi0+nRo344+VVfUc/91PLvD9YE22/A8RKlD9b
qdoMZb0PNicqpWT/QsT/i5c5qquC9NO5MJ4F9ujJJZM+WgxnTIwm7m+o5K0ImMDfeOg/hIEC4Fl6
P8471ta5zs+N30uzW6Ny4NH1skz/JLtH5lb5/uIPlGUunqnPTrgHj+X/qZhU70zHlrlHI7FxXq/l
BTaJCWeebxAA1fPoWKS5VNejlRwNgmUZmGoLLNEeDR9xo60m82o9suhvnEUULxnFQQDPtJAMeBzq
pTaDt/OEGoo1RVW7UyhZuTY2wGXettX4zu//yEC4RgYorQ8Ja4fnMu/ZWwDMXqGdLEtSwqOemaRD
Zu9U3YlxTi9sfW2tkUNLJRBoT+F1NNevoNBi04ZEJQ1mZapx6GJGDmCYLAa4M3L7LbhasM3EGYbG
/dV2V6vAYQ2JtGdozh5guKiWMWaiRvyJO1ezv4cPE2aEnPSdANT0du+NfzNg6mSSeuqBz3puDIe2
J6iU2yWwVNV6wlBeGEKZbnrfs57EgDul8YvYu4YperaA6U6686hLSu1eIXybKmi23NrOg2l2ZVPI
3r9cay65WJ9eBWjTTF/ASi0DShwKZjgqrWvExgyRbMfztyWsRphbIabLdddG/iw8f8u2bhDK81a9
H7WascJbsAhyRx6ZMlBPkTMxdfA3JzXQckxf0F8D++bNdd/ItZ6jcm3xWR9z6oLQuuOw7w2UvPhT
X71hByln4QwKv6FNHmkDWSdYCTSorXka+Yevl7Lvpo9ctsw4NIP/FQ8gDJJv3O3gSTV4P2x90uIY
zzk0/NKwUqGG4a0ss+VDwWU2P4Db7YVZ6a/kVxJbT+z445SoebhkyB0Zq0C7I/uushrAJWHZAgxs
8npNIAvxswylkP+uxRFYZUXJxgE1XKNU9HnZHhaXqWKUFNeLmSPe9qjRGVcNKMCbq+1cDq250ska
zneHatkCv9laeF7AB62rEKKeu0ZzNpfnmO6y2pZ+eRpuNSP7QHDcWCgRdHJL1Z0C9GSLOQNT9P4J
uu3qnbbknQxdxoiN9h2JUjj/Qq4I5gO91t018Iw7FxG1cSmNWXa3toT2U343+gSsMEXn95ly0llI
Li7psqr5qFask34Gs7g=
`protect end_protected
