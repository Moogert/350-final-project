��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.hq>dT?����
�6�+Pj�---��÷����o��7��soz[��ψ'8,I���?)�;���On��^:٪v�6�3U�nRz��q	�ϛ^��u�!�ZP�-��JxqKy#I�д+�fe��"�e �Eن$ �d��7�ͮ���!K����z�Lf���~a	+����^	�aq�����8�����ӎ���4�U���/���`׭?�V:���2��!O�������,jC2��{���`�
���w�����S�n�C�j�9^��8fd� }��91�,4ӦT(C�3����G��3}B�������L!2��}=oUI�� =^��qs��!�J(���1��׌�G������o%-�c�e��[����%�����Υƪn����4X����#�;i��E�cq,�t�gq�*�R�oh����V�7�޺��2ٟ·_;!�(OǑr#�Ȭ�tߘ�d7��6�!D;�F���-<k�{Ώޥ�W)zs�$Gk�V�.�t����'��ٕѶ�JK7�R�B����x�B��(rbW��֢�\ș~����<X`f���鏂� �[[gq[g�~x��K�B����/��0�;�/y`�b�6��H�RTO�=����3^��R��ª�T�s��I̼�H�\�g���L�2��s�޹�*���&�_��LI�*jiC�TPC�����!�Vˣ֢���|��.f�^Z߸ès�]*<d�A�j�n�?����\4�ٶ�V�:�ا>�݊�͈�w��,�����O3�ɿ�8�st��)���~�
��W�
��q��8	ѿ@';�=$���H�d��\
�����g�>���v1���В*�'�����=?}ty����X6�3���%�K4�!)m�F��	;c��S#H��?�kX�ڹ���C��F*�>�d�����>��w���>��7�bD����AI\�I���_6/� ��X!�s���y�v�v�w�����x&XT'���J{2�۰�����`�݂� %R+jZ���h7�X����ݙ�ќxI�դ}$�g;�C���t.��屫��-?����N�s:E��J�5H���-�����!�<�j���R�,T�ږG
���,Y7=P\i�#{/շ���s���h'�!V�����c��S�2dS1k@�g8� "$�	�&��Fu�fk|����^���wϴ�m�8Ň��`�?Z�f>�� Z�K�$M4��W�Vd�}7�x~i�:�}KK�?uyu�׶|qW����Xq���
#8x��[��H�ݩ��?$�v�U�ߣ{�q9N�q��ٺ�(�Ý~����OKz#H�/ _M�C����$��f�"�m��gTP���o�)'��Vӆʆ���:�����w�W>�=q`³�Ɍ!n���M�d+�X�5�(�݀�8z&@)�I�t2l�t�_.
�wm9�Y����Nv�2�ߘ���]\$���@�q�OfD�m�Y�xB2�v��@q��ݦ�wf���T�k}�]��A��ae�֒��f�Gf�;ߞ�n_���{ G�<C����n}I�_�쩭o�	wI��p�$��L�d2�9��ն�4��b�G<�M���s�%c�u���fy�N{_g���A;O�S����&W�Q�~��x�0����_ϓ��'�${��R�����a��(:�(X/��@�m'`k�4O�a
JQ�V���W^�^��� }��pe:2���q#�`�H̽e�<n!���"�ĦC�n$�,Y���/��6x�%�a'j�v�Q$RuƧ��C=���zw�1�A諞�!f�
�]H�c�[�1�K�Ƣ'j�T*�)~�o�M4O
���� �9>��>4��Ūi8��������N@���>���e��8o�l�����ޞek�pM�\W��3t����"�X�&J�K��	�E����!��1@O��@���_4��$xɴ�����Y�,���|�"�9�o=�yi~}8Ei9����0Uw��:�O\7�N�f�gxU�qB�3z^f!�o��5��f$���?D0Ƹ7��_΃̅�%��J��8$�
��-4�;���5�M��]�={��y\ʗWǁ4����Ŗ�;���8!�a�Gy5��+��.��Ǯ��$9�,��)3�? ��P��֢S4R����SGdۥ� ����"�0Q㣣�� �FؐTY��gXi��ןkb��&*��o����k��ߺ�")��]KA�n��F�ϕ���T�&�~�*�Bqv!��
��61S�kܤ�����Ρ2��y�(����� ��H�@"W޷8���z�|�$�P��7��4Ͻ8�V��$�q6'?Ϯ>��!�{$�K��g�1�K^�T-�|8�..Y��H��rm��G�.;0�*�ՄMs�GU��i����V] ��=R�]�"�>��������:0��%SHݐ���h����kf�X��.�`���Uиj�������Z�������F�4�0y&B�g{��#U���?�.�ʪ�[���i�mn/�>&��%�>�HƘT���|j,�|e�s�����.m���� 	�х�O��d�B�����^��(��ol�q�A3���l4w��F�#JE����Y<��f��]�<i�<,��"�- C��맿;m+z��u��L��|�ȫeFL���H��)#5���ܝ�A�Uڅ-��V2�/�T_*<S7�ay��a r;q[<�NL;������}�� C�ȀP�(K�90L0���YA�|����d5?��1�Z4����;s��u̍$;k��(k�I�ڏ��n���sZ�0���՗$C�� ӍJxQr�?��BVUrl�um_�M����XG�{O����O:biP�����EW(JvWZ2 #o�S:X�243�L�����w��A��:�� ��_�����a��7�6
����/�?�oꤚ��>%-\�C$Q�����8j@ݘ#|�a�W�v�b24�N���9!�:��slǛ1����h�	�����c���i(��P#���@�[��+�3Ϭ;��5�:�/0"\
��`]����d�zM���+Z�j�v������O�>&X��lfL+Z���{�Mf��(��Mw�Jx��i�B��� ����e./�>X�)��6K��S��2m|ݎ��c ���H�@�2���!��v;��h8k��,�Y�u���C����G�GM#�AR�;S��F^�<�^�yk�*K�N��@�=EiJ F��� ���Fg���fi|���(#wCe�١\��m�W�Pؐ����`A��)�#�X�=�%�����
">��9�1k��`�ٗ��8�y����T	fuw7����o{�?>ۙN�����C���|��A��p��躩@'�4�?dp�m�V��5���7�W9f+4�[�۱��M�y�Z�ڄ gy�g8����/�q��G$^�����T�)#^�_69tU��3�G|&a�{�z(v��ɍ��g*,h���bv 
Xx3�w���B*iC�$�d����I ���Z-o��|
�%�-œP֑(�(j
�L����� �s�0v��"�n��>�HdBC���E�,i���ڃ��L��sG�Z��{�xs�1���ɛFtoa�&b���A���g�8�l���������s���
m}�(�%q퀪�lB�-��H�X�9������x���B��L�}�l��֭e�b��#x40�l�b��FŏNVD�Z�I����ۈ_V�Q�\�ȶ���x��k��/�LkX��r��`#��-�8�F5����dR����Pɿ������d9!l��KW��j���%_v�3y�d���Z�J����ob��͛��0o�ܿ��تX_mR«p�$ �_�*�h�j}m�\��-��z�cWv�$�d���w��}������y����0�rO����|=�P%(��Z��՘=xi�&��LrSF�ͯ\tq��H]�X6T���h8|1�+t��a�`"������iЙr�gM5��ۭM;~�o���	Uͪ����h��/�;F��4�X��-�=�;BAm���|t����T�|2�ſ1��LA�TE��fxU��<0˷��Wk�(�c�z�]n<�>��W���HJk��k���2�=F�ב	��[�b�ם+zGr[+�j{������d�c��p�
y���EQB���h��3�Θ�H'x���H�ZJH�^ ����%�?�iĳ�%�z5�Y��35����IlqJ�'��k���Qk҄�{�IQioÄ��B���e��ו���m��FE�"b邖΢d)l�rz��NU.��~8<�;��#ܸ�� a>�����5S������R���e��(n�Tѥ݂�S���wo�2�z�����zuah�i�CҚ���_w/+��*�oIg�XZ0���}��&e�ʦ�Ȱ�K�t�gS��._����ѿ��~�&:ݶ�V���C���U.�]�`U�L���]���ՠ�C>L����!�Rd�x⼮�$�JTe�n�y��y�����쾮���@�<GO�v�����W�y�aJ��ӟ�����7w����W�>����H�T7X���Z8-��x�Q����
�������y\N��iNzܻ�cn�(j�xO�e鴅��|�A����Ǭ[y���WԼ���6o�?y�U��*c3��M���L&�|�$�U�g#y�GW�P��)���_M~2�<9��h��e��v�L�W�;ZP�{���($�e`p��@˙y��&�QوT?1��9����%%t��:��<�=LV��T3�J��7�Թ��D��uW�ä��9��b����u�Y��<�Q��Ck��z5�j����!��q��Үv"ǋ�'�I)���&�{���Mno�J�0���+u�������҇�� =�{�d*2!��)����[��c𽿭=��㹧�ݨu�����;�8�W�-�!e3�?��~���e�t��E�o8y�b�Kw���EB%x_��"�
��zm!���������'�
�1�\��+��4))�R�_��izҺh���")iP����<*�w^���ҙ�_Z�)V�?�^�	<�Ys�z3�qx�	Mk�m�'֦^İ��q��u �-{t+��L���D8Xz鉺@MWIO�g��9� �G����騽Ё���R�_C��5�^�"�1V\���9�cC���@�����t8���W��н%=�HA�om+Pt�ȗ�{v�)����mx��9�L��qn�y��1�m;����^+��x��܁�_m�+�x@�T��ɚ����-<�;W�h*��F�m9P�|Jn��{�X(�q'��זI�mY_���h^����z�D��$�Oْ>�������:��c�iwo�5m�~D��덿� �q�n�4�T��i���8�����Q��]���
gM�׼�����@0F����3��<Gz�� �n�4�[]�{�6ۼ�	�n�C�����Ǥ.��,��2ŀ7��7�8So�*L'��n�q '�?��j
�+Ñ����?�t�H�`Yɯ��dѠ��+��t�N5�w�2ŉ-�i�	�hh��e>D�=[lπ;A��t�
��D��O��X�hd��z��e0=���_�L� �G$��4�T�vh�h��ŷ�T�D�i_����4ŎV;��Cd���m���.c����ի5�r�d�\��J�s���ݙ�dLYQ��O'(}�Ҕrh�}�af⮧���ۖ�.sk��VV�������,��1l3W�Q��c�T5O�t���t�����ApΞ�V���)����'l��Z���Zd��R���
�1�݊WG��K�X�K�3vOt9)Ҥ�y>�+A�Y�+���GMF�8~9J�p�s��>�d�� ���Z�a6��38ss\;�μ:�N��U$�zأx5�f��DDs�9� n��#:�� (�r����Iz{~�;��C_���޳�:Y	_Sm}VB:��w3@Z��$hy(��@1�pkQ@O䗗 �dN���h����Z���tZKH��	�!2a'�J�˽�F��t6J�� p�=qqz؉n%��M�X��ƸvĀӋ)
����Fꂴ�<���P2`;���$�wy� !E;5��)a�!��/��;,ތpSy7} �DY�=��r�k�]6:��f��5VCKa��C �\�
��C:�4���:o멭�
J�%@(��T�;{X�Gh#���d�081V`2�l�Va�Un�����9�a��w[|�rG�{D'��}����[�=�á������N$8ၠ��t�w16$���u`���θ�������ʚ�(R�it�~C�K�xdʚ�9��V��%�?ed,1o��۞�)�s�ɜ���<�Č����{6HW������|�Q1��j$JĀ��e�i[�2��G��4u��q�h�Vc;��:"�.,��uTɲLz���E��Z�Z��Q�����.��N�ں��\�k�M�s�u%wV��dn���k�irr׶�w�>��}���#E�Q��5�K������Ԧ��߸A�!��A���N5�؎�A�t{��ƭE?}�h�G������8��C�������`z���ۦٲx�Z<O0fs��[!2oF��4��:]`f�q�I�5��,9���@�Śn1���Bb�B���l���6!RI.��l�-~a���(��7pD4s}��յ��V�8ZH�����E���; ���r�jK-��4�Ζ<���sj��+�~S9Vt�פ��$��"%'�}��6G]�uG�j�bqK�!YO��v�BM��V?�!��K��j)d����OCp�m>�(���s�Ԏ7mu7�V��A�3���
�,$�bd�4܄Q|w<��q�e�[���f����h�D������v���^�l�&��98L̈́�u�����( ��3f!#=��G㇖����3��9���V2��r�)�QU-����L_��29��RܭC˾&��S��'6+��������-�k&�Վv�l	�-Ѷ�j��'K�F4+F��,�Ώ6�p ��["�9w���+����'���i�>�^�ا?F4GE*�S�V���e���U8�_��f�$s׋
�?��\��R�1}�&��3��H�9�(�x)]�8~��c��<���r�Lf�6��q�E`YdҺ+�n�.����(�2��Yl��:���xx?�K�UPv��4�'o�Z��q
��=h�[7�'�c�
����C��v�I�߼gm�p���5��U5�7�IOu+{,u	pK������r@���j�� �[�$m�.	���8!fCg�0@ھ���	��3��=��6X|:L�8�v#{`߬����+Tn%9���*��vcd�eg�/��Y	w���^Բ��_�<qN>�,#X.�d)��R�Z�lߩeJ�䏓ț�S�ĵe ��yX3s��:=�H���C��;���\�%�Z��g���ǂuZ��Qn�N�7J��R+��[M��������P�=��"m�-�ɭS}�N���A�b�n�	8����E'G�W�3�-�a��������\�����"�/��\O};l^��-�p�r1���'Aв\Rp���@/�{z�T[�6�ϴ,��r�h�;�MZ��9�X
a\���Z!�X:�[Oi��h+���	�kg
Hv�h��H��/YrjsP)�"]�`SY��qg`���%��휽�� �ˬb�)�buw�s�&"�=%�H���r.î���u�����vL:ؐ�*��Ф-9�}:T��X#����KE��P��P�:��U��ٷ+��j���&i3����'H%�+��]��ÜЕ�.�����w��L�S�c��4�0�J8��&��8g���d"��%0��)�ݓ<��r�d3���p��N�ϯ7o�+=�gJ�'=�nm���@'�&ݲ�T��e6�a����.�M?Y��K:�"�o����Vj��	��/^t�I[�`������=(�@�;p����c��ڰ\	b�N��g�HuG�C毨>�b�����T�� c��y�W4�͉�&ы`wP��"��=)i�m]<T��L���	���Z n�G����9w��~�ױp0���J4��&�N0@<��,�1�E�����z�g��q�>R���'H���.0��8��$����pv`�����
%|��[��È�2��]r�HMK)t��u3q��ɭUj(�d�׎�)"��/\�j�n�}��E%����;+����X��W���c_W�w�!P^��k���c��܂�I?w��2��l#k�L_XO�1�������q�k�[aR(d���F��C �R�P����pӅ^�n���3�:MN�`��3�%���zٰ��{�vD9pH��@<B�^h>_�r���`���Q���z�H�i�Ǚ��ґ����v�F�}v�U�<��)7�5��̪f�)��K���X���
R�%�\��)�o5�i�Bh�W@y�Q\��R�� ���B�dxuA�E�v�K�N�g�>*,�Y&r�:ʠ���6�npU7kyX{����.\��5J���^��Rǟ��Fpgz�Ȥ�py��ߴ�qm�m]T(5����Dg����5V��]�m��"Ɠz� �-�ꞔYP��:��t~��3��4S]�iˁ���Э�,��)�~�TλQO��kC�+u�}Hɐ���ݼ$Ɨ��߀��R�ul���((�0��Q�;��Cxs���+��ْ��!eҟ���a�k{d��s�u݅��O|?��\�n&�V��.�����칦���A���ć
�Cӿ��;�*�2��HU���>xW��;wt�*��rXGV�p�ж.[��@U�&��{Hb���	)gmF�jS��ߢY�.`9�˷��Nl��ա�����Nm���)�o�d>}�eh4)k�C1��nt�H�e�)�L�H=����J�܇u�7:*l	td��I
M����q�r��~��l5���a�=�M�0������g����FP�|�	�h�}�L˛�3�'��#�w鏔uP���oQp���ö��r4#��*�N��c�/?�p"4�Y���t��úk U�&��V�q����FҀ�rg�{��T����8��S���pt	��i�Yz��Ϩ%g"��&:��@��S�{/F������W�O�AI��D�Lsk����7?�H#�|f�1������˙�\���#���"�rc�Y����j~w�-݁zOK�;��z6:��@(�����]G꼨�r�b�2�T�ႜN�IE;�G��ъ��5�$��r(�;�tTu�1��Q��D]Gyk'	˘�P�A����Y/K-���t���3bt����+��*Mti��В��9c�9�Ƌ�j��f�����3��RI%c�٥��'��p�<��_�9s�cē(&пB9\mD!I���*A�Q��ł���e����->�"
t�:üe���j�9I��o��l%��/��܂����_	@j<���Q��z�o�q�?Jݫ�dg��Ct��z����K�"V�p<Іpzgs���j1$�^lܲ�Oz�a�R��.F�,!~:�4�N"�P}��_4��Xԓ0Z:��Di<rzşWT�$~O���N$Q"[n��-잖��톉Gx�/�Y�h�-����};����)������������S[�ȋ��r�,;��^�D�z.x��P���?{�Jh�Ʉ�]�-��v����m{�<�ܣ���M�d�1��A���C>����<�E_�����c��3����
:D0C"偯��It���F�k��1u�쮷�� �L��.U���[noČm�Gظ��a~@���-i�dJ��t�� �"h($��@�0��f<̨��$#���.�	q/�?�f��vƳZ��ïd;y������p�+�	-�'�e�5��_�}9�z�ꛧ�N���ˌL����G�W�.��-�����۽.�9~����f-��ܭ|?����[�x�vM�Df^�y���tA�����r0?�.�;6��:�ݜ����յ��,�tw����o�v�H?����*?�:�l���쇄�)'ؿ1�=�t�l
ρ�s22��a�2�/8yX^��G9���Rs�	�Y�N�.ꒉ�Df$~Re,_���Ic�&��ʦ��u�`B��Z�?����2��.�A������A����p���[�2���g�L�=����W��?eG�\��[��|�����4�ʍ�ܝ5?��=}��@�;Rh4���Z��U�4�����s��d3
63����9̂٩>�\h�!j��bi0��GZ��b����`T{����e�M�I���i�bۥ=�[�Q�ҩm���`�x �̶��I��_��%��,��4�JƎ������{ǭk����vZ=pvJM�F@���O�K�Z%�y+$�/*WY�)��ȁ-��M�{`~hU��f^�~l��u|2�ة�	E��	�*P��9V�+�70��B��/��(\�N��yM����� ���O��xA����{#��({�]i'��8h�A��tt�TK�W^~�/�(��d�-�t(�<����/;W@�%*`�g�۾"֦��p��V�&�-�j	b i��H�g �v}�@6x����6أ.��@�~.�[:(��P;jP13y�x�F0�u�HB#erH�Cq���������E��b�P�E��=�"�68�_P�~����x�çR���!��ۇ$z\0���jX7"�$�2H�X`}�j4IF����vt��������N6��ړ��X8%~��ߞ�l�������N�5l�ܮ�(�z�ݨu�(���Ƕ�t�(u�W���������鬔��7a�i��T��.�F!��\`�͡���:A	@.�*�e��Aj�C͗��=.��K+�� ŏj|�e�m��m9бŞ�����
��R4��%��m/�+pirHޟ���:)eQ�W�ր��|{�M�! A����y����
�;���Q�^q� _p�)�u��I���_9���̬3g����j�]�$�:0Jø�"B�@��8i0B�l+5ភ�"�,T�LчpEr��{��Q��a���$l.�M�`Mr?V�'�֮��\x�+�wq���Hj�<�1^[�o��0rR!V��ϔ����<�Vf7Ȁ�$��]��Oq�ͧk,iE�xS��V�%t"� �af�-R�t�p49R6-L\�anR��^|6h��=�Y�����s\��`ˎj,�[��(��A�&�����q��"I �$�OQ�'\���'���f�/���L-��b�GY�O�!�����*���~��нI�+FN|S	�Ʌp�W0�������k��rߚrɺ�2�T��~.@VG�ŧ�ىr�'M�N��Im;��`���W���N�n�W&BrgB>ڃ��'�
�*|�=��]�j�nAE��uS��T�n��t�^�Jw}���3�q��w�Y;t��Ǽ��Ფ�X�Vp5)�8�&�,r���edr�[x�]r�+�w�1܍ux�+i�Fe��r��P`�bm}� �u��w�	Λ�3�~�0½1���80���OaE���C\XPA�~j��|�OXK���Tҿ�r��r7�b C_�hԡ�/�_�>��S��;�v�+�zgg���ls�S\���:D0��Ɏ�E��@�TkX�<���Q�ǔ������U�_���V�4��V[[����:����	��v��I`*R]�(IM� 7�N���a�]��x{�?c0`�W��fO�a#ݵR~q=�^>MC� \��k�0C��2��M�U&���Kg*�g���<�PՍ�q�"
��'8�sｓNT�^�lƥ8� ��,��#�3z˙hOW�GWS���)Ρ��o�p=�kr3�_$�8X�v� �ՕQw�#OR4|������1��-Ċ��(!O޾��bMIMK1,���ö�3۹6��Q���6��fW'1v�m��֣iV2-߅=}M���U�&o�+����RGvh��H�i��gȸ�����F�ӯCSu�{�c_h���0k<P��L�Ŋ��.eW�qr��t�$�"u"�J̓��r��ۗ\��ܼ��Г��LM�yרN7*�aK��{�|��`q������yˏ�E����]��^�Yt�m���	 [�H�N�:]�*���,����?�d3'&H�G �"���4�x�q�>	�w��K���E*8��BO /�<���D�J6��q�����"/O�4L�i�a�O�Y�/�t��Y�td��&.m|E"fZ�?���fw<E�\�����h���~K&���ZbŹ��g������&nZD^ $$�fh�
/��g:����It`R���nAoE{+��) &SS$]V)��Q�P>�ء�$���*t��Y�'5�b:�dR�&E7�C�#�eH)y;��-�{���Ӡ��Jw���Z|cz�?��j2��;{��>v�lr7����	/U\�HJ�H�r�"�	b���|��
�;��� �5	PP�n+=�)���( ���2��g�=�mb���B�7�-��]�K@�pO�J>��LIs�D�,�aR�D��=9��t�<����(�ާl�6J�|	%�P��2k ���� ���[ʾ��ۙ`�pF2��%�ß\�窚d`��E9�2U�r��I/�?��|�k�����Z�q�>�f�mrc�규���/C�xp���X���"H����C�ZCV�Q�����$���NfcR���U=��lzb�%5��;�uH'z�u�EƗ����Oh����L:�s`xM�;�З��ĒAu��B,�I;�쵒�"Gi�L����,C�� λ����4N���|�\���?з�&70��BJޢw_d�
*ͤ�=�8��{���2�'��=�o�yY�)��|P�����lK����%W.�� m��*�J?_�@���%���4WB&��t[���6Ȝ�X|B��6�r��yi2�b~8ŅW�Ѐ��H�Mh�՜<|��ʗn>c�}�MMkE���n��1�H�ڳj�#�$A���e��Ի�GB�+�ה�1��
z��'M�L"��� ���r��F��3�
9%i������u��Ns�Ĵ�ۯ�s�1(��'[�l�J.f������vg<�t���ʿ�W.��C��N� ��˼�H���}u������8v�6�����0���|�E0{����  %�;X�Hu�'��	Gt�����1P��K'�Ʃ����t �����8����ގn4]�و#�b*7r!H���d���4�J/P�݈�-�>bY-��,�vFg0�q���LWu~Wm�6"�B�C���|��:��7�����Z���I�O��q�{�N3��n�G��!��ue!o��G�_J?��m����c�f��Ζ,�r�Vh���\�O+ȅ�iӀ��fu!�~0i�A�	�"�}���*����qG�C��u�<7n�Х?,�#>H ̕x6�d7Y�g�����zr5�J�#N���5��viQ�Ma���νş(��q�'z8��6n�;mct�}�,��t����m������~&a��1E�|Q�r���0
$C�p��>��+�̃��eh���jc��,�4:sd���Ս�B|�N�l!������Z��b;���^c�����M�ѐ�`;�V2��a��%7"R}��Z��(D����]j7ӊ=~���A�-�8�h�Qs !+�$�PH�ڬ��tW�Yx_�ӝ�"��iP���Z!�ѷf�rd���e"<�h���)�^a���#��1����'�&,Zxu����X���7]j_X��9L>�;G	�h����;!����7ڣ�=�p��y�s#���
\)���6�f��z�qE����{Л����h��-q��e�_B��6;����a���*� �d��[�2KDL��)	��*�c�N��@����^�<�kI~|=������VDS�������pt���?0� Tmr�С�"� ��e+����'L�r(t]��5��/�Z3�&�P�Xa�$���t�t�>���t�^����r�ҵ��
���r�WP��R���%w�ƚ/��Y���h��)���������uɍ3��V����n'��9���%Z��vN ��t���|ȿ$Lݸ�ee����#6Q���ͣ�ѣV�(�c'q�@�E�wŽ�^a��kA�5<���K�oWM,ĒE���M�;=d �ji�UO
�#� ���F?��Bl�����Չ�2|��O�fHlK�U��A�8�����oTC��h''����a��n�6.���wqhT�2�1��##�CGbc�Z��m�X��~ L�c��7�+�j��}�6�����^k ����(\q�_`g�����J�
���Pr&z�q�����	��t��a��������9�b���1rN`(-"�nI��/0
kb���4r��\bf7��?���}:��.ς�n�����~��^�8L�f�Ȃ�+^˗P0q�弆H|�dp���˙f쪎D���"�w&�i�W�Gf$���x�p�Ȍ,�{���W)�\����G���7�0BXB�϶o�����\�u�Ņ���Nn޽�Ht"�~���F:�Q
��5�1�Iv�϶� /����S�)��ݸ�����5u��C�?
�6�8�=SK�?�t0��Ʋ�̒�rYvFp�K��?���a%�l��N��E)5�w>�B�ʺ�zۄ��������7�Mo�1�VsN,��C������#�v�hFz�3ܩ!�����Ԁ�4ϝH_-Az&Q'z]Uų'Y��Q�YV�������%�|u��~��/8ZK\XjM�}�j��:eo�sgb�a�0!iBC cEPMt��<�\���F��%��<��z�~�9EU�l��ċ�]]9@������ο�I+$z�NZq��mom���;:�9��m��^�*� l����}d�/��(������boR�d���B�{<�������7�Ϥ<�$K����Q�L�z/��u��yN�@��&<_���B)��pN�[]��&yrXB�6Y��ڄ�oӑ��q2��ָ�����b��{���~>�(��P?P-]�u_A���.�5�S2���Ũ�u�Z_;G��	�SfA�'X�b�KV�HU���H3s�>�Ж�ϙ{�4f�b��p{8S��:�5�䖳�'�7*F��R��Ma�RS�Η"-�
g`�z�T�I�K����Ko�
�����=�f2�R��9��_l��{[n�����;�S�����\I�5:�՚}�� �<7�����;ĉN�[��I_�M�'�*���b̟�{3(GN&���N���H+���\����6ŊH������PEST�GO��(6G|���M��W/�l{�?���~Pt�Gt0@ �ڣ����iDz*��E��$D<��R�{IQ��iv|]�a]Y#��ֱ�z�p;�`��j�o�K�]˄�����[�u�,4�	M�_6�x��h�7��-S�"|�)�&!�uP�UJ��Jܲ���ʩ��PW�4�3r�)+���N&��&5/���a�ל�D�֕��6�竎�	]ź��7Z�|h]L�'@o�ط��)N+,��>-��f�T��1���lS��^����甮߁	�1�h�h'?�ʮ��Ħ�� �"�,Qk1W�rA0��{=���Qy^if�*�<��K��^~G��0�d��S@۶u�|x� �{�hk_J>Ui#�פ])��J���"t�pQS���eʷ�q��$�
���_i�S��e��F�-^��e�(ؿ�����d� G��֏v�t�6�7�TNߦ&���c)��ML|i}lI�A��j�tAi��)?�>z	Ļ��ʅ���Џ]�QQ>w_�ĸ�����6��6�OKn?6���/mO�,5Y�X��D��>me	#�A�*s����������6�)py�/�:�g���И��W��*��; �Y߂�yt��"�Y4ؓ1ش����ʀ�Y���7?��S�Y/��U=���O��l@��g��$h� �s�SX����1��Q{��#�t!��X|"�6+��z�1����ٺ��Xfd2�ğ]�\���?;������׻��aCخ���m��Q0��1:�C㫃�4'�s��ʰ� ������0Uv�Y��1�|��:������b&�m�
�p�Һ������Zg�0��7j��f��l�I���ǮH��E�8.�Ē%㲆&�Ah�t�#�-��#q����|�x ��_��)4j�eye��-Xh�TA[9p���7��������7)h��XRl��RB�a�4,����
878H�u�pϹ�����g_���0�Q<#K�_O�@PHRI%)�Qh����~'��z����t0���#yfә�E�W��bE�,ֺo�d��;���G�:���/�?�v�mf��ݰ����s�����çD&�	�/<������1���B�d�a�
Z��O��z$�s7R�)@�e�gfs��\�E���$�\�D�Ƅ�kp�l�`O����k�4̵��?n(��]����p���@�R%&yQ9�<w$c,K������b{�zW���r����r��wii�P�Vq��ʡ1z�ރ�cH[�����#ث
��	Ӛ�%!�u�7A����6?��L)��/*Y~��	�a���B V�+����Z/����?Rq[˭�"�$H�z�7����P�Иs6���&�Ǆ� �4Q����-oD�+��▪�
~��q7h�ȏTó�?�)��Ou���EgJ��c�f����K&r��.%Kk�8Ѳ+XD)K���h���� 5ȳ��e%��/H�ۋw�Ԭ?ME첍;-bZOlm�h�i>�8 컩,��q�XZ6�lYK�!��듊��
LD�h�<T��m:J�`���x���nA�����}�U��;�,
n쵠/�m��_,����(4��f$MdI��>���
�$�Q�ҙB���Ƞ.�Ԕ��8�Ʀմ���}S�Y(l!2�^	���Mw��u�q���t.3���ݯt�t8ȥb�>�p�Ո�֑���/̸�&���vQ.��L�q�+��A����U`� {�5�n�y/��A<�i�bg�e�p7:h8k�\0˺2�JI T��H���+6��X$�1?���?�#v�&��N��e�9�k��Nw�	wԃ��$��(Q�]�)	A'�\�79�������&��.ۃAIк�r���؉���ax[��j╟���3�Oh��-�?IY�;/�MU~�e�$��Z���*@V<R`2�5��]��F��@���Q3�� ��܀���૔ ���t����Cl�!�����8��Q���~5�y�8\1��=W��$�[,�^��}��dO����Z��Y"�a��[Q�N��E}��E�e�������,2,`"�� A��#��!������bS��Q��6���5��,��L8�ԺmÉ��
�p�h=t&+d�������a�����㯄ϜK�H��0�/'e��L}��?��N��k�&�fzB��7�U�O��3MO��S�g�RU���!�r�h�<.a�5���&ϋ���7U�E��/jj^�6l�p�{�S�=����`�T-T�V$OߖZ�8��P�oR�����nx��{�;��rh�T@�#vhZ�I���6��(l�tdn��O��HF%�!����ą`m{�1{��m�,2�dX��݅�%���5H�ե�C��N���8|��Bl�V�52ݾ?�ln0���W^�	B�j�/w�hMP�W�c/&p?_Ω貊�Q�o����R<<�+/�˝n���e*���
 �4&�}^�z�`�5צrܮ���L�ҎV������b�����H)����z����o~��+�Zg'=ɞh6�����d�٧�ɪU��|������P6"�D�2Ps�=Md?���//qӸV�m��? lu�h�2�N�O�;��I`!��v�_>%L2�!���kJ���_(8qsTu��{։�x<+�~�S��>��D�W����n�aD�5�B1Ntv60�V��t5�R%���Y�ۭ�e? �������v�dIoԷ�v��5��q�� �{勥�Z��{�X��"<t��)�#20��-'[l���q����@�3�� z��,s�[�Ļ�~�����yl��h�}����l#�Ke�p� f��dn��A�b�\Ƣ3�[99v5Q�E�L�>S�W�)�y��$��tpko	�[M.qɍ�����,=j`\���N�1;�°�TE�w/�`�ZR��Ă΋��'�G���"}�w�`����?)�u�ͺ�'��(���Ƴ�g
�W����,�\��M߾o%3�=��Pv/���~KA��k�d%C�t�C�t���vO�`-tҡ�����yWq8�My��N@�RV�w��j8���}�Mm�kn��Q����3n�df؍�G���>!�a�xl��j��]��ɥ)���&�O�_ۖ
I��L*�R�ΰ�w�<�?�Rqf.&5W��<�/�%�$4~�6��\´"T��.�ؑX�ka˞�%�[T���9��a�d�$n�4d��JYl{�����]z�9�!��(�*]<v| ��=��C#~m��-Wl���y�[�ц\n¸>V'~/gD��������0]�l(3gגKJ����Ƅ�/]�^�";��(�~!�����W�S,�"H�=ܾ!�7mV��Qʼ<�+�B�Rg���q�(i���C>L5S�%.�K�5\�a]M^�vy�)���xS�Qj7�k���F	�JW�E�B	p�F��`�������h�oK��PB�FP���,ǡG��ۻ w>���U� tڒHV�ӮG�3�Ȕ��,\��Fg7���I�6�3w�B�p-v��0�~P қ�ù�m�p`Nf�:���3J1b!�f�ql&4�Y�`xG����"f�o+<sI�������O<���gR�|ϰ|.�v��C2HK����-:�U�$U-�4ԁu�GQ�d�-�f���Id�6��!���>D������,����=d2&'�{���  Ig��~�=�z�n%��w,C.�q���d-M�V��R����f��հ"����~԰c��1� ����%�,��sˀ�����V���'8�CV�P�n�T*|:	�}������Ï�����)�q�2Q������C$�(��}X'�&c�ɏ���{�|�=o�bC���D���Y3�	V���FTu{��߰��4����-�Z�I_}�$��H��������4h��`���-�H�0]��g'���o@�CY( ���h��Jiw9�f���}���B���e���Zw����h��k#�-n�M|ӫ�і>cڼ�K�q�!o�`��-ƻ��|m'����-h�L���6m��:�c	��z�*PU�I���)����w��%�Q�`Y�b�*�49_Ś��ʏZ�L�F��i���x	��y����D� |�ջV,%��d��~񞱬�VtĂ-��jk���^5Z�=;�����'R=8^�?cnz:��r�錞7��A{�F��m�����T�?�&c;�Q6��f���5��Сyu�go�F�PO1����W����f����3�h��J]G�̷;��.~���	l8g�lqw��ݢ�z[���bp���Kg:����4?�ǀ�<��6��\�`LO�A���c(.�n�cl�MZ!Q!B6��>R��<uMD��'j6G܂�rZ�b��cx�|~tSX}G�<����I�,���[V�;:����󙼤ڶIc)�"�%f%�7"���ݒ��������q���5��2ltQ���:�'ԣ�Q%p�U��~�8�#!Y�ΦD�63����R��m�F�3�4����r�P���	<+	�5&W���`6A�F�w�q�t�ۊ�} V'V��M�^�
�D�+,y�O�>l�jm-�Ɠ&��/V�;��n�l���>�4NuȄn��(	sͲ�f����з�&78�l��B@y/�a篵�Q}#>�ٯ	��qwF7�z�-p앝���������a�Y��Z���\BD�p�ت�l�y��iU��W�S�Y���1�zM�y\�a_t��dg�06�4��w����n4q�����<�m���
GU�'�c����¢�(���4�"� �Y�^n9�rt�&+[��r�-������ޥ+f�I]P�nP���l��0rKp���CX%�АJC-��An�l?�V�WsG�'���>��$�F�n*Zδ(r�,�����B�*^��d"4MK�k/зn���Ә��е%	�j��Ș�su�o)�����:l%?��F⎾CB%#���ǉ����4��r��������';1�=	�8y|ڠSOla�'�����<����&�n:&�أ�c�\ЩQ�k/h�S��,�S��=���K;k{@Đ��ژ��N�+p�������4�\��k�UU����+ɻH��^M���V����2���(�#���k^�|]�YO�U�d"!��KQ��}�Y��?�����9»���a���o��w�c��@�j	xd;�;�A�Фߘ�l����
�v�����عVX]e���*�sM�k�E܀8�o��m������)�:*�Oj�Ȋߑ��R�|Ƹ�1�EiN˒a�ݥ����{��$��[T�eO�jcn��f9\#~e1ЬL6�'�֟��
�g�M�E�To�g^�;j�6���O��k�n��D�M,�Z�^�;��a���crgr�
&�0Ibd�-�9?����-���O��E<�05�ń$��[��51.�S�JT���c\��?�?��g�=$9l��:{5�S�	��r��ѯ�z�����}��S�h@9�E�fp�k>��?�ب�]"5	�Hn}���D옕6�ʣ��gp�����f[�����.aT�����v�~��Lo0���El0g
8����1 ݠw˫���op�������B����C��8�eӹ�H�(� ����UN#�2Ӟ�����%�<��-�J���ʳ���2�
Tm��J�t[X�T��炬j].1f���G��A���@ֻ�CTZ2-'J��e�PS}G���c����_%��޾%xT[�e��$&;t%���4B�g>���}?2�]�?��x�]@��'�g�uܳ2X�K����ͪ.�"f�RJ��@Ct��"20s�_��EB�G��� Σ=�,�t�&Ջ��2O�������1��/3q�0�?-���Y_
�}��y+
��j= _�s�Z��gn�ׁU��n��<�)r9c���B�ը&�n�n��yׂ	5��Q���v�6�۴�����A<�l����'�#���54���|$��ɒ���:̥/k(��Fd0^Y���V>Y��w��ꮋ�B+�#��t�8�*}�I�x�pP���V�}B����@��d�� Հ8"E��)�@��gF�Ӂ���h=Ӱ�p)�pnj���M��э?�wjLH�[����1d�viѺAost'D�O�>��i�r�5�P樨���悯4���ŉܱ�
R��iQ��?!�I~�����m%s2]j}��q�p��H2��SG����?�i��o�i_Esڠ�=��[��O
I�v��F�)ed&����*]H�i�M.�Ϥg{�fEa)��=S�%M~;k�Q��)NN��0��.ÈE@ǜ��ڈo'��ȋ���#�.*&�u�1;P?����x��pH3|��7t;5��vj��t�+ԍ��y_7�;����뇏�Xtۗp}aA9q��h�����[��z��ql����4�[�d�9	��������pYq�.��Gס��4&��K�S�YV��L�}iڛ��^m�%�� 툙#`��í;����/����4�/$r�k?>�x��,�(�%"��!*�)f������J��r�EI�`�̶w��Rg���옼葉�\�ʙ"���H3�:�O��r�"]_��c|{>�lԳT���H4{�����Õ+-�
ӟ���4QqSM^����n�+F��j2<�S;H����.|��0�o�T���4�j��G��9��c�@Q{Y�D���(�Q�����G��<���C��[��z��:q"Ư�J�&y�œL6����P��	�u4��>X9�t��q��ue�j������#X��/k�Ib���	c�ݿ�e����Ї�,� ����c�/�]�	d�~{��8v�T��o?�z$�kbm�6v���7,H���u��Ïhz��I��+K3)��{��Zy�`��'�a���7�)�R�@^�f���q�[%����1N�V��$�_J��Ν�`1g�`@K9>[��
55�����ܓ!P�z��w|k�)E������r�!��M@9EQ}���J6���a���.8�\���}unqOPu#�_�S%���	��l9Lά�4B]o]H�	I�f����(���𩟛 9j�	�Rհ���o��j���{Z]�w<�6e��6M.������q��G
�B���PbV�I�A�|�c!�}�^�ʔC.s��w���՘@"~���Sܬ��Y�8�>[��P�!"|m�d
��2�6˄@V�(�/͛6/�zS������<4�o �.wʨ鼲�!7��N��^t��md�-�.��!K����I��%4������L�yn�#JA���4����Q��Va��4�N�Z�E�Sr�z׈��^	=�	r�Y��zZ��KL
�2���� H�`5��8�}��ӷn�ۧ�IY��I(�`]�g�4_-L隶EZd7`͚m�,�JSD���/��������h����*���:'.�J� Y0?�J)Ze�Y+i��59����]*؟b��&"�����4����@��S5�q��½?I���_^�pÙ;����ƴ����~�'k&/��3"r:�}J#�D�<�,�Z2�+ӗ�n�W��	t4Wic�/<�ؘ�Jm��%.�%4k>%�5���k�ڡ�jy��;�@�+a�2)�@�(���d�(�L�l�W�药K��p��x ?P�,|�I��X�柊�C�eY�&"t��l7�|�q6��xI1�]�#ޭۣ�)F����E�#��7	����� �I_�����(%����1@O�xx&��7�w���9�y���7%�8�A���<}S��e������$5�D��κ����ʱh}'+/��J�5E�{3t3�W�g����.H�Z�˟bZ��B�P�Hb+�ƜA�Vkי��5�Jk6(�񷚟���U$��y^�Bܿ������W]+�=���o�zb��F򧊍%���5VnU�t�D�Alޠ�鴐!�)��{Pe��4�}D(���q-��O��\K[<[h��v�	y6��X����dGX麺�u����w"r2e�"u�����A�N�:�DU��'�A�H�cyV�$��
^� ��Hc6�2��3nE���-��s"0��7.�k�����uQ�_����r���D���1O�n����`��K���LpC3������-(��}�}籃����Y-�o�ΨL/
���Z*aa	�E,��bNX��Wˤ/ �?�ܷ�3[w���/~�m�Y�I�C���t����7TB ��[��=����������b�KM,壔�2Xl�b�S��X�X�o�t����Y��S\!c�^ �	&dbM��1\���Yk! �S+�;������^�{綪!��d���$��6
��9#�-s���J�;st{���ǈť�,·v���e�S�нt�y'\������*�5�H�5��Ѵ��c u���� �,����tx��I�BM3|:+R����W��&0�Ƞ�o��ھ�Ɣ�x�řŬD�9��,;�dl�F����[l5��R��M� ��2<xioV�-�Ҝ���.�dm�O��l�=[��
a[��c��\��������n]r!���� Ih��qJ"@��#��2a}[C�~�ݷȤ��o۩��'��o�Q����ߤE襎��3�q8;�էMr���y�B
�`/�y�+�5�s&�0㇮�&V��t�6�~���Z�8�}xD+����~���rj�p�2��VI��O����1���Tv�77�G�k����>�RQ���n�WW�VK5π�[Ƙ�}Ü��3q��s�J���^'3_=g5H����`#�=��{%*��5�S�/΃mR��:�C,}����e6�eV��U�V�U�i^�*�%�5bȹO�g�&yS��ׄ� ���.��.�����P�F��3#Nl�A"@��� ����|�X�o��w���؂O�L �u` ].��M��`�!bc���E��'~�yɁ�mT�f��g�5	�/��Rsn4mæ[�:k��#��^��hl����hF�Ǩ���|6`kY��n�>��u@���<&m��
�焒L��"Oa����;2FAq�XʕY�=�*Z�G��zGh�o�����&�	�c�E~BĸD��8g�b����).��߶d
p�f9K���:��a#t፩c�oT݀�)��0��,�=�.?�A"鲫�f[=�W��$!"���s%��VYQj�u1�:���Cz	�y���Wk��^w�����aBG\0�Q6� /-����gl���`�G�|�����k���ެ���U��u�b�'y���H�>��~����K��ld|��õeq ?ژ��S�N��m&C�����L-�Q�Y��>u[�O2Y���㶹)�OZ����� ����}yH�kSw2��-ɭ�p5S��/,������V����В�ɊJOs�]O�3����m�: m!�Ͼ��U	>����%6m�C�ិ'�9�,nmC�$�U-BxS�w�v��~5r�ᶔ=W�j/ �K���5� �@����i�}`Y#f��xˈx�=�z��tL�m3��.a���V�l�麏�iD�M�>��~��ҭ9�^v���)w!�Aɓ�n6 �ף����۴��"��D��6�F�&�h�0w��]���<��"2�GdK�^uT�`\+,����O�PfΕ��M�]�Qg;"�/�?G��Ǣ�6O�6[L��$�w�;/0��3*��#���)��0�tz�i��}�.����(T���CF[�R�軵i��%�p�C���U�� V2��x�*؉�D���ź�c�"�י�sѵ�����,�fd��N���}��9gk7t���E�8�W�����欭�>v��a�������/�U�y�;�h�Yj���ܩ�������UA�c�У��L_�	�"9�O@�J=§m��Fufw��B�ݽ���v�b2�pʦ�j��k�ϰ͕K���P3��#p�_�>���o�3������3��R"b����B�:�0vq%�n+nA�	|���x��#�Ƴ����yZP�R�b�Ynٞ��]J]tpѕlp�9V�/��j#��E���A��F��f13����avpr9�a�Р��ʠEZ���w�^�����G%qF� ��ȿ!��2Ⱥ�V,d�w�5qHҰ]�9��w<��R�6��J֢��<m����='b҉��!�;��tk�N�^� #�����d.�yġ�o�]χHJLr>�AJ��8�C����M=�Рl�j�����r�!xƿ��v�ޓY���Q[W�qF�;�G�g����0��^�D|�7�; ہ\`p߼1 �Sk�G��t �H���kY	��ރn�U����4���o�J)�@ ��9�#%�2�K�~4�kN��K��͸P�jSM(_Q�D),X�� %�5���X�:�k��zf�2��p�|>	�f�E�{t{�9��eˡ"�{��-aN��=ӫ�LlR��.�)(�M�U�fm�z�"����f<���|�4�ޘ8&�Ll�4�r��+�4��ք3(��J�9�z��ʯ�N.�[�y��U�7��@������?a:Li�t���bq���r�{~zB0a�?m���Ws����y��<��Q4�� ��U��H<�.�]���`5�s�(L���j��2�t�?���fԃ��[��yK��E��n�Pn�������Tj��WT;�M4�B9��#p��2ʘ�0. �g������¯RA�X!�_�E�Ŋ���/��R�+��΋xg�}w�`��o�&�M
b���ݕi5�� ���r%Ν/wc�C���FCte�����Q	�El�P�ά������H�r����{ɭ?�����/�'�QMQ�΃��W<������)<�BP�nxE<j&�H�Y�j=;�����!��0�UF���\p\�yyX�x)ղU��U��,_��j76
Vf�	=#�:�F�Ԏ ��0
hVk9����q��G
��x�9"����+�HON�zp*媢Qn��|����bi��
�Q�2I.�V��Kv��7��r�o�0�[��y��Ӗ��к�'��_�="���6��6�)Q��s;c5RR�ev(iQ�\�������᰿��������� �'M�������kO	���J>�3���f��,�}A
>y��?�1�=���`x�mXG��6؀u�WG�6٠�7Z�b�M�f�r�aXXn��wB�Q	Ҡ�d�h< �]Jh�mW��౎��k6���N�:Ӵ�a=�1/�����=������u�1�UJ���a��{���*y�9 D�j�E�2��	"���@5�ɚ"��������T� �i�7ּ��t�u��}�?�o� i��8��:����saKS/1}k��fQ��0f2븷�2-0��ӟm�|�����Ġ�Q�� x�U��u�&���fuJ��k�
́{� ���dE� nU�	SK^\1�*�L	YkuQ;g���RJe=�ԎƐ@�Hj�g���n�m$8�%��r0�ZƼ�g.m�ô#ziET�W��n9�9��c�K����+a�Ac�L�e��$A^0�#����p�~6/���Oט���, s��>�p�5Dl�?�C҄�=�v��R� ,6]��׀��!h����8��T�������bH�h�/�NC�����`f�D��SY"u��l��ՙXN�+]Sm޶Y`�ٖT����b����=۳�G��v�YF��ί?��X�z��J�oX��R���8���E����D����ح�!���-����A0}Z�)%�:�`m@����I7�������zBq&����pW荜�O.@4��x�WJbЌ�D�� ��*�R��~�����9S|��z�������ނb+Q�@s6�j�߃@(y>X�y�ėo�	_x^�;�����R�ֱ��M}b4U�1é^E5���Vi� �b��ۋ㦦
� ��IdUd
X%^��\�*F};d�Ԅ�B2|Y���]'쒸d֞�[���ygvV_��^�@ʁ̨�(�h&�?S�iJ%)B��<L|P��� ��x�Z���p���s�TmI<O��DJ�A���{� I�;RA�#�oRI4*�=��r������~�CR�(J�[���F�Z�nG�´uݯ ;������*��\O��?%N����!q� `�!n��ӗ�s���R
y��e��-��a/�r���w��`���B+Cx��������w�ؓ��NN�z�������铔d� ͻ~䗕�'��=D�}t�dT3dK���o~��Na��,��	N�I�L��T%nS12�/�c��T[�2��/�8^$R/�p-�zN��Zk=4�nb���%���:.;{�D���Ƞ��8�c���}�%���ы�In��7[���d.��X��:��	N^�)�����x`/�;��Ee=�o�� �W�T�l�zB8���rO\>��.�?uM[�\0v�Mj�8�|��"M���"İY�h��r�c���ҳ�����)m�0B�O5�`�RP�-`�UF���y�+�SgV����1�/
�N��}����*�$j��74�p��*&{K�K��W�@p
���e�՞LP�
�N��n�����#b��ƛkad&~��/�������y�/n끖�x+y�ys��췐= .O�.1UE9n�I����wK孋lX��Q�����P��>T����DG��F���!�;8�?Qj�c֒��:M��
�V�Q�b=�9ʓ18R��@*���#�ݳ��W�r�h������9�v�9ҏ#�"�x��x����U��5�I�TšѡfEO1�-{�&d�����jݩ_��X`�Џ�P��R�p;"1wv��4\QO�w�
F���ʟGu�ozM�~��Ť��+=o��y� v^va6 4ԗH�j�s8���O_�6�]�UJB�₡5�.eI��8�>*l�������rI�+��&0�$��'�}�0������zO+F���^�>ߢ�F0(m�����7Pe��D��^a w���i��nJ3�WU̱&ʍ�(19VQe�'q�
�u*O�*肼v���<w��0��?[��IOn@�ۺ��W�,���b�}�˻_ s�Aa=��
��o�?����b�h%�\.!}�~�+��k�-^5%��+���J窖��;׆[c |�h��o*��9�i���Ih����]j2��
2*^M��bq3�H�}�3������{���\1��XV�Z�7NQ�ޙ̒����� �Zy��9Xr�@��OCf:��������apQi:�a��ݱ�|����e��ϫ h�vu#��J��#n��Ã��͊>�cB-"�F��t�|�,�.��&x���4��cŪ�>ϸq+folB��ª��� ��u��~ε|_�#���$���l�]|N���A���V�c���o�&�z.Ծ�����li����l�&HL�� �(|��]ȑ�aȢ�E����xJp{���5�l���;�xke1�.��#J���o#��(�l�������po68��]�\���u�\y�/�o��λ̫��O*���)��z�{�	�"�؝��y��j+�
U.�K�_l�A<1��BiܚY4]9�T��?}y�{^��u.a���3���t�?/��σ0�J'<���s�{�f��2J��Kx�v����A����6e=3�J�:t���B���+]$���V��;P�Đb�h`�8��C)\����s�Kꁜ&�l���:�7����Rq5�%����q�Y$���V
w����[�X+�U��&�����������S��9�E�P)#e�佘�\�X��_|��d�݆v��I�s;�����=�-z�\AR_�U��J�AP����}x�Oj������e��6��,G��^׊ŒA�_���j��K� ��Ⰾ�|���>�*-9N�A�Qm$gu_q9��y�E>�ݎ�?t�����h�j��Ej>if�+���*'
���3{���(&s��t����4���ybj���ʗ��PF"�#Bn�L)ĩ��H*�6B���WM�m|��>j�LN�D�d�T�^:˓���U�J߉�A4��>���.F�<��ۀ���=�YW����B����f��Bޮ7?�7�4���.|��j���d-�e�{�Y�x�)�H��rƲ��bI�[���������ȋ�\�t{|6��g��|Z������l]��!m���4_���k�U��v���ըhk\���gy�� c��m�����Y`� �ٚ�:�B��݇s�oa!�y��\���%9�s�O���nPC'T��~,��
"�D���`l�o���u|.�"3uT/!��j#v��/[�z�Kq���o�dROp�q�ҵ4���926������%Y^ 
�ԋ6����� �Ju�
z�W��1���8kN�m���4�A/�]���تĩM��]U�yo�h.Y������,�&�2��]J�Y��b��z:�F������N�訐�7N.o��LG.Q��V�#�#d����Ai���Go���%�uTGw=D5f�3�Sϥ�ALRQʾ}��p��"d�,ǟ�)���[,�}ߢ��d̖������S趸�0n�=7�����"l�����`\�Tc^v�+�gVo�b4y}�]�@��]�5U����0��_+��C���R�X�A�������z����@d�	'��?7�Ľo0��ȑ��\f�sY�Oj4�|�����_X]��ذ2#��f����J���LԻ��h�]c�>9p��h��2����f� i}<���7&�X�t,^I"���J�����^UR�#^ɬ<�Y��l��l�@ڸ!k^�V�dK��͢���v:�#/�g��R�����'6�PG^�#;-��"��P�~���(UU�.k�䞽#��������ɦ@DM���F�<4�̪�<�nV[r2@
d	��Ǔ�����|�N-�4�w?���Ѽ�et�w��Ƹ����9F}��t�os�D���z3NK���0�H��$Qx�y^���E*�Z�U�}@awl�*V����@c��8��r8cH�qv�߳�T���ep�����\ ��rKp��Z�`�����	{�k�G�k�K�N-2�Ķ���u48J���f0����|mw�)+���y����}պ{#0M���錄���e-k3%���yl����Y��?�X窼=ƕm)eaqNS?�|�Ы�ĝ:��V�I�P63�7�F����k��t ;���SN(���|�k/@�26?���~*֋�0w`\�S+�<�c���c �����/�����.�^ӎ��uMh�^�M�2��#|�Q�@3�j��sC�I[W��xH���]����ׁ��`�'듐o��@�<� ���bA��[�kށ������8kG�|����;�� n7�~}��&��"�H��\7ms���!IP)8!����U}#F6��>��H��op��,�9�_2rл`��^��vê�?0���E���tK}:����B��"���+�����Oq-|F����{��e&��͌5�2�����S��Ȅ&>�@��rTl�Z|��ܮ]|뛰.5{�_~e���z:���p$F���?>X���������dW`Q?�(.��
�>��S�H
q�0��R�C��."��q0�mgXz�֕X�q~Ԍ�ɵ��H�w{\��U��$��7��Wo�4�#lqK��⨴���Bqo��g�9�6��Б��t��!�c��0#~r ���y-�U,�z�(B٪��xE��0��xdW�D$lG��ˡI�e�R��V�[ę���6��u#��(�y�Nb��1��4���؇��[�qm�I��H)I�p��q��
#�6Ȩ�����a1�&��o}<߰���:շנ���땍�onK�!
00�U�zy�<â�6�Tq��r|7��Wx4T*?.yfr��,�ܷ��� ��A�D1y&O1�??m7���qP�T�Ų�ƛ��|�q�_�Q��F��w�=J���z4F�A�T��P62o�NOK���\en�+Ӧ�sKu\4Y!D�1?h?�r�NI���I0���1��{�>?kn.xM��s�|��-<�l�BoO����,���N����9X6�x���<��ǿ�U9S�+]�S��g���]5��@F��Dt������KZ�r�[+vCC}���LC-��!���Ƀ�ŋ�C��̑�F{�Zc����n�OJ8r�7���kf���A$�F*�pv��j9cjD8�\^�s�qHli���+[�fdk2���f	\$��I��v2#�1`o�rk�(	"��ka8�s�k���EH���H���ɻc�W���M����Q����&J���y=	��?�7mԕi�^<�߫�L-��@�Hb�i��H��֨/J5F�`�00�hࣕ��p�z�Ft0n���Ʌ6����d�AZ�P�7B��+���|=oJ)o��۠x;�?l�Su�C=�?Ec'H�|{ Ba���P!�%6�����n��;�Z��xcX0a�!�B���R��V���Yc1�tJ�bG�&� ���`�M.���N�vO�Bk�^�ފ	y�yR�K��/(���	14��̹��ӝ��r'��LSW��*+6��猚��Ǩ�yni���jh��o��i�>R�%	Ղȝ/?�u��M�`��0V���K���vk��%P�(�w�q�}n$5��Sb����q����t�Q�7֘����`̽����!�\��R�)��=�H���4<�l����K`�δ$���ޅ���1�ve�n-�r�Ɲ����g(<�������I�	a%wR� �V�W �b^0�1H��� ,����p��E;��h~�N�C��'p#*��ð%�9L�X+7�5v���}N/b!Z(��b�-���ʃz�y���%p������d��Mn�ka��>�	Y��(�hr)<A��s)�qm�a[4&=��-Z�qQE��u��\�q��a�"G=�� �~���=(�ʀ�)!�y>9�iK��}��������y�P��U7_WX��跷�oq@�mN�*my6��B�����/��q