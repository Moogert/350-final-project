-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
m6vNtTsKexo5YrGal9KWJdzrfxjtJagRMtrxgV00WXnbfIvwfrhuxQT6M9f5CQlIvCg+SQCBJGdm
mxIKnKwCb2RJ5Nlnm+NbI83q6afCcbkg8giJU78q4GNemcOXmx8abEAiOp8HVSMLgPFsVxvAUJDL
FW33IJuYwhiS9+qiuoqGVkAWuiAXjJhKsMAksSPGxe3hfpwjA+bWJoDnq9XohgXnVMAuJiSByij8
bDnWQcuMx9PXCK2MXyRGj0rpzesWhatWxYcOXZy5+gdYtORTWnzhJPH/Tp9T9mJjBpPyCTDF0uO4
CDRnxD+yd5V1D4QCepjqrHvdGUVqRuVwgJBQjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
zgt4isOwWZvM/IeZ+yn+rpKsdqYaOufUda8F4ZYifMP0h1L583eCk2tDoIm+YPiNmjvSwdOebd2z
3EGnzajXD+xEVSm/jgvAs2ez6rmavrQXGrjIL7KZGap7JK0ZcJtOln3tzRhDy7Ugk9z8rnMd3l5o
bWy+85VgHg8JJBilvdrk2/GMPwNUImPDgy7mgPgLd4tUOmhF82sFKryoBODOT+7Ih+ICJ46oFQtE
3DgzfNoRNqZPYsqMXL6GI94BEx7WBz8+xVoz4Qf7eoU7fdHI2Rfvrs8iAQkQmLtykjNgl8Lu/iza
wvPwAEvPjqDxw36omqbM6eT6i/INUFcrzWnSjOgWYZlX6wXwvi43Ce85Qw7bqDiFICsf3gD/3DxO
gROeJUlSyLKyu53rsw/21+9AOp9HhF+7bqpuEI8d5uEu01EtJ9/awZIs9zn6E/e5Jb3+9Yav+gAN
G48vz38nmoPjTVPPCT66GMU+CD0YpkSXModx8fydubZhq9SHX7ow+8+8VZ+3WI6fiEXLPT855YJC
rkAH61YcFMEYCqfmQbT01TCYfB6gRlEL6F+vLBoUz8P2VapH2mxV3SVbTINAu/I7WwH1fmIQzTIg
mS6Dt67w1UDBGJZmiMVolLPHPPcjjN7LlX6iUY10tUCzioEF0WwZbm00BLTrUQyacceLvagv1InL
7DYhyIoGYAlk06ScmloxcofzO5v+oLE3A72N1hK6bJSmcXgyDx0R1N/aev0AQTaytU/QZhbwave7
kDkpbjbHl1IMsP+c0Zc1WtDsfgVr7S0PN+fprT3g34cFHprj05BsoiAXPtFlPWRs4SPcFVo9TgH9
vRr+IcIpCJEPk3QeNdUzmF+FpRBGIQZrCYK05dCV96EIC1fDNUXxW3Vfm5bP5eQ2RWmco1ScmYMC
xArPugEPRR+CEORzn8kdUq2N6xGLTQClKd6ChzZyolpB6+4YpmRd7rHokZcGHiP7HswSYI0r95nC
YlcvYl/uBwxcrJ2diYylwAUt6clhsiVx++fBVSydc24Xqom42HKJ1EuU383sjZYSXZ7I/06gyoCd
Hk53Sz8qNep6+7BAVsy92M/4vBv9M5JaRudrrsPrYYODbNw3+p9yzJueEBZTIXhBcLnyetwBwsQf
j2UwsVb4N/mfIfPzWUh5qa6YjUmLGGzonJHiq3TydQLAX5nTcQLLiPEXj3HyFoqIhGu41SS9EwaK
tmP0YYp4zDAZxuY4AaIn1w9xoxjCyzn8MAMrQAw0EqPvUD1I6nzVD++WxeCdjA1ZUsS1Tggit3N0
jg09R9UUnRXcblLxzHrPgFd+YmBGj3pbfqRbf1c1hDttCnGmIVhUrNQ9itCn4wWl06EnG9hHu2zr
vcT5K7R+ElPXOGBzQsCMsuDLzhm7q5hreg9C6li1On8FZ++2bJO8QyYcDy7ePK8n/NbV3J1JdDlQ
7dn3NU74HCV2DlxqPbVEOjbgObG3Xo6qstvuNhiSkAG14CbP1HN7eZ6wKYS/1ZOuYuYqXnD4O5ZE
XekyOaUR37SooBA8HtVYCYL8PmYpoU2cHdMJSvN/Hx8oQv9JzON8g2RrpXYML+MWxdtpUrJbHkUH
bqsbLrzaDyHrqgqd4VA+Evv/MKsOQ7UEZWAJNMci0CSRICVxBSA1Hu70okB3IAAAP9JbPRGWmPJP
x0vTTdrIKtVH1uD3ueTrn1AzdE3P0bifzZGf1Wn4o/6D78TGXkJTALUvPHFhQx3I+df8OHl1XYZn
wjhIiHXUFGUG3/cXy8ENwGUQs3EkB6FnnwajDzjXzfbn+j3Kt8uc28Brswx6ovCW8Onjb9wEHFPH
EmhA1NCmiG1HfdaUf0ZpcEGhmOVR0LZa52dXvB8UytjbpNBT/gqL2ZkGR/GhXrRrYUunXFIr0I1j
H79WaqZ110I6KZPmzL+VAh6hR1gXa7vvmZ7Z0N84pRR52BitjpJ3iI9X818SPibrlzrnrtpRa2mC
Gd4nKewlhg1DtYpw+ee12x9vfgrFBieDXtFxtmjNscJNgI1BIgLDFTEfRfNwOreIeoAh23/egDYZ
YI2dSaHV0CYgFvAh1NDYCadoChjQw9arXcPG80XQakx7RxjpZgyoRBjAAcI7i6f46pgPhgUY5lfQ
YJAyGlroyVGkdjWbdkMpPIjWqa0BAOlzpVFEc7TfiVrJcdjJFwtylDdj/V9qyCfWe5S6/tcCm0sI
edI17C9vlalAh04ikhJmNKUaD/jwg0O6z8odj2PVgfFyccjWMkvvht/b4JqUQtgjAW9ne+aUbYh7
oNZHR13prLwOyf3/6Tvbzgu4HzKsusSMjE5MBziMY4Z9np/ZyE5XDlfoqLmNumF8Nduin1Kzz/VE
GCvy0tV06lVzVYnk0Jb5ZS0VXFI5AOUbnICNvIeR/dyAa2XrpFpRj0K0oIeascRcEN/DdrmGcB7l
2FeirDxKwG/HbYNutv2UH/Ce2T1IN8z4mC83OUoaF0d2AHW/9gkPiVkvYCx0o9hbzcylDra4U5O2
e+QkClpvf1Qb90Coqy+7bKu5rx+YQYMQ4VCZ3w+ky8m+JwNRRV6cY0N5P1xYtYRHbxS1VaGtJKrQ
TOfdyNWhxRwr/5uWLf0Y12tEzcWRX0NNEVk3jB2QwkTRJ9QsXAx6turwMzoPIdMQfNqBsgJI8Lfo
K4JIqlc6ExkV3QabuLf0fkC3BAtGepWxoi70COA6Ak0GHFxlr/GZDi+zjPOKH/kZjChjUtv8F+9s
3ygVYpV6NqSS5pX0pmxp5Merb06gCOybFtWjoBF0Zs1TNccxrmjkN9Z4mov54jz47pUEK8yZTx//
csFWLE2MXa6RUc/YDCwPcKGyrZmXqzku1sHcqsVaU9mOp4IGgNZS/DAEAWb1QItjYzg9FjB0DmZ3
m1/e/GXJf8dwOVHOE+Ne/l5nSoKZPt45L9l0zG0uEzwNKt9/P1s64Y0zdo12kII7UOEruvP+oBou
j0Ad9oua7QDfIjAcRossNMV0grqN1FB0IHpr1XoesYZEcSX39ZWLkCOczAC3lEiBZGmXxONsJZ9v
32JK4rbCO2pI2Q4pxLvPXQ9ggpOvuclRTun2O33Jjaq5yBoWDjkJuZyFhoYHanmwV3QtBQcp/Zna
6k+aQj6e7Fq9/djLF4LDOwImFYp6TpOcoOgi4R4/ZAsNiG3L78bi/ddNPpmcOO6qUSY2BEToLci4
n/rd3xQvH41aEN+tF0SY9oV/D5UnD/w1EV40EQM5tko2oesUlmUHniggJ4+5U4SCt0wZadKrVW4H
20eSdJ1E4wAifFwmLKyeaLBw5ewOLuAIKOUm73O1JR17WnZpPwkH4W2U8/AUPKD99nO65kBsMobl
MxOVScUj3c6T/ma0jNhx3kKLrK9p1pmTJzfBnhT6GmLEyNA8DyQ/z0wecQ2tlOZPPqqpKXlQyIAt
rq9lheIzLuT528GsMrgzJZIVQbvLU4nv9T6dbyBdwU0NJwjr3NfuFcLdGVBWK3asQ++ZWegOnLTS
rzCSrrLxVTfDGAdyjJ49xNofdEy8U7HEP/00Ety9lrztHdj8/usEwD3yoLIfVpgKRuHxnBlNJkUt
1JsPTGy7RYtIIXj9Mi+NpF3xxUv0YCAGWJ6FF9JbVPI4lwpyTGSuq5K2qSuJOfP7AG7kw2b9Ip78
UvJdJtLk+C0GASRusvDsStnxedx2W2LT+qlbYrxBVlqOMW3ku46zRnPTvBJqIMqiMLJR+bIfCwRx
S1whBsfZSwuQXuZ8smLinxfFjBiBNE6GirffDDRRIrEUVCQ9t6XgSrf1nz8ymcWaaiVetLQW3yJ3
takfFqhr9Z/DNTmDT8amF1MJ9wVxnjJ5CE8JBUPStjhKuK6cxJhBcgi1fHeqqrBNDhK9UESF0dRn
IGlQ2lglCvsqiwA4+baw+GwGuk1aUkgHmBhRFgDldEyr2XAmozpKSWmwbNKibSJmDqJ0olB0szfX
a6N7tmt4sChC80GG95K/EHsurSRlrs+niKS9/0Q81ETtCBNz+nFQ3IzwB4h0tWwqmGK+znjnKQoD
V2DrCD7OvtQvEBTbSAnr6dE8cYst6Ugst+UQy4MdEesOg71dPcC1zguSay20kxx3iaybNaOQ5E1w
o2SXp9ROnMa3U5XS5p59DGj77JnJSCSr0iAMt+3uGkmDojr5N//8Or4o7S0vfrGXOkTHFJPvuv5A
NELl1hiBeHO4zguhp5rxsm+wwEu6S1Ocn2hkoPmVv+AYZT+whAxQB1SSYDqBSFW/ehEVTnIqi5KG
on9+un+cOA/pFWbcnmYg9dtqOGxdrU/b6J19iCcnV6jF1Doj2g+2wS769uot8XT9vsmLUjcA7g8B
vmR5/4dBAneB2Rn5GpY1dau2fDVmK7kMWYsPiEU8pNd7B+8QHXwLKfbqJ2O5NQcOyY8hStz4oqe2
cjXSSY7FQO0oQ6nwjj3tJPC8mBUhf5RGlKblOJetzs6xa6bYqp99mydDIhCkjAVRb95PKU8gzTjn
geY3UuCulQhM7Cy9gbh9cSkMwTQEvb7NYB9YZ975wqw2XAwc9y6kRwZDpQ8DwKSWxo/6b/MI9I0R
HX4n+38mPLbYs1Coac1InPtQIUH+plxmCNa8s1hb2E6wfwum3tr6Kf7ZzjS46Ytm4WnUxAOikcWs
M9HzFpmCkcr3It4AY7ThMqdGzTeRwm/t+6NkQj6G1ZowwxhzcjhPXdUajYng775cMnMMsvkCR7OJ
Ukl+e955gHurj+v7XymRc+g2ms+tKD5TdZVTghUDNUTTv4ndxFJZZCZegUh+hEvdSSHvjJfFxsV4
gYdqNFOLieeblVaeO/YhA7ITvfZpAt06SJZoN5kiivOlBNK0EKaEq1LCKrIc28/tT4XURWt4gais
kDxjKoGq7kzd9ISTZE9QsOOX87ShaZwRG7Suo/9yxXDlwsu0kkbDQlj+l7ADE93QX8TYIZHPO9lf
RaEiuWa0EYcxkgX93hAeovFA1uEgmCMocGqC1UMEODwQhx8fplLTLmSCcdXm5I7sC8occ2vNQ7FS
gbazY4eOrL2pu5EBlms1SZCeh9Yy8HwK9dHwy9JsiuWLKxCKyx6bPBasE1SaT5ruO05VGdVdwAqQ
QQySv9wpX/4a1Ndic3COgSFwY8u6leQr97MfKpv2jDJaXY+FVY47/icugYpKZQLajmtzgTyxNZUA
t156QZ/qkscN6anC+Ti/PmxgQJfzmZDX/G255k+YBxPbVjf3I2hGtp5gSkw6Jvn8IIsYbdTrnjcz
TDgm40JvK90pCzD4qjeOSh2mrBOTtV4+awyUlnAua8aQ+COvbMeMWubxbeHuagDXgaJ7Wy+WGO5d
+ry3lYAmj+ZehT/innxnJRUsQVxEIef8A7QySUPRJ+TAvDL/5/3N1DNbQaNi5A0rUW5kFAw5jF++
atF79G+gAPRGQNHMUNnGf8sm03CG8nYx5qentVJlbXlO4hx3d0sOK3Gxp+UNwyK/bGg1fCdVYXHy
jxQ5GIG6nHAHtUbkthF0b9Ym5LAOji0762ow/WCBufBHzc6NK/kCuLy40/TU2P6OhDS8ohxnNMZf
rLPp9vqax3p1CFlx9nINT+9z9m9ZZKvzDS2rqz2Nj11ZjZnxWzc1kaoSTAPBZgAtT1OlgxynrDse
950axsaSIFIO74Y4q25RG3sGtgNTaRWCo4RfVgYcntSquZoW9dN+Ey2kHHR726m6r8J3O0mk52zr
SXUvmkqZxQ99aUZNCWsfANpWDQr51WvGFHK70YvonEQ+PvVmV/YolD6KOamtPDy/Df+JgMBHI/HA
fn67cwGhLBwqIcCE+ISi9C/G0kTwYZAYZxJixyJ//VNHR3HH1AASrotE+jbPAAYul+CQPPKvJRwL
bsdUsaHYi5hyxAb1E9IO06Ru2Xl+q7SvLK0WQ5ISFhYYnyhKiVuuEXQ/+SoOsZGIvve8q5hSxZiG
il18UBwOAoZ5n8oSyw8T+cbvroVadqqf6a98E9qTuWtzUR9GE6e5jgDq9rIfQzq2+22O2hQOh9Us
d/vstH4Fu2pOfrdfPPkL5v6ZDNHoQgherto+hb6G6DWJpjCeqgWK6jHPnebjpERFFF3XhZY6UaLm
JE5AqF+oUaJpHjmEvpkeZhDJA2/+yEgXSUuxO4hJdHtXOHunS7rl9vYneNW1v97ITQ/SIiSutYav
+vozhFv22kKqUd3wFNAqVssT8sBKboktFkKoVxEUl8KiHM8a3q74Q8rAcBoGHDZZKKnzQyvh2kKH
vfmYFZWKIrroDUjSLXm/n4Pc4+Strxl/9yjdAmYQ0Z9SzY+Hhm2GCTcjMSaAmNetTXITqthehmmY
naOSDyOHYlbpcinwAimLDR6TVEqdI/fo2aWyjTTPkaltJqIu/847mk57vjcRbWVeKEAsp/qrUna6
MGtOrddrCSc8Gr0Z1ylg8hjTlGIUl66s7IgBxKILrA/ed+CNoWpgUSLjWPnOUhH2+NAiEAChEvLj
n+tNqWgOdyUV9UVvVy8bk5M4RHMDgdY01Dx2B6dhrRFgpRlvfHoPK5/iHYlcrj9c+kodLM2vKohR
luJ5yUdp7mc3wpMGZX0u5MsQofqhcE9l09DCT7sLFZ8V7SxNmkZ6uDsvqjMkh+2xVTjIrhWTbOD5
4eHdPsKjLCZFRmcTnkI6Qtg2/H08LdnkT2UjS7Hq6hPtzWe/YFxQhrTVK5WrLJ2PTE5Z7avW8ehB
xGdGft0CWX/OuiXAAcyNlmadq+BuceOsB+txb1Uv4NFXdKmAUsmgKKxJb7YXrbgTPyjcFDocnGsp
si/yvAGv59Skk+kI8AlOPzaB1qJhOT1p+iH37KJuldWdUAJ3y8uS1DK/ZXwl8fWiV8SkIW/b21sU
c5fA6SQti+SfECjqyWF/fjoTUFCfU7BDEaYxJadyYD3RdAqYnujE+sS/6dDD1clI0Rqdg/5DqeoM
eviIGDmSgWfbAB/sgTKxesjXvEUy8/KIk9j6G8AQI50npEczjrH8y2F2FJe3DYlhtkVIcSjnoxYj
sJIxotoYm/Q6ZxF8NbHGVJSGrkmHCVoEumU8tBsOY2wbqSNdC9uXvadyT1lgYqlbGzKilzM4/Lch
8/GqGR4cYAFWuvGCgePB+x6mH1Psgh0lBtifjJeJfUet8b3E+n6bre517+yvpUFbQy0Y149IxuSY
bi6WlMRtB778KRixMLtvqYk4vmcVFQKV4gJo1w3RMEdaIvhFC1U6uJwZZEwRzDYUrhQrRzKaBY2W
H01lQ8BFLZOEEQ1k5swhYbheIYrNxgLu0j28LjuWM/WXPsTPvUMh1X0wGjEj3oX+uNWVo0Pn0M5Y
nC+QZJqFh+mFGqrWBxD/kIDEKFAaDlo7Pd5R3EIub/d+2cASoClvs0WV0f+YGtMcHmBaE1Dtw5DB
Z4quSbp//bFZ9MZE27TqFnQCYPS5shJ9ZWoW9LyIVEWQbls3CLc+MzKKxmLDwOOdN7CTEHkhXXVK
0lO1VYIxA/mbjmL2IrAQUgjlLpsJcJHVa20P8GJ6saKZZ2Pz83RrHOvbWCnNhNEyDarZKjoUA1Mt
5d/4qFwtbuJ6BhCSMj+chlaBenP081tTiZwSpTGQ2UZM31p0LHd6S1YIxZ4+SrHmsafk99ZNQhqn
fPn9zrneyN8bUYAlr7pZw59I2CSpE5LvumPsvuyreGdwLQ7c0Ih3sXhECkMXNRUCN1hteLovViyd
VdJ/QvCoEBXLH/QXUMjLugA4M9TST2drt+sVeAmLpJzz74AmVgjIXsYY6wRnMuJLf4yOj3S6jltV
yU47ISyTVRobNrQqS+hiDVLrXesQYbOnlL2Y3kvB9BQ+znrywzfQuCNdbxQJIJUf21Z32GAUJJQa
/1AqXImHC/MrimUnYlx814QjHaj+9ye5HZIW72NOsX22alzOfi+Ah/K2+fnabqmsfz36PFLPVUKA
CZqxpIosOb5YddhN6Wf/K/2HFYvwLjCarO7VTRCRtp+KXUbu9ZNFbNtlgmDKgVsV6HzMhWPhncnM
Az0ogd1kC0H3Jk9hO9Tfrj3INDU//GG9fUjHpy6X8dPAdyez4WACjm0eH2EpfUJ8edpaOil19FRo
3qDKKdmRP+ao9Iul+OQ93dbN5hQ58yr3G7N1Kh+1WSW+87E3mVeePGPo+rkCRWySOqqRyuNPitUF
i+K6VtQM5YiLXAuWlZwvH8Bv4my1f1cOOjQVQ5CmfmQpliNEXYIh9ZPogPVHwgJAB0pNVlqVtzaW
MtxfeUKk2zrtj0fV/GDJR/f0+uEQ2Yb24D1p9ZkzcW08Xt0XiaUH/xmAGXW1lJegNcFyz5HpuCow
u/4fZPWNmoBoeUGoq8fO4OfZgOxowkdUQyPui6Ozj3Q9j8OUJMDK0aaHK9vJb6iUZp/Zv4ctE3p/
niom6UFpAzQ9o6mqIPOyeocn5qQuT65WeJHkJljkHqiPd3tUpDk/tZq8J80e3QMwsP1na2wPKFJ3
b97atKWmwOiYrug5k3PcmqJmq688O6H+5VhKD24zzGQhGIopZ9L0Heb+cIE5sxdo2fhMh28CcXLw
0AbSPlp3PZfxYhKBtr18fOhBWZyEXRkfa3EU1CLfBaQn8TkcRaj1tTrFSTlt44DjENEc47snYDgK
a4byMf71nWxQtJKNOIMUwRhSpK9KyfvOmE8EvYl9z3XSHYaMY9WdXjqIX0IV5ZLJaBOea+PMxxGZ
2G3ANMk8+Q5TW2KjW9RKlM1TPoT3q6SHh29kZved+jGNZs1OPvuM8jmdGhGG7ASfUfjw5JpNM6QV
6zl2bdTvhzbugIBDwRZyVjrDxuJuSyi65XPLhi8jHtxtIUjbA/U+qFnvZmMkKlGNV2WHYzM6wmzN
dPBr+THVHgkIw83P0e+iwZzNllnHmSKHDt445R53PuJ8zSOyJTbR6DvD4eWVEYgoYf8KSbFEaXIE
4HyHF8cRDGhHhqTfRiRYG96Hjc8xzojViLSaTbTnby894h0FtQdXqLNhtIowhMJYxDWi/TU0TBgu
80UHxCAhZgm8Y1QIscW4Hm0faipxztmCfAonhd7UXi84g5khQoh4RH5HbhOhs/60Ip7gnoXOVGG7
0s82cqvyC5K33k29Hi4rAWTFxwElEusXhnf+IjcBQGcWfL8moSyUMtOXBgfnFjzf5ovIRn5/kxuZ
HuSfmeYOXHSnpxPm/aUDMvXpiiaa4Rl0O7q35r1FlxuEAZ/9bH+5t0pBFUxfsUrmfbIuRckGu6hq
HDvFlZbPsHzZrT7LWbGVltxnOiV5l9KHotxrrrx9qwji/GKDJEwlG+pX76IXu9cIFn/E58L6DhxM
6SdtvHnWkQSODVd4GYCH8116oE5FCMJYSU75H7EiK22V/2xz+zAon0sIsU7q2B2bCEXmwfaBN3v6
Fj+ZDXUQwEL2a4UoHzPTkqiM6hWH08z34IkVuteWQvtg+k5zYgV8fV+Lf9ak1961WMY/LrydV5az
jRyshvGWYeNqkNYuCN26QawfeL/FZQTNcc3jzL4fFM3/JPXBr+GXB6kibhlRcArUtexgl2MgDZPw
QOPmaDV4MLmrphD3OrOhXwDu82d1+tbAF9l8fUd9xAQVrq5CFWMinZW6vmJ9HVcprgi32e649ncC
Fi+he+nu/hLtMYFJJide9+o5abRwEObM5ql0KbhPtd2DKbOLEYcCp4ysQm3ikWbgisWK8izIqVzF
LfYg2VOhTVWbSPVCFn/bGJGYOg3xY/G7hqw+qmRlgeLZYy0VkHYrZRESxA2Fu75+JZ9ps694UllD
aPbmpjOm1Hm/dAHQGK86duHD6ciCUz1AY6Uo73X2wnWNQAwvpOdh56e1aN3rpMVD6Im9P4IWJNKU
Eh17EjTDzjb7CDbY84OOFUp8cMp13dw3Eh7uk2g/xygAUl59tlYUpn8rW1WoFXtF7uxgcvwGZK/a
7FOPjYh1kMZot54UyVQkQK+aKiPABbyEvs5FOZ+5Cj5fcOGr7TUPT9An8mA48b9VWvYyZgFvvcnt
msBGvQR9R12ogpLeWDPmTC4qZEvWz4GvUgTeHaIxsSqflq1T9nU3IwjmS+j0h2ep5y2g7XXsdJuF
/iKLD0T8X2acH118/n9YJvwnaBhL/nionj3CvtSKn89oHZXLwbQb5Zr+52cBZIRuUXsgXmwMfYFW
WqNmlkcBRsiV3fJv9WXlZNjJCRfE7XQ+rLJnDy1aD8RYTQ7f0AHbTk/MAQWmLwR3ZISIe487cuII
YWc6/XmTFOo9W9BqTzFJNOLh4GOnF86U2PhsY3p+GMndC5YQZayZPh98OBm7Ow1WH4rxBbr5PMOX
WO9pQkcUecufvV4PDbOJl///ADRb4xwnJbekI7UtFQrPz+Sx/aW/lEojl8CQJgN7K5MkrVDkjXrW
zuewy3+otm2BpwWXnZv0tudvOBWikqpH2zo2kACtHnZDzOKc1iwFur/SynqPrYrEYmKWQQWU+sTT
5px9MMfR4fpN6AiKxBXF7xDnXYQXxvQ5Ks3Y87JuibZcYSzcC7V8qN2bPwUsVP0n3u48mDk3A1kA
G8NASnZnpNboUrggVj/cSlcEgAyEw1YnHAYwFef1fIuC68PHDj+URIyakIcRFxN1Bl7ZHDFqwaDv
//WyFIwPCKhuTG9E3NbZKEEiBDx801V1x5AIWpEWh+cAxJkYaGk5sJ+5w7rPrFIrOWGMKmdet6O/
f/07XzXW7IpgZho+ZcFFlZSRQ7dDcS63wPw1zIJ7H19XidxGRT6J14BYy2WAnu/wYOnoqThJEejI
MOPQ6n/mQ6Nks5k7/z1b2kVpGoUM+4rys+gjGNB8bYjovtHT6YeG3niDX3xJ1hAXlbaCE1Ybj5vE
PRkTrj7rS7Eq+5TghMknhMjoX1flgllO/CnykKp2mpRULpDeDOy7hsq8pgtxrB4hfZRb/LF4Gn3o
yc/IoZJ2G9w696c3aGICBjdafmJuxJB7kFjq6/g2f45uE5J+w6uRE+Zl5G+4yzjtFEH5n/UQQFDa
cFTUa+6jIGkxinGd0Czkc7c1hEr8TdxG7a4OwzJ9SP0uMctw17+MeehyjsuSLN0BlmtPp/8ZO4EV
2rdaJJJONIJ4r1agBUjbzZCPn+efTa4w37042IY9lWrbXKm8lS6736NQJScDZF32ZWsQgwIc1YIE
39GwcxxRQafSv5cZX2BbwvkzJFK0/7vYyQjf29vweOLsFLHpq8s/orG1E8I25B32BO+M2mVj9lXo
bFfb9Cy4M/1kwl59Hs3w9lJwIaLP9i+bSk0V0nmclFaH1jXWrpPPJe8ImMmJg8Eprfl+wEzLeSHA
BNl9P98K8lnxmWiP4FNzPr/sRbMVV7ja26/Dpsi3zt7IxNcEP3P2MeOLGbGHg00y8RoB4QCjxhFF
UPG1KUxjdqY3Il7pZah8OAyDt4WSa80zXUMvpD89b2A2nJQ/V0Lm46kRCuq5rm7/rCy4OeRAwXG3
EyQDfs9fC/GZ098GrxdykOTNkuVOlPkGBAUugWCa95Xyqmvmcet2tC50GXIBE94RW5j16WtIlusX
CuBcwyjlafb+qMOvNROpYdlA6DPlkH0I64EgRGAzDS2vaHcfCvAZ5RNUJJLPtUhZixFrMElucllg
qCr6RJOGqZxSvbf6W72qvOuLzRbzHuaxcwiCaCSWE8uLSSeQCMxKZhFHTNGeZc2bQvOTdgrw0Lhm
+B1Mn1D3hKMRzB6V8sSZdaARlIomTdQngazC/ZiCDgG3XG3wd74MnBN3JhroJknASyZgr9Tv667Y
fMyYBz62Q/YAnBZktdgQmbgB5FGh7TPKLTn/pgfaYKx6VweRHucwRIdXBM45CiS/yyGS3iqeD6h4
1N7K9Qw/IbYiTOwzwnEgRwgANbPcRzC9UE7a+XxQlRnDaGoi5p5vOlB5beXBavCzSAhGRd1AYhYn
YknGiiQW8PDemcjhb/GCwNulST6qm0oPYK0LaZgfRNsmqCFUSNLPixfzHu7G4adKFLssIoZrcz9x
jo5PuPGpNn4/Tu9fkKq0FsT7aUWFcT2WYeOdoCeppea39TVx10g5y48JDCw8+sAvp/1HrX/5W7sz
90x8jHdO78+42lyBZ7tCyvoZDz3wiiIHVK32DDlPQErqaRVIg0LkeOXFRdiptPd2wm6YnGe85H+C
ushAGLvyUexq+Hm6H0HxdsNbvdQT08q24VyJnsC1OVTZEzw93H6Kkkdx5xyQ7nMjN2t01FuI6lFl
p6MOa2M42/b+l8oUD4tJJ8VSkI2jzG06a73jhybUgUmbrKSFcbbl13uMNrBc9j8+JpJAYSyz8c5F
8zjOrveI5Mk2Ka89WpvvVw3BBa3N2CvZr6HKFqcMod7zrDuMWPha1Aux/J1JowHxiD5K/55EmOpM
c7AuTk5J85EG3DTwFg1NL2YWVDxI65JUNp7Gd40qxaSpnVqFSkioLaNDBcOIeNDn2bVK0fuA2oxu
KhyapGkixMKvNzSmoOuiJGGSG79+9flfiw/lurfJ0vD9NgpOI5zSWUTkq1tpdqrw8xAT4XUdWPDy
XvUnTWXPQiJ7iJIwPIoPi3UW3rAiZ3obvEoFyyiU6F5HxujgIFv1N2ZJa9nffr/34VVVYUaBgbLE
NH0PIrcouAt9iIP5Gknq9gUbuhPxpWLji3vA5S5t9+xhx7F5ZmRPY2yZRpCi95+nXSOQ5oG+U1Zo
mHvbDUuo5ong1Hc3F7F9Gxdw7wMusL8h0pxVVRs9K09SjHN6FKMzgppnaiU6Qdzle2oN511KtsNb
W7I/kKWpiAM0500ZoJWULzhaT08kE3qSYFv3NRG5KRNLN+/R+XkyxWDeP3x3TJOktSc3/XxdHo5j
FDoMlHBkGAma5MyJg9GT278Vz9XRywAQYXVE7Y49n8KlVZK2PWqJLHIR9V4ig6eyUCViPu3PPYT8
V2nNK6v1YNyG+OPCf4TBuN1dKiO2bvY5rrNTk+GfR/FUis18JxpNmPv6iogMhjNyGzLCXc9u9VsO
Ad1pJcoYiYHXP3q7sFsqG9H4j4ktY5gKD6cbpZHM7uXkYbB6MUM2UmwJ5kNXVE9YNELwec9/xlnH
VJKtcfhtnVSKTnipytq3afPkERHfOyLNdArYopkCCLK124UgqQp7A3vPtUPdzNwkL1bp9RGqtppR
Bqf+rAOC9hGa+sInpU113XZdzvgeiHR+rvDY/osCJTv8KErJPNbFu+4ncxuFhvRtJLOBSWF4NDs4
HUhvYsUKG8wqP+v6et0W3uO6J1rg5D06hp1bIkQJh3fHpynEmeg+H4DosQsgHnDLosvWBcPDfmwG
5L6EaYE/l8DG+RdX7kHK6EpKKWO6aIdIX3VV1nLMOHmdIV9on9qw9SAUeD6aU0CwMEGpJFUKo/Kx
+H1iG81RMjEiCjO/FYff9tWH4Fim8eaBpnmayJzlkwB2HRPayG/ZWoHJxQ6HB3SsBFv0/mBawoq9
8FIyBLm74XtVwbIXx9nhlO6DVQbfgoenJvRK/6bX0fGd2uH4tOhDuDLeCfc5Pj14TVxZ+W1WeK5Y
z1gZy57KQJbxMhQlYpkZuICPpEpLU5Pz29eRXgzrv32rp7qtrrvdGLXFiz9nSZIRrQ4EzeR+wrNV
4+HfPx3xHagle7pi38/2jsmDoz0SI5CdjCY6+/gYXfFJkrBOXkWFkDpCae5BivDNPMQYGYxCwDnN
ra6PjpR7invYwcKkkuY7jf58RjesNgW1JBqFrW7Jox53kJ9TWZb/dBcLmQGzAgdrH4vmvRR6JOZ3
+e5Qo4MJADZZ7UIrx2SRnI+JvLkkR0Razr30uXF7RAqMiafdCigOvvPeChQKFB+mDpovC1usQ1mr
XBTSO+zTAyq/BBY9h0fSAMe611QwpYTrlQEsXP4q+wtccR4AU5vw8x+PhPtD9xxsNTNbKeh2IVZm
zyYsgc4pljHTW1R6hvkpvcEP03jMffHfOozhAyKmkDoe8R/YnMsFU7fVsOr89mONHZ9vqsUV23kT
DleRS6vHG0GctX2uu+x7qr3qsU4GTEZCKYdiY2U4bK7FjMGmiletS9WDaw/5gaFIavWQsAT+aVxz
QZe3CzyRFIUAdBuWaM/Wng8JrEJZZmPEKU5B0OK3dS03V74pH5Gr7nJmnu2S6ZrQ7Yd1hz+qBi2e
IkswWNt7wd6L7FWxrA6mIHoGTjzRBK4JCxEWGnpj0aSrbj+H1xFc3xPDJ5pa1fpyBZSE8YbpnLJD
uAIxj9wyN14KxxD7qCVvPHB1dMihiYgnWegBf0gekW+KRj7zntwWDNGEuBsAheYK8Rhugn6klAwH
458Ab0dzFhYhHkRZFY/RArHA3uDR8Lho5rpsSk+ABRWB07QLG6DkH82DtG2wc8pJ6cBofzcFXnUK
QheBVfpMXF1sSFjjSTuNsmNtMx5IZbyJR7+OAVoDfrMq3WhHQDmdOcSWni0/0JMMxRmmBkoYvVRf
zcP29RJ6/3mZMsPBjj/HINtvpgEUjqAEEzHg6iJaB4Bl3VaHTRXTkzX8bjrLiLxFXZmMokcvlOUv
vQXH0orWbfdu0e7bS7DGGS6RepY+HEQXYNArBM8Inni1GKCX0wSg0f3NZIjX5OapcfD2o1peG3oc
uRD/PSpGoLDGpT0+WMgJG21NovYMS6CXWVL1t6vWsUg4PUUXQbkoYK6SxRbM3Z2ugyL9DW0E4O/C
oW7CWedI1umyASWP4U2CNJRpo6BN4WNecl29u1e0WA2S7GxQDuDEEYCaHcwq/zdGzmX0Fgs6i6vl
3lS7lWDg76YOgWpEH7p8+W+pGPRPbwZwail81ltM4Aaw6kHLrkULDGNQlF/dxh6xMkcIVzgV9E1z
EnvluczMdv76PuYOZnabHsa1Fhvwlv/tuSfQDyRisfyvLDhSYRBg0s8qsdrowZcmkuPk9tGH8tSF
C0oI15pEHmry8YgBmyMdjakhAwZMLAdmTgcH9VcP1Mr5F0sXTel7EtoFCarpjzObZm3TU5RKVHNZ
WJmI+Pu5P2ZVTqTr7qS3yLn6HX1LNJC5Np+Jl3NhYG7uysY1AKmg+aaMS4xsiqpOU8Ao+Oo0IchZ
1iNrf+7AB8LZJrUbXNDWLVLz5d81NaWrDhxYozx6cltG/sHIxBDgEBzoruiNGW3TeYUzQ0JqV2rQ
bPD8azDL9kaI+6ueFDUjsyF7339cPxkaI+wmGxcnJViEmV8YZ0qHuj90rlh3HPT7cRSRHvg4bgSk
Sci8xVEIBqPDLeObUr384J3kmitIt2ClV9X1GwM8KkPyQ8nhVyu3fqgMnG73qxW2IQntfrLKBMhT
H+aPzshbzQzye/o7RbyqKwyhQipm3NJ2RWhZXXeffiDuOvjaPsxtI9ma/PCZnM3ZrcEZBoa11oid
GXn3gXhYF97wxdZmR5/JyyX3piQZZl1CwQbwFDgYlmBTLb72PhgS2CyB7xChVQG5NGMnSjtTOdTV
ib49tDxHH2B9XfoIpiC4/GnzKX1OTHITPY78j8iipKOOb7WsUzvMeY1Dib8uK5wTBt5kXF6uw8NB
Fkde2JdqmQNwczee1R5FeLgHqo8oOdYSpZE28yoNkZEd358zH8uftOTiwOi80hYgdLt4ZsHPV2Oh
ckAK6UmHAnfyHyboeF2LEIrUrVbld9GfRFRk38mnUC8kfEuoinXaLn4Q4F19qrqRh4hFoluJb+DA
ba6amPCAowXZlmMW+ch/6KwROOn49+n4XxJmSL9yBLyYsPAwGzun48OvZTX3tlJgVRzVpfqmrwB1
AFCczL2+daJJ9TROSvfWMbcVWq+5itSflOMsNQvk9X+w9iMGwSswqvpF2naNtCOcJxKsdm5aGCbR
8bPHktNFuN9cN8pd/xPyMlnmNgkz6vhSDxQeikKGslnwbxSg33NGuk4avdHp2nfxoLrp7KqVMmBg
Ek4jJIIUuJ3yIt9tVcLLbLhbha8rY8IbyRQIhaClM/3xrmtF0egSmIhrcK388encEfwqHUu17CiB
vXZKCMZU4Dl6HfFQE2c8syqXRb5yvCosIXzi6jjzwaZChuHDE0bdcv8T+iJ4Tz5dEtXHeXBq4mre
quPnYuBzbbuoy750iyBlGlmUZZ8qlU4CH5qykKD5MCd3KGTlR4oRHXD6y5Ls+mjeUJ3/wix+buUP
jsJUkSJuv5abJSq8uQnnZkM+QnKtvKtue/euDODkgxYiM9v+MSfdurxhdVt8n4XgYTRcHc62cutk
t446Dcj5iQzdHO5U3bVep4rIDbv8XtJfppS9UYTFTJkQRDulp0VaQ92n8l1Rr1Xo8cnfWgXuqXaA
HQ+YNxkmPArTNz++Fc7kGJzwQtiLAHtGCjDED2fSf4/eR1HxgwJGcAOVJMHXacfClSrSmEYHHoG+
DucsTSQve0YjH1MoAvEEOWyd/WskPVgvPoSlo5y4q8PGjLdXHa6K1WV5evWYCEXA124dEGwJuaDL
1MCDKMVfy1aMXc2jmUi3MSXhIjbGdchSSuM2YgtqUXgafKJrrX00vhKbkTrdf1/uvKAbYEtzSuqv
ngXKs2ynFKLRTQQcAtruB5ptGksyrIOmjQdynjVVzIzai2Qy0FRjxHQp88SSwsGjxnkr/yJyCi/b
FWW7+TgG7oUIiho6TkprcdcGxcZlluh0HsO/LfLwjjtuQw8n/596z8qZ6NaempVyhcebqlJNDR6A
kKwqSNunR8VuwZFeMF1bZq25i2r8OQRHBnHviBS42zTKjTLmBjw2rr26tmbBdrMy2fKHI0HUGQB+
OaHxYJXHB3R5CIpJLFiqe+bTIjpxZ9oqPjYM7Ob1Vr4w6ZuaSBwU1YMTxKJsslfHcShodsh9yK4C
B5HxuvFSETRqQ/O9EouMogJrD6QvedObj/4/eoleGYXmfLmm9V9KYU0NZIimcBAensmHrCcVTCt7
NFXCpK7h+5ffCgQIOqvfuz72tV3wNAlvm5t7N+t9Ztaht0DCCovWZCohk2uaO/OaBI6qdXz1Vc/v
HhLIQFKOlvJc+O1yIXkXiPDlHzpj0GwFJxztbjpIxeJwlLBrDRY8VCDsM9qg8NICDsH7pIGshYtr
DW42eIAASePNGqx5rDUsByz7fjKJjQOP9e5hqjXPREpnAC7loI3O2yFDIz8t3FUmWtdqzxbyRcKH
dF4lXdsdJVvjmpaWJkpHPKb9PANJc+fprJjj7HmZTDaSMQ6VKKV4pGk+g03cTndacNJXFy446GqV
ONRuYYgakZBo1yZIukPDcf5+BH2xj8/xfFoOTaalyLHBb6nMipnJ6vEj8mhC5f8ved8A2VDKt9MJ
K6r1cEWz7sVISAAVCNy+SupZGbS5TvUe+83TTMNwwZLhIObgaBY3JbWB+u6UUGGS52X2XgtaAEhT
1VBAjt0b2hN0pNeTzyLO4xVw0q/WQTMXzHQhrUS+Ob0ZI4DMTYcbuf98Y5y1X/Nuf1HUn7S/zEld
tEGA0CYWdDMPW3dIJxtRaRcYc1+vkrsq3xuX7k+2UZNZIjcw8+EBXlH4TuVwV8tzz7tMU44m4UDw
RiFgwVDNdJ7SiyUkqr4iKZrS99HHuDET9UgTPZqNq0IAXq0NkYlYB550nMpMWlsISAkotflBEVqf
VdpynY7DhQhzzfBNTJIltYLT2+hezmgmagRmWQJjT0ygh1wUI/+rd0hznHyahBcMaWLQih9LTUsE
WrSw+513zmyq6L5QWt8EkDrwSUQvJl0W/RcxljKJkM1ZB376WdyyBCJi643bxHzXIcvUOEdIaHnM
fB7ekANsgqTHas7kG20geVC8+xjvQTx6YSdzXURNiEqiDt2ZOdir0K+UWgAi4f1RrJD1gCTzTpuW
oszhCwTqIn5BpfCxo+AArwTe5+pO7N6K2u8y7zXNZCelDCH1xnnItDm4C0uz2116j2Yf+wOrfgfH
QgETNaMnflAANJPmC5gY2F1/PimlQFPMc8yj8zopTFWsDY8RqOqc0De/RTyVQJJDsvc8OHy7tZsE
K08aNd0AhpHhd5+UbTt6dX3UbKZjHOh6SJqfxrzZwuTpdSOlEs40/gHH4tga8qI1UgdHq1BEcR4l
5kPN+lIDFP2cBNa5yNt+b+ygyzsqtJFWIJR28ulR3KzkxZG6a6OsYVCf8A9rqp9fTknZURZxyiou
++IIZU3RANmOn4pjZnfi96bVPtRuR38vAnHNxv5635IGf7kRJTp7KWU+QRD5FKQAdC8HpoNaBfuQ
HRMZfigKVEdSuu8gQj+fhZVpX/ioOMwlYdGGe/YcmJ5xtm73cmXKjbKFtMl/SpAMzyo4kvDhXTyC
8pEujoNq6IgzS3Vzbe20I4H2iX+p8Mh7xy88A1sqD+tx6x7SSLSmCqQc4M+PklK/ZPw8H6MofVia
kVRfTfZamTxWhzrvExEggYilFAKpneHfxbcfYLSM8IdY1Ez38+WSPHXW1xnqWB4o5JrJ8xbut1OL
Qbv+5WLe+7bUcoWE8XGNvoy3NwNs7rTwWvEOCI7C/1DzVz94/wOUiITaleoNfRIQhtLGSam4pq4t
GjN06DiciRym7b6gIq/dtPwkvYI3S9JgFs8EoITibrXSyb+IAdAPmjDmd9Nk0egZbB1mYPvjOXVB
XBfEvTvm96v1KloV/wOLvXuOhDeMQPT+aZZF42mOZGzdZPyqMe68zcYQ4QoObI6Me3T4MgBO1A8W
tUZX0e9HRc9teAQP4tB8eKC7JHJME5bPyJs3NmjdVvfB2ygZvgxwQDKxgrSNy4sWiXFfkY485gLj
NTFifC5/eKoZVPnXTTFVgV7+7vvYzDi02/QTlvQ3LgydNtNq3YgLfkMNylMrKf6UJbNtRxapTRxJ
WfQygr9KLJCsEZ6aOwPKuhGTBnIHDQwImWFUcpBcIUdn3rRH8qbW0nNwR749QuHwyyZzFTTdA3aC
7O7UkjD/Q/bCvm8kmEg/7eYbAIs3DI6C24xoRM7YLpoqfqmjeb1DkW3loH9e1nCPefg74gfFR5Eb
jJp6tfs+bXzNObYX+RQm9Bt8D93g98/YtPwozz6cqP5517UH/yzI0W7bba2bAlQhHlsalo2f8bOK
EnM+hgm89DLBkB8Bp5nhVqbrI2DBFX1MN6FbT+ieOgARcC7lQ+IOlgW5PC+sw6RkmEhlF4597wCv
EhL5F/4GghiOEvQygj40mYXwcRKiyGze+7QHxVEiSgp8e4l3Ra+h6QJsfw87Fo6MmTyak5BTqcDE
WSgOlsgZlBPDDhwM5Ap1Mw4tcRL6WHGV68rKKEJXW4BIMv79UNV5ToAjSZsZv2OJQv2WJ9CEhice
boyixMuE82g5kNePCi3CC2C0DJD4c2+BuIRZk417Pl2KZYgML0MAgJ9onzuUbVpXpHxXTyYwuwfu
T1s0cLXR0Am1LX/frpBxSMm1Im25gPkUdV22isPS8XqhS+cihmHCJLffShjdVyvfuj7djYCqg7CY
2b7jMAzMYs+qYrl0D6/xEmvhLYgYj8jC139oeNMjB5H1Du1Q1ihwze83ATy+UXHNXFa3TODKujyh
kFvZBTsBEP5vlNPSB2KPDwsAvub+QDWHNh4A5aM/jSAlYSZpzT5kYF6ra3BCJI1T4t05UghTS+6p
KxzITeFVthIUd+HbPvaW9PJffrvvIRrm4IITLxSFFv7k/ClVdgVXbhCAeUXzcWfMrut1OXqe94/1
L0XgZPEyIyTG+BUF5WpHiIh95AMZiRqONGDTxcHtGi0Ck71eTEFvXjfeqK34SxUb7LMakEHLejVn
i/8II0KDKycA/Rv0rVUDa2ar73dHDkys/0oio9mscyVtt78HG67hXSoKQuCBsME9z4+THHV4DrFa
zmvqDAdLG7qqbUO+SxTFDsKrf1ZIJOY61RaUop+msPqReCXLH5OXQTQ+FJqMhT11R+kuLfaMxeg4
xYhJAWJLOP2OIVMz59kcA7GPIDc+j7i2LCgwXnVYCyHbCsbE8MzBsOzWgT3y81QW3TBGH1sWA97J
NLcFT73IuDnFCXJedCof8y06JqtZcC+Nf4hk+MiXPFoqnio/9ORe1cG0OXn2DitzkMdSimzDRgkf
TGxJG6AamyXj5Cw0PWITMrRyVicPmWT1hcoMXPAehAqVYVn2ou0D22EAKAakcZy2O938J3AvSL4I
HkhPJDRAkTqgptjGZOtVRng3vDPxSqQ4tJnIf/ij4V//vSi1ZQlrXgWdnpOisqt8gTso/PHUcfzX
wOSAJQKjgFDQRUhGM88QKWdhNEJ7EXfrowihoHpKX9xpvfmJoA9o2xnQf7oPNBRxNdsqaw8bbUGd
/HbzWEBZVkb5IHD43bscGBHZ3zoLraUYzb7theIRczxnPLDMDZpJGMwJmw4TQ5UgXKERoc5RR84I
He9E5jl0bOaiPaF0DWlC4cnwTNWnzqcK2HJBwHrJpP/wzdpG0enM+6IjvQ+IK8BbZsXb/VGsnoW7
/2JYwZwo3mEYAimOQoVPHHWnBENIUsEe+1abuOFtylIfSF2hIvaHbr4vfh5ahTwKJss9+X1xDd/u
W/6ggecdynXbieZW+Uf0NB8A9dBPN/CGzmBGFchoJbVP+EecjhEt1J4UnMY43JWHyioi5nrIapHh
w49jvOUkoKKy0mdNw4PtjUQldrDVLXFvtVpr7X6FM5YXWRJzwCAOLHUzh//DiKi6ougGMLip8odQ
KaRRSmIZmk7DK8DKCXAROTW69d2Z2WyMycH5KffyQKGGauWy40M4nFYcoK3Ho/iQzlhVsOuRPlEz
jAfLEcTq/Lsnw78x4p7vjY9JXoS+MPvyrVAzfwj2h3pVdUqpsW6JC8BvJSHqDgA2tumth40s/tK1
1HsHBYHPOg3xiX6V6Uq0bckqaR1H8+JKpEGXVBl6aAYi/5ttRaR4ikfVp8mRqB+o6mhYNXh0nwh+
RxE7+jrkS5Qma1fd/TI1VdAqpYJSuPMizXY4/S9kLL5djvGYZZlSTZf6pcdm1UYFJyOo9dXY+Eu7
Z1sXazwEEKAcFlKFyEm9I4H748JVsALLiNAl0ePVIrfD7YASQPUy0weZx3v7fS19IXVaS6ugehHE
d+vsK03XWltuHAuAvdl1XD4kbwpi6an69dLeYUzrAFGQb9yWou1r7K7NbZR4tEGd9BQ81AaqvlEU
VbJ6VdTAZJaW2AfKHozQvgVNI65XIWlv2CsP96AbF2HernQOG6HTZj26bwZN0GH4MV9KulIE5fUe
3rJcGj0UuY9H2/wbzTGsZj9V3yNeePOBoBKMrKJck4aPl/5bTMRTzxau2YKveze6JhKdJcsDUCAF
IZfx0NJx1bmRuPIste/ZjS1G8lny6B95AZt5GFTmqlSGgd4VctE75JNejyADjvCXvBRZCnwSKrQB
JTMTbHjnPJ+C/hopVVSPLil6pVI/V12mK6JEdh4kO7Qr8L28LAnUDZgrRZNSzL5E8zLj3cI73IF7
6uxrrojcbUfP788StC8QbbpsUgTjopDVtejpXEjXlDB7ykCwnUl0KUa6HcW6X/YDLxKhrgRFa6Uu
85jSa9IMhVMhJ9uDA4uF9kuFshMYDqNeXfJxk/POR7wbldTIA64XdgCTVw1CxL1uTDccw26jY8ls
PSobymEsocZEho7gGdiitNVaXclTpGxWhGRwuzmLvE/2s/EdfSRKzKJ06+PP735BXYI2azpz/e/Y
zWffAOJ3kU7u9qF5tTX9OAgYGrfiUQj207zBBo5hy7/x833NKWhCqct/zBVzfuy4Wl5FDp3j9Utn
SHe65Q6ElI5U7Twi1d3Qnnr0C3Th/FWZxJArNSKjGF+Bx5mqAFx9sMRLYxekl1O+U5+ki3faNz+W
DK4DL1CIZ1xNaUyscXEkf9mpV60+kCiyTdOU08blCAdYGQ7RKG0qDp0xwb7v2YX3eWWIea2g4iVM
YeoSy+MKkUG1qNQLQRukLVM1I9ngWx4oW/T0KXDpgmuOeYaowAmlp4Eixo+Tn8Hy+GoicDpHSlyh
eftY00hK9B+9pU0Imas7x8bOE5G8LT6VkV78N9J2lUH5lyRtVBYOkTsZC3OC6uTvZHYHVjYqTod0
cV31NdUWJML0Xt7t+6TVCviGuEKC6pJGFiv04bZ+dk7EKi29op/wHFX8JrWqfZzlOmIySMrtc6Sq
Vmj1FznQ4NiYoBTVD4PZPVCcishk4f//5DO2USO2YvGAao2aGfg4jPDQy0UEgoIHVvxgU+eLe7kb
MlrapmtCXNeh61mleLYiRx2iX1tPyqw3g+LkhqOtG6neWg+/tWKN7InEIjzIicyofkzz8x9ZO0w9
r4DIrzTveD+L4F4Iu1WIoRycGoeQDKLz4+lbe03OO3a6ClqufBCNXwLNTuS9Ak8mX+aSfbziadxC
C2kHVXPIBTTxsZX2WJniUY4vnxePo7cMmFIlO2Y1YYql9LQJh4vmyRDRUgQUowPEzgNk4UN8tXIW
UHxVExgj50/17YVVAkuSB0r9LPl5tJzD62n2vP+elC65WTFz3qBpvepCbIPM+aFEnqvuY4TGgWLT
XB0O/CtKk/Ybs98BjPhdkPc6AHbV3YH4mK1im2j0FEiu8DmCLTK+WVkmsgjff5mnfovAE9v4HKYF
zpWvE6XVnNxunpKUjI4AfdGisMqVI5X7FRAu/3/ttA/dws0VT8Kxp/PNEtiTizeKEheq8C7vy0M6
D6q3la2hPFaDyeTsTQ1ScGccMWQi9wakXXXIA00SfjIzG+ojN6QMRxgJ/UjB0V1jIlYE0ZmEcebc
qv0Pdy35jTYqbS6ieMo3uBkOTPCb8DWDDSXjPcaWWVe4cOIibm7YeXbiUEOf0hAsSaySd4FI4tIc
l6Isg3iQ+i8wkBxVIiwB10sY98vSI1p0JUufEj9RRP6YJLU6mJfFbYAYjhmeCyrCEIjmAfbXHy7p
cLkzYSK4pLt1WBPxK0ZkmkV1qZYpeaNcgM8i91BBr+e+3ZpWp0mYh7xqT8TTjbSK2pReWbIJcNP4
iFd+DSpOjj4xsIfMA9RWzCDpbxr+M45vXMplDFeERI0rMX1D8SCHO3xDCv76PZXlPAYFm1Q8AJ7k
ddKioNGzbFdqu5QIH95HgR+LqYJsrT5WkgiXxhSn6P49EQ7vdpT3AltQ/bko6bhbnQB/fSguvI9J
Jk2s7k71FD83JUi9QrtsHHBF16KIoIxI+qRyLo8nVGjunBavvKkrCD3U5ObFGdxYgtd+cv4qdZNp
fv0oONejCTs+n/KIVeV6XR046d0YdfPNhYhFs5blGO7fGcXz1TtL1a9PhigIMoeW5oGlTfHoEedm
YbPynqF+hQjy/gfUXDgHz8xcLsOlQUvBU/6x/W8f1pm5ed3ed04hUlxkYgatwqSPt8c3Cgbzrzml
qcA+lH/Id0IaH7FOUXb9e4ss8mrbDzltbHI8Z/+snexyOjFdp2cL7UM/3XwyjEIJpughvxoNfqiQ
nFoRklDmAZgrNjyT4fCtDEQptBvJ4MzzOcXRc3lkCPmlOHfVJT4DGo7TFGrNbsS5Y4dyKJA/Gwmg
zf1GRa2j6WsHquaj32hUujtniSD1q+w5Ip/lWiUJFT2qRtW2cQkcklVbueG9SHJOmYKjPl/ADumz
OdyUOprrhy/VhpBNtFVtAc+cCWNhwZJIHN2RPGnhqA2rR32B3jS//KCZdYNTJrls90w5NkJf8BLq
omEXmRs7SNKTDvms2wno14RYeh4IJ0Wo2xF+cvNmXEAUBhYFPZ5diG/Mn5e5XwZ6mT+FFzNJdcv2
sivqG1em+sSZeQu0htqUFbIiuTSSPySLF7LF4V8eHC8i+aXykSTuXaRC9awk8sknFLfLqH/JIiJ/
b299MN57vW0mflwp6fMmi4OL4yPIqP3jgiemGOuGJCpUz36S9ZhN+wCC2CLgwwpWqzAQmqnN4Ful
p+wgi3dpbXZL8t7OXl8xJQnyzoaNUfZqkHEPiQlo+15yjiV36HqGMD1iNJny3CxnhaukkLhI2YnO
H+ulowr4bLBUMY/qwfv/ESbYRZVhCx+4AAFLOgb/Tq+YbVEF8JAg1vxA3J9MJtM4eLftNjt2yzX+
3STA2dLLhFvh60yHoSGFm2rn7WoLzymwRo1AGRaP2xNlvpBhrLKAImRwA3Yb8fUUgDHfwiBeN7T9
+THxfYVIuD36PH203WRW+bmpItCli+cRFi5kZv16GmVP7MPw/EXzjmbMxf+gydi+vg5Jqw6qjQqz
DTd03txTSaKdsD+/lqGyuR8+vo7pyAr2Mio1Jdm3rLw8GwR3sNf5uSnWZgmbquSLqAULsGabGOYN
mtIduCnnNlrcYDWqGswb+PXqVUY97vg+6noxORkbblw2wd3K4KF0aU9iFX8mQzhNtogiCmwrrqYE
XEx/XppuAFO8cUhUJhhiMCl4MRmxxNHTdB3SQGH/JYfrgj88THY/kXVpEEGHwAa2eM870rIRqJ6k
X8QeVBvLIoZZBpLXekxcr+Su4VjL3TQWHEqP/P7li89Ik2U5tXqv2BOrkv7PnwAJGEih8StjieIc
6xjocdLQul+KP4FF2dGh1w96HNJCE5KcrzBFd+jjxTBs/6SX0Pc+DvYiluqNx1LqL+7XIOhY234W
i4vuvCIUTQollmxnPVS1/l0D3ObW3ocVsnLbfqJoc46JvwEVQrwD/d1Vkg7/PxRGB07bNp9le8UG
YW+P7dBLVJyeXxqe98ogBwZMhcjsdUi4rVT/k0H2DoJTxp8TaA5JHkBNWT9x45gm+T/TE5NuY89d
9wQ9BXeNpCoXrW+bQY7C0avkeIEs4IG8RR5eROnyhnMnMc5+yF3H2dcaOAT3OsqXGg8LoHTKRNpW
BABaxtJbmv6HL25lNO+f8M4A3PI1CtXR8AkiSo4CKpGdpII9xZIAObJUZnX9upneQzwxC4NFpbOR
grtSGRquQU9su46phmejIdDZmaSb7OOLkU1ekF/xC9lwtw+DGPcSU2WB4Gm5HfQR8e9sxBuyTk51
4Zwm4I+5THN8G1qTAc1nwItuvpZ1klML/4GwLH5MIfzNphqRMCGFtaTxGDssYDTMC8oKfIRk7HiB
V5U+903fSQuZVkfFSjx1yYveCRsmx6zCL9+nT4hJFThxcgMGrH85sjD0XRFesakGGJVQtnqKgHIv
yesjOVggd3335wy5DxmJ0uHUi7GY5trpVmabFca1bX/BWm0ldkAEheaD4nmr8g/eFVa5Kq8pxHLZ
yoVSwCos7vvBkNNJlwNHiQGOvIr3zbjCTZAyIsmV2vZA1wZKI5WvccVctLJ2kU/ShUOdhgAU/y5U
KlzkcD/ZV3729PvbwUlNSz2narXhOTnv6a3PiA3v+DyJdsqa68zAhLtvPk4Tf6xc3jsOQ0J6F/6e
jXPJd5z+TCy4HU1tMmlRilaio6VjWefrmYFE3OH2AGWGeTFg2PXPOhzZntQfLV7vHAvEi9jHvrXP
OqtOmldjU8yFtA5pT7tljSp+HGLZGUNwca1tV7r+3Bk0Lab9/sMCF+QiHv5WHQKl8EGQRg7C7mA0
GxAmetF9xBemhVo2Lox9ebw3ZUHUpY3fTTZiTCcWY02/zDeWF4fLzwnvbVh54qNzvOIM9WlmOyfS
8qxBuGz5nZUjXhpkG0Xc/f3gc/iOqlwsenPkiPgE0CAv44HffqoZre3AiqoJGbQRXMXV/aCh5hE8
UeKFiU7GjQSu1ocI8UPRal8vO0hUrLyLCCjo8P8nt8Un7n9eyUouf3xySVgv6AijwtmqBD7pf6U+
vgAUReGx7GIMEDiq3m8+a/su3WYCBtpaI1i/LBVVwkViu15gYdH3eACfMbr0lPJ9T2h/roHK0/Wq
C+pQjp9aE6W/tNZwMr2Oz0L/mpSIetTpe5yfSicewZyd/UXKgC663rVv/seRkzUCozVvNLu2DG3k
7L0b5CixBR0ellwzimuiGj7MvhbNWaRlHUXsCHLCQzLqAx/pjbJJaeMcr9qIL/fTq8VtdyHU+3Ya
0hsNbBZuY4i1UCiUnEyjNZUHwrKzZRVPRVigfXtoMgp9VS3gLGOAXhNZLHA+6CsLITwL2aol97ht
f+F7TyvGCfQ9edx2Lxp3l+WZg/tyzWoDtbtX4gbcyAKCUgYZqJXNXdHWGTSURIUDZ7aPbcXYWf46
0NkONvLLH7FHstwB6yfiaUDe9UXnS0cABXjLNxoCds80s8j+AkT4MOd4eM8qgohc11tzZl9plg29
aGSMb477ZKxJfF12H5+4Gj3ulLJr+lFRYistBrgu1jnkpzp24ETGsRxdC2gZB6gxRt32SUA9eynK
DgB4Bgkcjy+YYbiTYNW1G4t0RdJ5XzPF+rB9OaYFSatx8fgfYBKS9HOW/80hlG3YT8I8C+tUHJ5x
rfo4CQKPafP3UWEUhpmR/fW1ZtGJS1TY7rP7DxLD0Md6i+1ixTPuOIFzoT8fN+2S7LiGDzVTJ4y4
l9vfR2v5hl4b9nVDCGp8UsdusJCfgOvkcDwVqokhGETTkBavzBah5egto7pLPy9evxFfZJR7zwoN
Agc6CIb6rILQjTUkI6mDJDcj1GZloHjoQ65MOoyaobsokHQmlICNzi7ZJUYwWqMbVbYSTBhUrvB+
Ehv7vEyEvi98kLdc2yqcoaWUvAfDn8toIoLaV9BVD1qlOYJVLqprtvsua84rdsDEmb5giP72l1vu
6CFUehnb6iViILbHef6e5mxmtR/GpK8k+RuneVqPX2UlfwXRn7jOLwBJZakTASsz9fnnIfpSpXbv
BVs096mwk/pDDJZ4T6MNAMXcgYOxt3kIw0fyxw3B47G7ThIB8DE91Ux4mKwF51oWZxE1m/LIZDCS
VeW9h31EybzmfFa+KqUGExIMYvLKgNqC8L7KwShIOMSCxGZTogL3wh3Q+vJkwvPV7JDM5kbgUJg3
4ShE5e3iYLHW8boXquY71R2y8vCNuxqfXplRzp8wlKma+tE8eZOLJ7w2PR8M1gJNtlbVuAwIR8DH
MzHexmUKvBYbrkkOMNYr0A3EXA4n9XIKVcXTsJnc0Qam2em9J+AbUNp0gHNms5AE65h2va5HzV+j
TtNEB4U83IlPCi3PPagpyOUG0yrSAA3+S6SLJZJ4gldTdcU4YS1v9L3umnHUf10uEz3EpCn/LGCM
gPXBm1lo0ekyya622DQGuNng/w0pZOMmN6SaxdoTBxuA8pCTkqbEAKaC0xt+tKiB5FmLhyGqaZSE
up0qvp7ik6MAHX2PlVMqrrTWCkZKvT3YGUSCgY6abBQMg8O/kN5QooIUWmdx1k4oSJEBKNb6C46s
L4g04/Ae4dMxEY/szTUgADpxO0uds4G7I7JzbyxAMMPMWHivHSGgviwb0WGtVkGwVKahFl4P5H8x
/pCDF4a+xkG3GrEbzMCdquCji0ci4p9/IJpCKcsiIGFaQ1rI7nrfwp7VdXB6ifTsXo/NR9AYUB0b
2d/3607MiwhewanqaG13VLedVE7A+buVNB+nYsgzLS2Bwft53rjPCw2SDlvhofdSLNkBYekvRDOq
da6huCTwPL3h0KHZU4F/sXWMY8icx0nK0GKCoc518eF9msaMFTdTC4n6QFiueT39lU1UkLWRDTRV
G0Su3XiDRCWpnipEZ27VEqrfMMOHzH0IPbCAEtCxd0eREo4z0oBBa6kdOh013HaAdvI9hP/mAW+s
z9tF5ySTAE/k9J8Vd5sVeurK1FEsA3iEGpW4tWCV8O8oNjD3gybYR6/VHgCklxlepCjEDoSAvfid
AVowvBNm5iM9miy3d7NzsRsnmm3jR6Vv6evLBrL4nJCtzzg0VLusw82pSIPQSpjRWTUhCGp0HWwv
rgDdd7sOvYS5VoKPHNMHM8iUAEnCl4k+8CfEhijx2/n0Yf56oiQ7FME904ObNe5pEn+n2ywQw/3/
/L7HzcjJFtoQaAYuHpCK+OQpgxJeX3lEgUzkdU+q6fe0xXJ0z1Yv7yXQLnQKCRfCNLG2eQZfJpEd
Y111RiePfi6kVlZ+rn2jcvEt1D+nO6VT4TrgvCRlFOPAXv11BZwOuWVMo70zQ2hnmmR7ZiGCaZig
0QcPW8Q3Aq0TGJ3onCEbu0vLtOHncWNNJVQdCqsPT+YefoWaEqaISic4bXIt14OVoRRUQWlrBR9z
ZrixDlOMm9fikL8qtC12U2VahAe/aVuUFON7ACIFeH/1KgtIM1wpwO2Wac5QTag8li8wgW1tkzkm
YY6C/as91Yn31iYuWgaY1td4ESC+yhJIocUv/RVet1n1P1aU/E0WOMvuKZVfsGGuT+tAK+mzxQSa
Vu2NGXg+emrP724VAWeKIJEmbxsy9VkhBGTcy5cx8lBf5mMGLM5VpdBKrMB5y3MA8e8F8IPcfuLp
Oz/AnfxCmazs3JeU4kLBN2lXScrb1Tz+kbiGGA0yJ81XdAlllAVudp+2pWZHkssm71WCvbF476Op
3zFQlhqfP3RHAEotSSneuRPNLLjS7ZLKaBYcv6hfJZnM7USvAki6Bnc4gYuU7fTS10c2APhFqq27
0r0tZGz0HT/doPdxuVFFD+bapzlC9uHtBADIOlzvRxBWrOTObxs4jJr/Mu6qiVoWapK7xCiiNFwn
AccXavkrLYdc4p+6zUi5hutpI4i3jdZvhaEMM4dA9YffmbVJcjV5H4bgvfkPmY+ILE3VMgdHHDe1
VOCTAYfYHcBQ1/uy/YpSb97joKN2WAw/XwgFSK8S+lwydGVz7XhquJIDA/8GWz74GhyfIh5aYyKK
UOBx0Ss9BJudkb41RjXgGs35PeZ26MLvGETRvCYljAPYoQTBSO7NvtyXmLeyEjW9DiiEgRGKXHHI
NyfWf71fhr7pC8YPz4N9qmAlXEh1Uvoz2OeYgER5wR7RUoA1NSi7/NlQOXMj9nWCy7GOK2SjkqyD
px1T6B6W6Oqf+opL7YBnRlAs6Cv28hreT5Q5AJQB0OZ5RQzV8OchyWA101AtU23Dwtr5OSCbEPC7
2Jx8uhj8U9fj/F4S0sAE765Cdh2FBAoSGV6vfe/9kZ6bFfuDPUQrmguZrKHkbcD9QO9eYia/4SYC
XHh3DQ+zxgBUmW5KMvFoedq61Q6duxTBvHCIMwefVLAkqAq3Le4XcVhcZ36OZEzJdFnazYEkUnSF
po+Km0TjIaIU7Wutf2Kkt8GQQG7XRVJGOn/LP2VYS3xAQWmdW8sqHc4WjLruSNpc8C9Aq26xAl1L
Ce71rwnVDM7Salr+c6xTbF/shWeZMGqtCHBdwQ+XxpS6VQs+BUKMJGHMNGMxxtfKmty61dIRhotj
TdbNe6NmIAr/P3yP8oe1GjNnVl7521g4c07o7svWpcnlSU1+HzDh89TpybM4j5zt20hfwUDmsCyE
KAdacnYuX6PCE18n1G9kIJsf9H8z2uLaTH+77iVtFkRfjk4nqVVadWVBaQPhGKeJAH5FVr+I8pMc
uukbM3Syr0j8HvMdfnIqFL9iwYDuXEQOrLIVQyvOnzCEeXdMVMLMy0BPKCzkOwkrBRubwBer/QaD
dAG6bAIaF8x+ZC5heXghqJEYO/WjJ8USfAGQJsph559QntjIexdXtFJskh8SjjhJUvVe7R21Azlh
iM0WEQ/j1sWAUuAcWu6a6LSM4gHShgkNNMfofTyDVWbNob4oFkEYy4kEV1bilae5sQCTJW7Mhhi3
RTl7qHrG50XldC9phqEhPzRpmmd52dd6OViIzdJ8QyxPcV4tn0qOzfALmbA5NtLe3KXuXbiZlqr/
ChVF8MjM3poSET6XRv3toFLoTGxAwv+D+0J5TBmav2sc91jz/XZCyKr5c9V2DEh7cgAbHNIGvzqj
uF7o50EJCsTXFCVVu/TDNqd2PSA8KGTNXPTDhZvarBovChHALBrMe7mmcy0YLI3bD73TeIkvuQmR
dqE5A2d9+Ma4Dg+5Q1m1mwOXLvDhZChI5hQdxbjrumF72aL6A0G1oijknlyZeFy8llVQFK9oGQTd
TGpqNfXBA49KczPz7X7lsaiblujzHgKflawEmfTtB8oRkdkogJtbPZoSUNWTT/MFAaJ/kV7e5aUt
O2rZgFy2pftghK8pk88Mr6BdgvfFpmbnHsakmsVnGWSQbazHQS/tgJQ6CJV++dboRS0N/KI2YpF+
I0tjfVVx2xtDGAuLk7y8qsfnl23UcuvHndWl32vmH3YDfh3CIunfIAXcodZ1mOajDAWI5W02L46c
/JxXgbd7u5tY0RzPFfMAz8JlrIqIxW9ZXDsPCBP2UwRbK0ucG+O3FbZCYWpyxWK8mzlqwQFuOTRx
0wedacWGZHQ/X0ZlfM3JW7MEZUJzY1EULW8cYN2KjeMnHfV8wCfWmaLTMcbI+c6j256ovQr6Ztkg
SWPNXO4L0+eP4eCqO3kQSb3T/J7ttXu2pHSIPzNvM7ldgEKom35YMp9pxxT7zbAwi4m376uEmn9O
01Obu0SW3K9IMLf6ubIF54D0dG5BmIgZXyXY5PFDKitBHDfJrQGWGIst0NZt27TW1aWCidvUvNVg
wZRjHwxqa+YwuJm0CzayuazwozcMQGgS3lzSSem1Z3rI+ib24apZkMVWkdIQ8oez6eR/ZLuvbbA2
UN886rnni+fZw6sRbm4YEhMeTiGkWoR0k59o5OlF+N2W3hLjVRKgmLCI1jvcitgk70XfZ/5XA9LI
iIFxs3SBDGCTUaGJIJehU9pd05hCU0X1TcMVcVqGeXkHp2Uo4CzaBBtnsY85/ySByb8ztSekdT62
BT9/a+y8z8K7eEAF/BO6ehXoNWi6iG+THEf9zFZKEIlQlVNf+WBRWn59whoC4fa15xaARdiSUNv0
UJvBzzzmODT9D/iZMI7NTtdUhkd9my9S+5RsGWjZBBPjVmIHPGzq/aekE8lgBgYEEbpY/Qx5niVd
jC/ZkUZaE6zdi0h46xh6JqFRW9ic52w8JQZfOJ3EQ49CwgUZQELiLyuLhdAT8NKH5svGc3Tdm+Bn
jRBo5kfvN+nr3N4JnkY1V3ihE+nYuXbjp5NGAx3amY0LT9paJL/1sl9MYXnyS0BOce2HeCsxx21L
KHgKM1YHHP61e2WetXCM5hwHa/CdvArVnDMCAWPpH/2Wabyfa678fAVfEHA5mm6P1m1byz8/UeQ8
gSO7ueH5OGUU9Zwm86yTuwwoAaONJNH0D3PRV7+8il2B0pFyeQlSNDOZIQ0uDUWVwRQy2KKkBqXv
Zms0W7UAVqmSuYg5cNhjSmf372hZ74fhrRIrWdjW2PO4SV/hTsop0Ofg4sX7kjTUYoEUpJMeD3OE
4fjKSVko4qlTOtr7Fd58LXVoJItMMW/Rchuw/Xj+tEoaKco0vjhB4SWf0N56/+/+bq+6rR6h1QXm
4jfKiPbUFAT2I6aiudJQRvDNugPGVFeabzfBG144Rq98B2fy22K+mPhARGvqEXSbAd9yO4bxL/Vu
yUqYf+rBjJdXeWtwJhm1qW1llbw+2RaTySLve74et5BYYA4PnqshD2S3fgEvqgF/9JamAyaEWplY
NkbBH5OPbArwpcMdeMY5j4F0MDtCSBfsLcpSWisjROUKeUUnqU6MFJ7sBIfJDqBg4cGOSrHXPLuH
uJge840QUFysRLHHHCVrS5gLDCebNCKV0TqmYMXVSRNYhuYoiB76+b6E6wY9GE7gBvZmqO2WVFT+
36rgYDQ9NdThBFSb6Gq+KtGfXpiz2Dj9u/PUXZAfwVX8fyy3Zb7djzoHCZleqWa2oZ9Jp6TTTjkQ
AeEZ/B9guWNwpYSiCirhXGsWsFyoffb9yHybYzA+/8nI3Y+3xoPIQMylfHTjOMGHng7ljqhrC1vt
uFdOsHC/026hmse/t+gWjhTNNE16qHjHzJp11yOeAhj/R1PKqU1RDw8No5d4Dsj54Y7TSQy6J/5m
v4d7N1bUk0y1o1pep72fSmTVGHR6SYfHvMfk8c9VpCkJRBFIgQHf2EhVXyiLbRSu6v0RId0I9BxK
RZgZWV/CnnybYWFuT8fU8ZI0uDIlLjWJygP66IPOgzBbIhouV9TXldg/mg6MMBEaTVouGOSx2BuA
N9C0J/3MJoMm4X26Bc7dTL3l6T/d3fC0u9FXpT3ZsadmxNpB/OuN6v5/l9BmZyMq9RkY59VZS/H9
bq90jHEYN2s9D+Jfa8iw7SM4E6xSyanhCSKWe7Bh5XzXr0TkooPrVUo2ENF3TDh1kTxT9lsgrbj3
CmxmbAaKbu0yjgYIxlTWVA8tYFbNNFWRs6tExzcRHGhgIqajO/2A+0a6E81VqLMGgJMF8WbyiWQj
Lcb3tpVUrCitUL5o/L6MqK9KSW2Zr+Qdrm0aWXEGb+i1Hg7tKamLPOBa6OOH++vY4qQNL9T8RXtu
Dyl5gPqhtH2ejXyb1NlyjDZdgyAZ/kDdY5yLPsworLe3tYi8dn7AB8sbIx81ka0cUMrcsdYF/O66
/6030jW2HIz0cAp5TUTMiOFN1WaN48cJmaOK7riC9BYSfzGzAbrBB55soqv9z+llbi6b99mfhMCt
ygmDmqNG9s87bFKDMBcrrVmvt3+337IuhRKlm4/VtHylwLqR+g+7UOw/jfcM80UBXg/2Rq31FLyv
GwZZFeUFeVZ3GmNHuauEomN0sfWWvyirXMyiW3jt+ddD7F6RBt5kLgmOteNPc1a3OYGrZ45cE59+
oPjDI2oeFQwW7Y7e0UEEcBSrS80ghkTRwu8eI6nYvt7IP4mhCbESOkFkq8EwSROx8JJMsF4FAP+L
n+Gs8UVGCT+ZrcXmflnl2PwfaiidPwRW6PVetdWBHqo5kGdjiSBoPHeDSrvPk2wFbdMKptl7CdoC
jYNbFFXgezdRr376jjw4d57TtOb6UFKxlqWZCwkMr0gQhyE+36bfGecpgzJs33tw4WPoi0Y1Pssk
ALpKVXZZC83u4lJY3WQK5vWHhcSU2OAbnFiD4U38eOVn1t0MuwGTp8QnMnV8h1wblqpkSauC9aMQ
4JO5/OHKD2UGQyJg5zvLYaZrjkB7DyfURaIAAdE7kx9Oy3JstiWVVCpdMWex0Cxi4tRJVeW56BM8
8tPrJeuM0Oidl9HYF4ifgPtbEAK7KuDTyf7SCWwVeH7/1GjZB8CwA2EY0SzEhzm/eQZkmfPSxu80
cC9P4Kal98A3WjZcO6Z9ilh8PLnWypgGqnjBxI5q4DD0Qymsl4ACaIPFIRQpnnVjBk5LtHhdSP6x
ye4iviu/CHTFCCbOtQjO1UFVGqdETOwWafnRTisyGunIRoI7MXQiaR4RFzwxlHdkn5rHoSDbMPZF
MCRjLhwAauN5+3TAUol1peNeoJxLF0ZigkB6QCsyUSMA9KTZ2VGX2+NMNShwVS1mYRa+cBRbEBUB
Fk0pqawBFLbBwORxMuXpup4rftEbfDdWC8/oohYMLaefq5EL2vBSzstgpW5S4+tI1usQI9bUGLje
3e0rr0bswyuppQz9anCLZ4hO5R7umZjEC2FkiXtrBXNkym79v1ODwdePV116G/KmSuGEvF9ymsAU
ps1UF5bbJjwDXCKzjZNZUGwxssuwUDHzmhWDvy7bNFz4xU6v6g4vFWbeO1vmL/QR2X2sH56xz0BR
eq8YKBB9NzImSvKrB19YpZKps2r1zgaVUdP5s7K4XtQj/XvWepjGwhMPPMpSZrKCbP0wpNxHDY3U
u3ZFL7qN6lpL7JL1VTo3JNxfptrZqhLNQXFUxjRoG0BsHlVzqX/EFG4vXV0AZBJhzDnpswpCzERY
ldobM8+4xSdzNGs7Bedv+s9I0xUVi7us0pUU7rmcfPbCpKVqJFEdFd5lziomrQBRd4WQ5posaezF
UAxLRDAv5aUkS5R+3pE2vIVAlJEhrgYFX7O2kPMul+ntSzzgExV5vLurZ4blStbPdChxkaLiuQtv
qufvywsO6MNPla/cLTU8zCROWOxzJliHL9SpAjeo/l9zQ0u6dXSWG02mfGDWCVPyHf5Hmx1bDfPq
QuyvylsZl0tHtJ0q+ZrD7B8c14y2pPiPdlIb8vLqoCegFelNmhtL31bJtO3d9XWtepd3v5xZuegQ
4/qFyd4SZT1G5Tlup1T/j9N3pVS7vD/DPRxOWK0O8C3PBvQD07OjDL4CBi/HtT3R9/0PvfO9wAFW
Wm0Xu1eHTeFogL2Baqz9Y5JFGitsTj94sDdPvqLWittMjLtKHuUlGepVjh15Z7VI5wdTS3uSpiTb
Qrfe9ue5gueRTkdz+wZzjdAPMzg8YhfpMoxeaqoucUyi6+/+uUnPeOzFEYmjGGzi4mcGzIpMmkPQ
0S5kAQ7rFOPogrBDaoBdDPSdCsuqNQlkYN56w419p2jyY/JVLSHQHIezm+v4sbTAP5sxkTzZEjzz
S1yusppO53tJi0t+qF9fzxq1/iawy4DZc1BJoPqsy6AuwhmMbeXV7KS7TSXjNie5GV2zNaUbWOGz
VcrizAq2NeoWNXm3kJ0+lZfr6lzav0FsG9RMNdx2U7fS5s4t+jAfJ1hksGt6XVbbIlW7rmL4fgjK
e2YBLY8qIC1whHpdZx0UAG+2d83UON7UjwbbZT9Q1joNe179mVFPpKDoen6cGO2dPUZGq3p9kZo9
E7xsN0OS7KPwFG++E3jXXks7oakjqbWcz2uoWCyXKwaTDitmKISg1M4y+5ynBofvUzf2yqjEB4ew
1qsKZRMbGnA5S+BUkMcNcbaESK6DgzV1+tzrZ8GMmKTjrE9sr18ttAkkmybSVF56e9nnoTm2x67L
f6T1nCLfmnawPrBdA1E1cGWC4zZJSwV6vpXYn7DegeCR2CZJyYZqkIK0mk808o2Hj0T/AmIdDNa+
re/ICfzucVgIfhsDtsHyYFz4APVlzex/mrhsv9jtoJLAT0Tz7cMBmYQI8MuY3aw/oI4FE1eEdrCa
Rc9vCpA/tr50ujArdRczZm+r4l/16R+eilv3zvVGw4KTD+7A8lkwMm2BiqS8B6viRwBLsk/ZVSnb
HG7VBsvpE/3+Dkcv4kZDe5pn6+v6JtSFZ0YSEaLsFZIg6qlcUk00CpKnse406ZgYlVxD7LgLbrXu
Q2yQel/wECAxj87RcS0DjdBAuGBRPTv9+cW6ujKS7cd0TSYaTeL/6cv0HA+TjpHCr2tLaYS4V6Vk
cvFLp3FNEvRRbE8c+zXAL/D1xDvzwjfNEq3wCoydSKsbk6VyZac0Zevq+ZfJLwbgGULrOf2jlWt8
Ks3Jh3Dcv1Z67VgdrtRkpctHRDNwi5h2DiR5OAtLL9wE8iOf4+xOhVgp+4JMP31C+ULMHFQ6jM14
I/oeewRqONpyRAjyLWR3n12CFlGLJd2pY6Sr8grYOMp4zucD3q540A7sSwW/STEavzzbcASW54ei
liI2ilR1gJ7sYmY88JkjAqyXzjXCy9CbtHZgbjtXDwcJw4xMPFkfxUtOwIhuo9q2cA+TOT3nsHWf
6nzZfXn9LHMzZF3OzTilmXHWvLHT8xCSr9FIWmHh1yOExkV25iEXll7zrIq9RgdPd0/tugbVTygO
Vcnf8g4OJtnXIliNV4gzPgE6r1CaHbeU+LLcd11q7bCKjX/ULoStFp3FPu1mZRIuM9yMkgc74Une
RDCYHqQ+XA3RH81udxY+BSPfHRWcKgzH8gWsX8wLmp0w+pvlo2m+CN5+tm3ba81RidPrTrfVjZd1
UvroXPMro9yRQMEYgAVuB/p2z8VT6/eW3KeYE2VRwKVAMGty580WCNhhI8+tQ6gglOt9ztvVKX8J
Xviz0T8t0OpN5WN1ENFt9z9Sl3LjDsk4goqclsZ/vR+QNiQ9l1Xpw+vaIA5nISpL83DB4qx0ToDp
ui0XOF3UJ57xhp33DnF2N4jl6M50bX4jwZoMCPx+z1STjcLsxkFXTPiQ4wkGb1fOMxOD9Dyyh8dD
Uy9JvPr9RkmBjg5iyiusH3mcwP5giCMcBvfNi167cXtJ+vbnEN2BWGAgxsXLH6bWhnCRThit96n4
6tX4VYRWoqXqzEwG/0xuQ4L/TmVRdrA5ydoxe06lP8HuGhitoWjYdV9FaRptijGBaWLz+tUHU7VK
sH+1XHMPuRDGX8jWUXVVc5lmeXFi05goGU0oUVoC4uzD/sDrtLTxgjZMtxIZvlHZK3IMjhAgQjZq
Cn/XmcF7uRCjNzyVS77LUJjye8yk++CHC6K6xE9QC+lrNQH98xpKl/pAAlcWfFm8Su6l8eCR3cDe
B+AvgI1FFpOKpnbAZQBk81li2pf0AJKqDXT9EzhSUYTIE6aPQoHmWbIwF4pKGxxsH69Dl2CPFYyj
hcNI238H9IcnYhi6+y+GxV3fkaalzdEGy1itaGsNJDpYO75vUNuCnX3RSUvlvWk/mJ36Yvx/FNHo
zGo1lIDdBGvuvc+PyE1BwVlgtdV1S2XBP6dMYv5TlovNmbDr2eKtSB8BFiT/oPD/59oi5FrnWBPx
sT86sURcerf3bQ74gl15NANmyNQS7SW3g4BvAD3DxSlg2ALEGFY+g8P9OQNOtX6UQY3WSOlSYJv9
9q93UocPzuFqgoyT4oM4bY8HaBHqrZOXGhrqeX22R2OeiQYXMm5A2edSmcar/AnBGaQYPT4eLyrG
t0LPOgvJepQhOdUboQlkjF6KKWwNRR5dIqD33isDuOP1pDIHcZKu7XhFJ2pejMYKLBlN2mtbtfHa
Wjeu16RYH92TkPxcnp+387GcuJ48C9lG/3qd0Wjw42bQ23oxVVtHZENFkjTnRW8z5rwYH2uA4hII
fF+03SwwBDSBv9VxnW1g/wa/ugBUSZqXoEjAzdWBRboNnBe7ed1L05kW2u1+bC2wxGyjwW5bG+sv
hpg0wI32EzOrPJLzVHwZJxaqvgGQ3Azl09ParislqIEcp+2TTiFhnaTrguoiVAzrTz3xyfBluLp+
map+jRvGrsC6r8luG2WriC8BdFTqXNMQx48k+cEXZ1kWIERY8+L9jylb0pO6JuHD2GriykJZcR7C
xoSqIZAv1ROzNZRyK6LMGSCEsa6HSAs8xftSXIICLqKTRxpbUx1ra7iOgBNsuJevB3GHOzTt1iIg
HolgQGC3PHVQixkwXNMgudlTuECIvFL4pD+jGx53OJnAYGO8NNd7zNgi4xpCSzr0FNHgCFIdVd8O
tcRBG7f+nfv5dERKYpC4/b2lEVighMgcTk9tlLSElcMkRAryj94EjgB5BABtfe8BOT/4OOhFFHZ8
1KK4qMqg1zrlEiIFzZhWRrpFuzVpmNWAKEuOBjCguvTySt+DlNKTWd+pTwD1DvkUU6/EZ4Z0ws4D
UfMM6C2/cMa3DP8cFFcJ8KHU62Hwwhr3p3VqhbhbpNFfJU7aEJJmUcNqhhPnDDknJnK0qxzFqvlh
ea9XdEnfiMyQ568gPAVzpy3sx6/Xb50AR20pvswVp6y40yx+1FfMdmwkY5QTqSLnbYBbx/UbzZ8A
2BPhGe9E+iEF5VAOoyhoO+CAtv8NpcPOrjxvnSueXG16JXLCe488u74Szv5kEprU7+FFFeigw0SQ
1Co0nOw3pvQeLh3nCIhOWHwUjVKe1rr3rHRxN4/Li4DrpC8rf513mHP76wAeEV0ITTtAJKhNBQdq
YEVmkiWzofPEP+LUKfYeBFA9uog4mnAtiKpB0q63rDDFlb3gimIVlr3bDePvvwtZ8Cse4oUWavlI
gY1a1akhVOcygqGseBd3o81A6m2fDqicO9EPJG85NO+2FU50cxwdIMz1q9MqXJAWRd7OTuPRpdRh
0dv0P8R65ouHa+vrSqcs+OjmLHLF+CxGBHI4hgOktjgbRCWREnMu7KlqyENcjnPABfNzaC/ERebk
F2RIw8S2gbN/M72q+XMqW3bFSF4VeYWgDJ5LS2JvF4pTDZA8k9ceHWqc2Yaw0LokbMI1JI0wzAYB
/2Ye21nB/AJERasIiHBBaoL9eKstxkTrnNahl84ZiFlqA32YT8yuEnc6dE0u1BPfWI9K+4w8Zf6n
bbtuF5UKif0utbuyLHOK8jWAuJ2XwHKrj7I98T2YnHtIMRtY2AfP8/EYiU0WZhw0CJ7OVNfvgYUg
wHr07mCx7VWrQDqptomXBWKQXrLbjLC49ILv6Wh1dN7YCJyT/Ojnky/t6g3ftSoRv+v1mvsk0oJ2
auu2MU2YHZKr3Z/n8aZVANM8xJxuQCCThDu5uHi0niqwUNIl1lMaYIdQsMkpKYmuX5uWQYIaeQlk
vYXCAE+MSbIe7F1/AC97k8A1phUCt7ISATVsi+azPpMX3kWSbgpxjjK3jInXndiEiItsD1ovw5ls
Xk2emHl2Nbz7oTWUAMu9TFHeLmYQZnTRWsZ1D7niodga5Z6IsCv91aficW/fo/PfOuar1X2yl611
aOpUHLO64SH5X4iZUxTttn2QRXFw8bjyquGd4Rc9a46ITgZbyWS+lrdWnODPlpehAr71N6sEco1X
REoYiXlERCTTpm0fmS8Fp3dWctr+NDey0SB/GMguZpRH2Zz/sZhz9Pf4Vw3wKZ2bw5Vhx6e83nFX
h1GBn71OgTqRtrbD0akTa6LrWKsBFatlXzFwdo2n8gUIkfgObNpEnyUmIh6uyTzMFn1pKAFuM0p9
rmznzOjnEsJtFRu9YVASKZFYj/ylO2v3PqaqVSxCbLA4mFtpscKViHoCmc5pXX1RrPMwU9r0CvcH
Q5CwbqzFAXFVpzr6H1oc9TVatpNJp+P+5cR9CLkVcA+LO3hBv5sbvgQwjWXOpv3EZJIle5CygSS/
XNcdNAv+/FuuJcG4srCDJH4UCaB/fvlHxzHPPph0qTWhioOcIiyDzLcclbxsPsymwErrjMFmBv1r
7iqPGyn8KYcD0gk2m01I9fqu46zfIjeiBPVSfkVIpPRAZ7Ked4DRTAMo94wPfri2p+46fxCQOLGf
00gl6jPUTZGkb4PcEOukyW69SDHCPzAbq/X+I8zmLm9J57aBmFU7Z3jRjmA9PQVdY/NhoKbiLJhl
tgIr675r17lNM5roz6dLlSj/9hchInrYRdVU/W6InzO+66t8Iq49eBiVeFlWDmAJ5Z1HniG/iIFq
72LWi4gwCxcw4Y2WXN95AXFZVyuKPjXh1uxWqkyhthuTIOg66qCE3aAHJvHfm/bMliioEq5pvu0S
sNxwyjsiwprD7bPptFRGyPra1bKP4h8928Ap0aWzAe9FITtfi9o+ut42EPtAP6K/XOt49Lcxquw8
TmH4tpxZEKhmy8M/b+fFX6iCsxHStAD0nqLtoKK7BhTzRhLC10OrBSf5p3/XD8JMG9EKbav3Cl9u
R5c4P/IiBeb4ejV97prO/fRe6W/cZqLlL9fGRi9+vxb/0rPglvYA0NtfeNFaLLgEJOaS1nJCUiQ7
XUcZ3aCh+xwTRdjoZUmxyRCrMsT5RecV/9hqUAlRCwsfYcEG4z4IaCfiEZVDK+TQv/dJkF2KptoI
J7rcvvPBgRqOJLjsxUwlPvH4tFoTtJm5vIR1PosBufDDOhHhYfsQiFArxXCUFhhcmfilMCQFs6lb
DT6MCAetBZ0D/amr59c+VSD3gXgixuU1tKLw9GY3Ro5F626x4IAFWpasGm2xfRWMaBP6S1wE156s
y0esPqssZHtIClawWAmxfNK7nlqo4SVFLMfSbanM6Ld6yerMP80wt6gbFF8OcG/SeMD/GuOgt+4j
5zOUDSUI/q7mxtGwf3FYzKuS77ukThBHIDiQlmANg6r1cIqkp43LGfaQgjOAlQanwExmNLK0a+gs
uSzts2HssnAF3lPSh0+Z+suxKYz2PlyyixlLam/Oy1bz2meX2MFR2IQAdGLV9sDA7R3qit3kcNkc
YPSoXrCNnt9Cla7PoFaGVYXYNjLcW4CNDophR3+iVfLbvPEXCJjBr1FQdATd4lXbkJ3jaImY8ksH
hLaWOJYr5tS3k62J66Fari0PmAIVQcWpjkcIk4sxYsNIi3fkSioNrukgkHYMDjhG6EgZcqmdU7K4
Zg4Kg4PsZm04fZuVJqHN4hMLmWBAvMYnjGdWlrKhuMvXtEztQwaWV0tMRx4fNORv+HcL5Fn7C7DI
fOKMjKl2BqR0w1XaugsxuDPKW4eNGfkq9T3NuqEfbIkKzwV/YvXr13+UdIFfUAbquRJ4ExOAIC0e
DoqDoEIKqriMv9zu6rurNfpninbkICtBxfgEh2IEKK0jmfn40E0cWSryKRXpk1Azk2Qx68WMSU5k
A9i/q39Y0FF2/gfkl//oxnQTkz9p6k9qdMAaVNnSy/ywbKlII4nzaaKLMtnqv7hagl5sZHeNRFWN
gHI5vB4D8bIQqfUo5mAWTcJuusd2fGtxHsMgih51iCXCoj457cXv8VUCjk6UTaOmELE0hx5y4sns
3QH43a9u+bEK3teIw7/13jh/Ik/gqHJGzcQJgCWeV1IdUV2zKBndA3NWBpHUNtXJ3WsmH7+9hCZ4
6K72DIK3BmYd5FahcutV7uHDmvJe0prvRXhqxhFFCpWlnFJqc750j9mHv6MVDo9MU2jxzwafTszu
VkeLRi/pjnJTjwfIl4/HgsWtbCX7zn6VOyuK/IXYJRSh2ASx30HjanH2WUzc9iKORzqX5Anif8dq
1ZfeawvvdnkiFgCQuVzrBoZLFOIL0ZM7l7kmUTyyDP9YhqVsHyJ+DEROwN8U6mfLjImHhDGtg8Nj
ho66TzNsdnduLjUuq4l9IzzqvevnDMoZK+YytzmzJTePgw9/S+XdMuLJG+J+avGoh90IVXqcu8bt
eLqb/gu92JbjkpBuiHwgQJfWvF39gNxYRN6KmHqbvQlhsKMFLbJ5DUu3ys1+YAP7kW3n9mxfnnDg
93oGtW9/1YvDqPWDAR13WXAs5CROBx/vpI6RBPgW86lJxnfsL92n62S3iWa0CxLU4yMZmT3EtCbE
GOc4dFMN/8quC0A7kwF0CGso9s/CLwyETkaQ+qknGGsQyYxPsGeGkbC4/K2ezV7jjYi9ps+wr3Pb
aahgCai9E7/3RmpPjEu8up0R8BsXDg5wmAWhq2B1vjnQC9CjBiNa7LdjJi07XA52wXGVMqwU4eTN
P/+/pvFvpv6ywGAZ5ZVjZO5pobBE7/sUTt2D/a+HOwpR5faRisAFwume6ydMqJYlp4oUSdjU5/d9
XzxB/QrFHcJZPNWk/Kvq/zW/ui9kmyOSobzPS+3Kq9yHnOAmz430NdsM6YDRte8EbP1rrGMs/f2E
LHvCWwv5sHXFS0yh92Kna3o6zzvnJhrnYsYhVMIHQcqGvJ0qerbksVyvdR6NcmoSGQY/fmqDpy5P
rfM07vuUMG4Y0H89kvy/mPdyCw+BI0dU/aAL0TjtZgzGpxunpnnY098CawRt6sIzPjPOpJNjsjIY
t36mjAXZOakCmSGM2CflEd4MrcQsZkXm8fCin2PS/bkzrEK6gW4vAGiX03iuuKUxKsjqlE6AO6SB
k/qMQAYQGsK/tFbBmuaSpqjxiaJX7R1v6dbSPzA50qY1hEV/OGpPG9uV05dZmtQH5FlXwChKgMbW
DDzTPp86odHnx+Aa/P9RzIHB4grKH9I33SMocjjVIrAQWTXVIIrwKmaFTDMYnIZK+xDXE9esYcFn
qND8paS09E4MU24C/GF6Z6uRMqhXcAE8lYmcrrBB4JVtRaZZTQ8GVxxsDFOv+woI2MlQW/ayNQIJ
y9IYJmArW8rCZPeIluIzTQlg8X6oqyM7f8o1nW4xttt4r6or6aBuxtnnnj/O7FbUqUUUC1Gj8Aoi
2jyYRwpthgUrbD5cX8/mSv2lUcnyJ/t+s+eMAs9D+QeH0JUEbQ4oXkbxtRXZzSxI5c4zq5Fl/exH
V08sDNT910L+/J569pOFV2MS9daYl67LqAPphjdRAOTEisiC0QTv7tHBVGc2n/5y7+sui1r93KFO
tdNVUru9BuRQBgO62bqpATpOWON5DmzW+7ItaU93Lrwx/kxHBM13EjnX0czXrs+hXut8BjgQ17yv
siFIO9KTzSmpl+bXoE5UC4LBXlu2R7wUKnAoJE3krK2PPTwJXPqRXpgQY6J2pwekNolmj5X9HNgk
w7jJP/viEVekpdKHKsbRxnJSbxeA/qhVsEfadkW/n5uT/F2Z7W8LzIKHTnVzEfv+SlUATTnsSQgN
xLBXAhgOm3cLYwNoj7rVE+lReCmwuutg/juKIyR6w8OFOtxgLSfcp6S0kFh4bCyVlJFsv8YCRYpZ
z3lSTepQZWlBCTKnI3asorM2Jugav6u1OJQR5rAIuFOg7Y1gdVyMr/wikabYq6u8bdbXaoXAA4iu
yvOoHLmaw7yXD+FXiGXpKVOQDk/uZf5IpImtIGm3UeNmnXxAE7bEoIGN8xDl7CPBRIZLnRj0Dxnj
64CnqshKuajXWgET51pDjYbvivvjgZsxaIYhoVlolnxk7xpK7Gfh/EO77cWyZll7zVlTr3Ajx/8u
b9Y6XUPL7go+b56lKLCBrcobD/EWptgPF/IzQGmxN2ulOciVr6D4LfytYpq9gZnVrCCRJpPeHlM8
YstKoymTgGjcZ0jDR6wQ86jikNaWbNc/2B+a5FRMByGJXnj9/ojOeBneOi6CBN9I5yv9pyayjNHu
f+XiyEZiQnQ7PrisNEm4bkdzILYp7FVgyUBoHMLiZz7jD5Bx5mOy757JT/CjF+MNCulioHcsskvL
545rv7imLkEFZ8A9y/9ENxKzlBFRAnD1ShYMhEOoXMTTaSYvmHB2lDqPRfv/+sugGH0Fs9H8nlP2
eIXvedl/HWhISh6oVXQZiDuBPQhtC0pra2lUzRS/0TJECUwgMX+jxFjoxGrq1cjMAmGA5CvjAG2u
Q5Ch2M7xjUHxUO3hrbHGS4BqHCbOTKzBREvj2et7tp11UzLc4AR5KOAoQxehwlUnnzAYgo2ekt4r
T97hatKHFAOz5uFLCVXXmCZYIw3rvwVIlfgoq0u+gfTYnwzbgX7havGJElvBbtUZmjl2WyIwWn8g
+u9MS4kCrxWaKZGu43nQXdFXbTDJEZmDZU6XGiVBU90oqwesERU+GsYzelhH/D8q2rbwgussLvm2
1+3b+K+Zj+Rj14GsXtH26hhtVa+A1YRiFSiGqe0oWfLENYXpV7JgeaOkllNpqp8HAtOkXy2MneQM
mySu7WAhQibj9DfjF6Gxvp88YTunPmDaFukgm4HR2UixP/vmOVNPsERFqdJkro483IaqL7kwMp2o
9lh5KO/bOHEYzpeHXUOPpnwoGG66siR7sJ/0HKyZUT4wwgVS2A2U11FNrHY3KLgI0FcCLCKvyOTu
NxDa2FMYSzcizXhcN5y83YAgd/EEGrNvJ3mX//vs0qpKr2IiVtw50JOP5GIUvqqBtOHIhIr6+eZC
BTJ7JhsOs9E3fFWdVIxPoC69ydzeDHidCa0OPYmcOuoRSrlCZpSOhjb8HIoLbr6rho8KVh3mxkRK
C0ufZFv+B2PNljiY45USliYJxVtj3tykKpaahipbY1DIMizrFFunQB7vsvpO1tyyfVyrXEnN6fqT
QIWUzyCLb3SULvNpW7TRvm/+0lvZgAIOvZflQw+ZPUGUkVMnJjyZ7FeSB7TH2O7T/3TC4le92QFk
F1XZb9cfoP9D2YGEuAJH4F71e2w5cSTqw2VJkbJFn6XI2lcNc402fHKaYRd48qlXrVeIRKX+0/4H
dwPk1iPBSuyqPBmV2JrXJT7p2tPlp0oukrLhM1879KS7DoxhYI0cWfEfzOCaAxIUPrwGcSqcwkGK
DQXmKlORU+N2g5rlENIr7y2U0iv1AZ8lZ5vO6bDXgoAVUj2HcCxO3S+Kd9+78yiLkJWN39V2kMid
icyEAAS9gEZJpqdfxxZ0sXpAfo2c2LLxIyaocmHnhfah7t9++jZ2GVTCmGRSwxmPm0igE88y/EnH
8sQXoUgxSacPb8eCK3W9OCnQkE2mxQTbxADLVHN82QFNnK/f2vqvVe1cHuuaAOO8EF8yY/6PCQ/5
bJrRqG/tIc7U77McqnTxDrbCd0lmgKKTcq0aW1cWZZujQwBPJCfzleb7JrpMq3TSqiAuLU8VtZbZ
edXNd+SY2GOazh/KsiVUvyKLGP48eEYYX/qpaEnWICwW585emkS/6PSjXZxr1bpnqm2P0c1ZVlck
ZUit8nBwcyNvuZ85TO2IaPuhPDkM7jBc5sublPS9goGF4WTSEc12CC1TBywXHG65Tpl4AXyZhmIx
C8F+wDBRZgHuwThdB87lJRfzaML7NuCd3c3QbWN+aUkXq2bxbwcGqi7B9eLWg/Ig6EJepTNPnP6Q
u8MS7cOgxCEUZ2Bob1dVtpeKZegm+JME55FimPdygyXj/zdhW6oPRpHUO4pBS4DT6k06qdPfQehp
yGb49Yz8EIjsmkBWb2ZUtFDhQFQbCV2It8rjbXx5SoMwm2kMhC+gO3QlohY1XjHAKxLM5Yb813q7
HaJm0HI0kZmyvrERm2f1tWR8DIzjNlJIB3URdgV6LwAfrcIr9/yIOen9EWtCVTuuV1ZCbw8VZz6P
IZvZxTB0dJSw8tfWNUR60WXam5beo0oSb9kuyrVNbXv7zdCpdQmbySzIIs24oEUM265hXzRtTbFq
WeJjhseFyJuXwWORPna+ApCTv9LzazrLSD7oH0E0ut1QoflWnWlMSyrbfViKDhcEdkqJaA0CIY6k
+HFqqiolmq/ZpVJThJquI8wWayDRZXa8tl3a8saAsNIo5RiGHV+7qzhU3kJq3HYBbnjvkXKGmata
ty3RcqQyzGbNvwweCbRLSlrjZjdcfnRrQvsgUw96gbtLIBGG4SG35NMb/mx3qAfg5YJPLfny6ViD
6MucWadloB/7r00KcjrgruP6GSblQCwra8dmnvcTLO3C6XwTMeZTtJeaNQZuB2Uirtkd86aS5tG9
Ph3wSxVyV5XdJM5gTIWrg72K3RiL0v1/Iu4xlV68weoR9otaB7Pjm8T0GSQOVsV/R3ccT1sSqewG
q7f/ohB1Zu3jZqVRjOUrbvC2bEs0iQUmfUlqPCSuS6/t2v9a7uFPUzxN8fCmWiXQrJgU2WgxbP2E
WLrhXxjZyp/s4XMLwdx0cGbdbO6G8PXNd9huULaDswj/xTJVFXzCjyt6FK0MP+3jii/iKVBf9lvT
SGwAf4f0e9DJf2eueVLBzC2kOz5pbqSjBTu5bTJ+htHA77Z+IURkq8CTDaJcLVVIay3z2VnEOSdf
Aj4dGh2UiPnbD5SW7DzyofkOp4cw6RgCHabD96HynQxdDVl3j2sRnGRQp9acOn7RsC2pCFEkNYJm
OTqDzwh9xfVshhdsixLm+FYiSonGJz3XLyYQRrlPiHOyXy6Q1qyh+OUR+chC2S6AdxevF1WcVYP8
CNfuF4tbYCbreECBVobKLvw1+MzBlReL6I6lEL1Kbus+VN/Ki0EjYHqeumfZIcy1P6SYoDja7yIy
B5P0iMl4G5VLgjUgl4gpXAVJ754mERfGrW+BbreYl8EAFTmD/XYl43NlGCbgz9ZnEANzK5BDOknv
g2tARS18Jmfv3mhm4GxaYUBjAb7K6fpdk2i0vCMR0fsvDEeIq2QlGxno0Gzg2Ghl9OYYE2wSzxNu
hcpUaRBWy9GNw6WPPHd5CeEkfh5BUWnS7B1F3H4EvXIiL5MqFexPri6FI8Z55+7utd4HQE7re/AS
fgf7BtpYJmNimQU77gzN2hyHRrXsHlDyaJAaBIVQha/kSbFHPwe3VgOKrhsIg9BHgyatqZGioIEM
nWCGafYYUD6/lYT4T9Yxv8/ofoIPsDCLrEHWpvy1CDkuTvgacc9+YUhtVsXnopD8gs4n1mQpAcB1
ruJhTS5Ny9rpdqSsawOvMwkzXplJyRgVDmSFL8uQrHb4KVm+PdU4JfiB0yySSQcex08rf3zFPGvw
nVyqTlNmNNz7LyrLnSS5uog1ajLpxG1j4SurUPm2lPmhQM7KnQcGU3jN3JBGPkMZwE+91URX0S16
vIIFE6gvvNX5RqThmgFyLE90A6udgRwW6Kj7hCAr0sNMUt7Ce4a4B/KBiMrvwNiVuBafFNQT4/OE
9YnGEu1y581oF7lPgHkku87vVUT+UlHCwIVyfHpiDyvC5R7eg6rxQXjtStVlhNjtxHBE1acWOIKy
tdqGK380DhsEA0tRCn4hGyEMrH8JQTm0DULZQT1WijuN5EvpAVHdQDLrk/3iySBCsfUNlClXFXOP
wq6f8RLfMsgOtmwxrbuxna8xf2TXCLA86S9pNdA9ex+taIrDeb8mlyYv82isJYWLccXlJNZ9XoPZ
GjV+uJ5JC+XjzqV8d8VGk3iMx4tXkEjOzDPyE9j0b+MnkfJOHsiS/EZjPQcgdl3pKFlGIfWpN6u5
iwQex9WyUkq8HrGhgqpkR6Ig2sN4RP1eBYLqSLHiWGYkzrZdPz9E78dQCyxqYx9L7pewXDyERTPl
pAkO5h+CJlcctJv7v6aiHhA2MrIj6q0VxjD1/hQCpWhWYoBDalxtzNV44U5qiSRY+2OWpJ+thlIG
u/Ya8SixHHoId4LRCCjKk/zkC3mnUWUOxF5rqxQ8A2Bw3CERvGV1RREC7zYTwwo1RlbI54faNihU
vLyGYS1cjs8FRhThdy8JN1xzPBZDzK9qr7OeVaQL+XVbvITnA2LbCncszPyVMTiPFEdeisCCPmzj
K6OLHGjbfyC422XgzAyNkyjF0pFxSIsuOdfyt/k7Sr8t5z94mQkMYt2gd84FbeLjS6PxPmADMw4L
dPAXa21mCjp7/3IvR+yVB6Pj1rEgd+KZGw5z4/GZAkUKMd7bRx5jxNwBUKYXthaSh0cTVfLfq8YF
WWHn+gy632AGctT9gDny4jLCvsYIUUqtEwWg9iaOuOQpY28/8akMekB5O4psqWn30qYqlT0hGQRp
jAF0UFouHW+DKOXriy5w9eRlCTHjOyaZ9WSd5YLRDxMLBoFsxlBWH6An3585ZBKuAF3ELqlJ4Jds
t//oYq/HfL93y0lAdjk+Smy6UELyzlyAuF2FJU1sI491wTDqzVNExJ7P1Vjw9ZKGI6Zy4+i+CqjT
+3hj0fjQqi3zXbJaw2bsui4Hgbu5aSowfVEqkGOxRuVwld8AL7gvLiTO/y2mxHTiZhK5LoALwq9O
VgIOhKXWeAKxbk01w677QqVqex4r38jIYQ6j3Q+BFIiU8s5uoDAKKmYWeFsjju0M8WNMBzGZpOjZ
EsyTMsztf5dN98vNWOaC/BbguwVFcIP7x2/hFUTzeSwXec51nvWDU8mvhcC/AUqj5x2tU+exlgK8
6UYoIiPNgw4rnAXNyl3XOaoKG7z5bJ6aHxKHjNbdv/LYojB+cnjqLZx7GockCUzZAWEPpCcg3BEl
ReDYEhv2yHHDBM5CHvb67JH24XnvvcJgqgm0DyOpCY1F51iqC9JHF06a8xaiplf5TqJ3ymDA/q2W
hUSmdVZkQTaXU/gQlpfPePFJHQDS8JA6OqA1w7tcFhY76JR0Kdf/8vso0zzTnr/Oj3ZrI5eF/fPD
9VpbyXWN/034VFxUMKdqkjm+mW12zpeCLOcElv6tP6SwZbkffB6GMYYIFCemUw+fhmRnp2z4xfkp
02bANYZStmZXeiTEBmZywie6pQNww0jQYUsfsF8jEtchFMYyHrGb2OZj1CGIjNeH+Ar6y11FEYCk
dfM3BK5iSQSNipi/vRY3r3ceX65OPt42TEmoDbp/TKlCVQJ1GCbL7hidXOyT33EcPVw065zS6oe3
mEiZkXHvV8nONsylwd7oY5w6ofiGblWL4EakTOd/4afMEG/SozGwvQA+PrvAONeZQPdxY3Hk11S5
pH/cgP0beYl5EvJUqormVXNF7UL3923zTt7YhKdjeqb2KpYgRWaX5lIw7/s5t9QlTF0WFnF9KNoq
1A2FgrvHYK15FI+lNrmUdUdZPauTpSZvmFr2rR60h1peFWAOJgShxsbl936sFLftnPsMCurrnFum
uJwnAW6uqFI+gbS2PLldaKWy7YBI7L2RgrWMG6uGdRfyJb5/3IO1WlVfKlIi3s0GXBdXnMD3Jjmo
awH/z0axfbz67Z2WNfQjuFjkn0TmWC8BpWju9zcRoNVUf9qGKIXUDEdntJVjrAbuvckVv020I6/Z
Ik67dCNCEUxA7L/5HPFGxrUw2TKqc9htIDaScPXZZrCKS8KiHejtDTDJj0M/mzyEMsFbg9ckAIis
+B7Ivui4gIIeMuJvqPD6SHtiag4QdyUkzBw42/t6XprT02EDm+pmcW2LDjIanx5Ct1eeFETdL/uc
XssewiT8drCei759NcJLTcGPGCttKIva94RCJ1rYvghOkAyfEIqdjR4d16NFKCxf7An+bh2o2d++
lpEJk+qy15Kq7SUgSJDPhPeSpwig37bfpIPZ6/z9odiJvXkam89lHGMtMCKNccCdoFHZbI6ckJHo
xRW67CWDU1bStkZLVrI5yM6JqXM0hk7rAtNr50dziLrvrNRi8z9vRaCm0hZhiQRP43wNngXbq8+P
a71FyoFD9vfQCXQJSgvO7X+k0mR1yL2Ve0t1YjB2sR0Cynr1x2umgs8GalOdj6W7ui4LZJ22bApi
8SnzM5NpaISmZFdj5j22r424IfvF15AUTmWotCuo2DhsCakC5MWn+Rmyjq+Wcj/6L+EIJNz0u7nz
ovQo2zx+4roKD0Ozpnvsw38OeaK9LalKZYDcpUJ8Gs/qiW7coUvJChNaOeubV9b9m/Xkiub7Kkkm
zJ2k8NREsuhMXe5iUncZHHSdx9EcgSBRXFi1ByDfRRLmdJFt4naebGfBMrldaplQAFE4teO+hhSy
whB453JtxUNltEiXETcl8q2g5v5iv9X0vL4S3qq0QURW4xe5W5rKgC3D85KUurNrfuBq/j4atPtt
/4O5ZVGE9VGFIKmclYki369TPaWfUhwSfVRUB082L+rWOR+DNF2Uw3fSblx0MLAc4QseFyOng51Q
d8mfiTOZS66HFWnyS0P7VQSnq202csE89Qf97UP5CZ179GKi0lyy4h4B2/oYTWqWwjE8aete0KHB
sTupq3Ay7/gEZKn7rMScFU6ecJNdRGnnr8h1FAUCgM8Pu7/VFufaW6PFQuPbztay9ZghEjdRv22t
BN46zFC6be18tVcyib3PFpQYQ/8uKp4Q/CZxfuX/MBGqWAsNqVIJdf9uudA2I5sirgn4U0YzjmKS
Hrme/70zNdgfRLhF/t/0DpMbSxYQiTwbFbAY9JLgM3x5Fcm2zvKL4o5YIBMS3zMHaWyVLjMf0aRH
AVZfuQ8x7w+eSKX9D7qysiggI2Z2oCf+ynh8APOUth6xjXoFIReIE/A3D3R6oBAvMNmgLSiocFxq
UzD0M8OQ47+lwStiuAZ1+2UrYzEIzm/jHOX5YCNkWWNXkheVNTTV3wn5mKsTNN6K48FDk73QFI/7
By5WlRtYr78nampzGWZ7Buuar81gMSymbHZbUJ2nlEqC3qcuLkTer19piHcxzlnznS5oaWlzgRjR
e0ZC0X3lS+b3L8HVM/LL6iIR5UbNpkivYF+mXW8LI9czG/A30Y1MqcJTnmLWuqpCzV2D5/PtrzYb
4z+ieznDgz9ZssMyC7bXwnSNvuFYk5knknr5XE52hBjuzZkOleilOCd03Ekya8TPYTylXBEBr4CC
ERLIAeSDKlA93lmAwCr1H4Re10Q6MSOCgeYKKdEhZ8ytQRT9XBCy2Tievouf2pAGr9Jd/9Th4cJv
9F1Y6J1oRqZg5rM/ThjMQ9i2q5lduW+qwhJXTD3EHlYWVl9YT1y45QVLipUj4lzZZOiho06aiI9E
4OW0RJh7DITheWqNm5PDDOoEdVLQ54WiPABfBVu4UdJONW2NdR4B9RIXmdWhLtbOx764/5jsJGxT
JuTtEOwHfa8Zik9uPs2huRhPAw+hM2DFG5J3OsUYAWRqLKIjPpB6/I1wxVWGSFy2f2ILkngcdxma
Rd6cJ1lePdYZ6S1/9SRalB+DoKWojx8DsO8w+Golyup00pBuEKEq9yIgbSH2cCi3UH/nhdclxgyn
T8SEwogT3V6TUWfUJeL7sezTUG8+t8DlJoAO5cEG3GWH8nsEluSD3LAu4PMNTX0TPQKQ7ERR11by
/UKFXou+GyXxjvI6oyOH5bZekVDffMlpsgIc1kMpYjXpIzW8u+ijvVZBMVTXtzZW3gWuw6+DAeJ/
9o8VaC2uv1t1BefYfDR5Nfr+P3o4O4N99OrZwHnZaUYMwYVb+pnKDXpB1VE2zp3WjAX97ajerFu4
oFoay+tds6Myg0S/w78Wxq2qANpKPmj6fkvB0fbCLl+1x4NwMnkm5wzIjhj5cmnEW1f9cFLF/qB+
HN16IaC6FYXE07XU/8wy4oCWHUxSA2/mGt80XfTHqujt5l1it8QP1+hnd3ntlQStz+CGsk5pcqV3
Ebsa6//UIXfoq4eO8aeaUWvbCVTLLJH4UeR6CuqRsxZPGkK3HWT7LJmFNH0hy1UQVa79EEIJOtFT
91w1EfJvr59Ce2GFAQ+NEMBnczFItF/FOEeEyC3ZxbmD6cFGSc3HOB8XJg+omHnyDSJG1pn+EazQ
zgrm6avnEsgLTnlCxFx1dX79zihRW0/TYi9DVqiz+pI7yTsj2NLkoE2fHP914EsC/okNb0jj2WR6
J/O+i9KgpUCWKsG09nAF4yPwNAFeL1ki35Dj+hQyJkSJcMN0Cs+E/NdxFGdxMByYRHHcnGERz0Nu
eaHI7qaq42oezrIMtIfoCBbjRKsS9HuLSg/NLd4wNU7+/8uurhCvnESAeydpPGondR/3Z+3Z+cRt
csI+F1sbKwQa7dcnmGWDiMHKA9pQDMBQT04OieXKhsjNyrHi62rGAHhjFK6mrGJ+zEISc+d1kRaH
2eZ8eStfA2UOwB3spyna3u2cVIMaHW495HMN4jV71ua8l6h+31z0i7VGF1vRIrEN0fqzXShnXUwg
J63ewEIwMr+LR2zjghzpfaXlRd2KnizS8eV7NLNThI4X4pVqk9vgAh3G/yl+6gfkn60QpxQDozyI
kNXCyZtPgrfT/b2wiA8s1fgYWeY5FHe+98XfO4+36VtGCSc+qySFYIWsZgJWgjCPTX+iQdeGMdpD
V4nVH4bsCquCvCNxgXN+plGqTBj30HgB/QDGvr4jeic7dthk6fsn7vLakvKEJLjuJiCCM9Zyk73a
rbIle3V0XahfEOhkw09E/9/bkeM7vuITtC077WTkQIAGMUWRFh80q5JXshSENnqXvvdy0dge+Z2C
Q8XNyAJueEvmEO8WboogR4U3R0kUa+P7H+5n6+RMuhNKuscphYJXv/ahtk+OgqIzhqjDo5Hdpm6B
RqqbuYYvD8A5ZuEXAysEjWHcu8t8N5zwGW0/Ie9KRkewu5be0/rH/4vW9gw44AidSzdr4laQZr/N
ihMkJrxbwnbkls3qYrXW0GmEkdgD7xaqV3tN+IY5YJ3PEcMJ6dcyuN+7H6hbChGyXcIsaDnPEeiA
s1H3fgcxT+Wel0uIHyFGTKX0ycEJ51/Xb7YuYOXiA/dEact2mNmfptUu5lPOBImnudqb+1Dnkvya
HxI/MtSS18KjK68W7J5kbofqOW5pS8C35MI18en9M9xPzIggemjmTkPs/eiYN7LX0ffJNbj6TLmS
39nlX5eIBWATMOv8sObojkswOuqke1GuyPIAvKDNTHPRHiOYJqDtaQEbo22VQTwrpB/EIptc31sn
ZAIE+pcN0k8Nxm3Oc+FwhWU1sGWmTayzlrNbj3AV845fXmYUWC2cEE/2TWKPcKodCSapZkvD3Qnc
1aAwhnpgJNngNnZvuOSpUXFvDzXzuhzPYP5O8dUdOgd3CBP+ppUmpmx43Wkc9RX5v1/8zUV4s21x
x3fkgVth6l7RKOkTmXM/JW0Uat0oiRihn72WfHR513tHKXSGL+d+f/vH54i1DqV4Mm5dY6zyvSkm
P4GrPZMn7cl9+CR9igs8znNHpGxBuLH0kAA+pX4ps20EwmkhKVawwT9GP7/wcm/QYhRbXPxkUmkK
58KTJrcZiEyjK6nqqjkcTs8iTZrADfTpzb7YdJ7Wf5QKEoAHMggemTIYrCxXhdkeRsPgix5wZrtN
p9MhkoZpB7W/eQ0qToRuTjqxyQM7+WlulwIj4HtaoDIzPfJakhaYFUuYqHMtdmW1vnU4sPOQvQ1N
/ZunpUC5U+de9MEP7W4sUl7WU9MqremB5lyfRZJEYME84QXEoq80UdrONeeEMKpTx8b9IITmTEiD
j9tPrIsg1WAoJ55I4MxAGVT1uKlRiRrce+hIoeYToN1lCc7rDP/gSAG0V5iavqtfxwwpR4avCPFz
ccLCILc9WXlbMWdwikNzl6b6TbKQmUwSS6PNlWnn1xa1avZGjAXi2L9/t8VwYLy71J4PpkU0vmyJ
kAFsahMa5FftTd+WaeS8KEAKGcnnPhXMFq2cA1+n1/oUjbohwrF2A7CEo/k4Gx5FoH8wWHYC4rwM
9WryQsNPGBVtyW1sbYFlKVRw8DLTuvMUCsbiqFbjT2WYbw4gwAZ/ReiAcFd2P/LDyOJ8/xZwMvGR
rnNrX8dnbpcAlsiU5iZNz44IP6pVSO4d37LfpzalmyIQdT8Cd1EEZT0SeYcGPeXLSAeliB1caxNJ
8D5ElNRiGCYTZEYCi8ul5Tp8chnjI6QaK+ZQRLkgKwNp4CM/AmzWSNLwI23Tc3JZFhvCw9Xf42JC
1lhGCTW3MN2tUuND6+Gx6whSHolGbzobr7H0zT/xCBaNv8SDOsyZRFsj2AShUadyP80vuQFfDi1Z
TYld8RVChMjMKfyYTfcHUrshYTYXlyLp37G/eot3q9UFhLcZz9n07jfsTNJ2J42RTFB5k7+IodbJ
mlAx9WCDUQP2UjwKGxR1Q2cr6WvnKdxCRlhmEIuudUz7bNt/cveN8MGu4/N7CQbSFVt4O10vGBOt
tC10anGuAVamwnhLYiRtB42rnk1ts6Re9CmM5Yk21R/zsDT2pCwOEH/2OcsXcq/puZjLkaqH/Ms5
amwxmvQ/hvonNPFQnLZmk67LyA6kdEUt93ggEui2lRDD8Xw0Ed61Dly/9tWuzxvmDvCXmmak7z6v
KE28z4myqL+atYskHGQqRLUmdosWPatEtZYn50i32k+omPnE8Ub6Qa4DdLn49DpYB6q8F+ukNlr8
Rvhyv+AExwPbCrp14XvT6N9S4hXSYQIrGJLz7WO2CJ0nwVsnHchXZ4TVE4mJpMX1wosYCB7Iu6gC
bf+nWewq3ct+iVrsbkRZyXNn4hdRsc86VC1GcGpsvMdUhdrRF2O+hO5y6dy7L5+MLfYzkPFt+2ld
ejedW6S7searhXyptGmJvM4L9Yg5uTyI2hDIAeFGsLbDeYc6Op/cnSZQiGLFm//BjeaHD4+YfR5T
5hkJm+3u6qoIkiJr7TFxxncNIRLAhYNMuTIjZn0L8+JLhfGgm7Hw78FWtoZzae9Xxsot9+o6Pm/S
WeSxggtHxqfeircYJRPaHxTvNfZz3dywdBTtk09gOK2DTLPLBg+0A+lLRhD5XbvvbsH1DItFXf+J
oChcR2omF/mZZxcFr1lzg3LPHyBM5lpFOiOgyCOQuLpVbqqmDl2Ccc3yDGQj0chCXTApMdEZPSkD
uGRzIK/NxVjesTlyS3+dDdqbmeW4L6KLNBaKpTepJWOOuZHIE29cukJaUUEGh2YleHK18O7XFH8+
hRzjqKdw9hyVc5cJR83U+GlDaAYuLkaHog3tBVRRG498/8ywKOW0xBWdI1uXubIXhMHw03FlSJ26
0ya6UwZQVu2w1YWAJDSOJhYbLmIkd+Kn0m/QhXE5xjnEiZadCXHUxeOSV0QjB8iWwTqNsIbhVJbQ
qO5AGqNsyiNupfrHLbOhObuBE6BeRNTT6uiHYLiUrn+dqhpbup6GsTlUQMigfzkk6qoxAKONrkm1
B1+WjfhTo1Ozm+ED+nrxMsvOUdU+ow7nt0UoyfEOL7QHSs/X8DTGA6IozvSUdwP8e2lG/HIqE03Q
8ES2Wqidsru9O/N/jIt7vkUMWyXzIV8BBWcW1adyDv0mQm8P5REgIA5TXYGzi/wItS7DuWYIjYWF
14V8XhNrGQaS7IUvUIyA6W1WbyzNEW1+q+4hinDgIuQw0NeBlJylbRJ0EQbZ/fjmv+Ri9AwqXnSV
Ed5QF0VlQDeu9wbizFLs7w0O2dkSzpq+9ux3tu4+NGzYKOAQwdkcNN2TAmsG7ZfAOQT8WwefPfF4
LDEtpYo+4ll63Ov2zv3OwW6jGNZejxL2tMaAWQCi6jM0Xc/Zo4GHL/YcbwxAB+3Pe43xMmYsBoNv
p57/LosDZm0VV3n7DMhtPSMcXDAbGUmYgimyEEn+StHM3gefOmx9LkKX9S9bVq8YB16ngM98dkkk
+qCRebyi+2fv8X3PeTzBaiI6XWlGDmY4aQDJmw6uDEVOEdZEtkcs9IIsfOv17yb5qYn0uTlmzgBU
+R0gzZ33nYAT37YQlzys12BOgqt5GhqkjDZht/U3JoHmt4df68dxuzlvKyfthNzIUmtOv6uHKOk5
DZkXzxSr4N72Sq37+J+6rs08d+HcCXX8fnulGijxj//qF+exxHCSsuOFJ9C+RT5Df9h8sWTb/uls
mN4u5v9wXuNFp2onXEACBxxfwV8hRQSbtt+ukpHXe1U6NzeRgZfj8W6w5LPmuUESN6TJ9jO5mqf5
1GaNjeFYvxHASEoUxlMdsqPASBcssEYCSAT9gg9xxnkoMtl2ZS6FEH2XDKkU8plu8dkdzufbe3wR
iXS9cTzCbtug5mFM07mQBC5+Gfri+gD54S0YIegt7sbvbkXkBV984i461bL/M4BFsQ1GN1iUL9zB
hudO3Z/QZkKyq8z7neEeWFU1f0Z4FOWdr3+FFyb5wIPFNZsh0PdZ4I+XBmiJS9wxEUcjQEDZw/n6
uYtGlG19HVH+S+W+cBwNeL8t245k8bntCSZJWDmY4ntIpVsCJ0Pw8m+gZ33o4OfLTdKIWQGlPjBE
1tfO4ZwIBPf8R89dyfEhtqKsb2atxZrsb+RgPwJ39GNG4D+GY4SDA0VJnLwRksUtXdp1dcGLhkza
vPjl9KnadxRE7ua5RFZWTXjOPm0ozjgIOJlkAUuGcSXJQdpsPMujJ/0JHpab19/hHOWlCFT5AXP2
8FinljP5AkLBR7OSgzVPT4pRPk9Ftj1fFtpgkF7jJv8d42yCPCDUoTt8wnyDHSWDGHNULQJoD6AJ
KCIRdBV86HxDFbrUwchH2GbJgC4sZX8tuo10TJ9+w/fzT14tLmBeawajJSeD5yfZIzaJkNO9xiEs
5AVojo/Jq6aZ3YvF1U3TRO3yjEYJMHgFSwGraTfh07kyShAd3FnHOwFYgQit0PMzlFYPaMwrb+Cj
KZoWbD8T0wcidHaYrEBdrEgoUYTyNs49Tc04IJHHAYyoZ+4O0CP9seuNnxzBZfmsIAsPZ7WgV1Rm
TpWR8M8LjowWi/TXlzF4qVmxW2S3XqHYWS54RhxUWr1RBuVXXy4TvZFh4KiztKWzzY8zZ5HZvU2B
jnUaEGsvJQ1+nqFGb3COdt7jb+g8iSg/y4PFap3UvPK5Kk38BaTe+6TsvlI8wz4WfzM4zHbB6tnR
q/6KFWngvOOcLUN5hcdorUgcLB2XMNda1qxr4J+8HCcA5XzTmgAxKAb4nfIrOutJEOjerWTi82AG
QqdNJZrJKw7RaztjLa1YMbN/JdmVnVks6FOU9ZC/n1CA/SlTQ3TWW2AXZTlqEmS88Fqe+rEBI7VT
Tmys0S2mjXRG/ZlN8AgP5u8GmlkOS3rygPrduIaLlHliuazVSj2SRiL9unOi23olUFjd3D9drd1z
mu7axO5+i7Q0DR0iakBJ7LzGnPmFKPLHrV+UfRMykYMKj93/566zQ1zhzjGO8TlzVLSRrzHrodnn
RkQMjDOMK4Ht6XcIL0v9lUFRc1CUB43AgVJJUsBGleM9kNWRoX3a+YETdbKAmAg01ANIdK1etGhs
YWJyAWaQ4sZ1NTC+TDN8ckxpb/2Kkhh1w0Ow3/yz+GQYIqy5RMPmSRJIw2ZPxSUx8Fuwlp9EZJ00
6px8DQk9R/DSKAy9gyOGXlpMS7Vkswdi0kJN8cybhNbEEV6giI67pPGhzgeycEWFLFePUoZV6nRR
g5V6Vg4jIhntlOtRbV49cEkLHCb0bCdhdNtxLyGToT2+faK3ymoFwBNGNMoqHxVqcYzZTlB41Fu/
y1wqTYeHdSTltloY7awRdtFuHgK9ETUDGu0qnWwoQX6/6sxAfZddWdoh/cCPnHwOEVmTyoO57y+n
BCPcx2XYuNnoo4ZsUOW0vcsQRq7IpyO2JX+7P+zLmiSno79Xo8yUepSyWFz4LgVZHXJd2dOcuxBA
h3R+he0J01JHNVswlUvnkeMrJ7xTtZwL7Z0LY9XMJ14UBU8rofwHufZ0RfaTy3UanwxHY27IMB/3
BQnuSlMdeorJUV+nee9yqanAqP5AscQy9sj3n1/Q/ggmrSx8c/0wsmRCgp1scjxdLChazlGbIjXd
rKdjbZnWeeHVntaQHoiOm/mUULmaNartb5ia8TMCp1y+ttIkHMw/PvARq+EE8XrshOqoNOcMFb23
6byzUnqu64EAGnVQmAmVtdQRhTas+lomyrCSuP3Xsr3amH+sFQsopvprH5mFIJtEU5sVnCShgVB2
c1ib4L7ptc27SBxDrl2IavpC3XG1OOEWve5u606CAcH8/158WKGRUQxJYrtIDDSQTDh6DZJxN4+g
z0umTRKXTAhJkN2rYAeVeM2dyc7K+Y0uLCGIGtChVdU5KMCUlF9m4IglS504LdgTlePoiAjFSr67
sZpNSI3Mq/ah59iXa7oovwlwUZXFXnZSF9UEC24skzh83f4HILClr1qruqAlBkPoRK8mpg6BWHmU
zCNj5lmWpyfou/1AmlwahWaZolI9WoI3/Satp++XxRkNHUbMBQWwMH6XqytLw9/qyzUGFiIuy58F
6HBX65hV4cOYDyxz8T0R+4kz59YnX2jyg0XOHo/bGm6m4014o3B9Yd+zU/ODIVRBBuXSErl5vt04
T9hTPyZ70vaU+SUEkSeiUKPAnS8RlGpFs8SdFZJSOmKkZSzpcHHKJk/rd1G4m7cASHGeA+kfcxHr
9vrjY49evqVBZbjV+uFZSkVGR6yR1FhlSJXBlQi04CyWy6kc+qiulk/sfLcsowgzxxmLBWIVwYl3
erj5GL+aGB2PXZJmkiGOpCHqaBV66o0/patm0uzL9wFy69yxVX7orEnPmgdislewJPswFupLPgFZ
hn2f9FAz1C33QVc6+miMoFiPDtI9jU7IO3Wu6FIsCAkxZ/3wyhjSLl2BQDrIYY4V9BJSg8bJ2O6+
ExFqoNXLnRRjWlQmBF0N9ob/ZVrWS84Y8STOpKjZ+n2j7nzO5TW663gnu5oCQwt1HE19rHev0DCO
ZCXbpWJnXJuZVAWfwGG7vveAamWURSCl0mxCHq/jtxzpbbwP3s4cbaWZq6TEdiWpsqps2XGD+KSx
wk7sxQXXLSpdOP7DT2iPQ5D8IOf+CQ3Ej6FrvVpJuzDI76BUeuYN/EKi/MhtphYbf4rnrPPV5Qj+
Yzc4ZQ3DNh0wyJwmBotDvAQJzB9YZGq7GptqdFv1/TXpMeEpSqRW0gYZfILmazE13tkdOvQE9jle
TqZJrFhxYprJbV3YRIRqfVuqFWs2PWFeZ5XCOQNn7029sD7PaCewuOqjC1iIP4nwABtFimgKC4vi
O81Gwu80d2HaUt9d3Jrvlf2VHgW8Tw6mVXKnUfGZ6+e0J6k/AhUYroxIEC1NylNBFXI6ix34NCTt
s3Ten+WARISploK0wXU4tPqJPtAFN2hqoR8rmBw+LDkNxiZNhVPybxySfDpdufmfrIobdO+Rkte+
7XCkxU3eZBE+CO80HP7L+dkJihb0+gJJuRl6NmeLZa1l18ftQ6i/OIrtpzVOvfCOct655vNu+qaQ
YY8+SJz91QZGywZGE4DjRaGxHAmlEuhXeheacFuqRqlXksYCG8JLYO3axVF3l4OJe8g9domOH9bq
JmbAKB9pViE7bARfCnodLYjZma65P75ieENOqpxIRyhyRS9m+ajH65FQNKu8jnQBdOadLCb5l1fR
3kzujLOSETCUBYF7GKnCUZspojgP00NvE0t7s6XhD1WV34FtOwxCF6IEfOA2mqgYzwYnw8bRnFOt
XNpm69o47eOh2TbIa/qOcA6OmjAHR1ehVz5Bwb4gAkL3tuHqy40Yo5UShssaQzxA3bYI8QvJTYU7
FdLUee3PgnGd/mcB5BaGMO7gi37VH/BhCRLLm4n9b8064wTe8ZfF4+cZOrVrSyBrR53thFLQ1U9q
2WV0OPSsqR6VEgER0GPdOCZF68lCVQRgcvZ7UmHlMjdpjeTky3qBQqsgqEwtnEoOaQ5zlB4Gfd57
R1n7lhZYvtlEuLMOY+bcsVXRL8eVgYxQ/rttPrUMDO1xB2AVhW7Oa1KEczzHxzCvlh5CZiIaqs/q
1uus9aL7Guf8z9/9VbuRN2ys1Sk6LKCEWh6gdyVKL1lZKZlbqcZuwbxamkA8lq4eRqXGqHpIAAcP
4Cu7Uf1fd2M+6Xp5hDxOLjcPfS19YS/3EKhaGJ6DJkgJL/07YVPRPEiaHgjfdme2oO8OQbElww4l
KH1JlHpaWu+hfe3rnHB4dH1fJOYjiK9e5vUjE/DR2b82YKesY/ZGJZ2ehdHTMDaPJwd0yqz3KfrY
j6OjcY9bEsYzz/WDWaodvU+gmK6AECUsH4vli6N9ccCkubFipsUg3onrs+vxmYagOdV4KAZvf4JK
8E69yfvHUhYP7O4UyD3n/3Bj8SWTFgOlh+KkCdBXEXRn+dGkyEqIN4vaQbr4azQKZAYTQ6dT1yN6
sBEvaxE2ngRL/v7FCRCkNIi81inS3f+hnWX9PM9/svOHVeRa1ajmX5ylIy/GcRK5OuPUFquABJp7
ux1eUL8HuOqyiioS8G9wcY+EDR2IqC64AQKVkHCR5l0sa51SyjtCI6JESxAVkXGDvkOEgkMd42Iz
+2ZfqZu/qFV6AvS9ED5D8DttzVm2BcUPT20SB9ZbbJN5Bm2W1x5KygAI+1SZ9cSh2JWgsUMJF6WO
I1vo/Z//mW0ViOP/B9MEXDIL88okhCzs0lObMTfV2G3JpxgtTFsZGw+7k89qbj2g9F9TCGDQhkIo
Tk/MSoS1Zyw8N1+4NR+A4Cu+BhuZowiw0pmmvQQul1hg1b//2D0hhFR3fqMNzA99z6enJlyF1QRU
7Zt1/Qx9qmKFsYvSqeJBb59vZl2fMiITuciq8xo/eo1E+1Q2k+CoI3CYj3gsNTE5Bdl4Cr5tzydu
FVl/dNN4Cy4s/eFWmsZuKH+QKgFOx+8z/hI+j8ZSgs+fy9T7ngr7TBymNREA9K/GsK1yVg/zybCF
jlBmL/zrItEfWQI8yc+q9iOAkb9VznkjUkOSN5CGEIBqp+w0UDzkgBqg+lQwuFvbWWLi9zFp7IMQ
UqxrjmmpplFp4GDE3TyY0Opl4KcrP+82crpRVjpWwUBvAzjviDzIE8/ZRu54jJIB5t8vPX78OR/W
0YZJBrSiLuNzrzzDAOZbbz4dfbpig+5V5afLD28xPXgyBD5a36IGgqF764q2h4zuXcySbztXKdrL
staZClf/Z+zA9WuDwMeOWCIZz3hSB4dBOAp1koXjyZKgwbGNa0jirC5ahE7YecbhiA7XABITUFHc
1CwTsuxBcO4dC5HZ/Z12k3gyojzN4gmrfa1N79FGEInnbUn0RyIW6ilH8DyYtAYqUjygtRCOnfcW
ERkJnXryE/L8jDxHoWVqFgjJudICQhHV7wgPG2H1jfebyqo54i/Ors3aR0Y/I32JexSNjYzU2zPo
QyYGb7gRTe0VfDVRes27Ls5CHPcYfJhtV0Jhz8HB3eRB/TU4ZdwLtOoQKaVAm3bdoxTS9MC0D/Rb
XsAigDAQAI0jvqDDLxJeldFK+UmyDB90oeUHV64FDVZFdS17JfHWdVz97mo9aO+6au7tPQ1ufeBJ
w+B2B2zxwdjbFFCIQ5KRI2prGoBclXk5tUOKdNWzrbetPF0fqrffEn8odyjoTL7fPEi/zJRtSuTy
LIU8JrxZuIu9OTWYJHTybEOXfO2aS2u50YJN/7Zh7uGhPgInxBhKGuqfeE5zKmxPNBtBjKJ+BQvr
RDEjWed1sECEq5Xu6kM63U438i9IO0gFcoNt95H4v6u/1fy9JnQBy9wcT297XHy0MYX7GrCmK+GW
NdFwz7gLUX9QeiK6Q4JwPXbIboGV+l312qCTt7rrnWfYb9GMqCf3vW43C6O6tAkwJnIcgxYxSiUb
6aR7F/hRGmKNKZvtcmvN/+fvIRGamUJLLxmTq0F5KYhWi3riNl790+9d9ZKGdPYFaON1MaEhONtP
69nMEj7yF8Tci4DdPddYk5CsejuJncyu4qY0zd8WJU2Veke4NCzxH9DIwiNh5dxQKuX5jqxw7BlI
yIkUy8s+KX4RpqCvSu1fqBWCwY9ugBjnPSU0SbttFLCHz5eos/gP4lRW27BKg4+uI1D2jdxeZN2O
mBfle0jsPwfAaDGNBdHCyGyk/yajz9bjBqkoZ4sZY/1EfmrZOqx1YcW3iRuZX+eW8JvxHLKSbbQn
ajFwWAIxVZd23DxvnHsIHE6kpuPU9UukPj+ZAvosoCQ5BeNGL6XUuJaVtOsvFP103zICm9ddEXjA
AFSb+KwKXjqftcXr2t2rOKVMAoVKf9B70YkyD8mdubqgtMWO5jYiPI+59a4VBSj/vJSb97OXVRQD
nXc7D/9QZVfkhcqxURA13zBfC0ojPgQJZqUKNj0CbOPCDpYTpMsZpM1hcFNOPCvhQsu82PMeLOsQ
jNTeJQetULpZLSpGV/BaFI+YVyKsLpymoAjTjOsgPJjGswcFE9Od+OVVl8dJYLzbhDDAOrcrv6Cl
P31tN88Y1R9niRh+VoPgcJUOTc/xxuu6DUvHZ6IfRYFRAt1q9hR+oVpMsN/4PVT0Q5GNe7VqwCOn
JFtTW5a9ubCSIVclwh+jqIwWnXtXu4zWzhMYL5CE0D1fyVXIw3XGLEWGzr9stBr1egYhYR/23cR/
CxQUmIoTf9Dmu3fKz/mDbWW/lC+WohYYZBDFeen/4cW9pB7dGocqOISZ5srf6ezNws+IxSYopRS9
+tWj07AIM3LyBAQ0KwsQvowCvBpMlD6myEWaTDSrplbZBz9P5Ge0472OEfSMKn7Tq7yvaNW67WNP
uH6aljBAxgDqM98P/utkaUMRbc4kqaX6BEk2aNeOIqHY3cNlMqd3OK6RhiJ/+V0aI8oUIh1vFC0i
6wyisIhLK+eh6u+SPDocsICFVYxNZRo1wks9g7uyTesRJ7J6FX7OdncQnlrP6tGi2OMuBbzPVWpt
fvQgs9ZgzZ8hNLBek3rZ9/SwqbbvK+Bqh5OsfxeyPlhGzwOCt3s7qLiw1zpH9AvNYIbszbARoUx1
MbGycdoe3yzY2I7dmY7b7cFoK7EhlGS7wSRDv3wNTkO7BNbkBLXpt7Ls10DSNaEF1xtdmNRnO3uN
x7lKFMcdpVW5mBpXETrSIBfwJrRCI/uIClh9aCAqISYkhaosjMTETLxBAcekE4Qjw8SPAi7tNa6T
IV/p5hDiCSmKOG35PUeJbQ+5mR/H3rOXIDx2tOOfA8qOxNkRdABKejxo4Dsgy1/ISfZ9uici5Xtb
TfaDYlRhhrJVG4uboFdcDxxICMROMXR0XUlZKW14vGzXhLkRqvuCrt/gBycwQjCsnK6J34hEr41m
+GJUfqSfV3WPnuSMvRkkPL4nSg2tSjkkhrMiVkwYsll3kgtsy6wvnNNPVXKxY2j5D4keUEsPbWAR
R2P0bBngOVNHYUkMEVE0LZQkd/0+T0fXDplwtCfigdnpl6cdBLstcRLeZWVWSL//Vt7AvzTD0YUY
5ipxTWjVb1NjRgSY6Tc2+qGpbsfIuX8IUgiEMzuA0pP2YIR4sgS2XwR9fsH0PZU4lIa/brigQknl
P36EH3H70fYoqi+QRseOTVbbfTMiNlLIgp/sCOzU6qsr/0pv7bAgLJq5g3bz5eV0KAlYZOJyS+e3
Q8cQbwQarsA0fz+2+FnOQG60RIQ3twr6Vf/+Z2hXl4dZu8sBmiE+bD+lGKtIVolsAiT1mua+s44+
2cMOfBYzcemj/aKoPtt7u9F+C0UaMpHc3R5QMUdaRJBKT2tDASnKVXyJXMry7C8fRZAi5kKfRSnK
aJx6RSjYExFxeaYY10z3l9teeW9uoKcD6tzQTrKzvpQUQR0sS/MYX3i4N5S/NS5sJTGOitoy0ya4
1aVTA3IrL+z9pHLecE/uFq2BEPOmergnXK7hgl5CyC6qIY5AnzmgVq6owUjWIFUAYs2IwoF8AB9c
mReGY6xQgsofOAjsaN87iY5LeG9D3K5Gg8rt1cbTtpye5zY+1r/4R72NidhSiIucmz05UVQGHkKJ
BxXWuKjwzOTQHS3rz71JV66A4KCcOGlyTBRgyLEzUXYWJXHlmqSxf0TeeuE+ZfJ/VE/XNc/Th+wz
xNXt9m754RmU5gYZUFhk8LrKGVSvOtyKRYcM+J9k4n+LYR3I1Dsx/l/Gl76ruo8pjr2f9ix//R/Z
NtTAQ9p3S97vOlIV/se1XN/4dI/MdYHhhKUE01XeONQChyiZRKQ24T3Udsy0K8Lrcx5nFV7UaPsu
F+fl0ySb0mv75j7Ctfh0uD5wx/e66l2QYPzCmG8GVaF7tiekSAnRy7rMOicUl5YP7KmaqMBQLM5z
99EY5TS2hd/U+vZSrI5vDQ+5/tnD3Mi1zk7Q+LwNj/D6uNbF4bQvMY4IC/3rfPMGbZ7Su8J+/Wx4
vyfwRS2y6mjsD5IA1saXan5Zan4Cz+Qv3HEXoWNngcN3xQQrDyubCR///ZV8+npoMH5fFjee5avX
CPwPOYWUIZLm6tGauLHR41rpRREq0orIddKWqweI/zXtYelrEm+CyPPtscE1kQCNF847n2cZV5db
4E5Ne7JE8tf7wNX6Nu8ZhBDzBGiAG/4/nwitrDMac8QsCsWmYot1bBrexMpz1vc/emWlolBtK/45
OwlMnfXxvIiKqt3dje4fAtFBOoxy+c/2kFLnOIxBVGp4y56Sg4PAslkso2ZRQoO0R3MB3QMDYiD1
SNgly/oKMNashAMUpPsUWMqL7o+KtDn2Cr5p87OKVoW0AdP29alDU6Bqh68Vfdfoc0dghB4bIUCR
rM2dJhHXUt1yf6aQGOSDhZRZ8K4brIQLWjx5ZmVfuGCDSePfXtRlrMoB//EyTuwmzRE9tZv4cFBP
Oyh+xrhxtAvW+MqgO0s+rOfT250ChBpbd86sEJuiOYgbiTszFQddxkUhy7Qx9DD0B6R7r8uGEr5f
6kSC6ZuxcSgL9sp/RqKrzYKm/+NYJ2xzhiv1jCh3sO0YJ/Wu4yPvNpgMjp0XkomNC05ewLjtiyw/
kXCJsIQQ9YfoKNcerOMvXVe18+LiwBQiZhH4j3/g008flRQFUk+aPQjHtGrl22xKlwDeP/St9kk8
Fi1U/9B8UrwGQv7gJZf5igKV3iCSSfjrWtAyfMDC2BQEtQ97UZjQhbTpSznTjtr9t69Es8qnT/RR
9EgpcOA70qfXH3w44KeBpzlVPC5FL8ab4NkzcYucP59Ra7kpQyfhGOG2oIJmSElN3u4vFZI7natP
f/mFmy2YfTeXsNgHjOoMhsub2b6EPAcvwPOrfu4uK4Xvxiierxo6EZIDf/0aYyVSffKayQf6KB6i
NDt5n8Uy+a0ndUQg9MtvpGoZp65gOwJen0MAcK21TOwJYIJx1PQz0nTe6ZQtvCrvolxViv5CogFD
Rj+0JTG1y+bL5IWR35wRK3Ujk7K/y91yOcRC4dflTV/8EGOonqr3Nr6oBx6Z8c71L6+zlywsUL2X
HDhH4/Pt5UmLJ4Yhr0FB36M0SC1NWWmXcLzgVcsvrKTC17VuO4PUkSGOHjVE37yqrxNDFmZRk1kP
pUtIWfb3uVWjvMkSgNQtbyHyhnnNe+L4HRaEj+nEvY2CP2rgTeYrMx09B2pFJFdt94P9T0DEHBXS
5g5KOhuw3Rxr8CHkX2GFyfbLeVASxOY8b34dx0uTJ48rKGrfdDtNgtHIqpsnzB7D9y5SuJencJNI
tPXR6TqNJfXfoA5qCC29e6zyLYvKZldtgOqdJSLE+cGD40t41CzJc7I20QQX3AKMOnq5CUrDeWBE
ReiFv8HPIViPUXZhELKKHgQWIw+QlyRGYjSO4fIA7hZ8qV2M8XNtYabijfCoHRLm0ejBc1zYzsLf
XKQoZcDfrnFnTCqt1kh1648uNEV30BqKRSP9JRkAqHbvJdHkqJJMjFDrBizQkKq/lQzUzFfNLVwd
4OI5CAl3kKb13fZmMR5kdRQOwfEUR8CVfR//8B6doS9yGNrhQMxSCOBVa2+IzSMDnVxEG90Uc7C2
acHsrkLD7aiYWc6tFOuZOHR87vUZkBmZWTJ4K8ActnN+TfHNnFVi4BJFWXAsXXdXW9AOhWFHpLdc
Y9g8UpKKbCA1Se5IsCSbYwv6KIZjyUF6gfdXZRSQry08CPDcKb3mze1Q++xgUQF/wrz4iJ5Ms6lv
tC53/At4oQxQxA4ZDX5lZt9GrdalVNN6l1H2mPP2MsHGYlX2rb1RC7LOFSZwiW6lMvW1NyWFTYnA
3TLrAH47f3swL4yoVWjxy0D1+rRfznOZAIacD9As+l1r/kh6SvOsKi/nPv9rKCgQxMFHjHv1lDK2
OtkFBGCw4n07ZXNUSgFkIHYtFFwENhUroMUnLHbcNL2Z4FmkwSLpZCFxMBsJwboRpnGRQ1sFXOxl
JCq2f2CTLcA8o34UcaEhHSrhuzjdjlPaG57f5MYkeQYhMZbW+110RbexK1nzy4CzDHspD+fAvc/Z
lMUYzhrdG05Hxe8j/fcgVuKvwPet/O8wXtJhYLH++lGmUtWcgzg0VC9M1ZUogD1hALMSyU88qv7X
NvEVJjtL5H63VMeaguA8sHeqxP0w4Oqr8xPr6rbo+P3772LTQGu/PskIAsxOGSHIzfAu2E27heXl
sqdu8CIusEVC+Z+nnQ4x9Y1VS5ZszQD/Gx5GYwVyQOrSLWlNCmRbDVc8M0HuZ8B7BbgjZcVdsM2d
wBMsqvWFTSIQUwFntRxncBZGhy/VMUH8cczBwKLoMPt2Uze73P9jb4nJVzYoquS94IDV+b2CZLR3
6EIxq/8OVJrI5QWKi80zOovU7CFZHVTKpCRL+tOfAkFVdHSacMYMP/2PyZX5jbB23xoqNDUb31oI
oDOcF61FU0Ist5GBTMmU3eTQO+xcqhH2UZWK1bWjHRq1AY4ysn18jH58I1Xt9QKiu/RFyVzIgUJB
dCAdX7Lra9EUqlyIKuDLZGbgYmiagqDtEWiBK8p+cQtFTN7rcZPzorF1+UertqW2duEeVUKMguia
jaIC81J29h5kjhbGYrbiWVoPml2hue5kIfVKWSV4x22SR+v+ITXejC3v4AeP6/0tJR8CdIwqJEvd
txEDFrMzBrTXE6CIA5pa/JxEGapqdKFWOXPK2MReHVEwpX4go52+rYIZo4aqJzwSKnLqn1vPm1oA
J1DhvQbFRo18ys+ZqMBicsOL0vV2vJ1F2rm37Yt/9llcmnrJ8owZR/cB97gT5WsLrqwrnnZ70DyA
m8YR4EGnAoQpzu687eVPi0ynTcVLX4yLQfwQYTs+9Z7E/3Jr5t3cGuRjzTAiiO6hryG7pN16NCOd
N224H9D9HTKGJBQ9cC1SpWnRFAr2YPHjZvRwnZMyB6IA1eXJVrMUsqQBv3obb6nIQ8ZXZD7MtFu4
L+CErMfW5MYwzy9dq/2xVKMjmCwzGb12tDCYlb/dVFapoAB+osasgYnNsosI2rxwJ9UHUkhIpwHV
p6Rm5un903iafzLKTBcQ7sC4ZG1TAQSZuaTx1/+91vV/h8rQUTn0/N30lb4oERWG2uw8vCk7fzDp
juQ0IevObjlaweeu2F8zgghNFxlAlUaSTjlvOpOAB0XZL7w9NkQGvM4qmKWMP6lLA7fEmhjH8y6P
VgWI0SwRqOYfhY0wsEWafQjvjTshrMc0p9ckLyvRmp36cIAA2Xaq2GADhcMrN+J724MQXdo5fSkj
ZnAcch2sLevMysLvW0+G8cjjFPzqURUtyyuBmIrJgLvqDWmpEXY7gUUT7sgkm6Fwci49ieHvvBk5
F4W9eJmOX1GjFZKJhQV0ykZj7aBbhJB0GnyaNxiytG/sIGDhbBOve6aHjD+HlsIOXEVbsfHZrTUu
fkK+mDSUH/Jq9ZADYEF3YGNdGNPcLC657SBOLGkKdG5qkdg2TW0DNxwy2DtyLI5Ig963Emd2nGs2
+D6dJZsuqz+cy+W4g0fDc/xVfYR5p1SnDID1zsYed00HhNYSr/UNVmlMs1MdrsCcI6B2Kj5A50+J
NyN2m07IMLDk+lKXS/shoDIZ6lsXdTztMvYNNj6e/9Z/S5EAPRmjU17x+uslTLQs5TD96I6DafMI
tPx2Dl8qcNt0SR5jp1R+Ni9P6GRqORTiwwdkCHR/zzpxAcKajC7ASNCBOtAlsY3/eTKZG02+f6De
ZcQh83W3bv3IIJeD2t7/1fmMyO1t7/kJltnr7275CRn3X0MsBtm1sU8gy3+wYOcShoSp5v8NzgLF
KpSkWTVlX6oYojZL96Dvy5NLqigxLaC0em0F1Ntd36NbYVmThKXygDT8Ln5dixC0ZXt+Sshh/l35
2UJK+7ENoAN80njrYPAufGedSzm1zHidpuqQ3+JbpftgNaiNDUEG9xcLsMRa8xJhI70doYy/v9gb
MeFTYyUY49SsO2Av8ngsq5+ZTrYhHTHvPGIlhHHa/J4wCjuG7h/nWoJIyOVtVsVZ+bu2Guy4Los8
VU7NJwypYZJR/Rj4hwRT/5v1I4cGjB7z2uTiNW0qoR685v0bHD17FcLV0CvRQan8Igylt3WWU67H
9UEvz+tMUPI7AcC3Pg0WlJwGubH+64cgZvSeDE3BMfCIyU3uN38UMAJyXWAQRLUjhdkWqXukpL1a
DWBLFYWiGAnT8UpJN42E+3oePzsRXKT9Mf8Gc7JJyyyzazTYrv2rbBBCzdwUyC5VzMZvX6102g46
sDmSKJOoh/q+MsE/DZ24I7ZzXgzGOTzUFo4HE+aCld/0zYjy6Yyki9q6IxdazvkST/eK3EDOIknn
BRgd4HoMy59tcMyC49g+aNDDSjzkIbNTYOUxbzk7JAtBiw5VoEKTJWcWP4ynl7LTMvHKB4CYrT+M
hG1hFaqyyfw7jtxtELPSPgX4F+aRo0mAGCjiWpiweNbntjb+YPg6fOpLJwHKnj7ua555NkeryPZt
80OyHm1ZeNxv//e7bL/BLvMBchdRTrDSqGn2SXUUvSb7qdoKiT8V4qctMG7rMQNpr7NzEsNOZxL8
M5IdcYHp3JzIRlLZ4+ybu/KL3XPINT6uNn2eqs7rkxGzg3xLYUxB4SQvD5pCtn1mdTx3fT+DWzOK
AV7zOKcXOn+X0nBJviCyPwIDsVh1kMNOwQV2sjUeJ6mowBkN/DDN3SdSI7oJKTAYo0OZr1iVzp47
BxWr/2Nd5fR7/7G0dC17SKxgGE6AsyAeZ3UVAkZ9GdhkpaqnxJJAKg7X0/I6h2wnMQPvEKAXCD/p
o7TwcFGaCnSMlF7PrO1gTsN9N5d00aD4nBkqUQEbIhMJ4Awtp/iPbtrpjaT72HzsBtHc3Ea/5TGj
cVxLGMuK9VZ7yBI6cnK6YMczwRZODx1lhrBEbvKxCkDOkFkBNppsz2clbwKrmtQeCxtkqhwSHa0J
7/lg3NNMPrUDvC5AJ4c2OWI+pCyBYdvqIRTuLg49Zt3Xa1qfnOtbCmc9P7sx7hme709NXG/v9aHn
y+MeGxg5cL2k/6npLuIeivBYHsQ30pptg1NqpFUQOJNpeatWh7G1Ahq2QwImZ05phAGngUAfnrYA
UYA/HU7aJvffXVDkAymtjEuc3mfj2szNuToypX1ARNPe4GfIkvS07gaYVX7JyQlvPpSZQO0m/luO
WWyiunYnrfSVRHmQEA+pTsJuufoC1FD31j3Pykwk59rQt9NQBpPHAY5gkhboMkJ8QHf2qKcj19+k
a6/yKDM1jnNdN81hXn+LycPgoyETak03uhbRkWumDfvXp+o6ljtmEVQhcw/IhI90PmSgU0xfT31k
2Y9DVL6furJiXhOVlmeqb6VRyfbcZ+c3B2fIjpe/k2jzxqoFiS6cQNw2UzN5H5h/SpzcMFk2QfOq
525hWDHVMvW8NvC68bqb3D4Fmy2d8MsfI/olrVk7kIF52fWRTuL6TAtZdFSaAg2bMh38xXXcF4k0
J7yQrOkEdRMZB5SSAjjeVvKisostKSPJC9ue3lzmwUcerYI+XUQFVFfbgvlprtzcQehJf9fgBrAu
u0QIyeAi1VC2z4b/kOmUOfsmBgKgtaYykgLCMMpT55qNioDAd8MWFJq0ee4uMoIjJML6EUgbDSSb
RvpseEYuNL5dwmVXPFx2yNfR5Y+1MFhyB5pJgNgUKmc1RIl7gBpv/wQ/edaBG/yJgfqxO90Z1PUb
55hsMCB0UIPVDnuh2B2Xm9PA05BqzLsS7lbDnjC7MkTJx6dO4+KLOlpIb6l5Ejekm5ydsU0LsdW/
Y2ACP6BO5bkS6la84/5CmFX8+4czYB8zcCymO0Uxs4lbJIp7QZ4OefeoxQO5eJUDbiaRSYPHDhh4
vJcNGhNkxPP9964UycWi8GFYtY4fGri2Bh2xebbgkWISlf0Q9nin4Xp67OnjPzIsLDnSifffcZiy
xxs9oVZLBS+jVHe3WHwFYAe3GtK+F7lRqTsPpoIbs9iBuapzYLbz7GXshoAmYGsFmC6m6M3LOpGV
k7RXXBfhwKKxgLIlcCtw08x9IwyCTbPGmRoM/rcKAGL2Z87UMe3bLlFMMGuw8VxN2cb5gtVtczD4
9+R0rBMlbWjemJJnqOmxNinVRN46gHiQYhXyR1o0m8Av7ciICIODbl5UEA3tmCyceJh7cOFkaU7y
Wqi8Lb+aeYsC6rIr/Tgaq9j3BwVyPClTyhz03kLr3p/RkGsaiSpD0yUvOVqn68qpu8CqeTxnViAf
0XcSxlO6EkDNJHxEiJIBuIYikRmOGj/bnY5UfOhiBBEthbtsyC7RaBPHduR0Mw/M9KthBHpOADuv
wGPdv281yGPYQKzwcfQlketLu4MD+oRobMWNWMfimrdE+wRGo2EukzEWN4y6qO/l8jgwEkvWVwQy
kteSd29+wv+s7RxLK42LKCPHAXr6LBjv5eL3WmlQ6jf2NlEUQwkFPpB2vee8m4ynWb8hFpXgj+56
8XDONpxtyN7EpxZ9ubqS5OWQbS+KznmNVz1kuo/sqNdSCaWIrb0jVRPamAjcInLfngXO+9ZNq7g6
fAOtgioRITzU+NyIRPzHD9khlLT3GCQrCWFBGQA8tI3t4VQvrco1DS16VaDJQZ5HwIu7MSrrgqGY
z3sP+lrrCbKDsMDdVgg/MEVehNZEH11nU0mGjfmupHrsx6ebBENNZI0NfbHKbbBeAb+oG2ssIhUS
ZqFqEErlwEvemKaf9wxocptMND6f4k4gEGp3A+8gC9/7cRJFmRfwrrTyKYckn3gMftCLxkLyWrXe
Eqf3/qB7Ghxgd+7MIr2uegEgI/9DawtQ6nH2phBecy/s7oKeqTgQE1uYpA8NtSpmfgl22JR11dQM
YOCXO26gz70XwuYdo4Yd84iAZQnJ4Hcnb/TRgxd8dakxKX/Lipa0+MozZRF2UF5yIi9fahdOhwa2
f0OEWbK1uHzL2EybKzbFBRrl6H/BZlAWMCBTvG38LEpn1BLxw2/YvqTa/wg1Wj+tIx7X7TgLawcn
2bYuRMxO6qMhbgJ24UqODJJGcU29hDVlEyUqrPYERA6BXsY/sqWIjd5gCBBdZwnEIup6wmj38sw4
OtYXe1zA8y4KCT/w+TzRxnLQ0+hKX28e+z9NDIy3C9ogoNJJJLXXZpWHQo1c/3cjx65JGivWl/e5
3pMyfFqwxHKFTtkH7hMpxuzQVycfeCB6LIY0WPANRDU7sla4rK41ZWUBpIZYTb3mZ8K4vDF+kmvw
4P66hXgUBo6CI8AbwmCITJ5hY1o3fYjfdeAztENarxEoFJyiji9fR2FuJLCzlgzmHq1zK9zCbIzJ
a/1aAi9GlWUvU4lm3pTC8gfFBUukAZXZyj78HbEAehoqZEq+R4wLE6sT/lhRcwkc6r7AIpTsVoop
NxHahwBFBTEnnzoPl3IjCnzEylDd7ej0ZJhkX89gHr/PWDh9MU9XdyanMmS059zypWCzC90kr9Fw
KoLfFFXbFYCqjOdT59eFCVJhQoy6TESlBjpxkg+UtOA6XzpOIgOki+EGAi005Z9nKmRCunGmn6v6
Upg8VYSLWzedQ2G8QXytZS+36Q3+9x+lBeBWEGC3x1rM5Cmra7Ng5K+Pnp6RnwrtpxsUvC0KO/mS
RQGTqmFFWTTyLPFaZ+c7LtEhrBSv4LdJajHshaXl3+W3keSgZyYFjYM6KymeHoXbm8/PvC0f3icW
gtpPzITWEtagqFsUm3RtR4B3sVvNjGZaMIoh48xFxdMyqpyGyrZEk3EgSj5rLCvChC1xHcG8Hydf
3OYi6cViD1K0Wf3JHNBzKyxd41yBQ17MZR4+dswPZAfPmYkyO/8OspLjJG33BVPnt5JcGtjBZued
JLlRW7r1uBwvyQJ6kPnz26mJmjAJogUj740bYkJFo6n8Z0JzCMXaBg7huzZSz8zljV/aYhOwwEzf
iHN8xZmKq+hDcxDrlwlmGqAuEhOYxX3yQ0y/h+xmu04ieSt74BxXAxWmda0Yoeh2Q6HbskRB8jQV
l0hF6AuXt2LbHSFPNE2sBW551vA0eXDYd9pIBkQBqDn8EfOlHypWxV56yzX0YlMIm5adkGDbrlxC
BtTQ0mVWk2PUt1Q7dgWhE1okhkoaaMHF09XLYeHZalmFyQZITT7ubr9kUilvZNlYZVraW/T7GoTT
2I0vVBC3bvWWuXB8bGJJB7hFBuLoRC6IIMyOzXgSQYFwpgx+/LBRt0wNkHnrzifduYHNwTo0YdRz
TaJRG9fngF1IFrEH3rF5q8zSNt4iiXvs8i8IcpPam4zA3RHGfPFifX+Ca8egjgDHnKZjOtCP1JGs
ytUZIE8N7pH0e02NjiO2MKWGJwR/yNDo+GjajnakZHr1Q+cKje0xdYwhqPN2cePs8G7RgRWrV44v
k9WxW4wcOqKG7x+B7sNRE+XYU1egQ4poqg3H6leIwDwR3Palj4UYeZOyH76W6tIA2th+N0ukg/YJ
r/GvZtGrepnRXASC23V+Gz5KtmTeCzuv9DRmP+C2UIq3QCiRxaYjwUSscD7Sm6dXfjGuN1YgxzuO
7156n3PPHeBQQqC86/slOblUTq3GXFKXkDXy3KoE692y4gjlUqKdJnUEk3jn5nmwm30KNYbyJZol
/nofHu0n9gEp/H4wioXVJP35dVQ8456BLMSfZFIooXBVs00YSt+1jEq1dE88NpLr98dcJ9qpM118
q0ModbLrLtuoIWz5yAsIGjulHJ878NVyO6rW60chszEC4Gi3k7WLI1FJBN5SqVcHDYxxHaptrFhB
ybnsIzJBxT3jjCin0fLx8PPY4klvH4NhrJcPcPSuXln9GnrDgcf2FHQ+OvIUXN/J7sAgQCWjXzJh
CaYaPHD0w5pampAhxR+XUaRfTuBI1p2EB+AdlTqEK3VF43zTIyfX3bs9lGmIbJFPrPlJ0mN9q9qX
c/CRkCtHMVdMSxBVHd5oNGUpam5ei8VGLoE8oZAKT3NQLNY3kwPuL0Z2QN5UkdHQTdnH9MiPPLZn
+lCijy+1pOppOqmX4U5rOaN6EqrHSW95Fx9dWzk2jwM1TpBEwz4NKP1O0fBJZ1913pHnfKOJAJt8
7raUfvMuOF8LhrpL6+r/TvUwequ+FUTZsnSuGHg88gY5Ute4ogfiXpekS6jHuHkSMuLzn1osfI9E
lHBRQKLd7Ji7VyxV4i6um7GPFczcKF/X/MX3Ir67OrM9GdAFFX+J0utcV1HA5WjIH6ld/e9j4kOX
qRnulRVuFtX2xVFHVKzeVCH3eUIMdfX8jq6yuSiOUqp+1+WerjYuf8+nsodTW6cuF2Y90awI3T/9
AhdpM6vNKfVKWgqHds02/CSNtMazk/dx3GIC1sl+JZIULYN2+UxKbhTtJlfV0ecifEynWDWgQ8zu
rqNtfd7z0UtCQBS+ew1TbpVI7jiiJcuqj1Ifv/MnZ9raioXHv/PGl/tedah1LMYGZkGlGOx8++1P
8A5x74PuTMpK4kP/kGvNBqHCUG9BekrXLujKOSaXH0AIYc+IaG4joCA4Q4R0WiguBLDxbBRQf2Fw
31wntSofm8Y5i5zVThN5XzX6wch3hmohhxBm0MMC7y0MTHlzF3DS8Tf/ovyBgBrg23WYCt1L9raS
QU6RadddIXxrnXXZ5mHjgr1rW+RqhY+RWUedbpp/TPZJD42oOk4thLj22sGR3F4fXW4ijYCWaOPy
SxiQOwloO/+bpN+n2Es/L8mRsS3rWmGOv0wfbjVwptp1BK0nn+wOXdt71FuAZatNIEJJEom6FQ1P
g/aEdwXwU/HC4SudIXyXiVllpvp/61qNF+YtYWo6DUbUm9UzMpYx4yWNcjeQndC8N0WPuD2qousJ
sEKPZTHbhel+brSmXUxzVj9pZCiDdmRlB/8MovBtSpIYo/HWmvq10OvUMlo0js8yirM65rRAwiNz
MlO3G71PCmOgZdUmabyutGv9LWVnK/ue40hdAVFmfB1F0NcpbUui9m/mqQYIgl2FyLSKzmhhdEZD
wWk4Nox5czmVo1+yhGgBiGJAIXVtM9S6E+beehDxHFqwy/Gi/J9ugJjCVWdhgb+bBguq0g1YH0wz
+MAqw4X6Dw8bzcJGDdi03Ad1eJQF3hvAzPW2pjWw6UXdh8a2ZzRPijcOZ7xnk3mDgnjE6ro17/D0
LYqPyJr267n3v3hnCfiT1EE7REddt5YCiCuzbjZc6hgeF6fKBtpJpU1p+RIr/iU1KDz6gysGeBRp
wHAssy32wIs1NI4+T17OO0ZmkfARDdU/A43xY3UWY0VOTnlHXN1XapZOj5BhcM5zW+K9FFAVANbR
mZWONghBsxX9xiHQPIqi/gFYLQSCmEnLrEiyiVcBpOjrXDLGli0GWGAUIpBQ51N2V3vK9027rjiz
tn/ZS8yusRUoGIjPL2TYZY4WcsXDUk/gzp+p2kE6v0cNgbxq+wlAAISzgZhaF1gxzp2DYAlVly9I
wh9V0a8nO9nn42xaQj5X5NW+rELsT4opl6jDQg1pvwmq+gHXCrPKrBDAEZ7pI3O1k3aZaS9mx2It
gREmPOcqMLN/igt96Jv11th5tKNkq+falUe9us8MYYbLqr71Nchi9bVW1tmQEPg+rjIKNo4oMYgQ
xsPa0dLeEp5PXXW9VTald1ZC1Gly1mtNvgRoDNrWXaiWpFE9QSCzUo/Th18XNXnlMRwycNEihGtJ
bA6cu/EvaJVEt0cOYnN0Lk8l/18jM9aqgM9VArCYupv+VL/bDd8szR5fiPZx8S++uvuYGnp3lAXj
xBptYsGmphsVaA2CA3V3jbuyBtwyNwiioBHsHTD0ZY+qz/Wzqc41PvHvXdGHln3aBGeqCe+4vJ+2
gIoXwzPojWKowCqEhLkZEzH8nmVgxoNfv48NYb+xDP4zBkrCw0SpM44epEv8nCqLXR/AGdyfAk91
D2QVYnXjz4Gmz0h7FiL4JgeM1Xctw+8tQSWj5yB81PVSKNvCl9nG/lQEp/4m6nCa9MCmf6cccU+t
QjcV33Sdb6rFOy2ugb/2BQ4IE6xVd0X1BY4mvl/brPWIUo8T+etsw1pgNUutAbxLqcuwHdeid4jr
FB1VUWOVnKLWb5I6fwOkXEdA+sHXOrIJ4rTuxNBZyOk3y4z3Xu6aHCiWyWc4s6lEJrgVvoYcbecp
8UAaQnF5D0Grrl6CI6cM45pseoHu/hhxrJxE44Djt9choBCmAlXb3CaObs+6lOyrK60wWHNskFKm
mCV+fozAqPuGMcQwkeK3h9X/rORCCE0P9wP5cVCdXDZS1Ikaru227w5b4CuZQ4FR6FVS3pDpsck3
sACLXVtzVi2Ol0iyhvaxx2v4Ekc5V0nJa6wHVA3EJW+zI/2AfzEYC8ZikvUsuutpOQHxTDH8VewQ
UxHBr9vUm2TNLHC5W9sosJRvYsHfjOD7I7GkBtDaQZ9BHHCVpfjrbOKSj5pv5fPIRoPHhBSw074z
Co2ueThfwLsWO8protPs20Pjzn5Ne+ZQumRCERbRn1Xser11Ut6LkHHOiDWlnEKEmaNQM13aOghF
Uzo6L8viDZBbST5icPt6G3ZOWXEx8/SqHJAoef8G9E9Ag3NNGBJ5IGXIsGtFcxJAr/MAM/I0e7aC
8QIZLmHspk0HR/Uncved1Ux8VgGsHhRGTHXHw5f9DoLkDCW6aySeyiVHhbV8btSMBL0TEIGuxTY8
C7kLvsbtHR0Da0oY8XdnJ3jnqydTeOSwTXLwUQ/t/H/p5N0No4o2ASDBAuZx51yo8cOSQstAVY0i
G38qmku8b+/XmTe8sS3Ye8Jk4vLsMpxZg1GKGD8biujExZ1JjiUFniwR1qowJSQqWAw5Rk1aOs5q
awdWkhzEwyyRaOwwNWQc6G5lUHD5ihGHSA7H5JtiPzCkK+NaidnGFo9yQfbmZSIt+Gm7DxFZTdnY
zPJ6J2bRYMhjbdl3uQwdfoMxHphISynfabfiuhbseI0NyC4AeOeBkXPu45z0l7weBhcr0ktfsHPu
nGdPHSj8VqYcj/MUqsnUf1DozpohJLgCFb5WTvh4xuRRAQPLrHj5CfJZEl3QYpLGPxU3F9/QiB5k
GB7jh+ni8gD1r1Xs6CaxepcuZJiMLDoKerlL58K1Lq4/Qj5JZryEOj/vt2+bmo20OrJznJ1H2Si4
+GiGwgpg3mbHoh600tuuDajmT804HzgTeFZLgJxlkSV0Zs1YiHXlUM4rm+Ik/kJ7Ee98HhWar57/
RC3ahnTVAMlM4/IXq33e9UmD5RGIIgrbPKRHA5t7GFJfMoTCnUjp8qkF3RUNAiKfEAyYwL6DJ3Tw
SG3IdrBNSv6MaTWHrYcosQdZHG1Kzs0XXMOq9oBnTkBizRlRH471mYPDIdQemmCEC+YuKEStSyyJ
AylEEgDrnhy/1RQ5GEu1E+N2Yt32oBBp4flsFSIzuvHqUjnMVzIdFUB9gIxYs7M3WIx9AHmoaFGZ
CEXVAZv+1nKzwMmMWaEfmMpwnbVf/8pdJ2oRXzNi0xJSqAr0P1KIjp0YHOVXxxDihJ6CjXJjbl9+
nKoNO106oFxMA3bv1hL62+mBbmiVsrK9Kuxzu+Uts0XBajRNgDqV0yE77IPv2c79BRIPwBKycUH8
nBmBG57efXiKjhoHNRZ8LnbF9HdKuWJJIaMgm6R8F180tu64MRAgkFdz1gB0W8fiDs2qC2CwOxug
cMu+qN4qSfSNp93aU0oxSlh/xe+ou4CgklKx6XlG2kLSP+QrULF87o/AZhQ+8ZC2og3OpufKBNjw
ed5pXgyYr46ZUsqAnCe2zueTSilfi0lDQqfyz4JZPaRPCsh3A119Qb9enDtu4qATemX9p9ElFDXG
lkZj04T/ESpRLT8HrU5Z6DgHhUluSVYaHIzuEeytoxnlUGrnee/4uxkd1Hf2VYFnCmc8eJIBR+03
yigzFahcp8/x0sL06N7eG8d64fMw7pmH3+/NFTxFuu2JYkz3JoEh9ZkAnDkV69bouaelOQF6cHTs
KGSU0NCnNdgoRP3j09T2HHStMotfQHsV9QyhtTKhhy9kSGWy8b9MGrar4FZ89SFOPQG68anK+fod
n9sEfME3X485oTH4x7qOUxLeQtdFIw0DQtbBV+qzMw1KHezXW6boFNjcx1auTJcdJ4Yigq8nRmvl
fzbC/rcbva+D98bgC5e+3018CPwhA3RRtjlzIzV1iIQMScN/8ed481jkHw0YPYvKEmoy2/NSP2k1
Ii8ar0pYykIo06etvofp7n4qjlmLNwXVSJrdIh4477WJy1/LNFQkDes4wveuv/uWgsaSB8OmoUNs
liJbSKrNW9mCo8udJW6vTRctKEBjx6rS/B+dEYrsxFOa5rt4X6zJmDi5ArpqlkqrtuT5qeuLQXZp
0F5hMDT2ZnyxrTyvYB8iEela2LpVwz4NPGfXQNEyvf+aR1updS41wu2X6bRRT7lo8Vl/mZJbH2du
ZFEc0wJuTeHalR3hY0X/JP4KZnhOwvb+KCbEth4ouOJDc+kDrTfAwJvDXMaUqgrURkcbpUW7JY6z
VB0oxjLb/A6g0zEsIh7gIGBSiCoFlJG770Jtz1AMkdjxxi9bX1k4YgFra9nfFUC8qyQwOtenzRaw
WLpdkdjtGByr8cKfuQkiZp67/L8zgMzu6LSLcR6G27g8yq+5NaOz1rpQfkYAUtrSD5qfaT++nRnV
rLjyzKtiJnNS9O63L9g3sJlTEDp3EDA6bGtjzCfbGYmqdyG20OqTAJRPoLN2OqVT97qsKB8mFie3
D3fQIxQJPAyfw45r3Y+uemNHQBMtI26wObyL0pNLStt4rQsS0gOs2VlB8L+/2wlvEOjtsl8IcNzW
9T5xPAjLoAhDHVY4PRVS7gJ0iSTgBJMSKBsGW5EaDtebh8b9IA8qKznkIzySBRbhwkpsgi0OHH5n
82Ijr3Auky7ITsCRwcSIlGlKnVSdF9T2yHtFNfQIt7M7U+5w0Ktf+q4xu8V2StkecoQ/oJyA5mAK
B/v6vMctM2D55KVV3bSQ3+v7Ej5giuzPjm1FQFxel2NxvaI7znutGiLLAQTimRDZc389Qo9V1ejB
37H+y4ifVjStqrR8iexWdCxci5gOCyTxss3ne8AFVt5d1nH3KXmnXc3m4CXZLPC2TbOh3/Vq6jPp
ZRdN7c2O3JUpJLnAF6fJ3tflmZ3JFitIJZ/agXz1fzwxTtz+UsvGCcjpQpbf91GVaJaiykg2E0PE
/3jhZpM3NRJU9PfsFvmgyNjkfFnV1CQR9flr3P/HN58CSUJwBbtvHPRTY46tfYdMa9OCbi0GJcH6
4huvy1z9qW4XMdBy4VEtXB7OrruW2AEAAYfbf0b80JuQF3RfBjvaSL9rUVXcZPw557M8Z89UY2c8
K5zbMWUlTooUb8DMHPi9z6xXFd5QnTzS9lex0EySSREAHRuEhocPJXh22i1OUIou+nOMg6GZZR2Y
MsJ1dQTJ8qOpqQFxrZ+wyayLsPIZcGhKD0iiEmvd5jznbGgBnOt30YJGZiE7xj2h3Y9GhmdinFkQ
6QDf0uJ/2hEX5gpZTwLR3mS1b/T23GQcLHRh5Z355Q1hNVreDXWFDbY4nsWoUe26QGCdex7gzt9j
hA2XVEZkS6JY89VYuSWnjtwPpt1qgKfQs3rmc4HfTPN2MmhV8wSCi57Uo1ooylG/pLeDPsnj/1JW
dHliQZIWTuh+AkZdPO2FSpohIDkCBIZPcgQVeaKMGKfn14YT2h4Mw4EBp1i/1cTnM1BbPRk5+ABL
jgqWl9KWvy3n1oRb5N/oVjz3l/z38PbDbtAtOGYApBgVHiova/bAW+uzQ+TTjCtcMoRJZJnZIil2
KivggKye2PKXii2FrgIDu+YxNQS7AfWJRO5iKb+E/Wdt7eOkAtxxpdVL9iO6rSQjyUTMBfASdOQU
8ChxFrFghWSDLgXT1O7PmIbWoPUZ3gzbzQAtay2oLpNG6TejS8xpYtQ33/bTUlyrSrn8OtGO2TAC
HqtoJlPD7wCq33oUEHeC3Ta2DiiyQyVJfyx2vOc4u6vAscEm8Q4sWim53WglPUR6n4AUvLZsVy0/
4nZ5PFdBzUjjd3KA/W2DcO54LC4NK9tNDt1INFqDuS6g6dgh83KdExUdphtzwvtJzu+Q9R4VonyH
DOFAb02q3qakoxbc5eFDl7nkNSFS09Ch7HdbT0qXJq27zgZqpvXn+tQhUx+UBWOL/upmvcgk/1+N
W6Bc8kDxr/gFWZ5faf6KG8xxC98Om1tvxbYJhlpK6Ijr9oGxgQAIQu9aC7oVRWek3MvyLv0KK+bl
WNh3GqptS4cE3KxPTJux0J7vVS4UpTNyvY24ShFm8OzBSpoY84+Sw0tSB/KUCTDN4n4QK/AVVYMo
rrYr08ULhjOgi0u7FF8Ozc/jouvacf1slWa476nVA9Pt2xPyg/4THLQcdBiDoU9v9M6f8UDRwiy3
Cb/0NkWdu+cz3hvMgIIyJhROlJdOP5w98QqIM4SLBnDVPBmh//rzrGHKxa+d7mSMISHj8A6tAH0O
N6GPw9WlUCFiuqO/BlMoip3Src5Dxiksnlk0yVb8yKWMqJQ+54DGJ3k+VrA9mamDNfh7rz0FWzQk
V7syHEKm2HmNoHbetqaHuXJk3MQTlFeTUqU0SovunnfwxwWAEMJls2Yh5DXaJ91XEWSeanGJknqc
VEjD+CRz/6evo4nurN4Vvzj98OX0c0UPxWaRE9WDoVcHgFi+9aAD/gHaooNChJoICqVfk6nJAF51
uk0wk7HUVdKzupt7DPjmq3xu2e13tFHTJPWVevGBSCjN0T0X8E5kIDoGzfp/kk9AdqcUQkB56OhN
FX36lJlLcu96fl3Qu3SoV37r/evfGTG6Qpc3WUkDrAhR4OkFKz9nngCDULAYpnJ8qzcNMgE2Hmap
b3ubLsqBLMOjurZHfDO2z44vJ8B2Bis5+vWA2ARCwZqgbxicV8nNH2XTV+LIrSEopY+JeNPwqSOm
aQen3QDT7pSFjvy0g70gu9985HjbuRsQ+qNdPkYuiFJW5ZSd7dLIPEC0BB8UUDfsX4BpU11emK1D
zi/FVgSEUyt3xLZsUjtCYjPxguiw8SHzpWSLthOYWZJmGNnL6xr41IH88t2qkKX6uIgPi/P4pCns
qz4u8/xEk0HyHjnx9E8A+SrlbZs/AJLwr513/QoSahkL/BtwUeBpp+VkFWH8ftuH208cNeJI1xKx
ZUHX0jKEATM2wnQtjEu0MIdCNZtDNv1N3TUgLtrPAO2i50+fUvsDZVmZCNXbJ8Vb7vAWg2AlazHe
y4qgArJpYC3YucR22sdCdWhpYbtH0T6y1R5Hg/ZQ8C8FXPxj6ha2x8nyvR42MSAiofVnpPMSZAsF
k5byWKgvJiyyCgbvxToNbwjxQRxHJLT5b0x81utXh5yBCP1r6Z/q/8uh6SuzbTUiE0U5cf2B9Ikp
7tlL+gz1E12xjO+iHInDs6iPJ37VJ8p4k3E9qQQ1UCAxFVJBcnTFmgxpOASLoifAAWO3JkfpQg+v
QUGIbFjH5KP/CI15B+nMu6hclswXffFWw3bxzMK0+auR4RzgkAbHUCXqxBx1C5fhZVLl81DGCzM7
EGQ+pEf9F03Fqomdyu6jUfgYsXGzN70f6oZgoQ5weL2z/l7b2HagcjyhPpSBC97sFT66Gji1Ur45
An7jS46GUxS2ao//px9KXCe3E+oLT2A0vrj+GSgkJ3gBPZ/iVMN0w7YEXyo7ZXzaENeOhUqtZIC6
KGPHW89u99aFCSyS72R6qUXn6wnTe5dNdmyVXyK2Yhu5b18irzrlwBQ1IzIcKHnR+TyJNnVYt0R1
dbzarrzSTmF2/EpSWDhhEPVgBiAUK5K1dG5rPwDVP/7tuic9blapDVxC3xykD75CzSOxbcYc0g4U
65u4hwdUub6EoVMoV8I0BeABpUQ5qN/cA/lF1LpYn2rM+7LLoXuG073C5/srgSZEnnvE6sqB3mX6
hYYrcnBVcuAljkDHOtvvXmqhDCOcwIRClhb4fCcPJ9oMBmpQ17Hh1n7G3rpFYKM28TEgpmbVnPVV
8UklO85/CCWBj60uEPhbGKiGdw3a3HaukFCjuH2ZqXRGZqmuPiZCC8KxXJPxHHmNKfq4J+98icf9
a5PFOMJG2oiG/g1anKPyMfI3359n2c4rbTSWjrySAmyjHEEPeu3i7XrINryodtk6iTKfLkFlvTI2
udMK8kvLzCJBfTUn7RJKkzC5F07sO+76hJLAxDqDHhuLArv7l42epqeV7KQv3hqQy8/FNNM0YGTM
0+cIHYhWBQY5Wmfs9foO8Qi9b6vsKhao0NZ+k5Mlj9CR+mIV5XGFvDiX2DLV3X++/UZ0a+ZrwXH9
E28F5hURgiEBAaD+RT/k9yPGuhjsfmgq4d/VmEBN9YRHi55xwQSueC3MOuqQNtq5NHLififSN5nb
haETXa/JUHTniyabQYWQ7SFAqpoGa99gYHk2PzfzWSle9sLO1QC1U/ZcF3FBoxWDdREdFUynR4AU
34P6m050pDvi5jJZoKxURWE6Wt6rhAUt7KKxyRgcuZKIGf3U6jG12q417HeBsZiVkaSUJYXPIGZ+
2yucGdOI3ijQ5e1NnNn0JgDfOaTxNdV+VdW9K5Vw83+k+crB+gzGTUoaDByPPhZhYf0XBmgjJjnG
+V0bGFF5S9PpUteyJLqSGxxT6rM2zOVssWVBRKwkluxhuehwo9xner9VxK/V6Sgdl1tVYaD7e/qX
HgpyfvawbgZrr66dEfke/Rw/j5wyqc8Z158FIuG2mel6BsAHkEHTsAYLvUc/R4U5/V5MmIGwUndG
AzUif56gOYy2wqbKFqFkUJ83PZP3A1o1qFokDRTkgOmOYxyAi0xN0RvtQM9butkH4P5X0aBMpi2V
KHh+OvhOezMuzdWTnWaH+ugj2GTssRhQIPEMvyaK9RNawxdsvex8n1fRKr/mqwfE0lCKfUKyPjDA
PoaksgOtoi//Z11BBHiug6KGk2XlTP1NLpGdbLPdZ69VXX0/czI1bEOa2oiHAZunKSv2WJzwZLR5
f61uaoDcyHG4VVtgmZgBTOH3CUks6h4ryB+0rN6RdY7cmaKSUOEpKcHljLP5P9Qkv/XfWFwRzewG
BlQZphWDPgYHG6QkNkVGM1kQYcbjvY5+9hX+lcg4FepbvUgqoX+XFQxUObpsbTyhqvZNOD8ZAv05
jWyf7HOTQ6GutuFdDAw4p0TPgdrUNtQXz6TUIitooYfBLu9s8/dN802ws7O64W0Ut1ou99X3jFub
4PiSfCMHVJY1EAY0PrrGGwlZ7eEijFOM2bytZAH4pBN9v0g1ceBnxhdY9+/O+HS+jjOw16Yk4l9+
Qufzm13OMy/xfq7PZ9Zrk5v0C/M/8KaRlpiQlIPDueT+G1DnwfOuhnjyy4yMmc+YL8HZAy4drkM2
k+QYN5/lGT2Ey11msR8lh8TOAKrlJ+Fm2cvGH7PGNxiaYNk21PAcSJbgUitVyZfoKqOL3nuJSmG3
M7QzO3CEO6VSXvEN0sLXyhhOa27i8m6X5Xl0oq65QpFC289olF7s0Y/BNQ+dTfURXL4gLf++3q2Y
BR6dfgqJwMcIdlFq4HngOt7wE/TsRjypGlPhflHoIvErfqGAIcdG1IEcOK+hcSKVkDd11jLqqPwz
pIeeR+lcpqhqH8nmXI0d4ML5VXC2XeKe526xVIoH21PO6vUc069LYT5fHNZUiUxrtUtEF75jfWA+
oKDLs9+8+UJME7htx4xeAiG95F7ZueugTcBZLKfHIrFVmjghXNJzuugwHrE1aGmQAA0Ae9rP9EZt
6SWVjjU0VKCW1XEEsuMXtVY38DRaCfOOPD10VXUjRt+amDtmWetC8sRbuGYW2h+SuQFZunLcKEX4
jCZsjvbFT+xR5pC78NU/EQ26ULzQX+xrEoLEDyczCA6Rem100XCVLuH/rO0aPcrLZtpHHlMbtxQi
ndnDmBcSSJ8VwT/AtK7C3gkC2HInxb0ZmzCZcSXiEKQFPuiuivtUsPZKeompP2no72dVffcGXpmH
OIUSEIYau5xX11WatqnOyFJH4rs2dO3DAZDnIToRjw5wUrWvJf3Bn5JBtJspfn4wFp3LO9GRSWLY
DeFpY4tYeVnEEwAYN/oXaK0tQUBZbUnt/N02ymK1JNXKOA/cEA2drWt+LsoyndC2ac1uz6zLtVY3
/VpT6e5PRpvpbbyp+0Uw76NMXxjJB9yA5K3inK4PLOSkV+89HdLANd9p6w/AjIwrs8jagBR6sI/o
zZ6LAcchgE6isW7LY1xytQsjceA0Z/D7iOmUf/TNxh4xDH/7K+703jyKbYa5QG0P7hiUOzDTfB11
5dirJ9NlHfSzPhHf7mLZ+XEr/5sKdPpH+Ov5XH06JRdKeotGVb2WTMqw78U6jRGdMkDOHl32Es1v
2xePaGFBANSqyLEBDsyhIyah5VmW12MH/CA38cBj6ZdMmI1JJwjV1S4BnQzD+SjAAoWAq35CjTP6
gB3oIkOxLHQJ8g4XY0QGYWQW2VpwahJlUv6tw8Kqgmo5lXHSJBEJMgaWBuxYj9J5Fw1RjIfNhk4W
0bG9Iq5fSKNKWInLQXpQtbE/mWuNfHdTyP/EpLZ4n8GKEXtiLkYyRS/0UbSiuRiv20AtDAnLn6NP
EWyC+qJ3fjOxEhv9LbtUIayx2TPPWG88iMdsO2m74mn/ityPL9BQKnDxPFQUwuYZeaMhTFWiBsEM
FWOEF4mtrg36DObI7HZaAXJaRWudS2rhTblAyb81yLgKRB/4mpcbGmWbAwca97MXmr+O4dzxzr4J
C+tOPJEmLRNDEibj8ROZf7RyVXtL/jI/KPZd6tVb8VzDlR6CKfMTmmWTk2yjXqvAAcsAnIiiTf4A
Da1VD3zZGabtXf0lLpYZ8hXqsQhv3QefWfpfB1R8ZQCCJBGQ4zmKrcamA6PqAD9E5F0Rwp8BSngR
ygRt0c2Li63CUWsHL1uLHK99Vu0hCEDdxVhyQqGn73KOSgsAGyb0QkYc22A6eBD4oCYdP5IpSfS8
2alXPMe6Po8pax8R/qI7StSXBJrS2WUCN1cBbONmYdJgbpkrnvgIDQTvp+o3YZCg6VX37p2k0OY2
VSZFAJMPOrIBNFNlDTIPkVZa16BbHT3ZawHvrLBAGfXoSvJB+Ru9Cwt+kBe4Y/e5WmfzGlAaUpe3
p8Cajei19vic88Nc+D7T6m0Jeijgl2N7ltlAfDy0VgBCK0Uei9ZUQrKlY2YYuoZ1/4JD22yMAhv/
rkza6fikFYsGe/EYI6rFqfBbLd/DyXUE7BfbBG0+kURSTgNxUKCk5BAw6OWv/mt+iMeGBwjSwYhy
sretYGA3+BLMTgNB7Z1ZVZtvPiWe9REYpYsfmzUScpG2tyWYunWwWsT6K1FzK6HHIkMH0UbcPfeM
uV+G/nsBAA/5m2u+90Eq2GHJuFtnHR6AY8j6IuoUxr4CykIJl2nJaDuIL50evS4XASFsaoqIrM2q
Kat77b4mmT2GYmd4fTvHEjpd/zhx+ffrBW0Nq0UpLXP+l2j2L8O3xYF1XYi16LrMsL7FH7dqhAGx
t3ZeSHwEiTVERJVvTtOan+Cqjz9qt02ytfArzFPlM+3Lex+r6tyFMUD6NUB5o11aZnjZ00AiPppq
S/s7wEA8GYmrp+wdJyAv30oDpUm1Ej/v+SfK4AJSWyPyLlDsj3/fxbrCG2anO1cx9PNoxNNvwOOl
MH+QUERmMTMtxtoKSNk+0H0CADqKHBijN04Yo6NR4nSpdEASzwp9+D7sfkJizL2pjRGQvALFv0qD
5yCxnGMS3gg56UH7ABI2jSsQtcQM5HKwhWooid1wOjQGxsW+hAHZuYnE2ctehdnl+ilSyKlPYN0m
Czr7F/1QJpazOJmtKvuh2cRx5BLAydyFEXLcZr4q1VQ7DI/hO2RM3FHlGCTYauWqheMoBnp320VT
0Ys7CNIvjmghhopYoeFe2o7Mqw3yjuWSXpKvnwjLlwrdnu0plMsuekO0GSq4Kt7vRickW/hwsYJm
7iH7w0FgMwqDTX000vMyWpQI3VuuI7Tvn3vSlzDRZBdlE1fukJCqcNGW3vkniEbEzcX7gv9efRg6
J808Ntx2qwm0f93jkp1ePsnJvgjlHJL7X6vZ5Mmbz0xM2Of64bjTRLhVs8v9elsuxrZc0+a1sZgM
wVGHls99LSxl1WyuWrFUaFl7+K2VNINUkRwDYwMvdotZKtuprlqjpJtcFK/ja/xM4f2LQZmhMGn6
6iCrFbK6bxJoOnHyWX1On6IJ52YSXtCh+41i701KS6cyz9HS6ZWszxZwfU6KSMtZvkC3LL4Ii4Z4
90yvih6XxbHw/m9z2gfj+k8S7pSov6HcNZ+wcEz3BD+t50X45eBkT92DSS/+AmMYiqA24AgNF+9g
gI6LqQQ5hidc3UjJlExWCAPHve5SsLoCTTaYKimEQa+984DLvvuGy+J0Yls+K4IQ7Q/jEGz/+JVn
4AFa6WKxNFRC+0m1zBamXc4FOAhiIkl6DXg2LCfj+dr1aerKI885KRmNxWIfwLEgz1lf/osdTHCx
csRp03oYd4c0MufwTcyI6Dn1SbHdaC/+tQrJKyjZw5a8b0in6RojC+7xSzHvjxFp40r5rQuhlPAf
TJyGOixMQF5zhbismLQulEsYGm/cc3RsdIFqRyEMSOY15OTWB5ZP86hjJwYn7bnVgrXOHrwwqBLA
/xNbtUpAhsIuOIH5T5T/FDaKUzYfUwfrgESLSOcqnsZClqV3CIKJ3UCnKRXUfuSw2H7XGI8xRDds
83RSiosK9mmPCMSI7JmjMHl4E4zEFqbisI1ceieTBrZ2VQxPWnVAyRXpF8xdwFVsI/GrusUzYL/d
2RKcsZ2tE/Y+XRKBCiFA9dGIECsK1gDvx6jQJcfbolTWw/EXfVIVyeWd+xVg3pXKbP2Koq8/f06O
4vXVK9u3XmeZDE67EKrPEQgNbIEL3RZSnOikNx3B99fiTu4QEL6u2waidT4UrxthPiu7mMxHE6L9
zkp/MJIiOCdmvNTE4QcAqEGDSJdPuL9AlloIhafYHUGzVFP/gl4EEb6+Q8Lld8JOW5gCoOSu7Vm6
yLnhsHkZcTg9JTI9MEkORnJN/950e0d44GEFuLHo+XbbUNWgX3MlgAeA5DExIDawUXfcfPnwEnMc
qWNZJpjHokWxpqbfw67SaweLGmGjQ9ZbAOhk1lftmiuC4pyrYHCS1QYACO5suG0o59JEr09z0qWn
TzfmiFHPgF4CXS2tQAdbsVQeJbP5jjfl9eIxKioCmjOqMsyUELhqF+IY2qz8YNrTwnpqvAhgQW5k
9+l0Q5FNa1Gk6ewJE8BFBIKQEBDL+fmbZPlGoq90iFTm5mrJQZq/+LOPkOAaUGOIbwnLPsHtwnQA
ZPIDG/Zlf1RpRHkX8SDWgbE/z6UOjOeugf1aH8yKfarwyupZU+9eNVjjc12LVVhRTzxGOhY95xHu
uBbH9AlXaNCNsWivPU1vmsDgeoJ1cjdZWEdeBtUJnhRjs5UtG/xhTAxQ2QQmW2DXoSE5p/uESh0F
cydf/GyEYlveyYzLVp9fJ2rIOpljA4IL4j6B+PEXfCHUg1M+mKs20rOhRLYhqx1vwLc5+CJDMBil
LQpsDU6cIG+/2JXSm4VtQIywGTrnz0wNfylyGzC15IrHW8Oa966y0Fg7DWKYllbPIHpL7ZyqMmpy
Lae8CBmrlVfL9wO5vRsI7ul2Wl8tlCc9blrJkoTa9afcP8c2lU1gU03Xa1V2OkmYGLWVZ2rmdETu
KhgMoTIcaMeuOIeeOSVNz25ckqXz+kGSwUxdpP7lEAqp+OR6mW3Bx4RY4xaVFYvo0KkqTICGzKLw
0JeSiAhSF30/1iWnzcQZoRfikmjAQlK4cxENUmOA+qdOAnqkrfjwTjf7mmcZ5uxSDdWb/cqMdJcq
mMRJbLTlHusqK9ei92Vqvn1L7kMICUiqEasIFv0cqNSx9VvACJvtVCEXHqDJ1I7oPVJNuy2mJuWo
1lmH+Tcdda374a4j+sqHeNSImMfKBe4lKHd7pPwUVFfFqmAV0wW91iMCpHFusE8ftVO6GI3oV7U5
JThOpHI3bGHmHq7YZuf1w6FRBU3MqjyG0UyVFm/yW1H23nLpR4dUMpkhgjF4AmEdnZYC+4DvJRDi
QDMgQH3JY6tHzWLZdHxDSp6BrvIJId/XkV/iro0uQO2UtFJU8uY/Rt8X97vP0iu6DjF7WiCzCxsO
S/b/V5nSxA3wHbghrKajaDyDemu5QDhqhM3bWHCb4LHSb+sVVTvwP2RU5SbUjb4WOkqks1btmiXV
Z1mk7//k8FX9Oj064MyLmQg6mASCjYomxe2mitCIdi+g4Hw7nTnPTPaFgDSE1/Kt+2CVE8tqpzeb
Bp01qRA5Qn8uCkiYTBPiwZM3liIR8bGvsWcFihXiyORaT9L2pJ4IgLBupwNmOSRRDvbV3KmFQIeO
omHLwjBhuYfvrHmjpGK81qEdMQVEC4gpxP/2/OM+1tJEZRhGkn1OFRU3APRNytNRlBS6jpSrEM+d
dqaHFdi1JeMWZ31bkSv4327CtytDi8yYyFdlAsVmTrtPGH4eQXT3F58BgJKDe69IpdTz6OP5BUAw
ywK2xVotldQQwlGPF0c2evKG4kYJV13rD2qVtuNbEwyioPUAcxWDnvGQHVfYGSUKzrK5VPrGHTj0
DpzubA/B2U3YEcH/xIGIZoHHr84T8GsXywwXzaFa7PMxCPpINKmVU/P4BIEz2Z6tKcXFYC7Ngmw3
t37OFkAlOG0uF9kDgl3xLvACEBv+vuFYnK5cvgNPQzgpO0blSa+tOmgh2A9wkuymxjq41Kc5xKi4
XWIZomc4W7d6sblFHnDNmbEccSIVKQQWPR4cTHGNXXAHSzjxsgzGCZfr0d4PNr3nLPP5ftLOh6Ti
pQDJGI+TbqT4cKoCh6p3fayNTa/6xXYFY2nijXIrNov3rXE06FCMr+C6kBBw8cik51+W3O/8X7qK
BkCFGiEr2Axm66+WVQQNE++EkW0FyOZ+7lrVesPIayXSY2BdQXMkDdx5opm+zF2WtCd3Nx1XYgH7
MQdLN5NmDUfaEkv5ZM1j1x+yG0izSMZzxiSDw666xDBXpKdViY0OPbK4Gop2wyrwfHoiEIuHCN8N
oG0+nRObP8XmrqsAu9nIgA6AGwQ/S5yuCq1S/UwA939GHYKHI9uTgE6A7aPcgllqXWAwbq3II9iK
LjW8GNUXIzcVB97wkbhv2QfUEe4xpNC7GG3X9/M+UB0lElIHmruCRnf3eLC49m1JcfdaX290sHkt
qGMFQDR969+5KrhU2ZXvz2D2pIErijXCVHVARiwqdaFBuPuo/0Ne/dpID2JbBSv2xsNdHi1f/uaH
NMQHv9+Pf5gFlVHkgVaiSTBtXiH37PebiNaABDZmn12p2/jo+sAinA7SEHAiZ7ZjEQiSqQ6w14fP
s//2kiS32anSbA6VAWXMd53onXU143P85SNB3snq64QHMHwfTXdYL8D3cX5aK0n6hM8eFUPIPFyJ
LWxvsWFoh4nN1roQia311V/qB7ir4sSoQWK+IoEu1BRUq0IPuyjNN7ZVs385Wi73ZJW3iOCriWew
BvTaANWaLP9MmJ9/UgGEP7PWIfj1KK12rt4GuPWm1eRmt1z1YZnqOGKpEOihp8SjEl6QHOTH+7fx
nQ0hzqk5PiLWC7TVkzUOxd42fRIuO9/v+OWIZrkXQnRAW8YP1U0BZ4PnVrGgwqYj1tIoiD00l+Fh
+6BrKuQAva4u8ljzryZGBMjPQEEQI2u4m8MOsUWGMlWah06E4+tvQTfqmTSYJGAYVNRfodJ+TXwO
teKsyKWeirUT1Kg2dqge06LVeLOARsSEYzoF+PEIz6FtmXYFhHhlE5pK0lGXqBeHWnTWweiXmZcR
sMM/g1bY1XXy5JW1USOpL4vd5DOdwJpzSXRSPEBiACgWEJAEtuHA2ZaNNhBaDvfTguisbeoL0nmm
QIWKC3jEiyW+B7b1i4EXXLyc6FJSnKk5aggjzUfg5GtKZpbss+Yqk9Gf1tbxr/XakkO6FTQLaKFf
leGwFjpjJ0uEgvsbJfHvQRr2aadbppR5rINQvbXa+8KnZPQPbOl0moJzNo/4RgEqSOLRZ6QW2+I9
kzk85/gqNDLkKKBrcn1FaZvVZ+5qOE0NAwmL6P2vFHFz1D7wBctmSbXXdWmXxZyzqr7zZryliXvH
yFveJg8F60LCsMOEfM7ap1gZ4hpbVUbUpaNtO1G7hpkKT/7ugubJsAyfhQwzCLI1+IKJSegh7hIx
+W6qUurqN7CMaGKi0jU93FQbzGBBZhv8O3rOtVAwDfol/I16cFNX4T20PtQ531CiW3oeZDF1q9lW
hXJAfGRyN6jIDiatJsdvH3Z7xlCF4sjiMv9T3KC+3bmumdet4eP/5ZC2GjfyZVd0XTa2kr6FVhtN
C6yveUOV+uCPxCoSYoeanJf2lBE96DQjIzKRKFt+lZpUDlG2nKKzJ14VxeuILaEO+mLBIyj1+LIe
1Tobtbs5LwWu5QKDGok48pEYZ2MZIfP/U/V5tdqUFFC1MPq+wFkL3OfGP7NBOSfl695S8c8F/+iN
fS4v6hzHlLiMFc3Sk4kd7+0bXs2zqzOokLfnu5wxkwsPQOklo14S6mvfUxtWnb66CAPF9UlcK2im
LiedHb945JA00ADTTE4yZ/ZN+yqyVaRva8hqBwY6kkAT8jSsYGqax2fpYA4oFGUnLQeoZoZ0A8uH
h5kpoQ05cajNnIjBEeTOKwNrPUpYaRyvxU/H0ZHv0WLXdaQOMeuHmWGdsUMn9XlEeku5AS1YrcPL
j7b8lu2NwR8ShTKeHArbHhx1uyBpR1zh3Akv92fCJdfhGEj943atTR9gPWciFYNKI2yBgRW4ZcGL
/km+fVE5NmCKqojuRLQUsQJ/oYNsvMePHby/hKEXLSUhVakwEvU9I0ssJRwukhnPKI+RYiElKpcs
rKrHmGxhBkNOJeymocPKPCrbYsKggbVLbitjsKxDTjL+m7Pp2bQQUw60BxVSzbUztw9bNekH+i9k
459dxZqk2HLoZCpTAFLQCTnMdQ+EJowuiDBjmW6j5TOmnoHpj+7Kz76zcVuWeDEv3jnYVR3mWu14
km/Dr2zI6V0tFrGXYkS4SPqsKdfyLfbJvcjWO5J3gw0ihbRurHsHUqHkGTYSBbLD4/wKP2RZzurs
SEFJKoEsp2Ee6Dxtw58XtcXm5wemGRiLQf8GdG5HpO44w4ulEUbXqMKqTQCDN4+N1m2Xz+Fcm6vf
6tpXDTB/m2C60pKHrdOVnWr2F2n/ozfgKpYo3+VGegg5u+glrf+e6hAV2DXTFHTyRPWhAv6NQ/rV
fcd+JiXeZagBzAaZ6a5KguWSTLgzK88htDRQzh1tQ6GauKarXQDBV2yiKkkWgdvFq/pbRG3A2E8B
zBV0xc3tnnP7y85piGW+5xd7/vKQIZTRAQ/gWtwMZiSRPwQSMJ+QI8G53im06BRGTBCcEx3arjws
UG4gj5k/SsL2J2ihfZIuL0nPuD4AU3vVnmNqVvQ2IRKmKiwp0v8+7sBpT6fnFM0OU+pkjBH6JLOB
0E7isEMnVwHjlbQ9TV/bH8OHOwwirGB28UNb+MAv9Oz8I2ZWxEBFkUCTPAtdwnfAfVK3n/+O16IY
eSaKKkX7NEO69ysJuAQI1Y1xtsdWECowecIutUcTe+yy/VEXVOa8mwFBDimzhtmiwmLbgmpchT8r
emO1dGqZId6N9wlCOe6NaTUx1sH7KJToag+N7aoVPrn0hnfleM+O1frAGwheYCFtWJEuXsefp4Oy
JgkpFlTlQwNBHu+2JSf7W+5B4Wsntw4iaMK+DUFH18Ik6QsN23LziQSz8bf1nq2XXF0stMlmF9KR
ivTzygCz2oMMa0RwUJTc2Q96UMb93htdkRQLxWWD05yllTHIef6+lWJdYSP/Fmn/zhvtV4BSOEYM
ZRkQYJG2mM5HNo1OWCO19XfxqIHRfrY/yvaiQV1P0MPkh3E22o+axbEY0a73X49nTS27UdSC2oEa
dfgXlGz4tEEQOgv1LE2WCSpWdE06nFrPVY/8XBs/pS4SXDergdooQJcAO6D5ZUs8rWaUG6UIH1rw
AXhUBetA5JW7+EMeNUdbZiyVRPqZcXaFOJ0iLhS0mo1r/e+/ZlQGKrlR9f67hLOurGrHRyperi2L
A728ngMX5gS54mzBp9/pJKe8lPsrBe6lTLsvpTjbLLPfT2hK5x83+1HCg9WTizUeU97h9k0Avaai
x9pQBMpC5PyOqDFZnVNqPxShgpFGuF6H+Ukrwu3B8uiWN7ineN8HuWgBnOcJApUV4ZkrsXBnAZdV
kqiLb13dP5n8DHrjEJX/rZYEpjr/1IRHcCzTiumNOH0D3BjKh5N3f6Rzq2moWRQIvj5KkBLdEAlh
/+9cDIvPHuRXbHcLCikljMK7RB+wcpwGqvjL5jDYgRE4GNOaiCBVk+BdO34bJUhPWNwIy7ls/+n3
CEZaO5wQqhstxSbWi9jpsPXE+D4hWKYIcvLvIp3g/Su7SKJfl28prgsrxEuz5gV5zTt5qCOVUBz6
Rl2OxB5Jwt+UbP60R7Vke9INpegXXruGZt5B5RGOKD/ZbmBrJ08DMmHfq24k51m0hO01EWCfhhps
DGDpfGNfNdK5gI84R5IJT+vdYu5ymC+OW01Ae6SYCWY1om1W1ykeGAzd/+oxMscr4xa9lhKy8bz1
ZMT2b9TZF8rH6xWM89TAeHflIMtzOq4PiWXvESl/RgevSlD7TBpDpEAyoELg3ZjO1BrmCKcax6YM
sB/Lg2YmPlkIuWNVRs5mavLGFxhDSiADeYY9RpLvbgsdBEd5gjFmF53WDF7DGv3q9aKpIRZZynh4
KQChGWcl7B1Uv1lMfz/Knb/U0SRqypwje9MfVzzK5PCkRhAAGJDXBVd9s8b9Y5H7RYD+WroAGwDF
9jve2FmXh2EKsMT+tyOa3fRi9m3NHkpQCnFhCW/BWknUoP2uXGcVqCv5A4FxRQCpwOYo5TPejXuK
tHozW3MiWt8QmgVNyPDKFB1n/C/mV2cE878JGcmV498V6xfJYcPCQXugEt8u/prFExxcmgfmkUCY
YjNhsmr7+DJpa7Z4NlGDARfgcTslrh1+fgI1Zc4hWwkLqIyr5pDGhN7gUWLhrrb4wHQjqjcH3c3c
Yw2lG0S4iKM55MXCH92rLUOp9LdehhPvZP2bgT5uyYr9iwR5egqA0euSx0k6d4lsM2y5RsMbZdsU
NaRVm1Ukzrn5/TCSXMKGINxZqtunWvNbIPEHPFAsRHrMgPWfaHBybQ4U6L1zrY+HwH7noQhTRiZw
GFHmeKnK/KalU6PyInB/vrGsJ++EZkaQUpBVhOoyPBzBvQ4Lgv3aGlsvS4JoBQC5fHoG0hj4gxR9
juLnjA/TUXnXuA2Nd7ucSF94rCq3UGWH5VLjfyyAZpQlJY8eEOnS3wZ0Kpxl5Ubp4Tg4LiGWHgYS
Rxv3KrGKxMpwzQs+KqrqommKVmlIAN7gV2JO2wmS2CtKlCV7ItUqPIrJ1Szfh1K2QZUS+6DafysJ
XhHXqOHxTVbn7hkZfyWhsLdRigWSit7YPhFkwfbqZpMFXPx0pySlx2ThtWJbqeBQyIQ7/Ay9Fn5X
1LeXV/uffNcIC3xmQ1lbVow6TuYoQE300n6abdOf6EOmfQf0skuTsT46Z+up1PosqlCMbsSffiUd
AziMrB+nFGhlUwdmteiDfJa0+65e7HRRyXvCMxUcFBaQA/63OIQiqeP2Dq3rrP3R9bO02ywG61v7
6UvIcWlLMCXlbM0bkqJSsqpHsfiadez/Y8IMdZFb105i27/4gMviWx7s33Y2evKrfzH0KwpHXhl6
3MtLM9qvn5NuaLiw0JWQaawVB7vNgUb0/Ace0bnpsSQ3Ri9vhQ64uC9cqbgla/oa8VUu589100Ky
wgoCuIQ+fGF08gSPnnv2vn5uAKVA3Pf6UtpFy+tEmLzhklKYvWycof1m6+S0FPw006ftjuVsQhtr
GsmjWUbxIwJG2fOvCFRBnPacAhhI2ow/nWNZU8ky7A2j2JuabC9h+RmauAkwYuQivNiYCZrVQIVb
kJB3kcjf2fGEW4Nezh5oIQoWuoNeouMy+5lncJ7op915dut7gjyV8Psr0v10H2bcDRZcC+JjB7ba
aM+xjahHyngwxuLGH1qWm0RY9nDUz2/caPboS2BSzYx5uDUSiUb96mbS4n0IHLGTTqYjLeBGqwFb
IOinQgqYvP7VEPEwetGFyhQMPtPKr4F9uz3FzU4LKoZlcR9nqJdLWsOZAV+mnFniw71g2R1JsTux
xnndzLSGoWq5iLcfjtKVEBJVkJsGqP5isv6BaWiN1Xv9MCV5jHMA1kl1JeotTyZtlfXxo+5p9Rz/
ty9WIhg4X1waFzmr3f4OtDUjph7li2L8GoVyyMybZe282D49HTLq8f0i2UZeHtGHK4Qywr8byFjJ
SP4pr798nyCwMODFzQ2noSHKPWN/qP4NxOipsXDQhtrLTgatf7MkBZA0iqVIyXjfFehSu6sGLC9r
PoR9X1+BetHgPz3ycaJH4SUqLNtAXDRVw02MUeXp4Ipz+GwIyll/6WlD1X69GYf0D0dPElQerCoa
Mw0sab5uup281RjIMwjqlIK272lIDCP8whAIWw66iF1oZBud2X+nTD7r3rocWjBcSjujDE+OOqWj
x6zaHf1Qu2F90HuQ7zWNYHKim7nkD22nw04mmVfoZCuxx0hFuM/UiVikfb27XDIpN2DBKIkzBk4o
lnSPhX+222hPF40JjURHWHpNjVuSeMH8TtN4NDRIUcVSsmYD1z950rQtFUEgBsdTYdvDcGc/ozbA
mLI3PYK09Mskm72rY7yU5XghEFeySehRwqN1xD7trB44oW8qAzQIw/cC0FqoIl6BLIns5mGYUw8y
W3vNauitDxuupSCGeDEJs6u/D/zzpNACAScr0ySptyxNe19cB0yzoYjB7mMOZDW1azvrOOshgM65
ZG2Fk2i6dwgJRwNJGQ+p8ycvb4ZjNP+YyjQ/RzvBk4CUD0Cw9WVK/M0G/tdtsuJ10PIxJS6c3YUW
EmZTl+EOu+HZdwl4wVJacCRpbrrCutM7rWzu0sNCn+u0598rGrkrO37naANa02aDlubfxJSVvm+D
Uqw50RKsCT0tszONnMNZOTSAUcGFtWA5PXPK1h6nh2ApXGGjThUFbP0yLhQxnFwhBI4E00FyWuDE
EkwJq6disQdYZVeED7StmjzyCBeZVj7Jdj8GH7P9xFqOP4yF0DoAEF1MXHnpnVKnK3QMdSOm0UYm
9Xq5cu10C+PYCXvyvnGd7KTLqD9GbEVJRojRep/9c8VXveMdNyH6Yn02TtayxVv9jE14Ywmz/tDQ
YHSnXVi6jpezAEJ+Jd9fu0KDyFFTgZT43UaZmOQOBLjvz1tCAGgsGwbLjnkNG3Sd5rZT0AW+W3Nh
4RjOSr3VX5tmOYJzuL/rbh2WAGm2Dqyh8D+NtJnkSJ7rNPL6qwr6nk/iLzocw7AdF/X9fKKtkKmy
Fx84jsOxPT+GVgbsyYb7QNiVg4nLQnPk4gBjdkduNfddZtBzCxG1bayWioSsZ83pQ719Cq3yNkhW
fvgUHAOkklQJyv5wpuCNt3dVlKpAa9J2KUqdYcsCYNSQj7yJ1omJBPSDhsozOho8+OkWYZAc6zsH
XoXv9AbNQEMYKeDpOGtu3pNOLQCiu3V4GROnxIHmQniTZXaNYwpuh+qsd0rFXUH2XWG0rEg/0EVv
gu1RxskI1IFzGtp6E4ylxR4zV/YokRXsTa62Hd8fgqdW7fQhs636eJiYGCRLFdu/WxBcDbJ0qU7m
Q2KTKrMPgYvQJ/YBBGiJTtsoArTOD6uBzKMwz8TqplAOqRB6rcEQhrjJ87LLNMVFFRjMFHZDmr+j
xUlSmyeYx08EcW4OQweDFZ2zitRsEdyG79C9g95132C/fUmUYjK1oeFtRMO4WdU//HgmSZS7E+f4
1cgLSqdWYRt3AZ0V23myqoGPg2+GWRb23xFm8W/sNc8acezVpbW22IxiXbYGLToLT0AxfF1Q032O
/3TZByMJS9m31yfOWc7ORmhCqFeiBcyEUMIN6j36an7V/DvwvvlGdAfKtJfm9kGnhNoORXWiXny2
RoHxeI8L3EPyksH3y3uiUxE/ta1r8ORzU/+DyVwQJB1E3GX8UAb7np1dp4GRRQgtfIhrRHJJl0eT
kg2cWmzRLTJGmCF6c13Gx0mNSXA1KVfhpBi8VBGfq/k/bl8iVmw5tUBKjkZ97CyN3ZQhaS25KPbi
WYmU8aoG4k0arP4xy7v0MegQyFz/JY+PZTF1sU7+cJPZm8v5K98eq0IE+Dv0OXiSQ+3I5FmLcfBN
cilphrsMm6nU978FG6sDlVKvkZxK33U8lsJgayevnn4yOLD9oKrE2jBB0AVmJ7ncWOyWI1e0h2Ty
L+EBmqCMvp69HsP5vQiBC2+BrNvOxB7n880+fdFJCewJiy9WU5a9BDZy8yQsmbsZHw8/BrvkNywf
m+QsxbLtGLPBLtLCFfZ6BX83TS4wHvnNs1TOQX86R0IK8nXQX0paQtJ9Dt1LbexpG71dx5h4wHQU
j2xlvmHtFGbkPKZmncKTNOs5kJ6bM6MPx/DCvg9Fwr/MVu6zER/3EOWIZ/L25DpDE2dY6nUlhG57
Zl5KdFITppl7a4mkw6yElvzL+cnOoRqq1PAPUugfC4RJNiLbEMRGe8m2+KRll+OgSYe9Z/hSWCEB
9NyIXAoNoStt7Z171LNLZAmO88U9vz5Sgg8svhUMxhTZY/OVmVaiCVLVUMXRpzck0AJAt1m6JYE/
gNv/DKyXVcInXyDpdSJKGbkXKyLT392c+vGNt+oNM7ObIs4O4p1pNON29Pp7gIvkAPa8b+xrH1mM
lagY3gZ3zTg95FnYyyH3BQu0y2cDwWozcJInSuA4h1c52HRGJU6uN4r+DMyLVdkGrPFQhjpXTHf3
KZTP67PWYWUruGvP4ddB7sWfLS9ZqUqbrRwJRSHAVYNsr7rQp5WVYNRtGmJl57JZTfVIqgYGtMVd
9iyMp9BkDqeU05bhE5fRNOggmsR22gom0v/CT+KzOSdDPwj9IXZRvy3o7ShBkrtYmhmdlRwy4zDL
A/FTJcxUzXPnP9SfrNnaFoTgunpON7Zq8ZheuilwD4C/oENi5szLQ4spOYsw1lkAnuDkeuXIJiYq
/ewQVzX3S+mq2pKcz9qrb2Jm7Lg4GQotcQVtLkzwBdHby58kwQycAwHfEBZe8VJDtd5WWDnjAN9k
9nxhcHJeZewLgAHhId8dw6Z2agkpTFNeHqgzRFIzSjurvrCgPns9qEKLYoYSOfAsu2DWxY+/TRXJ
U/8rdTDRPGH0inG3IPwybMBZegBlLnoafDCQZxFiCI0fZR0aEPDj4wUvyNh96XGgKhWkPn2V+LTc
+P8E2NcEhJlx0ho6/+5DObOxll6vZ4gyRkT+M9fZrDuVMUNJDl7yewTZP3a/RuezBhydKpM3Oo4y
qRVzIFhF1t69zhRr+iMyw0hDkHMtM7i7/L9vPVoBNK4MY+RqJlXgvibCC95A2GIrE4VTHT3Zs6fR
PEBRYPbOQZc8PxDRhJHJSKOzhE8A689x1WXnEACaaRTSk6ERhrOS9tsW6FVf+4cTpPVd5cWgqLUl
et9LtOmMyozo6//ugbu+5OkswOKuSqe8tnsOVuXjjbk8KmdxryobhtF1CoyZqFF0JId0l42KP260
3DQPX54nXrA7PEZsosO5XwmeYbF4SWJrBEzFee7ZvQLazqEWDn0lpI0Z9LliC9963nfugMjFwMY4
5nZ2ZC/gv0Xe2vumgkgo9IZDv5FjZ4zWs/68KKtf6zyccwjZRiC9huDPB0ssUJXZHux9JrTwdouK
8zkU/0u5LerNmhEPHR+u+ZXppHurh4/rlCQH5bWLNoRtQlsMyas/e0h8T4kJCVjCoCqcAa61W4kB
ZJmXqvpCOBxXckSnbM0oIqodOlfmb1zQ4q8poxOZ2CmNZgcxhg6cfWrOWHk8CKXMyHc4ATwIS3zF
Ho/qbA4eFcf5fMSIsTi704S8S1iSodORn9zYqc8B/9txG1+2OCghEVy0/arT2sqg+HCKrAlS/lrk
hzV1zDRzILJF0vw19yBeXhJSZQleg3x1qAipX7dNIETHkE+gPknhWdAQ9wfTUVwU4Krrghu7/QZS
XZHTdmNNe+syJAIngLoDBF8vvSxmDje5kn/IxnczpTfxxu/wZlwlfH69q1/53WAmCMBuwo35SsG3
EGWZFTJYmNDO5pnTMEzuZSQZF3riwttfRnke7wcyjg5tnWdem4A1RbrTreG06Qk8s4tK1HwBO2rA
VKrqvUFRNZQzBYh1JahdItavMGvrw/EBA86ujyrlWI5DYK05oAjf7H/y/7NTKVLgNyAaFpZDVYeW
QrZy6VJ/FDjraV/QgtC1CX7Jgm5ENko7McGxlF4y+0yqHZJ0qZ9A4ERGoMfyeKkILzZr5dc3ON8C
GgBja2wfu7b+EQJclVeaedLLbSPX8Q6LofJzuhz6MAHK3sNUz/rcn/UYK9Gc4kphIgqzae/5Yb8u
7ESKv2FiX2ckYCJoPyfTJZAtb42oSjpgddc4sKqik5386+A2NOpFsFDGdl80LgfBgxeGK+VWG4hB
m1UUmHHhZQy00J6bbxLomSgkFuQE03SDIY/So3JL9msfPKIxrJ7NC9V+elwoOuBafw4koIrmEVRw
kHqSdjw1yE6qo2DrYzscBRqtevv6tvJcRHBU1rcUMi8wK88/5fXtKUt/hixB2R7EGq+P/ymwSBm3
oCLKmo4XXWuzkbbpXOBqOAOy4I1TA9sBZ2gaylYCIiWgFcy2a8IZz1SELYQyoCZkuKka8HLou6oT
naC0NdMDMk6pe0E5PurUhGJC15ZxBN+TeRUr9dEfkiCAuCMo+BYioIisnVNSoCOYkPAXrvyefeiu
z1KGLvHDoWXRhTlK+lXP7DSE8GtXwFvGbKlR4fZO60dON3KzmlW03YyAnYn5LEKSrC1s5Kf+lQ2s
gcCxifrch+OcJs5Sp05T5Mdp4xfc9D03fl/3eTEyAOX42uk3Wv5YTJ7rpV6LYTUb/Smyq9aakzp+
Z6hNU32HDpkSOQ1BXXmGPfrNIdQIA+/BnItZZrGCxDKHiMToUHjO/CdCW/PZ+v2DY/ODnoNDasOL
zZaMbtCNruXX/LTX/u+EFZBHgUib0+Smr3ehVaxdaYqrjFT+N5aOYTsaDtiYzq79nZo8+qROfCaX
M9oo9UEMBsWwSPWaoqA/wD+KuCt3PZ5xpJTQSjqeLp3qsYA/AAQuw95FNzfuKdSRvJnkluEXwMP9
gkP0ZF7IgrTvWDHlOqwN/zkuP9gR2x/ZClDrZlSBxNMc+sJsLr0BFcUCT1j0wQ6w94euphlXu5R7
rLHECj9LOcP0sZ1u2ONe+4LeQBtN0p+HFosP+ft+8pQF8RKWz8Joq0t2xOVGBUTqPvP0gONDRFj9
D9QgDJuS+GiJRmXc+xtF/phG+ZVQp5BmuWoEzCiSSIebCNHrWaMddtsY/zWVZbdvGtOKktg8BuOr
WHrwDcf+NYfjPLrkZtYn4KcStnwV3/myxh2bk17hDU9YlRJ792arocV92ntVJrpoDC3zOQhOA7dN
r+hMrNVwNqS8GHtzszbLAUkf8D2NWb+dA7heEdvlFZVAj0yV6sEyU1mcBlby1qV357LzWebLW/+7
S24HyzB4aDBz5C5Sq+4lboeNK4OAGl6Q+UWe2m1YewdHBuw2Z+3KB61YESd6EjhFdLV8oDjuUxkP
/3qD5VrqFx4ANJnhzRp+KYigXgh+RrRg4OopO1+A5+1Bej/erlGueN9pdXyDiJWrNCsi8PGB75Hu
1BKWMovOxAmnt3Z9uKvWsnhkfUT2AZ19regSuG1vnNGBYT5VIeY1aIoO3FcwCdEHceWlQ4EsXNYk
haIZ74mXdSQXrMAN8wuNNe+d7V2RmATJ19C6/6VECyLwrO165+HXDnfwOaPcsw19kgrKeppf0u1/
RCjJjkXts/V42cOYs3eFno+5zVQkgvHDiLi00Qd7VMLj/rWpgch3Wes4oE5WjENC2t6+tTsUqbzd
v4a9cZzZtzxHfXoarTBh4P/IOIziRVgsQzdfi7cj78EF5QGt9r/F/luzPIGFZK2efgTPFVmCpZNr
LAvI/FTWsUx1tgfIEqD031uEr1Wis246uWljMXM6kipBhkhs2QWnxNy3i+ox0EjkcIXnJ/orxW2t
+rxbQCJHVJzmSckPPRf5vdBiy0zfDesGLI/MWjz1CeRruH8PUsTdUFghYKKLFtOR11KZCW/Cowmo
bLsPATXGNZrIMC1a4FvLSMlavVvh8v4sk0q3wDw4ogYWU6VkeJOr4Ydx10vGRRRH5F5LiMIiCUY2
pN8fp4u0OA5pKqycleVjzPEQcHCtC+hCpemZ8VdOmPmUoqcL4NlI9pEu1G0MIZOyy8EYG2YYX3c5
F93a0sw1S7/pYpsUzprGKeN64HIAGcB80h2KX6zpjHjPv3WvlWwyMLFObtSPhrKtLYZkUAfXzvLF
WeL7SuwbBybG/RmEA8ap7ky9o/pE+nAmDwYUfHPdK04B03bkZ9PHgPi5c7x2RpyW64ueOfAUqSEE
IHZoEMIOnhi/t3/USK2iPmPyTIl+vpVMz0sS0G64DTAfiXjDvWbDK5RQnah9xLx9sc7ApEyVf6Yj
GGzRiMo57uIQ8uNEmANQKyZmftqPk6mc/k2hcY2ssf76MsNDyv+B6ykT3n0hGLX+VOuvuDG7GdcE
HsRepPAmyvUhuMA2PS0K224HcN27KAQ5NWjbaof0NSexjfGukNGOgRKLrNFnQ7rMJns9DspGk0J2
q7tCjM0pJeiLb/A6xY809isI+69WlVP+WgORt5gSsFxMEhViuKA3VfPUfAbhYfTMirhqt2FU4Mu5
7Bl04bNlz9BpxOjW5qsKTVmlqkdgaHwxfWwBPI24jN5ZNeCLTArLhiCG/Wrcr0LORmZMv21A7ECu
eFM1BX+3Tj/ebyP1g7NCPw7CqfU000/cJ28kwcAZ6GhOQs2WD14oUhx/wb88Hhx/rzSDVqhX828f
Cm/u2/+yWgQdpZkOIPUPXLHY1WGG/rnBhZM7H7XfiEvdIbfi7hK7/Wj7ka3C8XcgDNxHmU8yx30b
CbwEPUlPQXEpNIVI0yfdLySAg6RWzYGFfgbREy6qmm+NdDT6D0RtqOhePQSXSAB5hhiNxxacQOGq
eWqogmBr2171NTth4puuHr0TwRmVBxDcI6LX8biKId+95TknEoWrH3pEZ1SFqXSA9FKX/rO12vvZ
fe/9VHgC5+08R+3s71P9LZDJZeQjvzmd1hSGjUI2LwXOVmqT/pZm3zrKFUEpf7GM+jSaCh4C/tP9
Vhw8He+zQ2YG9PzMRUYpwwggaYP+42w/6GLksIqOk64KliBR4MZ7ezqLJDzxUpgKMsYA3JWxrshE
ckzqePYpHv8tUCKs29qnm6bxFRvCmqn77gX7BvjTpsO2nFWnsjHqjax+2/ToCQAuOJQon7PiWdff
hnasov2kjJY2bE7N8qjqtrn61yp6w/88/2LeVGP5azCV9E722TLaxg8qMP0XClYIXow4DZToQLk+
rQTNPqj880/95s8irt0CosSraTOH60rSFf0pxMmxRBZYGb0ZvLM0Lx8hFAsToUCULpbGXfSlvP9/
4xE9d+VayHtXnqvnK1bG49tNusAcXil2hNk9KSia72Ms3G77BDVQG485FraFbj1zEEi7OICxk7yG
wfVxUtK/pAppFBxbZv8oVKeqt7415QJ47hsoAqs0oKbpaEeGsFW5BRHnl8aEmCjvAUxtXUBHCiWf
FprlN9fcr0MM6n6NQgLJoSvULaCbb/rsiLu7qW5xXCmNYvngcd7oJoq2Cg5xeNuFg3DwFQZKKq3x
wYYPvaG7QPXpIGJhFnvaIUya1cLgBeFbQIv2li2kLoinB9gZpP4782w8/NcPH0skreV4ZgSMHW3M
8ta1MIImVqCgXaw0jpbaftLkonstYXUMjDPjonmOOuRXLiyvFM5LlJwaApOfR4N4EMpprYUZCyy4
kG8VYQE1xXRfMXOB2Ec/aNP3mrI55aKbmwMwi14eHKh/lM1ZsDD0/RreOz9y9oBBWRKBXJXwLk76
X/H1ooTrqvUQm/leJ8itu5frgacXCgLD/QxZM2Jvw24q+cgw4uZAZtfr9ZNWLfQ7H6ag9iARuqTU
2CQrxHlC/ZfgH4BZ7RYM9yb6GTySDEwP/YIRTRHPNvh4mkp1aB4LlUUJZ0pnycIGQqVks5AB9Li5
/1OmHIPddo16sNpamPb9+gNK3fCUz3fmBnRl/oHiTV4ulU+K5XCA99iYxbrRps2FABYAE8eZ0VE9
a3/gP3GG7qmWB46HGYeKPL6DEID8nWKwF3n37pfPTiSJPZMuCbKXr0HhHwL5YhUbTmUtZHel2mG2
yX25diLZq5leeJgJcGM8qEn/DIDQ1+HVlkxH8y/swPNSc2YqUNpi5K6jk80Ye93ChMyPM/VugAH1
23EyAkZE+bJfh9rnY+K6Eh6V5UDY/Knhk8shA0a7SW/DSPbfbF86w+wJokSDriE07K7J8K/Gr29I
VlL8snyUIXWq5h+HtGT68WcMVS9VV2SSC6/sgXzvzX0yhMpycQx5Cinfn+uIty10L1fU3LE37TIe
eX1GGA7D7ueL/uemoqvWaIgefnD9Ba3S/XeBesVGtwVDAcFxl98YZ5ueMVJWa9Jc6qqCuRDfcKrM
NI9YLC1HYB6WnNKSgE4/XmAxQ0Md+6h34/duBNwn008y8XB7WDmiyR5Q2WsHfgCOdPvFXxmi420M
Dxmv9OKGdZ2F9Beyod8qjwlM6caGsZgifIIqgZsSa8VwA5ZFIIRoBArJGdCG71Pg9GogrIoI1gjy
QIpm4DI/kP/H6PYNLt7ulAO55WeClgXD658RAp6qdNZdj4fQv8jWKZqgUDm0n6W40mbp9VRwnI8N
PC9mSa4snO1/aAJUjjWZUeLnTmHpvDH+I8M4qlG8zQlNJHO4lDKJdsG5W7RC5fRSi4bKHivXQb/y
9FDmcwc9EnN3x9qq/0p819NyzAavwt7oEo7OuTkkV//YVr8R7dRL4YHu90F2f0ksL64pCXZqfCM/
hbTjW/kCISIldjXY9mBNqSzi3IIUb8ZqzHtgJv85t4BqRCfgRxZbQwXyZS1d3pP5xrlKjAqP0FH4
88OT5xSOHYg8DleUVdd5M1nUy36ZNVkLtTsbhsLSEp58WPO59pY6otEF7qW4PN7Vx7UqT6BWvasn
FpW/95G1PjHXT65Xzj/AE0nCOYwGwQggqO4MSqDSNchNVRJZ5vRcDseApZFp+m9czicB1MwqxonE
L/8u7TodRlArpyxX2m7yn/gc7ffWGif8cliTInDV10aKXPVwc3Qzxe1GCBBL6DdAiF0KhQzhbpl1
+mpngdjnBK5/YYktK1WrqgwfndnpbrgesfvFKtQVZFKSKRPRh1UdN9sQr0eVEDbmhrpJf4DpNcKQ
d75jVQwwa0KddWpLH8uX5dlpxO3HUkALyyNsh+xju8njvFNxtBAHe4TqXGwg7D3kC+lry2nSPrWw
hU5fDV1G5QFJMYxBpcS97Jzqrpykkn2otkjLZ5p+iyxwoPfHHxQYffy6J6headNyWm0sC9M0WMyu
xNTgk9rpvtIWRcNb1sFvzYJvo8BLgwpebPUxbTjr56uficGmTCpOyoUri9wC7DTW73idNXWmO9hd
ZdlP0xmzX+p5kMPQbFbJbZX3xbfLWljX+NNwuXdcgKhuVsnY8eAnFx1oncOnOMyuL0V8q4EmRdBL
7CRz+IBtjwWR89u8SyCCpilhJBNI48V0XUlRu1gUWnssJDDCz7zfS9DA69dwbbDu6CTz9VX2TSWa
n7UkHEReoxxghx7Yv0qfPf9m+0NA4234qHN+9mEJ0+BZAFoDtoFrFXLPqZzjFM8L6JlQx8FXjD5z
sJb1cnBvT8n9cD8rJIGXRqINoX5Ik0mWj+CuoBiiDB4hRmfZ6/WAopfsE3VphwwR9U5QI0qHNqxe
zvZP0H6bvwHxm0J31KzXj+b+nOVc1LLxShvGxY0N4pcr8oRx6xFNt6oh3lSHzB7fbgN9QduwRJsJ
MP6k5Bh8hbo+5IlPfKIISkjnoY6tNCBnq/lMPFKeuZWjNJubmshN9EK58gkRsLSIXSTg6E62s4DT
kXbMxuz9yL0HWhnsy4ocrZ1IGdIEucXKtdIqmaiDgZPaOsf6iWqyMzO8fXC7UXgS1K9lR0HujbXS
1+HdrXbPiBrM+Zq9GMaiVQvDQyjYSESUat3zPIPfxYIEueNpeDq/qhvpeS3tl5u2OuxgNnzfqMUI
JDdFNW6w+CfMXthQve10TjxxAY4RtLR3/KMV7EK5vVvduy/EhMrffuM1fCCgwjDf2XdK3mzYnJJ6
Z/3yNQZ8+eGEx8BswFkER1vBawniHtLTqIKI43pVoOD1Rut1lvCXe16nasFzrM9zG7XM/K2O7YzI
AnL/0zUkahOzeUO+AE/DkpZoRoFRkDoaAeTty+RETPHPVTFmPr7rD27seZT8EOSdIk1oGRXYSKVZ
khdvu5tZ70OSP0bpopf+cAtBipQ5L+q20MEYQY5zuqI170rNUu3vqkWBXN+zet+vxqLytsPeI+vE
CGujAbyK6zS7gK2preSgkqZe7PVg0ls+uzqJFZKXj417cB8lfc2M9QVvkyn7r00vMAXjg1ACkht5
8hTX2e4fbjIc/kFIPMMtDe3ssPPwYmRroYTQehtRsshlVA+DdgyruKkg6OyYB8T0+FxgfGvcHbxh
FjbxWxrBsPc1zoCZl4Vd5nqNsWnWjtQ3xfNxCdHIFABeiK88kEDN/EFsDR05C5IM9vtcwuri+D4e
XViEyED6Sna7H9/HnvrMhnbSOqQwmYLL7foOLfcSwTD4maGLjUNST5NUUz2hdx0ivfth2Kyx7DOY
kbuL3UZP/bMpaOCnFOQOUfszMhImSxZB7C0LPp5sSVoarxSyM+DM4TOGjrhXYz/1C6uUR5sV+hB2
hhDvMwhzdJshxGLf3i/HYGZbkQ7u1FSujFB3GYRdwjOZ5h0/ztFLxvKNAqlYtCBfzyU2eMLl5Bl1
MsSKERWY4Wa39/1oSUP22pi6Ninaggy8RQqdMFde3JA4wKZav5ENY8JlQjt82RnmDGnsDPXp0yHk
7F0rQKkmXreZwdx+Cd/RnAQQMYdxbYpI4qzZ+mAO77bPBv978dOcBdTpQnfJaC7Awa+pBGLGx7xT
vPBYa8CRSKxAnhBNSkGKK5G5/EHbnvIvEl8wJyt8DrA9QKbbxV/r/LekegzAMi25H7bnQ/oDfOk6
O7/tznpPaYRHc0mIxE44AYIGXmNEAhvawe0ldBV7yN7thlCyX0yuJeuJ4GrRSI739TUfthsfygTt
jta6Oz+7ACY/HwgkLsLP0p7cH7xbBg1F8461fhkzMbDHuMgI5078JXuMQaRLS87Blm8orU7aHFi2
qusk2mS8VYrf88fc4nXW0bb+Rv3XgI4q7O8jnMXTa2++e6ovghgk6irTAgvC5ft/HZfbTRVfA9wV
7aEefwO1FQvxTQW6wVUyCqYF4WWLAP6GEW3nHUnj6ar0ZyeLzuEt50nrdATn8Q0J37u375cEw6ld
lIsDhP9rFLk4xDsFJgJ1/VGToVYBj8JJXsgc8XZFqg3PuLDX2eQFNQFxkD5Urg7mFzYdOZvZyQDy
tJ3E1s+GQrz9GVwFnQOEMLTT/WFhO6pOl/08sTqPNmbQk9Ubcpk5duIZ8nqPzOv1YIrX1uNr2fVf
N7EdPR0GrvReMhvtiiNS7SLWnrd5x2PYmGFQjIsZi5aEJcXzs2DLoZdIKaEZbz52HaCCGJM6pNNq
RPeAfNx3+V8rL4Wmx9G4DKyXgw3vYniCB5jyRTwUKohUdmilMyMb8205fheQFWs8GTJ1qUD0bRms
e+lW0Cg/Woda9VPmfqSGPZDNiCmFJ9dBqfRcIewoPRBNuzPay7fThKMIWPF6rXkNrzYstEgN3rFd
OWzBQl6u9Yg/3EwCwUmnbJB1dSA0fsD/WK23t09/qCf+RhCKAezcJ0RhEKHBjHx8BpbYQRxR6mAN
TfMfi7V1YcVRCNzvZiU1ZHjlh+XWvM1nx1+7MkuNXA92g3zHu9k3fUXv7rP0i2qeAhebIaVnUa0Z
FMphIieT0oXI7CLrQd1AyG5vszbZWNPiwzi5HVoWGnTKebsiEIE3kdSR8buNoWmjjWBYC0wWEHIb
8Ff+8/xLypL8pJl7fJWwMBs14rJt1SJHY80yQc2JdI6FdiP9VXpMHym84tcZ/Nkn85ayWgLAIZ8H
m83vX7g/Qx1XPmbGjqTGmpmDtYabxZRRniC1iMfunpwZB5kNSq7AXXMKtKxdwbcWcMo27joGxDnU
DutxUrTp8sNCRxoXWz7RD+V61fkjnQiqHPCAfqRBOgc7w1rhsqtPxLCQXEGtR3Mus73mYaNflAsz
Bk/hHkr5+FnbZ2/zTwE5KoczuXp/F59VKBbSZsPDgpiJehcz6+kXiHVu1An86+IvfVa/TrfrAPYI
bBrCIC435yTYGYlS5mwUUd9n8YOlosg2tirRWiP3rVPwEaBd64DrNl7g53kwH7ZKM+Zr/LTONL6y
VdDOoL3kWl9y14yGz+MF+JhsjdgxXz0m/m/i7Ztv33djcwLUCZPhy3Mc4v9VgxSl96Nwaf1EkPJU
uDPL+XfD8mlFouslnlDcd+LR7pLs/hIYBgxPE1sK9a4JkSak0DztLdR+pgTuuE25Zi7l8tRr8hDO
pPKrC7NRuNiPZ53yhOHJufBJhWkSPo8yEIXdtPJfsL8mb6KjWHR1iKgtScwxpyAwuFxU7CShDdAq
FhuBNMpckstb4+ZVK9wYSG53HaTXXyauJIp3+Vna9UyD2Mbp4hizcG7hzWd04Rlwmk9xbCdsE/pz
Gsa3J8LH9UbSeMQSXTI/zyQlAqfxJk41ArK9u3Xg+KLQFd8RQl4oHtaIm/IBZwclK6eKC8zDoUbY
iPJ/M/NhH7XttZrFv7JxVd9wy3ZJZE8Uav0eWdBIZzLvxedMFlSzIRPTrvoVV6zdrD6BWSMUiBS2
c0HidLckQgYHTLXWLFr7LQdGdJYjcqSi9fIXgHrMFy2zI1+IWlVTnTuB5qfMeB2I8k8/tqj+pysz
KMzE3wRkPdBTzKfO2ez11Lwz7qGKYrwo+i2fugZZS4hyIqL434CiYDRwOZTixOLsDP+C3GscXzRX
ZvIMesRTpPcAWvtZ+k1V2FMMtO+vSPuITQMrmi9/Jd0LMJ4fai6deD/F+P9j+tnyzSeRbVC5Q5Jb
MIKzdW1rmM+MabYlvJCNQ7Zp3FWa5joc1sZ0T+Tvs8vxO8shVL+MvL4X3vgENYwQLr7Tx1cZTWJJ
7OCUFbAlO16UFVRW/xWS1riZOWo+EGS5K2YUnzRBDT0mLJDrHGPcbcrbBly0QKdb52xIwKmjfMCR
NjdzpCS82WpxG5t4+9UME8OKDcgc/JYZ5PV3m+enK2yGQ2G1QoiKMuY7NYY9TzKz07k7QPbA3M+0
0KefZveqPdOmMA5KgPxJfCNYhehHl9BiaJZKiO10brMBI7uHM5bgbXwyBBrb4hhyWMdR/V2x/lNj
XQnCeSfTOJ6sgmnltyYbuH++pTYsFj/Bj0nPZeoYRLy5EeRwZkNXRq8x+Hl6INrzPzLo8nfxQR6O
JFpkAghc2Y1lqOM8JOoPZAhgQ732c9qRjwgeQmKeM5xHW0hOVisg+hPKhi8FBkslG7bkStJ82stO
gH2Ct/678y/03QmRI7RahXB10F7wFCsYzPfZkyG7EXWjHqSOtd/f4gIkOi/BlVg42Nzaz5TSRkpc
yd/VVmC47wsqlV9AcguYXzzNFzkU33DkXnz0qFYfw4SFczJTFaMQ5C1YK/qk04haFuHhVPaJghKV
OG286UGWYH8JQm2MtkMT//ntZLBZYlBN+0AvVLVNSrdRUCvkiav85yVXsdw8PFv+63RyyeWPVoty
0meEv3ZTsqWsmY0TqIKD3Z3aUbxMi7XoWwhGpGgvTdkFFD0bs6LRWe6tAnYdp5gVo5rGxKUBDWmw
4C9rvmVAuVTy1F8W6vCtTCGYQi372JRApEaEDkHUzAbO90NC8B4pfekqJ+FAFqIiFLmenaXcXWRp
sz8bURS394XFLxADRvOHFqBugAJBfpOFt9ovSGJv9TcgAgY1Z+JIQvNV2iGYyUUlDKl5cIksWJTK
AKfhxFowLY5ViK1+PelDMI2WWron7vH3lStMPwuJLTTWa4f/7r6ls+D23/dqNAQw4f873AznvemA
xlvKw3Y172F61/sqYB23tfRIkeFHve4UePPZzTy64CThIVyi/qGeuL8VzQ8rK0jiSVSx5qyMCIni
S4y0+Rf7+YAhlads7eqoZthpG+njsZ3AKarRMyCzxTut8GUsLbmAc6lHdWPJVY+dPzVA/9vg9ppR
TK7SfbxEtRHJ2WjHRF1FQtmFeJ9/IEnu53htH4DfaLYWTRYZtl/bHUiF6eJIJw9c4IKgBoSN04+W
qNLywZ3gdI40JDOcXSprUqkbV54PVsZfADabWY3+tyOqdqf0SEy3pvGSUNWuIoqx38XPmfqBwFjJ
3ivzClgqjILQS/JRdZnIHGO7oy4K7QWkkhKm6puX5bDDdGpETEEUsBL0xLCFyrnqq57wHjk9R35c
ufVd33Q87NKGfzNoxts9WS6N4t5o+1V38cxaXZXLMdQwrn7bxYxwKR8MTgf/g30TYbk5iTBvaDTF
CG8Z61glKoUAh0+Z0Bcv6DL5SS5JTG8ptxg3ymr4l2AFzLEX99xaHq0blvHnuRye8HO6x1nOO+rI
ZpEqjtYApluxNSmMi92aWdDZPA6kF9oCczWB25riM7T3oRgx7QeytHfymAlTTRZM08qhUwo1CcKJ
r8XKKM+I4Lpl+No81Nw6lA09zGqRpMIO8TKUhpasV4LWpWsAFLvV/pKqBg/GGLluyKkyAFjEuZRG
9nN3yHfIthCmSEeoOLzGp1rs/ZopZKcyH4syoXRrQJB+CTBxUfhhNZ8aWGUVadK5FziD0rUGC2A/
rTsgt52We5Bsx24tLoCYbepK9BvqgfRDZ6R+Q5L/pMadNbWfMvdDoGRMMQYDX46R9WzWal5dMajf
czxDaxtzYeiD50ARjv2imp0WrDcoaawcZMCjJKPPQIpUfvILdOLSGSTSERFGQIB7J+fguPVLd4Qx
/1WB8xbwM2izWjO9rLId/Pjrzu4ilRg7dLSrwqVBohepLFT/QNVApaP3shf67WyaAU8+5jxOc0Oj
anl0TPD5ApyIA7qGu6FjIITdB/8c0XAKZUhISwYdwL450SitWuNBM5bVYxKdNtfPjMFsA0aYcPrE
L572YgjrHxdNamZpZNIK8KghcFlMjoHdJdtJVg+QqSu3hwtO6h/HRyu59TsFXacRh3vEpnBC9P/t
rOocApnfFdTWPXVPXs+cJfY7bB+jADglOaGpYlNPvIcmWPlMlUyDswZyDrcwF3CNtSCuyt30m3DD
bnKFOhm8WLabmi9CIsGb05jGr7KlyWM6D3j0BY8epIiTP1LW+HFMYsTgGx9CN4w4++ia1gddiBqP
c76+nQy7w+ugRTwiu95h0rEU+oH+JbaEeThcW2WVyMpi7b+BAcsU++uhV1M6/GcfnW5gy4Qdtly4
WbZIOkz8+YAMBFw9QxqzRAaCE9zA54hl6dp5tDAOfXlw4KKPsCgYGH1a4BKYSJ9khzu69T2FOmnk
7I75dOa9Av7aVMBjjs75JkQyGvEItcA6KZhQY0omXAwo9dt2FH+X97lMgDNNeoTkeKWeeUKSJrKX
mRhcLu3twpladlNknfytYb+c3lpKrVRKn4Xxeb+fRWiCRmS3svoqJJQ/gYkRWN4Rg2EtTZ8waKiX
pc+02QFT635Apz6dctKuddOR3U274Zi2CLLvPiWVPsgyupzwD46AC97b8N8BlS9lMloOApyx7hRf
ncOhRArUubHF5JCTA1IChj2EoGWS/7KXoxndi/HzOshRTnfaF2TPEm3G43XUMGTjFns+8CZG0+k3
sYKIN+pKMAbGphdTgaTIz8L+Ngg40dD6AF04dvpMvUfzf6DMq28spXtQf2LH042litRhfNs6MrTC
MC1yAaFRR1DYvMAWzCgCOEbBNUP093Vj73GHY7/lJF+RTOJN43MayuADAgaterdJJ8u08FAs0XQU
tT6RGLO83CJCbtiZzolI8yg0sTmTDfw81+L7+A22iL/Y7s6dVP95yFfzeCM3hW5lS3ybT6xGW7oV
FuTj++TMaOe8suVv9HJ8aq3KjvjV1CkAKmnS2LCIrqqVV0gtgkCCb2ZSdBHDx/oQzHYBVRQoRZCG
jwvBIaZO+VZBW3rAtrzSXkXXnD+83giC/Ih1kkwEP8RF3Pg8Vj6to/btyixCnUNvqcr3NG1W8E5f
sLxsESKOUsGoVysDpwwHsqexnrDMt5GZYCfXOlmkBiWFODryI6YafZ424ydmYeGJY0/OinaCDP2/
tjts50ybEEuwWVMaQqMKxjVOQufpu1+GaztkC0TUZMnKxVy+awqtidJXzU257kiedOUWY/UC+dND
dqOVOAIJf6hNuo9ayadg47dTMDEPmZuvTMZzYKM5l8WcBcFfHAlIgmzEEwwp87zVyaHtObgTa3Z2
65/HKJNdbs5PPCQdDQ3nYVu0PWbHaM3LwTqO763GiQyVyHkA7EHdoJUHYyiI/qEU6QA5PBtjqT2s
pRlGWcFJPZCZHP78MyC0FHPn3+4xCkz/wwrxQYUoQRmW2Ry7SYtkrHluWNx1F8jKNPBCBEEcgvWf
TveVKvRoXWFiSgrR9KNv8J8BdvyJ4WYsStmvJ5ljJIeYUSI4l9jDX5BZmtw4UIJx8At/k61vo9uB
BAHSxdq9c8b9+LzLTrU3wGpll0C+Nx0ZxuEO08uUwWAIZWPuCa4gYrRI9zU190SBAHeJtRQVLYgs
15D28Qh4GBkdMX0743khSk4myybop9cF5XexFG4qeI7ce4KMSHbHtMYv39ZEduQGHdIls9Pf4fux
nlLWiRAXGIOcHQFuEbjNdktba2fsjMjO4F0T+alXeKG8917hFd8Zw/u0A4p8tHVhdzqeUEGy6sGm
OsWfGXIxpQrc1orMbs053+vozYj21r0un34yRP+ZSoNyo9F9k5gL6w4UEX871mpOoR03DXcQtnEK
CKXh0v9ZpjUiudS2TZ60/J3wFFjwJHumjcIzpEW5apS+xZRdw2fBl9pdLX9eiyLU9Af9PxROVPHZ
p7+8Pzk7EY0mcITkbf6YCmry/7b63A4ufHlQRZXMwHpPI7hzV+ix8jy1JXIxTLvi0L7mV9iMOty6
lYAiPJEd/0ODwAUfWAb/MT+TK8gbkjx+x40BpAKF0EN+OjlW+oEPs/0GxK37TP17Up70I+RHlpTf
3jgfd2CCTFbPhsBiR+putK4gicZnjKMgVDTbl0FFsGC+CUF6/LHoK88hKYPz90SNiLkiBo2TzfGU
yPCt9c3Zjvmje7O5P+dWA3Tl6z+WVmp0u8lg4784OuoD8BPFTzyuzSE1vreRCuBYsiUSlDFic5t0
KXc7jRQ5rsLV+ikCGclSjlxSHZgJxGsOpIPvIxCv9gnp4EKeiblqDU8BCtcZqwq9BpJ9KRVpdIc9
JEXLdE7ihUxWixVv0SndGCnmtnz6zbclA8U0o0imOMtWgDz00MswHRhARIsxOQYJAJKKsruT4aFp
C0f4lFJ/9QSDt6v2qWTHtB1JfNr09Hlyg8fcyWYaRfxMlXTX+NOrlw/BIeqqS1273oRWFVTqqXNZ
Irpl6C339n8GUF4nZgYpCf1NvUYxUP0tE3DbzWfT5U+EQI24IfSyBB43OGZEjrhZr9WszZMI8AmV
VDNxEC3olj2EfWNcuTp4W86uTa/z4eBvWbK8hVgzbY9T0fDY31SRL7f1fBYZSg7nZRoplRJJ2jfi
fGiqGrmwlLyiiCII6YN3TP02+X6qFaFTMQvpXUPQCWYySjbYfNn7Ph8jTZVE6ysij+hTLuR+9tZw
jbSOzDPF0Ecbwd22R49+U3hP2TB5avpKdvF+ENu6+smNMCsQex6O2iZIdvgOfTAOZ4Rd9PSzt483
BN1qFMHWgSS2WiwjBuR3mVliwRhWhgV6xSDE8vmoWflmduUfNqrRkXfPzb3ZOuftSibL6bJnLKo9
0cJQU7n+JWiHmdSypXvtiZfVWTcPdNsqQ7Y0wCQzApRAyO2IB1XNPAUlHoXEUs2SwmO9C4vljOha
BJZeIO4hjxaTp4pLcyfCsDMb7EgsOz6GQg1pfPqFf1TlD9FYWkd7Ww6X5z7CLTyTkC12jRQApzX1
nckbRk3zJxsJ4JjOM/zwTrvPQf3bedbOSrYqDNRrzr2ds4xq80U4nE+5+Of90eyUz3JI/dQ80Lzj
RjnFGWeFHpA6BM6cZMNaqTryKuk0JVdRnq2XwXdPFewSX/RLChcPH6Av2hgLpj51W2DfNiYEvBM8
LgHKTbMi67OTQeN0ihPpePepinLlC8+1U4cLN44p7ny9WoRJnwGp5lLef/BRgGxrHZtotD4ayRow
K8SZEysKZieCIOamJw7P6gry+mDThtLa4qtqTyBIDpIVk4BQ2mvsmsP33BmplE0SzcS2eTsRGOM5
DXEDeQ6FWieQjGl13yTCItkpUVm+c89QvycEmi8TtSviQB1nZCylEbn5/LpdsFW/y4+Hdey0nyOd
Bd6Bpo7N+IGVJ3zVYnT5Dd0Lj30e6gbZcvGdYHYlbkY27+LOx68SKFo9EvzukmpDIVvTHNPOmeAl
6CJ6+tsEkpPaLdJOkT6Yi6EHoeBTEblSRUxH4dTycAoUEfjJE4Dr5eLFCZ9hrzgbUxnaJ6u7jaK1
5r8V8MtfFY1ZVYjTq4lhXasywYqjRxx+vgeuJt6jx/dDQOkHvgRii45+4r9ftXonBaNZC6Vwdo4M
waHXjdhbxi3kK4me53dDXJpJwUQKDkQJ10AzBVeykrtXH1GHT045jhyt4OjpgY2+GqJjS2dnuCod
RBPWysny3ZjqR4AM0Un1Ucm+KQ0CqrhO0IkFKlJmJGT+DhHxG26UvEHFNBoyJlIIfuwjk5+/rvVY
5n/ZYdBMplEXM+yDRKmuIRRUHfadbIFIZSQ/6U5KqqEZeLqa+ERzPHz+YZh42sTGW6Hy8XE/2pTD
EjwxlxTT/Fk53qrVpWzI+HzMaz8OKJZujZ2gEt+RkibO/pi85DJkyk1YVhfCfYBZ1YJuSRhgrfBf
3S0AKwkaSimUm5Tm1+KD/JzceG7rEID1fdSUgCNlrjQog0rIutpcpyA/J+9Km4fTtwXLfkylrYTp
LiiSUdgGhPL0dYYsxtpWPYacGlTqmYKGnIYQzQWhXiQz25HmEr59MFt9duio/MiWDENig8HkP5/F
L+Sl4b5hfocUHvuEyppxUw6q4HtBgpGgOkKvglcXqDTF0m0kIDJMgfAOpjBJ4uc2cTEh716kLaeT
IEe+RBIMsBSL3EupnThlHVDNhlUAwnRtxwKqEb2z0AeRN0Kurd/HqLn01xUM+Xm7VcP3+22BTZjc
XHzetIgP361unnslNA4EC8HFp7sFUDkbaE5kD9hQbOZrfz535whtGv4HiJPZp/jRoGeO+8E3VAra
jCbchL+j5IMDj0WZZriqSn3Jn4Q2KehDSOKTdZAIbWMrt3hCGE/07NBnC9r4SC+BaxfRSmtNBZqx
mLp6gzS34sl3mgnvQ9Fj9IABFMKYyl02uPMYpHM08IdA5P6+krufk0G+lVUs+9NGq3SC4PaEBmPj
TenfKLHD3Io1cDEiPTYCv8jsLQMk1JHbeK656WFfRMUPgr734kl4Sds2161trKQmNl2XfORoFtoX
PSeS2rDcmQ6/SvCbevmvTxx7cfc0O0CA5tZcZ5T2Ik41ArVL7eIQ7dJNTL0wax/yKvbfKPP2FLmZ
q6ZOmz1VsZPhWSaO866A6cWzcipC3o/N3QaWIgRj1MuUAHh5Mm5C3OcetfDW6uMDEtbyFGkJ7Bxc
7SXo3iJcTpZODIkqf7Etfwa3FC5REGTgRJuzNOc3n3lkv4IAzJkvX9LAEtCTSwltzHs0+ey6ldHP
EYMfwfw46v+L8CzpTom6aaAFFX2hePi4JLE1lJwQKbDVHGAxd37p/iEU+iQ7ADNlK5Z++fsml6Rf
wOdIFZ6nFfVaxItPToGuoXlcd1hBGwk11SCVyBj2RJJEWZgSv+mUEmT2dVzCgTHwstvotlHtUNo9
azOjTU8oFDVnUjWTvLEXGaw46OdrRDrplU6VshDKzp5f2VeBUY5djLR2qovCtjGWdnGxBx/uzqSS
wE/0hp/ZyBFEYJu41h3sGD/NkfxLAGdMGxD5TkkOaAcqWXmLkR2AE1R79Sekhj4/PuR6yz9z9Rdr
kVaVBsUZuk5vdQCevAkMujfhhEpJspYvdDwX6M09hDOJbA7baovQ/tbVobkIuG18t1X3IrOhpHoO
1twk7FbiKdUhMJbjkV4r46c1i9PD5N4O5GPMor32NUKkeYlsxkq93yGIea8WxYyM3sl2BC81qRIS
M5I8kpdoPDC5I1o6M2057kKokKN4UY+luYj5ndfkyETArPDem6kG0qn0WwAaMtkOR1T26Fpe0pWr
dSwa5hyl381O1RzpYImO3T+0J3Qq3iZ8/PykkdnzGlekmGTpdsCplQiDgUjmrBTt602xX2A5/g+V
RABz7RLaM3FDHtDhri+ds1AsrCGxy0O8TlVmNUt5cf/3N0dsz6VRDSFiYu8qj3RyllyAs1Niamqo
9OxL+RBYD9iz6TP49SGd2h6CxfzxgasKxfaxG0bJEonDA8Kpit5cyNMFTBAqglZL5rFetITyzBt+
BtwGfcgtLT315mJxyfwx7WgC49UqJz8Tg7CgQX9HCSAiC4fTpGLLWMsvdMDNZabRFSklof9njo/E
H237ClDyNYTO/YoqjfeRW5SU09WV/cQBygM2t2NbMD6e5nwn8NvC3eBWem2y4UqpHffbvBtHKp2X
wzA9aoMPELdTb8eQx2Xjj+0wWGlNtRuvoxOVfcwb6sDjm9SYig9Pwi7SuMk4OUPX3hzi11YXrKsy
XvLeSt1tD2uTDLVFNoVRv9HgNvLUANSPcjqYd6wyaQcY1Gbo/hTgaChtplMA+B3a2aiMCvJdmT2l
0pmSpJFmuSFSe346XOSDF/QYHhBSDAKZ/eTEPXREE+cxVRxaEr6X/X/xNNlgZXNa8NGRuXxNjE82
XIwr47+RwqDpBiEEqqR1LLOtf8D68sUf1t9/cZV43tNS/ymf2N/u+C+5k2VngUwE84zV8nRQ9pAu
WalEhKLwkMcHGECO49/ccdJjh4uKm+egwLP5bicSEBp4fEc1Z6VTL6SX6NzqF80xUjoN0mzZOkpS
MWedJZBROExwmUTOfyVVsb80F4gqn7NkF7Wi29C3x2rsrsMAILSBDSDZtiem1dHCBGbK4kHwzfYK
6Tlj+dd1Q6Scenpcgrtep4EN8O28N0TAekFUUluLYoJlsOA/yaY2OhjefUiKKCN9eKxn6Xg+/EC6
CHsbLxqMu5nACMveAghOA2oKc2qBZlw37CyhJKjg0yvPIZqhfyk60tuC6oEXB8wgwa3kJbZGy0B8
gjpNWL4fSyl2L7M7nyXIFSSEaeM6JQLjLSu63NQuxu9eTKw5U/4Dh7K+U+C+jhj/EArjHj6VLI72
miSz3pG58prPeL2D7AzyLXLVwBC6VKLbDUgt4DVQ5PsYkbJYwTwNwF3AJNoUJjQ3Da+U1nHTuj2j
8+OnbFPxKzDakHeV4H2Y67eW1+KjRJvPGmF6dH//soT6dydboLHST+5RppARGcB9gQdjCm3dHKAk
lTFRL0Fs9Aou2Wq5iKIAb9FePPW0bjdCbLohtyyZ9aGhu/eMt+qw6VdoqP3FRsW1+WZpIDotbZJw
A67Q9Q5iCCtn+M6n81soNkWDeizw7cSXmEn6O7c+csdK2RliKQKsZp0GHxcCZXaKFs3TC6G5QqVS
1smXMkRGV6GRU7LmqyufKp0gjyHQF7jqlrLVm4B9amDFBTicl11a4mLSH9fjgYLNAr+kIHGGDu5R
2Sy+awFbQ9MCc8iukUoKpUTAn6Sh82heTRPfIOqZtrP7LXSe34ybXQqpvhIsvGhzlZh4kICuaetH
XpB2jHIb1M4k7qxWBYfTXS+vFERjXjqM03YT8kaQSVuEh6J2623UREe+CixfrOkWTX4CElEwhbHL
PTbC9PvusycBReAkpvGtdG5O+o8e0mnQW5IFAKmF1QnddbHrz5UfPEaycZPx7uqsDBxSRoKQW08+
e8ucQ5RROcU+BVoAKCtPLcgqjOMvjsBY6ZZmvPH4Wliv+ay9JdM3YavSUKUqoRHKRX1clCscZ6VB
6X4MhCaV+6gvdjBMQTFhG8Cn3ZPB4CZbPj73+wao8J/cUBGF1zMhXFRjV7MCGnx+N+mA9PWnO2NJ
0FZ9AVl5RTeSoR9FXVvbH2X61LEJRpIEyWf4mOR7jbglZ32u5584hVK8UY8IMqN6bkIlAMwnLI4P
apDlG6cxkHJFIHbTWZIfpwlDidEf6W64eWcOngPe/XlZTtt8jgQAx6cWozgjTXlo/K2//UJeHcR5
O/ap6WvD/yphdLUGzXQ/9b0EpwmOlooAwrx0rza/miL3tVR4R4U90vFFEAT091dAqXT+1N5izlmw
pYVWBaepknlSdrf1rVbnw15oFPZrZd5LmzDSwCGM0BpN18otzXFrjACYJ0Axd/6c5yyfn2PUfTB1
Y/QQvzlDTfxwZhCvqvYkXp+gXb9Ei4x1De5b0JLD9C8N3B1cX46Q8obVN9w/vemW0ot/qrM+BD3+
mQw6fYUViX4NWVh2OWvUuW7xJCuXCAqt4mn3aHXUShpCFiKP+ORFDj/AGOv0OslKdFz12t6gmtqx
yPnIlE8fCE4tpSJDN/jyVmsF1ltME0YGlfddOpwUHWT94VEeR3VxxATq4AoNSQ8t6XvFernY20vE
VGQL1LCrnOHLP5xOxC3O7rN7ioKx64RdaYKRoq9K0ix4T8KgmyHoUKVfJQOjwfSedyEjws5yXaAx
snoUlpBlfPgLhm/8k1mfIgoM89hrxIq3ekYBcAFAK16PVenUD27ObX7WuU7gMqNgzg9Xff/0dlnJ
7J/I9HQZyWMfQJ+Cz05Ui19iojFIs4fuOaW2opz5lZcK4lNqPFzjNFPd0rh5jQ0J15Z8hhDCp/iU
111SxwuaY2Jqc9WNufoNeUg+5bJvsDwHsx/3KGY76iDBt995MltOnWIHryfTeOZQPeA9FjNM0szu
szEbkhXhkYcHq0wvghMe1msHyGsZyUSiG5DCSRrglf0B4X+SkwZWTGvFX/5CSIZWVqEpuJhmvAQX
Pyd862rLOnt6Gfp+TW01RmpXOLcel8pQXUeU/1yPEI5LIh5/a4cQ0m6KRrl3Tep3EOsOJbqIERwO
7yOX4SVCLhUbREH4aYJ/CYy82okAfxqL1BDHIOHZKkhHA3MNGZHo8mylRU2q/G7uwWCfmsX7OAA3
m13JVbd4wgwGVfpps+edM/fXiBbGZnxiLSb5gx5tN91fdOFz5qPfN5MRN4+8JGokuUw89I44NLeR
bTa0o9xjBYd4I8q80X/E9DLV2KSODdWNJCD5g8b3AO05xVtkPVvzbNkDpK+JYN0PHlrEGTdp/3l8
tINucAWmZ0RIV8BHOti5WNpldSU9p6KSpYdsu9ebS+J4L9dLpA95ecjVajQAP0Dti6MQGDjmtAAz
1yMSb75aSwq1G9/585sgJxUP/IcS9C6BoRepvsxAUZ3N8GuchePE29ijAHn2AYKWHQ8+Sm/b825W
Ut+O2VL2Woodx0Wq86HMRxiSoBzM7CDw/giUJKMnZao8Lc9uV5qCR8CWjZaNvnIieiQpAIwPxlQp
5DDdI6V2H/xZhCZ2zqmchrtiIvxZeLR84+rDQuwfmzfBV8ojgkK50xQ57ICIP9TsaGOQUk6n9Aww
Gy2fKsM6OFbIDkAPQTOrBrNiYpzLWIrJF0acSn4xDjVsNHVQHvLv0Ndkd4G4A82LMRqPrZ+GWLVA
7YZgvPaivYalS9EnAzx4VrmyS5TxNayRQNijKcf/SMYENr/wWP6woqHyr2SUzJyCemqd7OlpxXtr
Z2Tp1htk8OE5ht/wqw9qlb13RC9VL8x2PgXeOsxFnPla5hS9W+uYdYiiu5LTwH6kA53nFuaYJCBF
6Ug3/TtNqhTKqJZ18b9nc05/VxZ2qrLVTfRKX37YlVnkAn6PNNePWu1VxrcfYNVIZrdE1jqt5PSL
cPXd0qoVuGM4OnVlrY7Ac5agnonBV6VdlWP6ZqkAt9kcCM3GXBpFMJCwRwKhSJxLvV4U2mLwEe8x
x+d/3wFYj56QRMnk51NlnFU7pfXWUGFFG+LOw5JFtV4C3l2SBLpVv6FuNRXpmCyrtkxh7llzqbLV
AlQTINLAfAJTQ3gUuWdz5Yp817OfTzTreKlywG8bJGWYIF9WKyiuhht/vfQ65xOoM94kiOP7NpMi
pwuXa9coO/XvOJ3ixhEnkFVNs9uzEHplUift0EksJOb3kJC2Juwn3BsesrOdml3c/3nvCL8wxfvt
/PFhMC0Q8WtP81v4l/j+k7cpjkOAYQBKS/hX10ExlHA/ONy7RFiE5ks3FLOuJQQafNLh1cNAukJH
GDuJDH+4VK8hlJYeyQKyENO746J41WczGwKwBymjXft9vm744rmo71vxmrRxS2TaSVpCFtehRwY8
gzEkgsETukxR6GuhJErRQLRNIhhUvahqbvannG9G4hqcqigs6ugqbNeVl0eVLA0mHOyEmQnYO81+
iLiyKPwHve2Y7u8seTiTDFE4CT3y6nIM0AwaiirpH/Ru5WqkdUWGgl5c5gcJ/rLOwms1AY8o0qhb
hOHJDLcddIT/toHQeFdJSE6nFXSp9nX/Gi4Q/f0pJQYrUxZHLhCcrW7n7eduFofQVJoo+Zg0L4LR
GTpgHjXgFE1oK97kKpbnByT9CiPobDfwLWyIsXBAsspbtAPCFvYgTfwo06wJeoN7iN/VezaMKHEL
0cV5iOueuvLJAbEtEulyJSk4FTBSI9DUzCozEAzqp2Bd0pkk15ZcnZlTVkm35KpdvDuzcEvC/Y8g
IoCw/cBkf72zOmmbffdnWtrR4DAue+uu1nxDKWxKewYgHbKm1Vgfa5c8cr+n90Tisc69DJqr7pJo
Je8wk+vcKFip9rmiOma0DS9rdsxg0VJFeQVBD9762c9psE9Ftw42qtj+HPpGwdE1m8JKDT7MZkwq
i5sl5Ti8OqoOFSVaH+Zm1fuXaqOGt8lviJC3B1s5q6sD3MDrhBaGahVYTWTQtbgk8nE9Obml5eiZ
CRbVm7vVdf6FK/LCXZepTCsct2otirQjPu5ukoad9byO1D0hK7IMAwsWICBLygIS9Tr7M/12obn4
N31EOSTLiyjE5heMSuwAsA9nuxDgET/NEY57PAMcIkzQ2qV1T5/bHWEss4Zj1CqOaPLQ756+9ClB
lTXVjM2BXO+WNADyIotwfbJwfWwUTopJbgXHm6LO8UNpJ3duOkTuDoVn24WBw5YDNapOd+lUtbJ/
LYSV9pu7xVkcgR8zCtWoco1ZTAswnUgAjTfROZEsVNpyqlkcuUoVvIpnra3MifGwgP5ip8Rdh6fH
SiGH8wXYMDI/ibdKpUSpHlWYRNtk9ZT6TR1vnsmcse1HuD19kFdEOzve1pPM/TIvXEOImaq6kj/T
5hgbVysjI1G34tXKohXVbOSlTWnWlsy/3lOt4lY/FhxkeZk6dbi/xRCp2OoSmZHr0JFeAmFCnWBF
NyTXXlB9MG/nZkzIsOtifGAmgqmSnB03JoWHTWfpx9jZkU3lXbPyEXeZCo0BOLirC1k94b+UCQGk
DLU2w2dGNMPiUhm4+VdIJ8w6mgxOcb9aK+ZRbUrFBr/QfzhUk6wgBgKYIv4++56N7HT2cZ0/hWoM
StLuk8DnJYI2ydH85SREpp/phMEPGVvC+1Z08TGyhvtNdW8U+HfgQh05i95jSFtgVCS9sHmCAkvC
CiGvMyF4fvmrhlmv3bkeeJQ68nHQaeUACFUnrEbZr40UhyLFPMD42Dr569iW8XPCdX+EhNDGcYNK
42fNWwsVV4zq3MBoz5b7IMV9i7xD+v+3w/KXqj/nNNklTGH3kokA3+OVIrgQlMDMEGim04Uvvupz
CV6I0tVR3XpvJo6dM8gm+7fAYgtUHHjiTZCjCL9NnGwfWq5er0ek8KK1iLE2OQrtLZx1Mh6djDLi
9OjnYZXNlbdyXgjiPFGZCS6j+UxoW3k32xpVG3YNFHuXgM5BgKt7Y6CmjH0BmPbeflTihR/fzgbI
B+o1hRPyyiP5vrYMXs4Atha0Ru1HsG27LMggAhpIRZC2exlObLpS1WT2BWbbbJH5RBIWndeuv9BW
nXAygzygv98SlmORfrsDH9IfjhXunqsT58drfaKzyozp8Ovj92U2Palu2E1lExmeGi8KE+jmck4e
8JCkgypbzVSCvlXMOsCOEX3HcVVwu72OzSsN9RWxZZEyrGDIRwno/BOma2Fg+LaVdGNwYT8Rv/D0
IZxanFzFaKO7/RzxSEVS/J5gMtzVDYhdtTn99r8nhamR5jLFNhoPYxwSi7oQZXmE3rVMzCMq+9q1
8bG2VDGhDtrCuKgotoGqFLHqiRYwuPmUHXz5bN2tkWxp+MnDiBblqaU1UZ6z58GrAmHNNWwjYyKX
Lc2c57BLLacKtKJiNRf3DmZqqM71bYxs64+1KaLtHFe51Gg0hidC2CJlNSmUnoGPzy/MCJdycvy9
pNri8jAZK85JY0IIz3sQdzWUlBk3E92Xdt5eC4pvGqXKH0RXuEJhhRx5EcfdoPD0gbJOq5u52HwR
OcpMoABYEoo28rhBkB+KWIyiKNdFbNB6y0QtUQmYnlVeQv2CDxSJSxmxkD5sdquE+6NknSAsF2GF
QccuSB7HUwuebmhVK3LBiHyJyYLvkJolQOZ0ShUuqTz5/XxdGI1kn7J/QHKnQOUTZPrQljydDBSc
cC8warvX2Nk4f0f06GC1fI+p57MAnfWF8nN6yPmricEs8VBUK09usoKWo7aRVN/5l36cDwMPt8B/
GgIBhbO8IagIqY4qhdBZf7V8fF3M791IwAshRSsTqPe/AVw8wC0fmLFv9mqdt/SwEm5r82YjWNVv
O0x2Bm2xVGToQYPYIDdkr8dKyfLmNe4zqR+SY9VXbU3v99XbLPZGlUwcu+qlWgFNwsPiP6hIkndh
jd1brcEvhwOkyZFxrHqq24gsPdNZaJD8D210y17xgrlLkBrMXeWK2/Tt6MN1zdWTRvKDdUFuGq/W
2ir2sjcfVU8g4VDhD5gbj0elwwfqKzB5MHYzXz+W+Ib5R7TvMQQK/gIPFvfzgaZp0oCXvW6NbySq
kAbPv7CBnv28bOAeF+o/mRDIyNsJNpZqYuuYfqMWp4TXXOOklh6KIrEVpPzvzRiAmIDs8kotIuuJ
/8parvm3BVVfUBOug6qVVDGEnOoKNZw8sbTWqvn2FO6zJ3wlrUNvXt47o08KKSC7y+kfSLskHVy3
kttPhvhDJetL7hGyYRXnMMAYJJNNLSz5NG/VBa3hpioVKXZoy+2cFUfDVIt7mWkK2WtssGNIc/8r
eKskUb9efd9W7RLTyzHDwulpV824w4uLzGUVafMn0jGtO1+fWZNar8zLEo45WLM7g/+l9b/TR3zy
ZRsOVMyJaPLSOvzpseocduXwfxTLcwzXrObhI+qmKB5jhTCoB99t+Kpv3FaFIGvBH40a9H7Z2NE8
o0bPqFlRdneHOZNw+p+Esb1WZV9INobvFpJZssstuiZ94tLpn+OJf7jdISNFapp2eBSrYpX7n+Nw
ai8pchvtcpPwMv7u7Jhiw/y76AdmiDhmiESa0g1tDGtwmw5epx9mRsE5TkfVBTax/uFGulYtZZ2e
WY9BSD7t+oWOT3fnv3m+g+AKDzLjKU3CZi016eCK2R5VqdxR0zQfMZxhU8Y0LshA5zKUofjV/uX0
7SFgrSP9PNeYY7BQj0nzan/wZCmHZIy0QCDy2fHqS1AZQ3bGh2Wdmd+AVXHgmU3Pu+x2kZ9ti+0B
P0Jr0nBz7sAPGrIOmqj3+ujScYex53HchFy4ObrTZrczTNyU/1/pOEcYefXHFjlDl8o7T+qcP+hf
dCWZKcfzFVy+7VnQUnjvOT9ECqVp3rxNweF3TCNRkE/PKUQ/Pcie5j57pen6SMH3cmRjdo+f65Po
sCdd7e68VQuttYiVPAU9JoMWKWtJRWvpBixoBj8wmIw/ohwJS1iJlYQ0V3xRgpDCNwBhQA9pnZTZ
ucJh9Aj1t5MVN/5x0EKWnPu7+zC/hyAGMFsYdempyR3u69yqUzNqfTfIlcqsWAGHm3atgIUdzT+V
SC097NOa2bn8y5UozkO265As48dgWFKiAX53JBDndXIqR2c1PeY9maf9NXCjGbQpOn0z6f1yrYJo
iZssyL+4CVyPyyKWkrrA/kULmIfP1h4wXaSC+ARJrlFytmhVJ6rtgh3+Bn5uVrmlwPgl9ML6Z/1R
eX4g1LhBiv+U9+6kNDw8uAxoOUIIXGE8l0OVAhNHjDshpimJQGliDIwOYODjv6q9S+DE0Sl6z/RD
8ja602Mxi3R+OVzlt9SBuKsM8XYX2mLZb8swYSljyfMBV9+T8Z/jY8kAyiVS4AIzKe0PWwH2Td5C
YrT0JDc/597f8mxd8MGhXknYoRDVY4GvM5S9tOOB1UwoCZuQuqOzf8rR860lvH/sbun4K9gMFCLA
w7Y8PaJEfH0pXS3q4ohI/iWaWmBg4EyHfCkwrprQGi4hvJzuigAUt1FeOVk7VqEPWzPDVJBq1CYq
KwQI7c07sKnWh53auqASOPnXbCqrqZswoooiLeTJb0QMCmXYGkhuIM76jbH8WAkHAEfnzac/v4aQ
Pt16DnpR8Ws3iTxnzMl+OebhPaK3Zj1snSwfN8vo60rwiIG8HeyNk2M1RDc6F/ViHqk43WLgZsgn
aXmGdynfd4edEAwlXry7RNIAWkraNzQ2BEQkOdnrqYsP53JjOnRRSbnQ3gtdRbXxRbawjADgM3v1
4q7xg/3YuHKVEGcmvwokrKxh3bqq6uj0rfzuYH+g/UOGLCeo/JFp3le/MRQj3FiOWebDnrXv3m3u
g53DURl/p6SAuYiOC30z1JKeDl3zY/rlp0TyXAPIiR26shgU4qlHt7TVNJU4K1ijgqEAgti6DYkY
EUKwr4y6vWDAbJybFjF59tozxWj+rmfZyNKmme6P3+XEdpi/wbPXQeRNZBMcXg/IA+XlsyqGVQED
6xUCcUsN01L2v6jc8+Kqdc9tBbndWAwWmFVnY6NMw+r7hDl+YCQ6mGEq5ooHiVRc/kZSjbm2VCZk
BaKDriiXfqIe5yBG9mbNkIIfQbZarLV7ZsBYdOp9wxdgZweF7jQ5fXfBxBHnOPO+ivHG+qBEjMXr
cMBg6NKwKJ8ecIjUTinXVuU6n2jqqwyNN7CaQkUmIS7falaYaxfjYzVDFHcOLkADuXO+/d9ndckD
Sh9SqZLQv3+0PpBL4kNT4qCKYaBjWVbqJ14pkvk67GVKZ7ZgnqZO+VxGh3GgGEvQTbUmdb/9ENqg
ruAQxUV27MaMqEQaUu8dW7GtdVhvNI/f/hz5JB7BhE+2Z0Z5JjsVuPoaCWbUMwhw+yZuMcW4bW1/
phtzQnop6wBoxAh93KnEv0fNhoXDPmtPHi1ss0UGwg9Lx/92//bqmBNkOCbMSOy9dmWzXMUY6Rqp
iVekeSZqizUvlE/9ZHQxxlSwuuFbjuBFZsnkKOM09vUDew1rn6uho60c4TVKNOPW6GraSmQERyS2
uuE19kEY/MhdIQHRFVXnNHkoRGcHEGy7s3583nRAydc2XzfvdGEiswK2bGbOUmyp5vw6GZ3eOTsP
W6tuWS4vdVr6/w+s1XLYonYp+mP6irAwb9FAbuVGPsfO2R94e/gF0NG4/pnNAEzzmnPKvn6Klfd1
vIF0bqACBRsClbELVrt/hU6oCmfkRZfzWTZ6X2MxNqgq6RCeunXhBxT0eL5v0F1pmc/RnMV2XsdY
rtssg/uhe9FCrWrgYfArLh0lTtjM5IgsrkfUoT6j4uTMMuOGr6tKm2MDY4LJc3zuR31e3ZirJaZ1
Pv6Mtt/KKe9f8VnE4WgfbcbV8bCh6E/VcO8Zccz3Qp/23XOw0Erbs4JPaXzTuXiBwy8qJc9+FZeh
R5n2PWl5+84ileNnDWNJC7ExGRlSdmdqkyDM6mn6iOefZTcWcH1bnhuyPkn53bm1a52DpRQH24/4
MqraOaFnpl3a04E3WhLm8hJNR/XriJ+Mhwq+iIcu9cE76YUXn7ygckr/EXMOz184HaG1PV/Yabnw
BO9zUM6v+3jty32owxmPN3QtY2BCDDXiNN4jjqtzIGrQUnMZqkR+HBFug9UIDfSjlvXcimasBWh3
lDPSheb3M+sri6D/8JWK8t3fyx4In3FN/jDIK2rgwf0ORXi3EME9reJzt4Z+UfeDQIi1XmE9IBEW
8hlryBJLKJ69b0V0Wkgq+yU09qJlYCa5+sDNNXkdaN5aySK0oTcVHmQ4EUAZtBB6A5E49Tn5c1/j
9x1X1CrPlFIN9iH5EtV3FM6FytpAN7OSkC/XoJVHEYc02bAbuEJ269q31ecczuPQiMnfCCTbmwmx
WzrHHS9A4Xr4plLRDqzookZkGXy4S3zuaz4J60/cuRMvcxtppSfsd/MARBoulyhTIDOG9qBXXUg4
p0XPStIE1TEwwHfhEc640f+qvgxqvnIez2kq6ShM2RJo52QxssCOhpTMMw1RRteV5zOxxtVdSyl1
cDtwMiUgEBZJ7FccMowxhDZ559LhBLsoLMWE7+APOOm4hmRppXEfZSu/Ed7femXoIk+lmr2q56eJ
DmbyiREYSviVPataGO/K7jCBraqmGvtO0Lo0urRrvTzj1/XIrkaYDJrEUHYOVFtXaULheL6QrU3R
87CkQ+BjfYb9Vj4joiMtgL7IbjwoTDBPZkJNVI/S5tFK/coMf96xcMJ7xPk9B1TIoZHtnaLEYgQl
VUFLN65yMe64IFdmLl9SfbVQzSpHI/ubvfcNFApxG6E7iUNyXa1nCv7jcLdjZq5QuAFG2h/p7VA3
2EqLsetPSMt/LhrMlUMr7CPfmcxbJbTyhppVOnkkhwfUsMdZvQC1zAjgFjH0OcwIjjmchgxVnWJD
3mtxoKBTXTyYqZGwsPizLzLd75eggvCXlcR6h0+fZvsFG3jnLezt9w1Q6Jar2TmIPOxijvmGw2H5
LRnlw+g3q9n6OlJqFj3PYUTbUpZwOHmv4TPVUoEt2U1oBecBSTMG1om6AjF4DeidRhIqF7+Q0+R4
DD3uaRkffBEAv3hgmBoS603p1NfJ8R1sxEjoiMS77P70FItQcbQbyqIisB/Y+jyPLbF6fojUfAEs
Bb20YipCIzFbVFWUkdbapxtRwbbeGmbmUO2KV8iNBH+ZyUnnR2fAm1MQhJmFMqMU/Dp+Jh3XmjIO
nktDJ4I5VhPKsglbAPxkQBtL5w0DwYMi2jOdzOh2HBQBJwxtrXL5nONKFi22YpxrRqEP0Ot/bdem
XaYPxlaIM9dDvrAfVoPQLwM+dUnBk4JIsOD/qYCs6FW+PMaC2rMT0hA6Eq9Dk+dLAWZVYzGZJ0b1
VyqsFcfqmZlvXHKjdiIDpM4h00+6HBT9tf0l2eXB+5pc00ZnBQEhvhQslcwI+6zLSgo+fmps2llD
GAsyeN2fPgyCzUGrgcVVmzL9cEcL2zp4ixyXPTagCLkc5wlniQGkGpOOtdXa/4vAdKgYxfLB7dzw
vsREZbAfK/XKMubYWHilLH+380mSlpixswjSxycirY+FZ55C/52WLT5aboja0CuKptGYnvZREXIs
+8j34dbadSYJsf33EwumRVmLyNrGORBM7PQjAieeP7xebZdWV18lTM95COKnNxM/xwzEGfXDeO2c
xxXzNumEGNsRA56CxKlbjqkaDY4TKQJGItJplSYWn2rDDcqPslRrOwRVl4fDebTCIgGLndFcGfp4
u7H66EFR39ZSFDch0gi0y9KR+3hW+EuC9EKaVHHUb/AC4CkLJFwYs9mFN/U9TyChxT45tDHJRiey
rFFKX+ntjJ4EpzZcAX3rNAziYm2skHW4yGRaZo09a2yq9ZuEk206vPRwpYAmMPunzSB9Leho5gXX
8TiZA80CQjnYaxrVeuDC9PkqioNY16n1d6ooomuSY7RYebTwcvNnUi4rDwgcMhU8ItWghYWVsOds
fPrHI4DZhFZzUZuDmozG6nPDE+Zd0xhfBxV/Gb3w4Ey2i8H3FtmPuabhzAA3Gmk8EH5tloR8nDCs
Y1a50SrFgl4DDWb6vgAlU/WHbsFQ5hhkt24bzXmRYzhdxTdLHyOXtw0fL2PyRPbeb952ELXCOw5j
fhBwHKvH0wUawQhlzZNKcKt+suVPEDv0dAJLmejCfJtMUYAJw0+D9RwDV7suFogqYeIAkpXABFYV
OjLIjHr9BXWr0WPZd4J6T9UC0/kEtJ+sxE46u+6Rj+OcFFyW87Z2pDJgsiFeyJHBDfxbwrqK8ged
tREzLdi70WaFc+R89ATzREUu0wPH43xW7umxw3mM2kw/n3GKPIlvf4VZCXozZ2sG86cduHiynjRn
4aLKeP/gKgPQk0qB2VDdYVXs5wRbzZNmQcPyxp7An2Neje2z6/u48gIWAWnwBgylEB7WcEMIrE1q
8kzNXqWBWsQRZlGWwJIUSRu+QiW31i/uPdjZoKeCt1C+6gIwpt09Wa8pDVghw08jKGumauy4gCl0
ACspE7QQJagaeDWafvkSLz1NQC8LrnNJ9ddwkeRZdcnkm8SLFvEng/RSTYW7popiCw1cJOxnOeFA
/xB65oBf8ADyiSAwUOcp9XZ0HubsEuLFzCClljaloW1HoCzz8D+zP569EPrKLte9aF8tWS2NJ1io
dOUICIcY67noURhFMXDLcmHzHV5XbICddfLZmHTOoXNfi8iTVchTWYB3UkYfWYtKEhgL6uzZonxX
D2cFkMUOToTD6pwsfQ2sbpovR8uYSgrDYQtQJMl39MK1jHGc+T9hIsoRP8e6vuZ5a/62kDx/ICfC
+UPHbAhvwYLO85ikYTzJ8sUbyGaXplODRqpI7xQVD9f+q5wmmFJ3sIJ7uhNOrKTctXvYy+u3Ge1H
9WMSvbEqZKZ6alPrX7zV22/5jMQCViUDdqUNkIW9af71Wx6KgV/DrojSwqBE0NsnIk7vI4LO4lth
Iw7MYiCr0oP74xzNvURQynbK9tCbtcrumImeD8V9O5o9pOweELsR4CVaQVP24YsLsDLP/c5VjwY8
dotGUJI5cTK6grvFRLAFMalUZNammj+OdY/TTcnMIflkJHzsIlKSvF1V3yT07JgUTH3F36zGbBL1
l0AiSjCojA/kpqTT6Mw14WGpw12DkQtqyQ4y8riFXwzzp746sGiU6cYqjkNijw3O8fQ6Z0doI3xr
5PX97XesmhsTK7I/9wP0DJ5HZ0QMAdSOrVkg69pa7x01F8LeGBoiCHYV/XuAFF7Hmrx2x+SVNSb2
Kul9X02z0AZ9epOwqEd/zrSvXu7xe8gz7+W+Lp/nVej2YzIg9JUjZDlGn9PbNOtSsRk3es4pD6EI
Dyvx+uhJPe82q9Z/2bjpg+4G5V5/4FimO68GLBHbrTRbxrUw6bPR+ce4aNxGVINO2r1YBsheb6Q9
ol7kAbEuxHMNXnSidhgbDbBnWJv9QLe6AO2d4kI7D5U+M2yn4x+NDAlDtK9u/uQjIaPrgbeZhPDi
kufuE1PhAGVLvIjP3kq6I/g3+FpucQDsWi/ofA9BoezDZmr3+idmpSrAhDKzxUoX2yoYh4eznbYH
L0qLgI5b38bBmERgDMBOLkgpEPxWd1K0WAFN5k+37XgjguNzQkiS07SCwVqgu1cbTPORWcTyscxL
USBgBc/mR8vA226DYoyPWolbQgUQnX0f8AlYdPGXYuiGhwvNXLEezNBthgqwILuCIJ3p6uGaRACP
FKP35goY0yrdh53JCTkJH3OO5nQvi+J299zsEOhxXcd/rtqgZ7b7IDjds3KGcRWaVEoTrTiLFWTf
p9ZP6hVCpeaW3JjUQJeu1Em2VXdZAjpdyzoSzZZcM/2EFyI3Yvv5BaPLQrnsySvNiDjR2bN5Wqab
6HUAHXJI+v+zo19Kn7xAbboO6yI2VjFUZtRv3MPip+vvZjWVbeGxYBCVCeKF2THBQRMKzzI2gYxu
0+Muv2atFecTgZUapMO+8zUTw2DP40StmSagqyJKc+51KommXr/gh1Uuh21UeHbAxXEkYEaYAsjv
zojunk65chH9JhABgYTf+XYAuUo4gWtDhJT3a4dwqaGal8vfl3q3yBf7NG8GmkuHY0i6+m7GS/8J
RGVC2kfNOlUGaCx5c9RFk5MaD1vpxcAV88aeOS9rGIHfgH7EHmLhBiL/zODN31leRqXxJR+2YmOd
TpT/rBppCskRlhv0iKWfPV45zZa03Su4a/wOPeU4ZTXiMIS21N0nCznND0/AN9QHf9h4g26fI6aq
dgemNnNRaAgzlG5//8+tEnSR1dTtC8YzDAqgLb2KLTzfMDzHRdheMRISAw6X20X4xXkUMDdHXOYg
MPzJG16lEtjZBZS+azpDVr9G1EAILNucgU5yEo8XvSULObRyUbLDax8Kx/DC/05OUrWw7xQO4JmV
gbtxsYNh9VPvdR/dx5+9UqetxrLa98JbCimzyzOaJsYyuqKi0Wes5y6X5SL7P2NxMQIfvKObAC6E
52yCcj20wfqllk5wCnTSguPDVFiIpieyXnnWYAtqFiNLyOBbRnlKqesGXT8BiW5Ana4+0WHKqdN0
tec63xgSC8V4mVnEI6FwlishtIUVAi7cPOhtzrwHWzgzVdOdAtESL7zvvGR3+F/qFB278pHW8CUH
yaCv+CZk06LIzd2BV8WMLom/z7Hsk+NXVjhft63xW2+Xvbp3DmFjO6TnWbvYr5BDJjNOFjDQsIz7
NuAw++F6ardU8Kk/gAlCxn7557ocxyqSuXMjP5Uq5jbFf+sUNUbeY9gJGZIk9MiWFbl53+DDtGxC
Eus5tIOkybCY4Jo3zITdSyDNWsXQunpARnG5kgI6WMQa4t8rKGsR7Ix7GV8WcODAvHkV93mhiF0L
oe49i685523nVt/N+d9MYNCBY8aHuiMyIWQYpFFCB0ofcWdSGWT99fmhaxF0L53pNW96xYBSczp4
zCzfyOT5cIwxVctyuoAEQzqQMpMGCFvR8qkd37wqoyCnXMS2rbVI7NJ/y7aRZRUPlDnwu7PJHhAE
1XubVkoLAQyBoBu7VcEhm5ybWvy8heDeH5dqFulWTeszhPkpHBhkfZMUce3PyLHdHNv4qlbQUivA
rbDW01/GekDKsPedC2HPDOUOayhp2riobi41EB1dT7dTxix1g9blB/OrmFOMrHB3duq7T/kmotBj
tnhCeuPQhOybiNWJym23IAaWoBhV7TKz0kApDfRW+PcbXWGHuLBhbNdscxsW4vgP2zT+sN3XdshA
PLPCBMFad19Zi/XJ0VgnZr8b2E6sctQjvCVo68HvrJmuhcyQ/4T6Ym6za7cEMF7tMRjMrGCTFsfn
wYbni5YI9+NDdaQajvHPzphuPZpuEXO9dUcngJ19sdxz37D/H1uA5naUzJ4Ugt/XQ5F8K3cHONZu
uHyClX2P2CP8ePWCP8DiELmn5x17ABOfVaTkQqBNo99u6BE0MnJzrafqc5Vju+ntD2Umw5O0wjMw
YQ8ImFBnRNWg2QNI/ePcjBs64wDGbPuoHOQHUMrn2CXmpOkcExp1YH9YmK/zX6Qm0zoq+wqhjFaX
iTI2J0oDucQrAeQ/KnoIIXQNPNXxmoqi/1qM48Da28d1eFQ7sx4oHLvWiBNciyMdbiRgV7tE7sn4
BV2j3lEui7eEyoTMtK1lkfixPBrNsvYuK9ZXqNrBpEiJXa3Fk9IJSeXugnLZHFV3iKGOD/MJmMAn
/1k6f2ZmDlg4vxVi87OXzHWd/3h953YT9kcpo2bFI/jjyEEuIb+//poz1pYN61GaSV6dpuxPuyaL
uCmLEnUf/rgXzdO4OZt6mChJmrmOr8+/JEg/IAYc1JK51TzK0RSkpdp5XBAfoCvLYjFKG4Ddvo/r
Wp79alGyn7qDaqDuc4J9zvuYaElFKMDvDrKl20ykLiqpiLxsOEskoIdeP67QabBxvI6Pfn1x2nOw
6W1c2jn3KOYZ1FQbVuFbKmtYMJHW6lCvUXq37eXecYra819b7SKGSYH9gdibsFVhjUkBEeJ0+rKX
cSbxkmuih9dtWM4j9JS21zVso4gWu2PueYLmCZyiNxHyBz7Sq6ExPyVXhedrKBGo1+2n54p3BS2m
hM9ycCY5wqcVvyB/8/0pzQUIIJome19IaIDLSq7jKbjYKCOwt5hH2dO5HaG3yLZk3G62lA/74zLz
HnSQa6NtP8aMTaf5T6YL6KOlN3pdFQK+3TnfYUZAnFeM3j62DnVioeKD2yfg1rfJ7rBGRJzjzcE9
nfz3rPXZGunYVdCPjNCOnUH111gKtERnIS7rUuvZEzUF6hLussP99J8l6LIY7ZDv0z6l7DCVs6oP
abC8Gv1C+I0+qxpeRP+Pkwvcz7DcXc34J417/OBgE6NZU65xAOcq0w+rJbgVExsAk3eEXat81QCb
VUXUFE/UQ0xZKFjL1w5rV6wUqDEyrVTaaRzN3oYdAkw5uZw6smsWjWjZdMzzVhy8ccE6JhGAhRyJ
WxEZDGpI97hl6AGftSpA92cXepRrk5hzboZ67T3LH4RnjoKMYNe3FzAndnOQAg+5TkWHxkrxjcD1
pPL1Q6YKGbQXCe+E31zl7th1AZA0tQjM9qY1VitvU6jZQDiq16lhLgjFZZb8FUSK1yFGlIPiA3/K
rlalty0pWIjgFSH94z2WrYHHK5rpmlnR4xrOoFoh2zAXUdsGNQ4bcCRngube4kigkot+kBT05HWF
8heEscjrgvaB/tVdnKuiMM3uF7QJwd4ppgSxa+xE9AQ9tDruvhxWnIP2IhzZoNjiFTMfUKYw77fn
myinHSdbcgrUm5xM0B30SzUxItn08obGaWfF9fRX0Qv1Gbn9/EZAxsIVzOVWHQmluZ4TDFeISgfP
w6v0v0yCydZfmC5Z7BZNmv48Ix3g7ODFo5e3jxWSu+X1Ngw3hHYw/RAfabwq3pgaMsizH7WN5or2
KW0KdHaMGfdypS8JSmUtqny+1v/rydViBHSoWPf1U687+szbYZG3NWsVA3NCsCHUM8W/XgZmqJow
Zcythacq9xopmrbnkQLh9A1Xmisy4HRPXotgvuyYLjYUNPM3YTIG1C1hfvU/jM7h7ss6fvS33YtE
eSThdpj2+II6swSoZoxDVvMCU2sWVyT54epsqVCuI4gmXygcylLDyi03SrcCxjPBtolRSkMR7U29
4BuXe6pWu7r+NefwxQ5rbKaHMUtOB9BOoW4pKNIugzWnO41wCv5A3zO9hejqUkYK5/44NaymJGOf
zzBUVoRPK1CMRSP5PZBc8y2VedsqY1MXQR5XEdtI2u+8IDBquwkevyZNPX+MWQXvCvd9kcTByXof
6F3rFeC5wZ9osxUQU2a58LyKf3B+NsgG1IH8Zogd10/rdys98gygqr22MqUiKMcppnd+HyrI1PVK
lMD6tsS23v0UZ8rGlGqtu84cIHigBpVidxl5MxsTVr9EGq1LxKv1vlxhJU0tuyZOEWhyRjszdIuz
0xnExLpFOt5oRCOUGJMJdaVr3rrBz06UcePo3/bUy2nWHQT7HVOVjmm9gIlFP61hrbon1F40YP0l
zkT5LUa5UUZWSiQaL4JSkICNBEQquYkm1/0N8vanM/96gStpZ6csWZr8fTN1iIZhDUtEl15tPkwe
0TzFlv4yculOPVTVRJppyNUCD8cIzieQGS3911Ef3PD+w1Jzob1b8ML/G7sAVLmMW2NB4HZ2wkP5
W4DdcXdsr5lCzBSuJj3oCzGUN7PX1ept2kcFFvmdG9EfJddf6ytSW1o7WGXSGtzE+kD/0d28gq3a
6xlMKM3e6sWb3tgC9b927pXGaywn+w84URux2lMhTCG+JYRDK17aYF4kSRF5Fqt+Qc1e1SQHnjQR
MQKy4k3Jzsn9ek+mAmh0TRKytdOihZ+QyT2bIU7yttLoVm7HKNtmT1GlxhRZDYetlP/KR8yzxeZi
X8CwztGqpEPfMxUWZc9Q0wThAmtxGvmiWsxFWUKxLy9VNe2boy75hN3oEZEPeg3yM+etfEACk8/A
sQDaaY7psVS+FqOGW7ar759Fn+cevOOsMOUcKXsA1n7OTJLHPLl7cH74rl1jN6/pNO8eW9TyMnWi
TjaIwXqfdSjOKSxHT9RneCEt/UWomIqEm4AK307yk6BuuDYzMNIUZu3CTl9msnvJs+SMVR1bbu1p
RE3S4YKWFPk1Wydi3M/RQokRJpLoMnV0HPaTmud7DxaK550ZbyaOyVEAugFBSp+79UtU6SiD8wpd
S1d56IAin26CUKrBEYhi/oeF1UeoG+5m+OUV4zPVEdcyDaQmfRedSW3vTnxDc72sBFhY6xQCTZkr
791FnVbGTDuFPt4QwDJpK+un911objo/Ju5y/ACj5pAtBQhsoxAC6WRjaoaNLfY3DsmyoNXaFPbv
KD5GtlrXqAcEm4UHIVY+qyVD8LnoGuObWEBfJZ4kDKbzMLq3Pf6Bydz/s4TmqTS1Uh+y8lmDe8kE
YWbseqNM6IrDhnyJSUtqGPzDbUkbt4smtimA5rW87wWDgbawUvrtkLERBmUYUG6Qm0xgfxjsn9rE
gLfi6VzR/ASDus7Wclsjn1ZS30NcuGZZss6qinb18FO7r5dLF98PUvRXYt3uim+PS7NQIzftfvzA
aHN2Ke5gR5q/+2fafeYFbsbkHJqLmlqBDRMLeuGlskBjPhb0CztZ/zJJHa5jGvZRpNlllz9GnYq3
/ZXeBcxv6Le4sKqkDlge0kydxGkqBJyuHk0rBpW2ja6EcpI4lMx2tmw8RtCzwgysrwKMQzRD4tWn
NqYImspKoGUM0VNQcXHQbwDwm/leNvfzDKWxdL9kffDTyjprqrLjwoQvfOxd3mqkx5Zpk9OY84bE
UaxC4333E4dGNgDlmqy9LA7eaApexhCqxSYvT88CH4OVSCYX1qtqGPAL/kcKKq1N3tQ0Dhh0r6wc
L1aQ0SLb3gm/Jw/xpHA8zpU+jeG993WWok3YN2YOHnWqZu1vcVlmt1d0Gll9LYGAZ1Etv5MhlZdL
y7vxyz009PQlUxpEN2suXLDkwdemDhe2WY6WtWpZ9XuE9KNfX3yY5ndYjW8FSkfQzGUkj6pg9myG
OB2Io4vvylTP26+2pyayYzvIptHNV+E8MFbqYsJ6R2m3i+SuVhdYtEHhQj8gLraPcibJnYtOFAnn
HWsdUBMhyAy4GPjafbKzLw7XMST3l6d7/qzangUxEHwaodRDzugwJT0W/ADbVJRqWCaDZyGsDhWG
wr8jsy+yg4MuHnZ2U6HaqoU9CFkDpmLHy1Kz3iJr+Ss2QyyDrdwC8rVRB7Ef3r5ViQShlei/VajO
8JxtHMS9IK7mpWZBCONNAnHDztr8LOjva3GXefLOy2IbaG0onUq+uJxJBGdnqSgvPBfdLY1zatzZ
CGMOdmEeDu2dy3lZPWKm4W5lodAFVP6LovzWSLCWMFMhlYnfpid2n2VEunT3NKb+AOTCTQrtcPAj
SeisqgCpT0twqnotB3qxioAYKiXQQtFsUGZ6pv9aBhlQfXETUKKQevh3B11Vhw040PxS+vajro4j
GN9jCxBd33GXDUi+HW4D41JvU6HS2OUP1EWjgstHPtqehJkG6zPYzJN9s9QnRc4bs+WOmembsjpQ
S0mMaAq+RT/qiaP1Ah2MSZqzydFeIHGU0aCJtEMw0ciSYTxzTxguVxdLha65PGUFqfx2f2DLgJ9e
ngpn8APM6eIhS1xGOyL1/bhb0ZT32VBk3ZcX/fGReL4o5FKvsLfzJVOuBCjjQRuVGQNqifcPPDHT
1ItM3sCgw00BIaiYWYRnTxJ5yDIyJ9a8871oTMNnG8Fqi7darpZU04lZ5vPIsbBUiLrbumbXVSsw
orsq4rEdUr6ifzuA1Ooup+MPnPN6KSx/BE6oOsmOvWek2gxZCy1J7oHaUu83rUT5GexEJaI3qx2w
wE8Ccn94jscoC/VsfF+Lk8q/khijZE7PaEdhp/IlVDu4Lbtvs+wqL/AkibRUOrureQ8z5tS1j+TO
T8w5feJlU3kXkkprhK6/VAdeJ9Q9UeaXT0dCJQkfYpwnZ11SG9hkqwz5rRRlp+svY5WZJoBPeJxe
6hGtfVN3aRmsZnqsqWMwwkb4a5t7gqmiMiut2vj3HRuWPOlcc2jCHprRM6h8+XxQKnYMOHmSJgJ1
AsVYMr+uSgQedmWl9/54Vtz+tzN5pzFnnlBzf+5GBlsY9b03O2oupAz2gpBVY9aRIvgDbRi0aGon
vtgr9kCNt6OA7pv6w3xnm3YTVxU7yOMp76sfImxzetStGUNk8SgZ+D6lQYeDziOcKVtCt/deM6Xs
eFpNA4rQiRnHaSRI6OxgSMMK3LFezW/3UaVxYyFZSQHrxxfCaX5cWj2zPUvZQwkRTZbpL8RIc1T+
RjvV14Vlnduuzu7grZhCwBbYdfcnEEcE8E4dZ/AenadjXtSJ3C1N9UnXp6vKneBaHQOICBSNt7tx
jEQJ9kddX+HGOiKZ+oZhUO1Lm0I/YD+bRYpgSUncRwhGE2aaFaH5J5k4emtp5g8D9vaB1KqYypKS
xzp/67EJ21ZMZ4BFS93epQ+Cnwm7lisK/9MI1mdACthAjTpmxU67tv5MyRX/MFm1zO22QtzWW8g6
lPFoOuuHEtCP3PPL0MqPbcd/eRbRbh1DPzeaK3+cWrwYnTdO6W04sjaMimSMCMDG/soHRk3+h+N6
t8xTlyo6Gq39to8K8iK6FFiFAeGAMRXCEb0ld3abGJM6etvifUDyum3nZJQpvgjCXywEwMy0AKxX
IzemRpeizqB7M9um4UPx8u+oBofgcr8ht7NmuDeRTEp/g0bFP28PNSMVJDS168t0YJ+kXO6w96ki
CUsB/FrMgouHOIMcib0n3Rsg/QI86Ksjy52GT+bRbug7VEZRkA1kn+DXzDeHCIaMKNg1BxWEn05Q
rKDV7m8aNGji3DkqoBhTOEBvo9xaK0OaIylhG+vrXLmVUjNFslgcD3al1bZ7x/UxlJc+zd/N1+C1
Gby/sMmcwkieXI5JdLmp/z/XSDzuIbVcKZGgBiAaja3GyPVODraBaRLGZNQNutZx73dnfzyi5Yms
HO+/h9QcYt6a+6910+JbiCRSVr8XdsjBAOMfVDqp0RS9v+mZqswZNvb8JREVLQYi9POroabVQ2PP
fPE4OZdw3Sf0yMk6VnpljBoKBYbqQFnqQ3qTBWqByJDUDrilGGpnZZ4P9DCe0dYsK0x4KXKp4iX2
i6tS/BX3EJNgiqTVX26t3853w4iOOzXaZl0cAl/ncmHcePjavc6pvc9m4TpT0TWn8+xJqioD8Kt8
wBpT6xinf0rqm0iXhTV9iDCtfnPdMNkQLT+vzBHsF9oCVnX0sFqNTtHVb0qwEXOJ1df9JoOxweiO
ZKmC/WKHDXK+HIYtB19g4nBU6iR4T8YH9yiDkiH10ko465wmkP/hPo9adjQd6LFf1hcc6dV3AgHz
ssbhaEe6zO7JboQHhc4CXyOq0Ucqydle8SRs1Qkg8I2BV12XMkjBRSSKc2h1a+H50lCsgjXMPN4F
12ybRd9SPP2hBonkutAF9fBr6KLQhOoDyeJoF9vlN1OC89DB1oEdvtoZRwRohf/aAspUT6zjVJYf
v8CxGWjPoBZKgvxw8Ub6ooys6+uVJbA2MLRqUlLtsClrmmUqWs8cmSuSCZKHjKOszvHGVVbOi+F7
yajKc3RY5YvBhkj0lm07t8XkAWNTPr/K7v9EjU8bMhj2ABKsq5V+1b2EZLSkIBOBKC/L9Gtc7nnV
dKLJJQvinmPcQQby3Y5bSEPHq3wppX9b5I9TDigoo3QuFAYf/I8a1svHq8uAP+R7DLmpx5Vnojvj
TK2eYT6Z7l3kW8Yb73lHTITxU6u5AfXNgK3DeZ8zshP/nZ4xAJXfkOKir8YBOgmVF724/cj4LZqB
YkobOf2AHGBnWZDioYvcnfxy90oRWOZNlz5YPOyxf6PwFlUWE7ihVxylV57oqGz1VRcJ8MJzbHQ7
o1TXGOTq2oGYyyuSnoExyGALCKh1PE69Q6WnHU/a1cLBDsAYVSJ/ODEZWQeHt5dw/40coMtZrL8V
Ru5HHfPskjhLJkiIPAHMr66SfXbjntUI5Srs8bp8+fec8Z1Q6xBCsZF4TofTVqWK0T3yEQyG3Vj5
e8rnvhBR1+wn3ePM1mUanZn2xu9e0vDeB0cv4gpDoumDbcrPUGlF8sfGxh3niY/6essdKsxplH/B
kIfeNxDgWJkV129i0ogf2VaPbjMAqepp9xFokbzsbl0vKxsK12U1IXmR0MZWlUC2zTbIyjylQLQc
4e6SHYw+TZgQKYhb2EgX3DvfS3QaAuAExq8d2nY1hh891P04w+N5RLdmW5cLuGrxKQpvlIIvBqGD
pGP9fcSgCk9Zik+jUdiiNlLZOm0y5O5rFBVUpbjsHMuTtK4ELxaNzwZzyhkm/uOTiLAUdjiAtEyN
2cpAYGdp0T/7RZCQwFRo+XhutFBtYFRymyGsCMlXnBLzQ84o1VMQxAP7MF27bYZ+ylIv2b7zFfYK
6rCwbayKNHsjbijF647/XiZhvLivQF4hTqXG7yV0/EF5Aho7q9ZLH6GeErCDGAReezx1TprOVdyB
xc4Zo5dupHsbt3eNt/2jIvglD4Hh6hVDybLCPnttb5D2pJOdOXYR6vPAi6aLO8pl5Rrv8IF0Lb90
8HKVGrCx8wTifeIQ4mEebA1iW0FrmcF7DvGT1+GHmYOpJ3Jv2pSo6mk8Ez5wqWzdSeQrWuImyTcO
g10kMm4P/dhu0kD+gj4dp5xeiZkf0QTNLfx/GZAMXFfg7c4qiDmlKUcQ619jQv7xf717mQOvGKyg
Ae9CPCPLC8qhMALaY1U7kcUvvVvMLaLAqoCKPmDlSrjlvmECUZR/IpGVzY438Eh/o8G0kS2LA9PI
RDNLuURGvr1MEG3PFL9sONjbrmvNUH7sIUDScD6aAudCwdLoU1qaQAIqdVuglxYREN/qbKPUmers
p0eRztQFy0ukgff5d2VLut2FhXB7T1aobW4EqVOsHXIL1qnl3ymk9Trc1aAZUAP7tKxL232HwfN3
utVAjfqQ3vEWCsk/tSiXol0LazCjCPchsEDWb+lI1XqDGOFr2GhzdkxeM5djbHOHA2MQD/ymJQwE
r9lE8/h24wYTxwudTHZnfzhjWZyZG6pTo33KhOQN+EyBUWMAw00OSU5mUbLgCPeJawTCVXDhIT8j
zh0C67z3HuYQRAvY8NBLM2Vw2+xnV8g608e/QZTqgIwaDvdiKoe/oPFpKIInrn+l0F5yM+R93i13
CE+s8LuxfNunU7IUi0wn/w10/UDsFARkcqM3N7u40OBAtsfrehm2CpiasS6czLSRW4M+jsT3M2Fl
aN3v9mf/J+P0gKp5I1gQ5y7hYFZHR3RGeYODNhudtIDkARvDWxGc7PSO1pvr00AGNcdztk4l6xZn
xrMbQldvwLikcf971cXjI/jYOxpXrSSM1g0zvS48fYgeu6ygBwlqlr6BSVToKehV/6BDHrSYauM7
oOScUVfxKzZBz135RaoyvpZ1Ep3ZwyYIiDbIK5MDqOI4f3pvGdMCYdahs6FnFY/ULrGA4jy6UwbT
WhMHAoIPLpULlHiZ3IOirfCTniv6VBrI5eXcr/okW+tWoVjo8oXS7XqZv/hFVi+yG4z4kKHCfT7z
7NQggHGncVMn7U0LZC/KqZskp6VgAc7wAM9KHvvm8dcY2HHgc2yH2SlR5KGYATzE8F6VNLTF2eyj
UMQnDbC80HA/aMqd92wvPlDZVKbjy9SYD5Us4wlw72C8bhwj7NB/LXsKU2wTx/otBjt0mGKlJrmk
sOfAotfb1OyOf2k9BeSsS7nWPhRRFZa/AevT2ND3QRKBA6lmwlaFESkXDTEsMWuarliEr+xGYPiX
ck4lwI6fJEDqvTlXgkLQx2+OmbTg6mi0ELV+tN1Y8DPkDV7tTSA4r3G3R//gjMTt5k6CV6mlZmQE
mtgf1b58AoI65LCnfWbPYLGLe7POaLCUB2ZOSI8h26JSPTysVcty7ponvLSvyeTNQ6vxnDR71ILv
9mf7XZ3VU65ya5xizAZJEfQKGxftLj41PZ7nt40P+kEnT/y/OsUTejBlqgYVgs7S1ZCUPOg6yGax
mfhG4j81c1HouAhvV62BG4JuOFMJP/0dyF20PibEjCgYlxB/z4rTCB8WkmM3xiV9LtHYMsydXwqR
K38pweuHornbI6xmEOFwvkwWJBHgmre+tmzXNzwLqAd4LGZaZP0r6I0mlg5pMhVQ4If2ELqIq5eY
SXmMb16IVIl2Xi9JVIJj4yX1DkYNiCwcjsGAVgVhAiSinMdj5kVvywKtjA5ChXZdrqPNLEQu5WLU
Mdb07hcu2DP4elbjWdWlDGVN5W6cU1EcGklfh4tfKko8L4FXwx5R+kDqJPk/gT34U9UErsymDcfe
YrZtdLiQdNE7pt+qZidsgvvIlU5LqZ2oAcrHLhTt4tFr/FzkfWQNPRRTUy5FHSDH3mvxJ7fjVNHF
nZcyxZtS3MKD9nTU7ytuKQ2Rdt3/GpqE/lTeb/bEn465QXm7Ay+S7HKFExB9kaYFJtrlrQJOKSHE
CWVe1wcW19bvTrENeTSs942pp4g6BWQ2vjRSK4IaSoG8Q4R6r1PI1ezSpyBRoxpPg4OnVEIRySn7
JAsWhxHZkM551CzhzIyBVZlvoNaStUBkPn476A9SuthYRcfwrIIFbK3jefa3bVK+lefwmk3A1clv
qBkMQLFn97Qe4KAZOWdv+dMf/A+mz+AfxGWiJXEzKJGY6TWN5xmZtK6UN7SeOXZhc6/ka+UFScOn
I9ESp2LTD+njntfI6aoecI0PvuvOHrMrqhgjFVDwoU5F2x0veBsL6po2FBl1CtXvZzUHq7a8Qv/c
OJyiWDsCs8qWhtKTvQ7AnPqENQbz/u5VD17bMerklprxSrxCRtxCE4nI3eR9MtD7YFDw1Kn8h7Bb
VPmfjGuvrXmTSCYk+0VLkael3cbOKzuqA24tlsnPAOoYEN+HjNCpO9oYzJPrzk5s8uaG71WkpiU8
br0km59euaCZmSxn0Eu/FRQz3qwxh8u+E5JPBI89sMtl7ezoSytFCVNX+3ZQHrsxvCpj8YykucwI
siV6+6vhykKIWbyK
`protect end_protected
