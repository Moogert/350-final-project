-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tczflSz9lVQujNj+sIaVr+uK1N1zIr9o0I8xDhcaCT96QTDPCRL+0RSUM8WZgsShZn9bCiVZHFLI
KdY3h8DLO7SDzEQYpkVnORam/ml32XymTf32FS/YpcjLC7K8uhJXCnMzlDfw8r1v0/VFyn9VrUlr
Gne5GolpMI3KJxoXfEdgok7ECTGNF4TuaV07QR+5Qd4Hu0dyrblgqCjhBlVwu+v0AKWX4Ydnm1FN
+LDZoUV2i7HTh3q9sfSep5586o3cKsLEUq3GuefUmc9H3JeZ2pxG6bqY8cbIbugoNvKheGnMsw1N
6jS53Mc7PTNNrt4VQajAJdOVW2V8PoLVMhN2Mw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
ZC+6aR8NoFFlItGTc53gthpeRU0XPf8YSV8Kf6o6LZoHvZ2FY33zNlZ7+F1fbtfCIJlKHKf+U+y2
AB320DsMoulyyVs5zASWx5oWAy0UWwrZOUoZr/E23Ym+qcv46Q6kfkCfkVjk9CmAojZJ+Hn+MbGz
SbqXma2kNhSWNjMJB9Ldrj5/Cqvn080G4Qz7Y7TPkuHoD1YyYezhABnxH0zcmOfEPbiLdWYbjOaG
lIptMQHk1sRqVn2xv1dyNMMEtOYUCA6k7QGXTSxASvPfPJpXKQVEAb0XQdeX32vv/V2+zB9fGNml
8YXBx9MGGAvriVNn51fQY/lpfSV8h0FdF4b0QBKu8hprvHfQ9H3DxDD7HF7B3zTvnowYyb7XSoZ1
rza7EVPcvmgypQcrE4C5GRE9faODfK2h2GHG/LdOIYDiB97KTEdXzv9T19FySgnkFygiwawpcPpI
7j6SaRgi7ZKZaAAkUxOoNujrCH8xVMgCNak5r9n/kW2VFf+YTzohgwTgPWLc/UC2f4Aw3aIYx8HG
teWVC82ld8TON3uR+bs5f7xcueIFdRxXGDIRLhdCWGDQIGV80fOKUJSlsyI909piHQ/9voGFz4LI
j5SYsl8cz+qQ7JPOoN/ySTAc0IQapP/oD6QRc8h/j/EtscNGq8lZHUc699kWaG/3BPSLaYayUTVW
0SjrEpX0WuhgDwdzjg3zLwgKkfumES/O/sHj1S1lHSS9wIyC4rY/KBVRgo2aolFgqkLtxIlQpEAQ
H0WafNi30f8SLUdO4EkrgfiWFp0NAjFc/MSN901fqBLWkWhrZXStCwvyGjx1JaOIJgovs+vUWUms
+2p7SVb9JEf0Gc2YdY7iHXsuTG0pONGuHkcFvG8WG/7CBejbqn6tuMD8NJAjxkdRzjTHORpBt1Cs
iZhLQTjCWY8xrLKa/0/EEGoQwZPTtODB/gyofUKaM7mmuJ+6kMKwe5WUDin1XtqhwURoLh7g9OLB
izZjMV9z92KAliJjL5IKxcx5N11t9lVTMac/E1+lhE06vvr+8PBSZewRzoOKIqbGdE+WT+moEMJK
PiloQtfE1HNK7iSA5I2/6m+VLBWsqSoT0kwp2d8tFLtt7ZE9yFFkOV4LD3EDHYWelclehavr/uTL
ckR51CwtJeyuKMrdkvmOKcirt/769Mi7ukyrQY8lqPp6oncyr++owxyT5GWb6GB/rWzxgsUYyqRw
FaTxj9WsLjM0pzeRxXJCM4H3eOcfyzcWGQXuBC0/vST5R8nHg4yeT+cL7lVAGBFNZtvW4IXFDUEm
18RpbdiNoBTnykX9hAJpK9lK8G1w48FLG6kVxrWp8oCIxUfzJEpB2cdG+iIQ3xVkf+uWZ9ae0PYN
Ijun7oU8dzVMLuAHp8v5aYQvllHDj78orDye5E5D3M1RSoYVcbDwS0kTbztHgJgPuLBEBNLEtGM/
DPaG9eUsbL4iWn7KaLiP+nRhXhTvrwW6J9vVrqZAFJjhXKAfDPNQf3VbXW8M+nmj60Cqyu6tIn20
2cLbNLPPB3hHRfA87CqGyJ0UEnbLz6KdDNRB+S4SFX14/kuPrVYidPP1lbN1Kg07pGhJeDHTrm8/
62I2E80f++v6+af8Dw6phHqkUutKtHh/EU95NcnDlJOPi73GEH+QdA8y+Aap12DmOC1cqiqiTnWK
kGb2PDI7sFNRe61BtY9AjDNimtoAPeCETcE/djRiyIlgmeBP5Q2o4tPSxjepAqSymmDs+oBcERR2
1c4FhDbeq5HqUJtSlvCxlCygAlTvX37iThHNadfSfyqFUcVpO8DVM77+UHjYTSbgYE1KJryvrMAv
TWPfWHPiFu6u9Y2fKTrRJ/GGWOPiQmT7dhcBL3OTe/9HQXVmeTGYafUSHrTPwAwDB+Nqe0+GCiNX
Vie217VMNzkBga3tHpZu/HTT+qzKNfKofaUy2dWwUT5IZ4+lrN5MJt7qG/big2/hArSi8NCj27KI
Nj16anyaSNZNPVEZfV2BnzuM/VegcDDXsR3iAsq8UXwbISxKwRdViCSD43H+dtzsYPUP8tL4agY5
0e6r7bSZFz9EU6/83hExIBxtcGuSm0TWiVNVVBqhTY+BI2WhJnhaOvXOz2WnE+doIPBOUMoW4z/7
+TNQ7hrDBQawc4L3d2r+FW3e4pjt6yeVXftf/bm9y360DIXH+R30r0eut+et0q8Gds8tmDPYASLx
KoTRgaHejs5fRfnjviNKpuWev/B3LnQpFB3aLi1jmsACXLdaGG9TyYODN+brYn6dEDt8GJprzZMS
esAsfb/aNG3kbzBBZa8IrgXob2LXQw+AwgfnX2LPgqvj5ALZDKAiSwlJq/0bFK+uzVnEz35BYAeg
36NkDuZYA9r5at2WTdKJ56aSoAob5dyskUQ5mOSGVgI67msL0BO9C/Ortz2kiyuJ7aPBIzraSYxr
+uGgCJ/Wje0Y8WLHcCsSkaCv4JIk7OuaKsax29Y0sn3u/0ywXVMPUsLOAxSB2FWJjfbXSYy2IW/L
OIZRG8xaFk3yNBGqQEZm2dYl8IfsZ7dkj2s3gX/Qwso62lyNP2P/vPuJ8FphTvVT5JQgT3bVQndo
nlyLjOy2oCyNBXiZqm9NIwRcgyAti/h2TjSpsm1XtZJxErqF+JfyRws99O9Bb15VtEyNmpNQkUB2
JaZumbyFuoiFOxTobPw45Qsc5H1i5AoTTNhNjSzcGQg/uRfMcSWvyC0EuCsnBGbbVGjap1FjQf4X
GjBmO3b8SdCIn0SVKiePo2mhGO2yGEDBzJZCspnNELf3cOH3QEAhKq8RyZddfZjARJOvkRZ4vdxW
NrEInQyRmfgZkuIJslQrkCGCwNTzG10+3JP2bkZ8RZF25o0NVAkHwxGPs1jxKHzUiwp3XVC/wQaO
B/CRH7p0dDKuAx1xk2E83kGY2i+LdamcydlcitzrweWiFPuL/qIO+CQDSLZpg+m37cWMxodtyC82
2g71dyKZDW6Ten2usC8I01mb7tJuAoTFNlaxekO6Ig9lRERJL/Dyl9B+4kxkmVw/RynNtCXIhPPq
JzdSaxGsFC01I+/r+fcshXSY9hedWoDZP+YW9g7KDUaXSsbg7e8z1uxskI+SSaRhwtw1WnMcKXTe
vVtoziajj3iBMpW5zSBedw9x9y2mritwpNCpD+WnC/Jb8AmhQxOBvhalXAvKJq3vibFZfng1+n8Y
siv5ufUH1ggUE9F0ICbAbCuvKdnIAZ/rPQUEw/4cS5zlXEgO1NFoObKZzK8xanb/bA1BwSAjOGIJ
G45/A6TALlLhNuR+Ib49mnbEatY5NyUsKM41LLRmhE8ENd3e0p8i7R0uF1GUO1mhWHimz9xPKuVs
3+pwScYZOX4J9+ATI/zcUWF88Nq1tta5Bj5+M/sQszVvOW5bWqkzKrNSATNQvj2lvzY2/ucY1tDT
W4gGN+U9KI8pQJoZQUDGnsOLtHPCFjnGi9z62vhlwvv9Am7GRfKq5O2EaKy/9YNa/LxTC4EsP7hL
eb6NzPmi3paMYpw5ZZgRSe/Oj+wCGhCflu8xwt7w+X3lhWlR6DS3GPcjMXg9iDZJO/cSV36Lme1b
34iipCaiSR3GBNjjQyH5dMkdAZkMB8u27NQ8jY3l+8mpvz5OXzsjkLaJ4CLzaPvnwv319B6tHua4
jrmU39/EbEJgzqTjnhs20zuhR9A/FnL1qBp+DIdRYU3dVw9InTJbrxfuUBpxhx74J0afbNKDcL+y
OV1dG96a3keDWUP18ZnZKLyB2tfiViecK4FxC6gHcLV9rQQhPA8QQzTIlUjSnNU+FayPt+xvj0xW
H2EMO9sZTVUY20Cq+Si1UKZDUZUqmg03qwl9JSDAzQSpB9FK0VSUZD2FxP1RA/pBVDwsysURn/QM
rF5xcuAmKZyyPJSEjU7PzZjTfLVvuoqbaPth6wRxWv6MhX2Rpr9ZjSQJkvkVfX4CN+9hiCP5O5WU
A0N64C0BTIPQhYM2BY2B0sTx0q8GammCs8czIaU06e8FGitZsqtkzy0nePfpI1HmNLcLSaONJvPB
ws/n8QBUSnxy3kp4wSK4O0wtmHQN5lxKwX7qmpCSefuVZigFC8gkV/h6ZIagDYV01DQBvZkGxzCd
fCKAAH0GE+E+vCpaMLcH8iYfb2VoibhJ+WFSZ8PErNHxwcJnX+AbD3WTFaiuTY+79Z8690w9QnMR
uFa5dwuzRJsdCV02BsywbOeyW7qG1mffAGIpb0zpQn2PiWOOK8sE52kwJ8DPIKFiuYaM70T/v6H/
zE5/uOgMYCk5nqmhOq9fp4IxSPVSRLDblY6h0g3XlXFebPFBh4+ylzD532zkez2BS1DH4detdJyz
hRLnlHucWcijoTSewESByrj0oUWT4PESVWoST6UtdN49F2quOpGdsFubuHjYFfBV8PPVt8T7zoRl
Wz82xwIN7PW2Li0bLqUGBs+oMFoMJFSUk/qK0yMD7jBdOBGPVZUrSZnZydM105FpFtYncTIWenQp
PxBaVGx93ELujq7Mv36MqAnR0rNjU+nBCVvc4oSHott5qGUuRpzqgQp99zUsDVZXPRLjvTbteFAr
caf3EUFMbVEYY7ckv0KlJf5XX65b4iM1tes4fo73XYEUFr6WKefPhxftnlMdTR4j1eZClxik0m8o
TST4DyyTdMDYDZHWFIfxpWTL7m6yLIc+965CAElhnUfg7Pgm3/7MdDw16zp5qg1BqvsFoz1cFflO
n6lc+in2h/6UgAkRbdNfz93Dj54f8huyu+VSC/XP9yalDRftRtmT6iqTJj9h0JpzVUkyKhR+6/B2
MLsXYYnjExv3+xu7RCPAFpkhshS9nVh2zKKJXHlE8q6ujOIhwVQPTNe6YFrBJOp9p/yfIwY1xs7v
t2qfr+eKKDhbqXfi134IbwrJRcqvD5dVjT1F1y8NY7MV05QWanP9iG6bw4Ipwt/3LgZI5bIo3HNX
z7PezjaDNUeTqGQEAA1hAtB5pM54CF2bkYKskz34o6hHLi6+op4HSK/VHB79/DjYl4zf7+gOPHVn
D3ymfh71Ti+wVSYzAGKrgG/HRVX9nXg4GqnwkvQK5w1tZZypRcFlpoSJEIjga3U1GFzI8PgW+FSd
pHYBkCXLytTN5/jYC56uVxtA9wk1rplEXuuJI/qmKSXTn1WKXQ69KjElaW8/XEoYbwFe9RJ6oRcp
ROj/dZZyrDDGyWQXA3Kue7Kx3g7TBhJHP3EV1sdGRlmD777g+a6PSVCevcSeHuhbke1txtpu5og1
1C6HMmsAH56/qG7Q9/LTdpapCk37BpcBal3F+MK9hmp7pHLL2YkmpqrPGHdto0VVg1zfQJauCaXQ
HYOCOh74rOCBLORXx4zm6e5/+cL5bfI9uSkarVjT6oNlORua+cgVCixXh+YjdyRWlr0PGdb8ekB1
lL9ghBIscYgGYycEgkx75n16pfeZZy4rksOS6flY7Usj7vsat2s6fxgkwiikikiUfQeyL2zfds+L
plCaZY85Xftn+Ybj+QYOW2ZMaE7waOwciVOrjG6wOX0j8VSJMXJX370otP1HUXI8lphmpOfeJRAD
HHJ0ciuRjkswoH+UsJQpgPKBnf+uZTpyT565lZYRKWEM/FQaW82y9n78ORGlu1enlBc1JNPQjobT
jGYFOq0QxF0BVqlaZdYsgxZQ8CkgRKKJi0jmlwoNlbiG8X5yPb1yACkczqNBGLmVN84yhyO+zT6Y
9MR/igufsDr4VwlIXajqsjpAEkPMbMgTiVHVQ/9m0ewqj/6lWLWmEZuiC2r92g9IYSkvCNCT9+x+
AQhZ+7+CIFHoBdeUNyOUpznlNHgQIjcwvQ8Cwvt+a3MLUAUWdEQnzka4D7hmD0TM1dcRlQIq24CQ
zHc7u2xCLzR9NR+tVuz8OhQXutacsEysfs/XByERXaTrRBeVudoGihBoeP7v3iK6PEQHelTHM9BX
TjBQIiKhjtypIR4aduldof8X/aLO3i6rSVasdKxWpZqKYtUFCQgFwrYuefoDIbSsyQOq+BbCXd7E
zgBYJcqAF7JvMYB04DPFi505qWpmRIPcX2tlvxzS9H8VnN4A4HFPvqjYTJReIRKw/hPX+MA9lHdo
YNQ5GEK/t51eDm5VT0ezu23HCeOaynHETaOXVQftDCoBou+DxaTljSgI9qB7o1lyCVu2CNfVbEV3
9EjY6MunI9GgogVkILdXx/qJ+bJVjehknW+RSCHshGqBfpH/u584zgpN4M9AfWKABekiXy+onGGO
rkZuyY+88CWv8y6kw0Wy2Hbva+Co9ph7lT72olNf7W9rerk0viyB2cwYU2ald7cj32kdxk1pNOha
WnXbwziVyCYNmkuN8cicp3crLIFglj/6ptqvg2frh2RTwx6NIu+U8CnmpY1TyUVKPESQTjwnBN7E
julyPbeNpluAu+F3CPTJ82kKDLtjcw3IDcr9WUZ2IwlTTfKTtg2Xg2llUKPVh67MzwgX1Oe5w+vW
PnEeCHIpyFyMoVkjWqTXCAaEGIF4aZwhr86yR55Wa+AGHwLrzmMAnlUaCNwk5shyi5KLbVvZx4TY
fdi47NysyxSubqrR0THXhxk/9Y3W6yE2zDnaYB/BvjIrQisODJIySJoOJ6PP5pvSNjEsvTDg+rz7
EbijU9D/18rpXuSfh2X2hnE1uzkUlPkaqJtjatWwICaoEIbYUWA/GjnKq6CfxWH7ngOhYs+Fo4dA
ytsuFnFxU4dgf9+zDEFiRBFvlBgM4L+bwkWjQY8VFbQUv9gdJMGkWztrqrjsPJeDvucx4+KRADfC
/dAnVbN7JXQeMMvykEsQF+s4p5IGUQqrbzcBumQesbqK++c0wCxJobvWyT648Q13+ClfV5oLgzO1
lPhFwj8tQzSuK0CPj7rSed5aGzzJ0KWv7sY9iZhw6s7CuoRQifB2Gz0DKmAJIQinvdCDh4w7nKyl
krlwW2ZchrkdGDAvTiWsk0rPxtx4B6D58iwIfVgCJjVmZVGUgveFVHdB68kfHPRM3m/WxkUnoSpj
rmFtVlyhJcfh2y8KHeWZk1s8LM+10hwRRvoxmIMq/3Wi7KcMyqlgPW/MTiyNnFXgAk9iG1fPLv0m
H0CtFd3How0IV2g6Sp/ldC4Dwy8avGBdmJVowVYKYctnP4keRenf0XdzVvGaHoxT9G4z2QCEii9+
6Rm7n+uxHvAHYN9MbfPF7sglw8Lw53y1nmrhV/n+ysRQ6FjsmNiU4gG3DzxNKKpAz9IPIhr/r2Bn
6U60kd9oGK3ijqj+bQqp6A0QZZdTSzchoS/GHb1ZagP9u0M62UmenQk+ro97di9JEhYPtLHt/aDs
RHkGG3+enZQKXujB8FwIECDwafhG7mt/LlBuQxN+GJfus5o1RT0Vgng0ryLY4U45pBTjT9BI0DgE
J7O2FudwBG5538RsI/Aqf+foJNlnFASpicd9NpydFqpplYyBiKOdbyw8vmROvaYgJNm9OPrQaS1p
b2k3p5h+1G4PALoTnz7DEcEUNfZf3VBNP/NGJLsAfzIc7K7GtJenXplK6PLsOobUVx5hTwjbOHEF
a+jg/qUpO4O1pf9K5z7VQ9QyClzT3+M0Icu+FRX7ut8ephqgjp0qFUdfSDdm17Hmxuoh71dn3E8A
md33tg5iLyUOfjSD1kp63fg2PuZN3sCf6EPNST3Ab0A97KW2cQJJsOwHoqvHTFJ9S8PJa8ctQX2e
r617gWK4mHws1+wfE5QugE200zBpG4Lc5/zJrKjPvA7hiJBeyhOQi+og6FUXPm0MIqIkuckUlpI/
1Bkd4+vci9cwbbCH/12MgO7pUKqMHWzbbJMEU85OAu7oNWP7IXtgxN0xPl/6WM1cNHiEapD6IrB6
Xliz+LYJWd0irAjpIC/KYhjoWaaxMXzgY/dAtMq4iK26mecad4mjgkbr4/IzD0zDDtmq/RZlxKn8
pNSzMG2lJv+L76sJZi+gIluYI6VChml+72zxmJLQqwh0qaYqbd1uv9KWOXbwmwk4Ywf3y8I3BRko
pirickU8RAZSMyW/DHGMNkKNDjZK9f9SkmjMi+/idn5DoL/bjtvNgAsLzD/YXfw5s8xjvvbaqjZa
gMsGy5KoicZ1dstAunDngvTlt/qkZk0S7R3kjPVNcCM1soDxV2P9cz0GfBnNokueTE2bVXckdMvD
c9AiHPj5q8zh0QaMzSOKTETFSa//Dac3z5M3IS/NwWdTpFGlApX3qRT4UNmOQfqzVLdYLZpmPZgz
+j4FXLf5XhmcG7bBhqFTfDTo3WjmEQxCVzvR4RiaVk0tBNlRdxd+DWS+xeczgtONfyKoh5n6JRmx
vPn4G83vU+PvqlejHD1dLz8vh/tpkoxLMivjCwQ8i86nVURl3d6RfmCOSyd8jPAC4oRKnVImjlOv
kfxO9F8BqWzHHzs8P+I4B+yYiByB6JK9aCIJ/385OQSBTxCt7PFImpXSbaPYEy0mG+cee8vefrh4
1yBtrdSMAPNcKJEYPTtBsaovm1LECXFns1I1Nke5dYtn2uzcLxAoi0pHlGd/3I1cjmbrUWAQ99Cj
UT3Ko67+/XGudtyB05SjgRFA4v+h8mb1ykOAM+lIuVPG88QHvfJB9eZskke+Q9+z8CptkoLfg/pC
+T5SPZACcoyRWI67w17r+9Je9LqvVPv1kDZpSWX9LdDAWeYuXQ/lhhEVjRoiQNOVHisMXVVyhwhB
Z4592p6Yez2dGfy+PjWxKgJNLA/UDurvzddJy7EEd3wQTKLutZmbddBjQxQAcAgCRVCMu8ly3mVE
Lts2qKtb0al2UMHK4ZTXaXKmk2mDE/V9sNxwBmxpfk9prtlT52WGFFzEt1oi4sjqvgN9zE2k1sKm
XRmUbI+bj7mLngBGopC7uI2za2svrzhQ0odEQA51iF6C/v4zuIqDKyt4/c7xL/NkYbNQp1A20des
fZZutXhO2coJTG9x/z6takjYbxos+nSSPmdjh1MEYfql7XCZ2kbFlK+uziq6T0gfSdoe8cxJUEHV
N1LV8F30L86ffJWV59btIu/mQsiHbuCq0ImQb/h7L/B2n5BkjI7vK9/xf5wYodVhI7etrKCYXaFe
JnNZDe38Y6xCnvuHiuacsUv5zv9ZjQANH+tYF4+dUfYkF41zVg4SQChO23ZPzrklFIU2QeommHXp
KBkWG38D3PD7BGsOhpaKv4yLIeqhDvYtassG566VfBuLxPgjrYoBMnT1/dx9az2GzSKL8ezF5Uhb
m9NUKqI5cTPPnF9RSSXwUEPlKP2lGR86K4KLtPNxr1F37uzkPHjU+uecWp2xqHNToOgMKX5zfySJ
atPfU0fDdxxpxzoY25FcBrTP5P6qi90w6u6gY3LXNBNIzfaeCXbuGmcQ0vi/TeDC6kWbUArc3Wpn
TZjfKDvgE9+ZMIWMQIcucErYLP7044AfH4hdcOuTffxgPbv6DjNxJWj7jzLjlQohPu+/5OLzA0Vs
JnoOlKqCNZDDlDCRNBT5z1Yc3QH3E5Q5P8zcAs3FWM7eIIZtYlWa6XuzusYibgwCULCSQkwqRmGd
x+rYrNL0M7QmJDEDPI/cP8mO59//3dsEscyn1v21O87EzXO4SivgjHjtPIhg5+AlQ554kTiMYz3t
Smvv6A7qipG8ZrIpoFN32SOI5vxDj1xhb+U8B/L4PTjKseijeg+3NRsPFSoFm4E1rP0+2v+njgjA
Ma3gBXhcALkdY8olkpdwXZe81rFJcyTtd7OGPt3tK5UWP+Ed90a9R7CwdUD583v9niVeOjNZwi4/
b+sABz/UJd5hZJCrWisq/44qPde1i0IRErOD1Sb+nYRo73+wgVcGRO0f4SC9QdepJnqv8vIhqdm8
RrK7aG4lbD8/7/qMOsHWyaaV37RKGzfK/VphPK8NCwkWIG4mIkxHXAtoxkdU2Y4osGSxTwDQerOj
43u0FGP01gOJgwlo/2RkDUMptPY7ZpNUYougamE96X2bXcnq0Xu9qAnIHPSpQOBS8Tnqha8DocoA
snuC9NlqKamDuhNZAb8XzKjRGIUyqTwVLtdXVT9oPgeSuaeG9SSMmHiML3MoCksDE1RyDVTgX27m
o+z7maWlQgHXHegimAZ2EWNK/ZHL+C0zz5w63oRJcoEWi1DFvk4iWbpm0P93gAsVoQkQpbElVhyX
V303uSMS9r7wyAM3nYi32JsJF9qm5+7byKNtnczxd5H7xfMlTKma2HOhnjTh6MuT9lq4sVNDgj/S
emYycSIVvnbKh9jLJZUotHt+ygrQIfCl11mNJgNH1XYoM8lMtAnktswQmof4UMtkm4jBPRnLTki+
Vm0n6p0BWsQahnQb/VlSdxA=
`protect end_protected
