-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bZ2QZpBXDtZ53CyTH/hXgemgb8AGvAz5Xg4P1YyS5SWVF96X5hVluGCHaUk1nJI61az53njm9XGI
YRELeSbT1eG9Gi5VDFONkzBuN31voXuhORsSn/2oga+pYu/+QFM8c4Rwc1vctT4L/PR+UhHkTm66
ktl+Dow8w9DYKv/38wjkbnnqONzk3f5Jtcy4tukccwtKaQfTDFNnIhR5w3bwNY8ldkd7hEsGxEff
Fp2g9kDq5nj07Toi/clnRwAJiwcvSa3Ds2n4IHSZnkeItofGur3DAFzy+Kj+AvWTp05BFKGcSyVL
puNTlWNSPualLlU/IL58mEqx7XEfkCmQF4jOXg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124976)
`protect data_block
nwhZDcsdN5LiafZydjYEEBxYgTpHbkYhN1wQtxCMbiSI2lQWJ9vtSQe5PmRuNz19w03PHrB/ZK6g
TXLBTAWhdLY3OsxzkaBskgxVpkrdb21akZ1HWsuqwbVRTdVq6Dd4oR4AdF853bDZ2Lg1fU2aAkJB
7X48FhM0yjvCFXP8KRTYAY41OwcQJRo6w4sYDz6TQ/UOWye/nOh0iSE+/2BiL7REdzxswGOjJXHN
m8DWxB1dWYmb9clVlyc/abQkNzXwjd9r2hagYmhcUmTBRx88svG4Q/Xw1VTfmrxrwKc9+nFumZXC
2xYXUtrWm7gsgD2Jsax2mu0NFS9SzPt21l0Gqkz2D/Pl2N3f5H+CSRGTNxb5dfpSwd+Uc20/RPMi
8F68H871gPrkgNcpNe7w7CYEA7bJe0CeMkUmcU2/4M54VQm+SexL6VnXDOGoWYdawKnXpG+JLR6I
jZIBKCkJ/Oup1xDl9nAjE1Jrmggz1BuuMIHkRW/XhG3/iu7UN+0fnnOX/WuRPgGj4l920cZoRz2I
wPdcZZGqfRP66HzmhTmlaQ8YReB3qYbFxlo7DZcD5FJ/E0waH0dNozPD5J3/muJFz2O/pwVdpAd0
YqI3IIY9kAD/W4s9wiilfal2DP8aBOl48VrYIxcxPSzcYl+DM8vlETNlfQn+jXNmu40vaCJv+1zZ
T9n/DyqqDv9iehRh0JgUPtG73fI+vp7PjT1EhuJ8pFckPuW0wShs9wjOTNQUNZQUt799Ydk7GqY7
YQlgZlmWYjBVHTLSj3IF6ZrNcntMETbMdH4XGa4NmQxZDEAlZaDvSZ1+BzJzUBivkhG6x2Hu/AxX
p4QW3UxNyTDB7LordS79ArMdWpzpePpDI/xLkEIcKLs/v+X34GmUrjMvDFYmfU+3drQ4gMcBUqS6
FzRxgUj2CJ5wLCZAkJEM/znI1YV49olS52X8LWcZYUITuJBY/Z9fEQ8QUI/segdgt+UOTJcnv2Ze
QCxqkPTAmmKcd4aECvrReRqFjUM7QBYYxNmwYhAPDLfYqM2X5VbVLIdL3XL+35afpZ7k85FXFRga
xRGGYdl2qBHQEpvH+ix3ZHnQmJQhyD/EKqT8kiXaMltUgOILSAjM0h2tT//aZLVI6dWrK/tNWb5X
u+yvwY15llS+lMZxu3yNrV5MCRac6lur429eP/+YSUuoTnXEiP/auXqpeopO6idOcUEKQgRHSUAc
WS8k8H7LWm2R3kvOQUzzeONC64h1dnZlL4JS40QjPVWZSUmOIm9ZlZGOK4iDoKwNqzQH4RsKD9KJ
8+TDK9RJaQvYwVfVkCFD5lBqQ1iMggxtSBLf2PyeMg0UxRRoCJjdAbgowKubbeNGKIuBh2LUWao0
imGASubG3y3PdAsCZPwnNW8Ddwsr0s4IQlrcZ8sQJ2A4bGH2Uz1shc9qj2iMIIMS9efKG/4X423X
AMFMxrK6jb/3OiLbrUWKAyYFYp9Lk6ZcUiK0jMAQoih/g6Oe5WnJDoUTenH8Dns6SvEFcwVDPVSx
yktFXg05QbN8/NPWeVtZM4ErLhlHq/h0041z1+KuYjtAikleZdocF+e+CkQe00eUeovD5JjDYJLS
6VniVdZ8R/6Kon9zUlJRgdFuE8IkhXY/ymwVUAFTz1ueKEMqHJVTCuRTc9uzSePUmFA50D0Ty0Xw
N3pZaDIDwYsp1NmhmXSoR5OtnfRYjSitwtkX8ZAb/isutIg2DVBUL3PKv5EV3n/m8Xy2rrHHQpse
LWvw/iDiFPNSdK3Kbp9UychB6Z8b1qS5evOtp955WW+PQW09dWrYFEzD3Ej7XA2D1KqVR5jwntvP
YMugRK89q2RVWQQLw0HiOCvRRNTOt9usrlKFfWnaACkl82g4V1Z6SEuxMVROY7z+6qHQxw7OAdPz
h+O9bxrOh8RqnHdpVjakBGz1mUVe4zSjXx+ezN5tYb1e1p2hkogtnQ+NWh8EGxSi7W/abudJFQKf
R/YN4KXLP8Gj2iEDb2K1mnaE8v31ZHFNKR7JLab6x8CqymoAdZaPWvniKUpd0ntVW4+nZb5xbo/Q
jUI0iVrJ0R+8icTwE4Vq0n9QFY+0EvZ1ImetICNoXEh6QXrW3ywkZKaC5WpCgCw5aVbmBThj6DPG
AFz1O75o4rSx+45WEAZOr6Sm3GXSZ5jil+IlF6QhYPGFM8lh/DPKUdAJrKQfRnVGgVUL8QILJim8
055NmYNB6pzkrCDcrr08Q3xccdtHsJbaWaZGh/ixIhlwEdLETUbZUU/OQjV8TjxT/s6d4kfCb1P6
Pzn7HFfyAOeEMETsolmznrQbYfHBp0lLoiAYXYKJlsB+Fetyk9c8L5honajwfEutwPed42b9H+UE
LGQNxjnbcfcMlSBLpkiqo/Sd8gEWEHtup+/YwPSq7bvatqbChx5dBOsctkfBf8mJ0nEc/p/XD+Nc
TM80uy9Qlxcxo3rbMolQtzhNe0quN3f+8MkR3ICP/0PIlt11t6Ayuewvh+Ej2vV296E7Bgzsw/Rr
fLkz5Mt8QzPse19ClVhC3UWbE5v7VrzV2HB3m+NwaVYLqcTkZBWeLacrWe+Gd/jRaRd8yu0grsqB
kjg9mG68pVKB8dzucddbeyituc7AL5g8hzoP9j3FbjSmOMcwbiL53MIEhCcCUSLk51X6oEraIKHA
lvZsJC5QwoPxr/M0yS3hAqT4kS3uiJhk+No7mhH6zvF8kkKy/oxpfEQQ59ZHEcOUfSvnZSAnZ2Mh
gJX0+BaOH43pLy25BgVEPBOwJbi/G1qUX7ihhnRWPtaSbJRkFHLCkv4+LkhMhOngJtTLoIBB4kCy
WmuVdRwAs3CXi1wEDAfrSdyxDwNKtGhdYi6RbsgVHZShCsmxT7vVGsnYAz3eZWld+dn8wVdF9uBH
XwriZUMleNOgGrkNGpSi3OLoUFN7iNvhWUZ5M1TbnwXheF9DlUJ622Jb+Ta5XEjx2RKLJbiZg40H
SorOGl1/VXmGuWFUBXFXXOLWds2271ZSC09l2v7TyQjIpgqjZJl1uUGI2ZcFXlyL/5whCzFwaeLk
6lKURZMMOllrIlNDcBgLz4U+IKmSJ2MBZzk3ZPzdXq5+SpNSspcJdcL/W/sJTjeo2rk/iL2AVCIr
VSVdBecRDogACiSgPAgDe9/XU278Duzj7gGxV2iSmqy+tHChE/UvAm02X26AlDzbn4yqDaqsuV0B
OY5YVBnYGBpSUcuzWDyWZ0lx5Jbbo5i/xZLn58b10aGx5p169+2bVef/nb7svwkX50vYf6C2A92l
YA/FkfflUrRsjw0YEmmMo2oh7vYNGPgILhMXZj1/0ttZRVFDULc7qL1DsAE3/Cc0Ia30XTR/lw4P
g22GBdkV8nbuIBzcFh1K0I9TK1sZNi/TzWnSFW2+LeJNQPcGAIcP8lvV2XSHv2HINo0qWtwpmdyI
/1FnBmyai4Ih6kLV+GkXv9AAmDWO5SZL9+Y5NMZ8LNNf+ULz2ILE5O4qBdAJU3len2kykPjdAk79
YvHuktwWiuTpSc6dwSP/yiGc/cfEMRvoq7NCMRwVxdb+oITG2KmvuOmgtsOtNxgygjuKyb4iV2lZ
Xcy7EISy+ZLJafXfGvYQQRiZ9iZ1Lea+SdJIeLet9pBugYaOR8ieQnKW4UUf7LF8clpHyX5vHQtw
kSZPHxQTr0hIdU1egn0Fxb2Wus75U9GZoSNain2w76LD5WhLQkgzBCkrBh1W7icBKI+v/4JX2YSM
H+7SP9r7fdmy5913565znphHjIW3l8/46x39JfNO7sVClzAWRNP5JQ6gIlP8dv/jNtRwTEXkpRZX
xgNgs5yKHKBDiM90p4mf6MVOqTwLAmekcoPulSg6R2epofT9nlsQSIUWV1APeZvWgdO8vPuhmqU/
FcA6iQvLviRUvk46Lf7zZ7uhJQ1Xm31qf+GVhR8eWKy2QhT5njORP8HF1nHyhAcWzUx6uwvFIw9D
hXLHQHIq1YI/CVvIBfDzsxMjYsfhKYp9a1CF87xk748OAs4pqqWaWGHV3kGbLhedAe23/KYbVexl
laiXT51ij4IGGnmAi6P+qMsf2kL+miCct6fVUiNV5YuPTdxZUC/eg479smvrxZoJtpTySNQcCOtL
TBItS+uJM9TXzCPVzRnw1kfDY+ooYPs8efREJZ+wrtJZ1oRO5NEx6ASJbs53Cay1Im87/lmkkSEJ
0glrepuIhuBeQ9hgLkzCB9Oybx05iYJO+ueUrhAZmW9K3vIxoxoGofHcZKTU/AQzOQGKmPr7hN9N
qwA6tlUpNgT7vHRDOkWZsvn7vwwli+mIMF/IMFJtL+yuA2iwSW50qztdKPy8EKIhBLGpBUZ62ljR
Iy6KgjxL7+uVSBkUg2s3TYUcX6w/KHG8ufqsUGUHWWKcXWNUGpvSlANARFV1vyk4hc4t8DM0nAEW
kz52g98uc+t3TtD5tmXSHp+FXkIs+NRyOH06avcjZHaJFmTFQ50AYBEkYkWdxqkrm3VZr8oi7Om3
1RwcfCocP8E0yQAkEf7Ku1F2xJTW2XZVfRUnc4hBcAqXxyc8vzfWKMsCxZGVeK8mACVWx266Ox5T
Bao3DgtRtYVmtEdQLJ7NINL6/1q9/VHm1UqK9Z8R4trBNFtNAtWWHcQyE8UxUJ+anqa2ARIqDXju
pWx4CPzgncBAAPya1/36quJoyscfqKkYmoCRpKq2+RALfNBkHl8/HZq1ClvW6OksOHPy4nreNB5w
AnNj6nUR1cmeCyFKbYJlatDd6pIws6DkIpnO/0SoGbOWX1wEV7jbO6lgKIjwv/1rITuGBFfPIuaE
ca1cvOd5FIY8h3ORA+KS6tvAJ68H1z+sOh6/h7WkttKJEVSJ3jpUFMRdYUaCXE0++mTPSJslu/ah
6FQf5JNBbvwhXA6EmgaDmZKQP58WQ7rzsZCoDFVGRK+IW97aTiqzRWad5zwMD+Ufk3abrRLx+2Xp
BqtLP0JzEga1BJqOONqrHKqnjhNDCTSpeoQOpkETSNkbTYxTZIBeALhT20UMUTNaFuR4Yz7WJ7nk
BC9d3CW+uJE5P/YcfSVuj7YHR7Pl0sYuMzIoBg1MI79Td/c0sxdG4kmmyz7wEs1J7sl6ouJRtqmA
JLxMHr2sbFWxZ1Enha5BaRNj0gvScf0LoWEnT8xRewnVBilvZIh9+Xdo8zNFs/oaOuVKJF6+FZa4
34KPs1ERY10O6Q+rA9qyt4hAenM21jrk1PajOFjesQyqOskktLLWtKqpGG/BF7eZku2Lo/NO36ze
UbDHLWzKaLfaAet9GdaY0e04oQBguerAN7anqeTBccpaci2u+OZJFQKbj9Qp46WLTBBflko4Jahi
hKd1d9cbY+5d3rIXheGeDatRhXtgIDhZ8Qk/0CbLsYh6oArBXoG5wNze1qCLX0JGaggyRL9YEhcU
UNgA4Wku2NRxSwe6BIG109uLI4dXFKwPagrdyoRWc4Cpbfmz4wRi6/YkKVVZFXgM2bCpfzXS+5sL
Su/52XertZ4xujiHXLOizUtJlyH9nDEdvLx2zY0W+f6U+x5DlhN0GBeaR5H8rU/91veBDzcIY8C2
Uk6umGXETDt2HFumuYyxO3YVKCp0SuhAhJrxcjjrvJJRiOf3eTJCmSdVlbjbRqNHWhN+0RztDR7F
62dKgWWs+fa4V2gN/+gpfytik+qLjas7Iqy8uUC3byhSxe6AEA/axRG8ciZDDf2cf+wblqZ/qMGZ
zK1EakP6kTt3B/l0uRxZxWBC+XJ1UnK5+4REkp+wnsnVIB2iVKVKyonz+fQZzSkVa9KfsoQOHE4G
uJtk3BocaHWpFFuMvVn6nLImq1p6uIwsx/2EJ6IK4BEbr5MQw6EoCxgBjQ6G4G/dkkL2Vom14NbU
LnuOXQjXWtrIsrDWOMXWID1eOCXHDIVI2j5TCYzF/imGTMj0vlkj9AlvLMUQAqp5lh3n5mb8akTg
Hcgjb+uH+OdH4nUAjyuNn/IfTmKP451kJyW4kJcoF4t+iR5zEBF5pAhh01qaQPrE3BswJuePm4gi
+SLx/3za84/etK/9m1EFE6f+qPJwpISvBv6dJ99594BZnyOfSScPhAqnEger10HDSQepDkwPzN9M
pJ9FKbm2ysI4U6cErUeU0jiahjYfpesxc0f82bOwpJOs/OtP9JYitUK0RGwxZoeSoNgO858XL9Up
6KlKvJUu7mdZsLUydJr7gVIa72PvjV75yU4P6EnweRE4z4ddO6z8e36qmTZRbzHSgAsZI0Gv0QNy
7Zxwhkn8c6jYsN0G/jWZMhZt3MoHYBhRXDgpkvYLCVGBUdOO7kXWyQtO678D5XSeV18yGs/lG4ck
Q5xyI+i2qdRYZvLjlQZ7E3twK0uuGzUveLdzQYFCDRUV+U1Hy9aXp++EIHXKrGHFTPDUCvUMquRH
gltyT6LcC4nug5KFjZxJvClWJGzRRIFtmvE2RtPWOkP+TkNHMr6SPevIdBa4Yr4fsZMAa+6r1bps
tXTkFwdMQS5yEIXAzTZXarOQUXThTPrZF1lPPdOMljzeO9CbjsSfXEXrYcz0lNzIGQoCJ3iEwLtT
O25XXaVUrEtteXZ4oetLqc9A0gfvuZ78S5YGF/BUKszVXLUqQvPsC47EOLckGQRcRYnAEd0E/aA/
ToXcdIFk62TDFbZSK+Vko3nY4ff0/Hikj+nG5IGR2pH+DcmeNxANGXt+kN/J8YIE24ED6iMim1GC
98k1MsSKP3ekMII31fo3Xkwgbs9P0N7ZFe2eVbrprpkoG7bdbwxBchEtXoPcah+o3KHbnuipgzmP
qzMkO2XxgyWx1st6BFqi9ZND7D/DLE29tcICnIDq2XY+4vkXB2aok44QANUpO0xuazdtptMEQ56m
VDzBWHkg+gnvZQVpzlg5YQk0aRaXZ9sTI75Mqs6KnVWWoROS7hLcR9+SpfUspC5z3uvy3e1WqGMy
0Hy4aghF32BmscnroThru2w33ffkFnNHfL/WjIhXTbH7wnrVEQy8DZBo9dUc8CV47oAeGyzxbt3b
w8IiA8XCIISSrnAT73A6M0/nwzAhwylQgK5XezWWubHLHiKdr4FZBDV5AMaDIa9rK6aV8mWepMQu
JpaeoN553bhKW7OpLAsBrT4Got2dNS6f0RugpYrHgInXQs425iF26zFN3q4iy482ugOUE60E6eGx
vAE2GKud9pQP4pne2u7fcQLuUNmWs22W1aKwTLuJZJ//wbhfdNFpGu9MWb0bLnH9ub8q/Kl5cBcX
mjnyfud6aofcuYYNx10Nl3fQMVFHvuuksvnHJ85ARwUyHjcGE15FkWGd+8J+TEWQogVcEWxDuf+n
KAqW2EdD0+jUsAh+pSXmyA1WK4BbCt0dk1z3tVdEFmUnCrbjqA+1QHVNYAGF0fQWG+wB0zOCtMiA
IP2DdLmW5FRMjVO+V3V64yMLD/1t+Dl8Nay3mUq28Uylmjz5OgmcitioUw2cZWjggkuo827wJAS1
ybWCUa7s8c3wgKMyFrmY6B4pTiRFzEBkjjA0XoBLNkzQhsj7eEeTQKEr5ABc8zRxUwjGNZEBM1q/
BcUa02DYvLFnV8GVY4TijRdmaEWdS/EgCYi37mk/9/+M9wfsmdRBZDU0vqkzQjvTP1gcqRkr9/xC
IV4OqOA/iMe9jb5vuPxrtCEhOT7XpYV9BOPfijSZsN8Pp9o6VzB+UGrV6qnW32ZOoCQwPMjBLgI0
/7JNpsk0aTtoTyLqhdXYRj0/AIeS8+l+XO0vey2Bx6vVECdp2vdI+JFykWCusDLxHWYPnw0nKkEx
by0/zn9hdL4i+hKCCxc+30B6jQoe5VTk5f+EI3vTFq/X3sU8E6BPD6soM0WQ73SgrChAVjs3AN2P
UH8U1JtVDidM5Z1l1KGsJhTMEPbLdaw9fWGHlhBco/YPOFSgJ3W/dhpctQnKwsIfapbLRasykZxP
eq4GOhSVizBiOFeKxdnoI8WTLocdtWil4Q5E7wzDeBvPc6W93mQLNuKGnJB8zqXQwnAeEb1v2Gqv
+cRLPPND2weC18/zeU+LF8ZP6E3HytD2Wb6kwNAlIUf0efePYJzTwmn9FxR1/8NiSKU8BLK++XAK
1THNumfgxB/TtOxbcXFUtkCzvsD7P3kI/RzV5ca+k6ZnMXgweccHIQc3ivrqQuLGQy4XGOwUxnko
u2NJGnx+oiCSebMJX1XL0cJan9e8Qjco6dH47aBIMIsrRcmHVbiFPcEOzpDKx2i//0pIuG/jiUbr
ET4VNhJWjrofffSSUgciMmTYuabmAbeHOSsc+iI6vwwlBNOqq5qlrhzEJER1biXR+7KixbMZNh8a
B+k2klvaAy1rKX3cWVc33wrAygKe12RU13DhnkoHUVFIeB662LPtOWWTs1j0RjNWdTFQzyn1QgQS
keI7vOayjYAjNJZrc5wG+3h7yczD90GF6nwqXNbKQGIBRS405Ud4VzSrqC43J6SFW+O0KMpuZA2k
UnMbNytdo7JurQISer8E1nZtIfUME7aFx+j0pmtgiX/fIuuJTl4+88jNICgSWcMDCXtJ7NdQaHJl
69BRc5B9EezBt9/6AHvWcayLdR8z8mbNJSLjwzqtRAv3ctz5I1kmqRGnGSqfHoCTJr3diSaYwVzQ
YIX1gfGO5PWkOKd2wV6qMVmz71eth4oCP680SDlEfhLsXQdNwiFtCFo4fnN742xGOYIkiSkaeRA9
jZO7M+5wXUr+fEZpCktUsYDelpZen1E4fn9HS2Jxklh7/dqQ/wlU9QtzybHnmKgXWUq606+cIPub
FUqJZ84+dFoZY8OZDJtPsFj74LyThe/LXkzTEFy5iVJoSVFcmkGq7PBYmu1t8dGRRTrDXHoefSQd
LcaODW/rFItM+5Oq1UXEnA32Frtl7ZR5/YkZGkryJRAMa5P+8RKmAlDoI3mpwKdoQykmn8C9cTPO
HgjmbOurNqOKjL/XKjs4dCKOX1vniTIudB4wdje6l2x61UVEy6Wj98oyDBMtmtlK7epMVtPU2hdo
t9R6DEIWLsPFxHJ2ySZQsoJjFuOTZBfItoWQrOcIF1YQj+TXa9aZj1u3qAMBcO5/1/nu96F65TTg
mFLVfSzUQ9ISm4DRrh85J7S+kyqhQ1K8dChW63BkRwsVzaeBv2aencAt7HStJaUPXBSSkXFd2k6U
r7tJb7KUTyIX/U3ydllPnmtTB1CQhXpkg28kAIvd6nXNhZyfehX7vlDxdatE1t5sUNsDsSA0hPNc
STPEC2WJxkIgFdj83mMCUQGonqVIDZ8brK+/t4Rc4POXn1qiBUvgYNNiXWqCvCAP6j7YfYFhMHKx
Jz//gNEW9ypFfshPWLGTRWPcAeZIMN/AzosAN0pC0SkdmD900YqgUgfcX6dBkHaIVnZqK43SMgqO
dnQhc+Dy/jPtxZK4qmbIAlHUMYV3fHt+RB45OLtoYBUiJkiNBsJxvSNPEiPYG3zva2p4ALFO8juN
nNwJE5CVbonD8a6ztTS+3d01w7dPsrYv3qFT+JMGvlV86zylis3tGvDI2Lvt78AhsSvKUVznXb7H
S10X7Oppqm0ia6//oN8OvK5Yc0HjYnyXktPaYxN3+kIJ7YEdNiZuU45+l/NC4Vw3V4pasRglSGWa
pjFfWRUewQWNdzHadhqjeeCY2Sef+ssUaR1badYK5pgkWDVbbpDWBi+bVWP3ksCsP8JNyysshNyv
8gFyzzWSaPgOE6sf+XrREDM73CAQWi7ISk2keoi6EHxM37kxhvfx98pNg7/aSX93GGzq7G5+Xdbi
r2dsMWM/PFlJRcIiYLN2RSHgsOGKqwxgcocwmo/0UAVs5iX1mFLsNxxCgSQZjM/jw3QQvKAYQ32m
LNXCTby5sKmKbEZ3chCUOUsxHOz2Sz21xT33oZPT5Jj6ruESHU28kCXCi8+ys/yHFuSuj4jpl46f
ENCPheG2Npj7nnlG+3F/f8nMMEZCuUZTHT9N0xAjoQi4Om+gNSdvzr6QMyk7rsab/AoWJuN3oh3U
gD9VL/3T0Ac4V+WFHvH7+zVgAkzyg70i6jOBUGzhSlyFpiHf4Wp0Olf72fN3ialb2WrqWHFSh7Ay
R1jOkd74LTQfSrvRz+c+9izkg5Dy01yd0mS3HNsCVT9J+RfARKKrNGurLJsnHA9bs26TtcxTr+b5
81+k2+kLhtP4ITuzuQMmSBrGHNqbJQFTVFKjglxf8NtKlS8YUdbCIlMowsBPMYHyldPJOAMDO3El
l4aFXHPBDbTlPGaZdBPsOc4E3VZGxV0I+xV28BPUUoCyx1jQUtCWhjI1GTubevE98xDXYEYAqGRg
GlyXBNRcIJVWfHZEQ7nIiy/dzKMejYR4zqnL5+voQo2+9Nsmfx95ALl1LSi+09jnepz1+CdHkXpa
ZtvMwZrVrxSxPll3ryNVWzOo4fqD+penOPl7X8L2ZfhzCHQP+Z5bZA0ZH1lS/bBuYmaMCiL/10Mf
OxJfALWavacl9R+V3hbG4ZTBnG519iUeSe+45A4RP+m6avesVMIOTqtb1IykMJDtg6ZT5o/n3py7
o7Ky81cnApSN7T7I0fu1/MyFX5XWpXIKOrqGrPz5oCdKXGYPWBK1+PrMqNZ7tHlFfUoSfSQjz20k
NN7njDlVL/NSQTFmkOrBMNviURi9r/TCNI3T1vXTthzyyPQ4RF1PmC4AHdlT2i86CtwDjs2uO2bP
2GTydnqMFk7K2T2NBrrocfIVttKNKHinBz5ywhrPOspm7gZgGo3lPiImy1cjFHZ04bSObZPqF/50
lFW47mgdG9AJADR5a7FenF+0b308Z9a/2Pl+fU7vAqwU5j6/b7W5sigxmA+v2HUPKqnP+ArGfUyE
P3SEFN4NQ7VnY6LodEPVbIlhTk2C1vIjroTiYJnl8FWXOjNK7KcPrOXY3psXCfwPLfuGzk44Ab3B
h6gu6He/RiUupFhb5YMONgk7MhUn1+6ep8jnuj0RC5gM19F4ORkveas379BT3jyXgEKhehviXMxi
RIJS4/bQ5CEgLpPiXG39JZenqu4UoYka/I3byXr41UnfHzo3Q2HsBeRodeS76RQBIqzwamtvKKTH
fjIbjc6kvywxJoWloyj8MmYQ+P5x/lkmuStzhs4ME9NHqDcLaBMhPqqoJfcWm5FeSHGfJWPCVG13
KIWWVssMfLtboe5fFWRDak0wupZEkdKo5iedEwnwVXJWr2rpTHeZsOwk5RXY7+sVbBpC/JgYQ25T
sb1yncO1sNwPUTDTdaKPvgoia9IYcx/ZTvA4zuu6oGWnNjIeWEOLloO6NaNPkU0cWalMtSfhBfO2
9OhaNDURZ8xlJ80524UyGlq+apT/Hxab3EA5ZrbRITn51IfBMNbOL3WY1WxSnkfS/9ZNqup0anOT
NqfwefKY8ygk0Slt6aOBEopZorQgFfjYKSFtJRRGKq8y5WpmU6E/kpHXAr8UAK8sYQT9pKmeVMSa
k3DO28ipkZayCTmP9QV9HWdwT3GE8CX+VJUMc4FQL7vstS7Kb1vFWdb52zoCbOoRrbzYoEiShEhZ
vgAx4eaByRCLCTENlK/RF62+ngr2pHja0sqv2CdLuQ/XG2gsbibSe0CdQbD0ufymZQANJAjVzBTn
KgRIhVF1MXp4mVvxUP/ecL8J4zit55vuYkrZwGZxfFgL6qR8DvSqkEeZgOUUkptGW9tQ/vzHYqBm
+OL6grvdVLhu6eAEuQT7q40JX/WX3GQ361vuc1KP53NG4r5gHeaooUOqwp+Q8zGXJxpGt5j6tFAO
R9oaoDF5WKNLf0zu6m0sefMm/yoTHaOhzBT6qO+3uYJuNifTHt0VcBkFsz56CfSsNPMYZjp2nwSu
8W8uucI8+ThSh8JuBCjJGoviXDUV6jfNuKDegvqgJyl+DoExkUW7/brKY8M/ZOrcbp8C4R42uVu6
3d9+3gAZLlqWGydYcOVEBCR0VAxpGT7D3KR+jlPWEFE1K1O2AVre1bedrBMYT3NKy4MsNuDevndh
GE2bxt2dI7QS+YXHt7PQc7rMNUZJ80kmO1fcurETu54BqKmy+8QWxBIb9EA+DJvK+tWCs9oghpOi
1fe4U51EPVkfAeSVHz9UKszm8S1cv7WrDRMcNT7pfd5sQXMhf3X1wDakLatHaTJHUfz6SLMBLzr/
BzeIIo7TyKVbbcvOXUW0Dij34ulO9MovFYfodLb5inbYmYI7VjnzU/3wOIbpGBDYyhH4P61qbFNo
RqfQlkZWBQJZ8ZQIOMs5TwIyXKc7IIg+mgEu1o5Mbs/AhWMYMYW8HzU2xYBuvF3lsGwMXVUZQ/zW
o2ql8Cqp6rcyxBYwtaGU5srzRJAOWUVxpetzHyotnH6/1YljyclV4bca5MjrzBWknZw0JBiJUleu
S2YpEggcuE5s1oOBVwGugGPv7Mp8HJ77qoqL2E02ZCFxseEY/jah/BdmVzgT3n554b3K8l1LNOoI
fq6MxaTyoY2MS2fOf5IBOtFqhvWEzKe6el22fsRJsJfGHEacV1fcD6oybTTnRyk4El7kDFeSk/BH
eDcZV1QGv0CfHTweMM8sZiImABaeUpBYURXVdfYPjW2GWeZVWJIIK6jwIuS6kDeDWaLz3px0oy0c
1oiMeyAKW2XdgGPg1t+vWtz1nAvYNe0jj6RuEZGLTjGMRAMt84C2iPyetyK1eNSjHucZUjN5exFb
p4LrlZoY10lhv7fGJWEi7xPyxUq+G6E7FW0xFPquXOhEJDMqyQ9hUW289eFTLcEiuNZwPoYczTWP
9wFmY9RQWhX7qKMvzvMx9mMMjbiiUxsP6g5DFzGGsRsiAKMfOnGOotLxOlJIYDAZjM8A9T/HcDAZ
GMCLGy4jxx6ewYkkJ5OOQCoAruZMoSn1JHSRN51dXfX1DQaVr//LJvXIjxrQaxaZz+bhJ6c4zXgK
eRxT1EyLGC5WETSUseX7i6Q7EpCd0wO3JaWt7pnVnDz5s0E0gR72jZ1bwVmMLEkFDrU3PFipGNga
1LN//S8ZTTqIBRl56/QsuaMRrTKvygyvzVwTf2GiKjdjoKzFkoKKxefe1JxdsTk3CrmFOqajSU2i
26eEhkU+YJuyI4B5gTcVHOOuc1R8Y9WWVjZacvTieAlrZ8mhBSEkHfv9ZaNSrtep+iWVFbsyDFaf
vqLqPqF88438c387xOvlNmntykygIfAaO9MCRBWTvHfJXnsSJU+qHlK9/68fGGQstOKV1r4rUQmG
GQtcEXQV+zEd5SqHdCep2iaDgdJKayzQ6kzyWzwXWZPuTjZuH3VjhS81GQ62LayQi2wayCjCHaUp
aQ4XGYkdYyF2lpUJlWroyHS0AsQiownwB2oE5OL6ZS5DqbfV5e1mjz6SFiGftmFvRd5hdo9grazK
GBeyexPhtgHbOyXDaxVFbO4h2AIYo6mWFzu9pB6LmcaWBc0mKS970dU4qPykiqQuaofxQRQvmF8e
NBhdOmQec3wsSsYKy2Eb/JSXFftq6QpoEEODfWBa4ikgQNxvkDw86p0GiM7Wwa0mKL9EJOJEEzzJ
ohC1TCexOqjBHQ7kCWt4pbokufOUUR2mig31BH8CDmgLSBcZkduMUpZzfaMo3b3hWoQr9xRGodZl
SviwEwADH1Tt7GYEYqTK1UFnyQvw82V+RzyadVKobIqHr2rFwo8/Sm6ZFgRGG2dTsP/6DZVGvtpO
bWV7XsrEsZZ6qocgNruR74nD8CyDD6I4aSuFpWyzFX1Y2G0TmgpQcRHb5cdSkqmNISzU8elqq9qw
IGWO/EW6ds1xvd/IJoROEuZC2IqOpTTsq/9m3wP1eKTAEGoffPSQIu7eiNIW67mxW5Z2SxahXmmZ
W8QUtR429pFtkHAKGH1b76IcuoYcj5dOyDQCNEogr006a4EXAlj+/yTyWGThqysSC6O5o0JLq5+o
Rug2WU/tIIMUqahXdmGPHbSMbkCIcbHEfyI6k45hpdjsuPDVi1yM2UDSrO3YyW5s2iVcbXibb+vf
tUKIOqZQcbDe09MEwe7cwY4yzzmsUxwdoP7NADr4iNQApGJhGGB2OOH0SqKRugny0M/VgtKEMQ+v
+H12a6UzYjXgvr/WHg9DkY9Bx71yglEJXI7eL12yiG44ekkntBE7GIikz7tAAR4m7k0NwLNHDsCL
9U5lZiUo3BdsgJnbQTox1ZCRljAgYfyqM/gmJ8yD3tRp1R5A6f9/0Y+MznOWs61OtsGntJGy/plB
JOv9KO9yBwgfE6MGbXcbRpfQK2vG6km49EhX/wMpkS1yTY7wRLMBIAcKEMVopJ77F19M2cymx+uZ
ZLIwQ6HZIYWZNceF7rt/THyZ9vcwiERR7GpxDcmc4pGdZ+GSZAUHnb95Npe9W/qX/lU9u9Wiz/Qy
DzyCzsGAOmBjFt8LOfwW3j1yq+Hq7cxtIbx/gYT8L0qgZ45RnEsBjExTgMosoFvsiyV3aILZKe0b
WeuVsFyHxacCBmleX6FuvLZep/6TMLoGAqrBnpG2W6v8nCH6eP/pRzqPNpoJsnDTk7ymAmjMYZ1l
4o6Edwvjo3GA9BjIfSB2XVJT812OVbI4YKtIqSfrpp927z+CPVrhFmJ/rvITE8KmaRLwmv+6ULr/
0DynKf8P8W7VAJQlLYdQj7pEwQU50F/zY2uSUMWH2B2xplm3KpebvPWlabP799lkkfflBiGvoae8
tl5bVjOut/N13nqrVTzaPB4eHKjcykgYpIoMWavUsiUjEuv3tbJ82sOJNqYaUio+PQTajrgwDvXA
2kuWA8x+ZTYIaCZxF9bf0zzcw+ywD/ZE4XXS0iHTFnkMZeFO98VKy1WpCa9ALW1BGfQVgnQCrrbu
ow6F+iN2jAije1wceH/dP1tO8admz7KuGxeAriXe+M8+GpXK8U6ykARpzoGzmreRMyINvfi5f2p7
IKSJtdEwuEmVZkukEgnjoTqoEXnn1WUeJFEdocqzAKF55kpzQUMAAGNEqfsZXzMPC2QOPwMLgZdM
8wJKRY+vR+DAM/DEQxZ37m/c6Dnuy0cXKCaJVVytgUyNhzER0OEbd2UUzImXAj8wDQw68C+4qTpr
5JbTt4ceS6oKXDm8Iiswv58KS6OmNlnCMLQA3SgzZLHYzCgj9jpoQioQbPSt0r0hchodEv7/iW7E
y1MvoST/Apki9ikB6w+ur1LH5O4BAdqe9qdAbYyDd8TMLukWH+cA8Jp+Bh89RtnUZ0m/fy4H6vOi
k4f24COWQXfHs2B9M0MCnQUcCX3qFnWlMwm+Ji3cWKkPWr/EsbbluN031AaG9hg4noWsGipZCZcq
xaU0k+8r8DhvcudLDwinxuu5KDU8GG1yLEwfB6tnAaAwd07BDfqMQ6RRX1OYJ/GzBWwN0hgdbZpr
X+JwBycms8i+fRPWLN+tFEH8PFzLpYTmJ9EFx5cennWWHZiVO05yktvQJlhEszzfUj+xYUiYX87C
SURYmwQoABBQ0DPpvaHVVpJP3OW6uPkQuNkxF2d4s2/T/0OgozUMybWd9007CWVCnA49TBTekJ25
qOw1Ueq4QYqvpjrRC+1TVk5ORTg883kriOskvhAs8fJk1ZOX5406fDTEKMpF1g0Q4W36sKJ97ELA
TsluxJHQHS2bMhbNSgJfYm4CkQk2WUpSZEPXscnjn86f5CGEiuQ2ZFfIa5Dm0/BUzZRmkFRulyY2
32YliXt4X1YhejpWnQh7aauexAII1CCoqEGEVFr+FE84QSLOb4PlzQk+Kd2H7Zz4aRaTZ0inxzWN
3VaF0rFdE83ipwJDSleVpP4ZJARwu2DazXFid5S9ZuBvA4vD1N6ucbR/CNtNoYwPCcvVMdqjCfpo
/N3ct8G47fGpuriwFdMQDlpkTyBnx6NpdA/T1gzkeuF+rpYopWk4LdoOoqqw1F6L+FKrze7MwlJc
Gy3GLN7qgVquTVcPGBviCbeuHsmZYpKeLGAH28+JPow80ESwFEyo8uRg9Nxge6c13wqXHGk4fWMy
hHXqPnv1mqGYBAGX8moguD7n0HXgX7sczikHcVIdekn+DM9ATqeRUfGn6Py81oxYQb3sssoEWbNN
8rR9PSlUtS9qjxppsUpf7zBzr0HxFbzKcuCBH5UTGELzcR69pFxGCMo+u4R10OYN7m4UCuXgb+Qh
RB1/fxLrIje0UbJON3EExJsW/BV7gQz0zm477HBr8SqpZbTTlfjETx3JmEnG0rO5ov01YSXnOKWi
bYsl1uzwP7MyWJg6FhaIoun1hNrCG60wu19e2FsP5/t7WxErEnyIQX/+Ffiekp//y2wuNDumIUqW
Q5uxfiy9NWJWLKUpcXX+vkXBt5ciZoqNoGIyZVXlPSfZbsqD4z2gEG69b5IuNNFnd2rVJFo2h8r4
cg2ljl2Fo8hHrPWs2URdhTEO/1N27syV00cQjv09H7MINr2mObp7xl+ka03AHeOUJwgTvC5vx+E6
bHsCd0ObHdaUTKf/J7wQ2+zR6qrsIAPxGNMm+CHDMbk9sh9fVtXf5gX6vjmXucg+43SUce/yvuxz
rtxTMQmP2UDr9leLE3HZU4OZzW+68AnmoDVV/IuryY1EZmvbr7+c5+YrArQGSYbGLZdQyXKXoC5W
T5IvJiAi6dY0e8nFu6j1bPM6SA6p/D0DRYdasg36MVmQEYeelXbY4KuZcsJiLxJ0U7+0mbbDIvmR
iXXhXcAqFqxFnOAfSlARypLxuz9Vo8vrfHcSqziF5MnuSaYvkjUxolNKLFgw10kAG6PQivVrvC/y
x4Sn+TEXV/QFSIcemKsGN1lRXWFpka3AjNjzg1pXgapBzagSRIxK4bVgiGKYy1hp1IpW2+wFmswO
sPiIrV6/tW4a7s79LeGWEF0I9bh1XArkLeBzRqpW+jqMbFnRQkJrx6qki+URCb2hdEuR/1fCLT2T
Vyk/PY223qHGf9Ex/OYR5zcXDV/8lDwqtrUiFqkhRZACVyYFsx62174pz4fzLqtY/pSibP/slo8z
URvKywfj9jL5wycD7EiyGCGoWA19ySoakPXgFALIS3KPA/rtF1TfhCRA7nHGIpVto38qtTChT+5K
dmLd0DZVj1QLy2BGWuV9pqAvCT5ljktFVqh6pjebRekNvUGMd1AiAk3tcLfhoStImes1A88x91Fa
TaN0cCF0cMTeztgrSrzRZ3HFRU9+apkOHROw/ea0G9D2v2A6koXQ3NVPG8BuZBQ/VRRVYJT+5hbW
l7V2DkovOsQ8aVzfyN8+PCzGCDdSdE+55rbtqhxVq9NRS24qjAJTj++Q7ZO25oKg2GDxUq3gRYc3
iW1aPI0tuOBZj4AHEfkCSVg+nG/nXwTAseuUVRLIZ27giELTjvDXVrBieL4stCIe/sopU0l/dvuo
8mcChfOV6pgR7SUP/zjubIK1Z5ulkEPggjOS+11z8/Sl4hvzLZbyvRnmsd5+CgdUPnn2UhOQ1lPc
MYdNhl8qGgZAMGSayWoTH1rNUfeD/KxSLjAIbRlXj8xdUfQSbzHV5YCuaZJWZAkzMnJZo3wp/6iI
mJCx1PND/3UA8P1x57wZyDwlX/wAG5XbwRUslY3HSYpCNJNG1VsitSS60N9aQrcN0ScyZNsl/9rb
o4Pz0mDip45TdIs88uxo4hTQf42tToHNbWAKJssYRKXSCnpkv2gf/R16lnPy7Rw0gDlJGPBAKWXX
WRRd8osB5zXJBWq8iMIBpenhfcBI6URfA6pHoZYup1VrBz7nYowKxQCp/05RNVtJxQqR8i74Tayr
1kNiPmHhv/reV8zG8PwMBHG9T7jrBDHWpHCXaz9NEGzUo7AGtPP9zTu0GZzzKrYIAjHx1iv6f9WW
8ILUvJc+96BagplUHNgRCmw8nvnOc7hUpijIWuRC7jt1OTGCo5LsYNHunKHMfKMHaa2m7ZksqNah
yeJ64QRv/8wgjEXY54boLnEJIaM9xnbKFZfjeotndDtabO+4R7tYVFvn88lvpaAU5vZ8HpFj3h/K
bfxWs4sHkmBZCc8EPb6mDPhdevlECFGcH5bvDkirfZFLLu57yPYxdOuyAlQvPpfIvKQgz8l6JZ0k
CnFBejgrZYZsiK7sDr4KGV8UHOWQqMnbdlmENLT6pWPsUA8Ek/ZKHRmWXc8CrBB9sJgE5kDjEVcS
b0dARn0IFRDAkyen3OS9vAzfMyFlts4m0ytN4gbgCOYZ8fDFCi0NTqmBMDcRyVvg8gkM9K2wP1iP
dg2fAoCoYL3HrfFNRAtCvaT5slt70bYts4qSuwBfl8CPAfZjBfoD66u1LKJD2iAX9lCQ3xRB5FsZ
7TSRnJRgk03gkRT5CPXxcqhmY/GBWeP4FuQv3izEUplM+uD2qjof5hpubuTNpmecSGwr9kk2nPxT
uNbd1ijmS1yySq124bG0MDIwPDYbGtyPDg/YW55cajeFpPGpQRsTEnADU+8E0/+rKTpOf1nogc7t
ioEVRB7S8oFSSPPwuFSHr/VR51kexoSitZDUJRQVTGxp2sw4HfaVSM7J3cBYd4nMkFNenxgJu7Bf
2LVzhouV5+r2HmIowYxq8nezLHIegHCWnvmHwubgjTsXRr49NVbiahieZSXSCSB0UYmNfZPUF3HY
1LRqUzK7sVi6tBwPZLy+TY6fytNoS3MAcwQLr91MCwbnccnbTBPGxzGc3Va64YXmTCQU4/4fRtfT
VAWTe6/GmWJl35qSvGJ2PKtsKnb8Kf/V9kJTV8738SelGlArwSMDhjUMeAmySBCX/lwkIyYVSF2Z
mF1fpq5WDRgtUasGUOTP0ekfXPMqSMxgS9ltaF/AZmoHnMt8/69iZdIgoF9zK44Syemb7Bvl82LP
WjsfKdW3CLS+eibZfeeQSYJgm3m7X719j6gp1TSpOviIlL/i6dWv7cfWTFUkgQyh+VRvCvstrxfo
RDmWgN0GcTHHMaNlcltfUVy28YX3PtagwzV53/cSO7oYV7DlNQWRvVEc00CNs8WYEtGV7aF5tJH5
AptqtYA354uD5dV27fTWXoQvPPAiw3+OrVSyN5X9mRvyqX4susz8Rme1+9r9TSUWCDfv1vpc/jHf
uRh57fIqegIJIP366P0/qQyJfa30tocyFTwvXSbsgsMQmGRTUUy2qHoGkXdVPXn+f3zkwuJPPZ53
idOoP3xfg4QK/29xW4k1aVixV18e8UwoCwUKrUF0TsStcTiGtIiK4Kp5jn0VWAwUaW1i2woKfolX
9QJxwUvCckYiM/RztztDBQEvq7LSPDKfSm/MKSH03+Njluv8j4WuMUWUWP8Ln8lsUE+KmDaTvcpE
HgAtBOH3bCosCHfCnVfxYhnwyyeV64CsDRPbdYd5ofmOWNPHjYutjT0C9N4FsN2+P0Z+QXG+9o6m
X7GN4ACNIB1P3aTrjeiVsh05qn/BIkAYd71QojdKvXsbB6SvorL7T1yrcPtGQ33RRll+6VGe2Sa+
gw9mDaYLLm4F0M1wpe6FJek/yy7azquPse5P4bp14wZ4KslmVfDQGo+WF3M+MSWNckQJXI+G5uW1
r69EtOcTWgZwIwpb7b4N6zci+LkdKjPVZUxzj83hZq/17u/xA8eRZz/IDUI3wW9Xj50yvvwhTNDT
E2yYPTC6rL/LKeWv5evSAo7Gwn4HlvkThh08647Tf57sTU5XRx08Oy7QEDAuIeQ/aOZsuWAbOLIY
xu4qJ+twwpn14Y6IXiKpqbc7M6yN10x5VcWSxUs4yWH8T/SaC7CgZhxRoNg28IKm7LRMM2Vl+rcw
mUzxG/EaQm9yK7qIBzVDEVdA7gb8Ibd85Wp5Zjk3QMSFYQCmKtcbcj53WvXgbzYsXuWOkbGsquXi
sPpA3ujwXtEmojG9d7hmDHgzg7xEQNHtc0VGdMWs50pvyJ/vhgaLe7F+XPRgiYgpSEuTT27FG6K6
05qPtFR9XYGOeBU+LPg0NaLYgk8MPXMvRa4yGLf4lW0dnozaDmmMJV6qxoRk8rSh1oyYxmGgVCMM
MbPAbd6KfX0KVqneTUNlpZk0xThQQAeS1fybj2imT22zZnXFiwgcUU3I4sxs263flkTsHfnSvXqD
64h6NpZ2uG7ge1B1yvbLZEPxowQJ68sSr+0LirwhnGbvZypyteuD/XTbGuGNv/Z5ugcJymMs1aux
rMonNDfD/ZU5n1k4AC9fprjxPKMrzJ6+icLS70hVqusa4fg6OVGEJDMxUY0ZSsY1E52mznPnC54/
/bG4OZo8QyIkgqBrTEvk7Y09U7fy7o/+DAzGt2bAdOOjN684ZU7gMrT/iO4jrTdvAbrVdjUu59WR
0bAF4pHcUHvUuxb+zjw3GpEuZDJgJuNoxZz2FHLiKuzZRldX/hwt1EnNmymE/7vGLkHME0/zvuQ5
zavlHSbt2KCKaWU5Ei3fgv0vqYZ90KuK1Kx+9HG2cPYXy/fncsyGheKmSWl0HOgFCHVF+AfPbRgg
+fAME4vESuIrSA3IWwY9rZmSIZGrksgSB8NQtfYjaiMQETuj/roWQdw9fri2zn8ldHUcdBrAjdFD
iC0EBp5gXzHqgueAP8OxGIUBMa9gPGHZ/7iez/Uz7oKjgmE6evy2fy0mzQt4T54EjA5Y1kkV6EiP
2Xzi842UCT2TqS87DqXYozPWnPb1JWxaqxpPT3e1s42UJkS+nRCIRWVzZ1qoJU32jvYd+RBf6LuW
k7txS3B5uEg9w2VjJ2+5DVSyTnAbmg9iRqJ1gW+vTPX/qwEl2dI7b4VU4GMBtIBnYtwedlaiiF1L
gWB5buKJAsnU+QT7EDdWpR2V9b80MAn8RtaSesi+PZM9oOVIA5oS9jeyApduCrdRi/fQVlTfCVSa
TsxLhBVscNMILbmCgHUA2CAy2K97fLL45aw+MPWMKV39AcAmOpPfRsiWYeYlDF1iDslGwz/YM0uB
Em1JWTrU2eJNkctIvsB7WUFR2h/SU8aNXPvI44yOIcq+1ChFkUfETnC5tEb80NtDAbpcsOzzcRQc
VHYUQwkTOWl+K0ou165/fpIY8TgOplUKFBFsuFodzAmdnGZTQmkXesRRsbem0eK6bR5eZq+m7vbW
UQAxEdD3HgXKCUzCyw3yT4lXNcyD2+P0BCCzDnc4dyA5Dglp3ONRVC+syemQXdQXAXYjHlwdQV1D
CwGmiKteOKMCaVPsliPfeMCJJjU4TArOxSXAE2LxiQnUMgG+WIhCKOYcp5eiq9D02CDn/4uixMV6
BwrblICtJV9tZwi6Ld1gYlYsIXalDe67bDUa/apZDZFrlDBOHo7afwkz11Ag92SGeWQDcE3kTnqL
5TMdrLuYw6iZym05jKdpvXFNw/iLK4qIcbVUy0ZHg9k5rUOzyfqhu0tjKmq4lX2DLtSjJuxDqTBK
Ud28Jxmu/x7lkc5Z7l1sMS877bu0vLAaRMBwWRO87x8/8J/soaLxYUjYN7ByiexqGYxgAQm8W8eU
oJmd3nDFRNjfaUfBLSrKo6ELn3es/B0eMclR5wnNUrL2Ujytr+NXQQAGyKUt5vl6cW0svxWxqH6n
S86CaGCwel7FljUEtMuKlsgdANrr7x19sPPMaWkfTh3CQlTD6QEaZUzAKlBdByyHqzGFITTNMfdz
3BKlrHP8Y96IiY0UbOnu821jhFtVPjd8O/c6/rmhXXcf88BchIlYIl68qWxXKvDNNuU4lI9k/A+V
CmTR4LRiXqCSMFjez2Npn9Q0c5DHYBOajcQuureTndHhuwkHi+ocsNBzDFXC6nWgXyLnBTjXw5+V
ZUJ2z92Ku1WHAX8HqVtDC8TQHsXZPHWnKs83YAQTU6Q/7ozAoVLEfor56Rgvtye5FVtFFiIGVhhN
WDvf5Oq98uPEIBuNblhavqdZttRZY08HMJFNz9Fv5GBd0g7P1lVVLh/7lwigVm5/0YjSgmXjeff4
+Zs9jTF2sFAOqAoBx4FJ9Ae25pzT0sp2F+QQOeHfZBU5NlbflrhoyvkfQ4rBfuXygBLC1Eua/yY9
GYpsX0Bjr6cB2h8WZ5vdFfwmsH258qtU2hYuujDeo55TLQ6vf+XB8O4bbfpGhCGeix0tkRLHynwt
Pp4sSyPjY7A3/InD4aEE2afYlOLiNJgqwaY5az1o6gKSG6Na9BAWxNFm9Lm6fvLOFVJ8L2oiNAzY
PcTCAuKVtJlmfYivCQpAMVV1vtx0MoVEI2tG8cf7t6/YG4ru9TvRq+Y6KSkZgQd4ugPKRzDR6WF+
h1OQ9VdVrX7ypSJArujdtvWeT31uio+x/VUCqZRdrG1yCynjDDSvFnIDz2uEYxbfRS7GzbhEel4H
A5jrEPbCmYDSPNs7/KG68BtwG7VWYrqSAW8G0MHNGn/8brG9oiEIlJaYCsjCRZ6DnNjinlO3EY3P
mWe1LvMc7zaEQsGnxc2LwRvIB3w9axcty9L+YhqxtdXNMObDHiPV59lujW/3JyCKiCSxSy3e9p04
SaNfP9TE9bvzcvpwLloJWBN/do/a/9LdnevYTDHJ4zv4o1bPU7Bg+P+nVPYq/v3hpZCCnYHOvA6s
r5JuZaKH580J9wxISX2FHxfFGUExiUSqnUrOr9k1uhkGQWw1fXLmmr7rKif/MOHmXxYuYjbmb9Fg
/Hh//0KLod6gL6sGJJqDJt6jK0yp6VI9/NeUD69jY6L07gLIBNB1nhPZzFqRSXRBjxcbrZXh3nnu
e4Qait4vW69RFv19zlKfeYqK998iD0i0XdLNNHhkBXxMuie8rpFQMEm+7cqKEaoYq/aMzRrLl6/1
r5TN9uUeTdxh4VzzKK1XqxWhDMDggUCt6D5XIMhpeNERufFJxjF/zdPusEqz3pmA8Ta45joIe+cZ
XjAmwG+lpF+OQ+nKOrtQLbpNd3Z2wmK7Vmj15rmHwlnQknqQgnc7b3zzJQj3ZNJYLckkm9filovA
rjoJT5WBTlOh2Wf1lXd9Rj3nuTdlYXSG1YLf+aa1rx3p8maMle+LIiVLCZ4SSmkseua45Hu1DqHc
kvIXP3tBV4I5xLMyYs49Jt6e/1GQdtmS1Ik5ESq7XsTAvCHATY/ont3YqUipT1UwaKemDlLuqm74
TBIh1wJcl5G3n1fGcWcmlkK6xdgk9FzPvInBsI1oJQ9RihLf4XMHYmt+4S/VvCwttlZcDWTX47dn
XTTE1BdejTEB2Un4ANIMfZXR2GZucenvCtSR9Hea0oRJaonUApcScIWMKNWkHMxrvOaAJsHWABlA
+Hm7HljTQgLHnnPZkWptS88TiaIGb1rqIlNcJcPzclvBB52GvC2xfRUSU93f1lgBSyo98LFLye2f
MuESAnQK9BoWRhZrJWZXXlfzurLEjvnuUrCoftBIrAh4YQMhVFQHPmD7Sae0sMaTzF6b/LrLyp8P
np9tKdJRuMzuWnyaz8B7fPir0rKRI61nYh8A+ITlEApjSiyot+Mk4ZVE3BUUp0wkk3oGK6GZYXx5
17CPlXGo9oKQSVXf7Pl6pifmzbjCHwWtglx4CstP5cK57czN0uYGbjnkNqUvM0Qa6OczHS9XQkD6
YK39owi8yVuGDTOTOOWkZBVN3IV78b2ihYxkUhEjxOIf9mjz4bnqXGqGApUbZ1SJDdPM3wjrHzeR
DUXrwnesLFcC+/Zf/lW0dfPOFqIuEpavm2gSQymHXnkoXPo8yZH0R9Yv/6B5IzL9mh+rt7u3lxT2
gHmLBqZl1uSRdunS/XTwBSiHZvRjM2vXmbi9lhiR/5qqvxPlQAmQpdFBYN7kut0s4G5QFbR77s5R
/7AO2ZaBycGNdWSxqEuIili7eNKr+m+tspIl7Gndachai6ioTUVpdIqyvCDcl2FrfLIs98DulOWb
+TOM8JWPfpOHiZGJ96aGndXJjTnNLmcA6m9Ua+PDkeyeQw64kCMVcLhYRgO6uCd16Bd8+F2FkBFC
4wZeWswh88FAeWXF0Q0PPgrzmowFu3aC1FhYMLma/shnU9bVHwIsA6zS36NGwhdMzI/xArsqVxWU
3mJtecI7kUkefBc2AzltISV9tj8AExymghCs+aOPjbjyAugvP1Qo0rcisT7Mv+YxayTAeqLaK/Ix
xbQAF+3RSmAxRxoDmb5dP+MM28i3MtLFpAh9ar/tQN4dlo8NLqxyf+0CzPVkI5CoudxlkFBdRPf2
wDqVybYri9ZmHRnHzjoCdrdoABQwHwiFwJrIGj7tDhBOkNdKRQmts3tstXUDHJ+1/WITmwZaSvE/
kNke3o1VQQKBu9ryrpLpkh40hZ/G9AYGpivKFx6SSqBNOkf1jv+3Mzkx2Q+jszlec3EFvq7b6ohf
5NpQ9OkJamqlFEfhoHUBF/A7tUpO0b5Y2DlvOOQ/Mkz1NpteH8ose75yrNDUE8XnpYN6q6YWcMsS
B32EIXijBYCPZxgxp1Qqlie7zsMnjuOfHJoTxg904+18+uk2phLvHqVEzX0G+DQmPJcd1b1LiI/H
8JMv06p8eF3cKgXKCYP9J5yU/mtkyat/dSBozUAvizfAUihsh4hQk74SUsonORun+4Q8ifgH13is
ykdHEeS2yVT/ZSkbPbc3ilGSHXpmCUTk6xdCK3fQfCiNiQ500AYxoz8L8gYvoC427AyMdXqPqN7i
hXBtY6TAfb43eklZADJltGTn/HXrEGAFNHNpbk3ZKojIq7xKSD0yWdW39KU9R+aDkCbguxLnG65L
hRe3P4bj1ifW+NZ8pCcmDI2qEMSDtnxh5IEl9Sqtrb67mn4WJB4pt72menwtWAwlFnvSJZ9hRDUM
uV9YvAQfqqGq92t2eVa27YVfkBc3ztb7cr3lSu5hgzG3iCBJuQFSLSHb3fFBQ0kLDo5XtJcKpSO8
vd07QttzjoA9I0sHCcOtQF1aR0vClJbRCr1G8+tASCSWK84+VguMojWGt3EnQMIInrsznr1u/Gcg
ghcQsIEobkGPfonRDnqcLIHTHMA6nXmTPCZ1ijD0L6S6Zg7Rg86ma96GXsV3JVXsXtecxydDiqD8
3CM5Sd7419PndOCDqTSP3k+rFiffOQAjp1FoodrreUXtFpBkB01vFSFPnvAKRP/qpnjmePP9eIn9
XvXuaFb94YaI30GYEXnsjF3SSubLyIWY44lvkzCaP0+5EATP9lPZZXJcA16t8i/yCdUy4sauwVig
4ttamo2hH2GRwLTbbfFuepn9u9qLC/21KLxeJiaCWqSoCo/7lwegNb47UVk3QTBRO9elkOYrtf+g
hyXclENlp8xk4SWR7sH/vocS4ABiJsUNWzStB+QtZVoxrJHyWzqeNABnVLKkZIvLMt8XXcwpDCRY
7wHRnByTjn0N6KN5xunktGzTDjhvLB5lKfltL9L837uP9TmqUnHxhnzETSJcbRDwtuWWZzNvHdjD
oTy4KifxOWPvZ4aR4xEwIpJ1mST3TcHeD8LaYS7PlOQT2gzobw4FaA5O1Q63PXSbmpQkPw+Nfc0R
drvxJg7tL3GNKwu/w9dVV40I/oxHSvXbNIHya0RmK6BdWpOhj9PmwncrlxblXUBsB7VTDP2/uPwr
RXio+Ou89NGqzDof8gVlZrySL8TRF0FvImqaNkqTIJ+69Z/TzHLFMrfbta5Yyb1DQnRzuKNQu5xq
wBA3aZXzW8hXOe1KD5c+kkBV9/CLbi8IEA2YmSfmEfIb4pqFYPjwxufnd0XHmZYyp/Mm3H9RTdMm
xe2oUJIxMX02to3Q89nUBzYfIZahvrLLnybIIEjvN6flVPnnUIL9TNUIC9HlivXnRlxYJvsPYNn5
feXCua3w8c7q7luMyemdRdeYs40IXQHjfxrZt23lHKgqxy9miW9peULI1H5zn2L+eQ3tQ9Io9k51
XIRLm8nLJxelNz5W5weEpD5Dm/XCb/iUEXQflUvC9s60XZ6PE9y8DeSOfK0W4lYuW9wcQxakzggr
TkwCpD45VDStfOTTam7GY79J5A0b2PKRoEilV8viPBgQUVuH6QVYAL7xinpsiTTjNgifiB2TDD29
/U5QeMifnI3N1EP9L6oJAYit3I0QepDbUmes+N2RppHOrdab05dICIsCre2IpNNuNPnKSSEgm046
DvikDQzAHyX+mSOTTFBnPq3ZFgcsZNotdL+oizIEYeqETJZ2co4qb4aPrQqHV8OrGAcrrBtUHZHR
B+O++AaOggatSMLS2JF/nshulbk+PmdVa1AjVSzlBbZFCWlo8RjWRSb5RziBaURoxN29G+ZSeFZO
gyt2VWv3wbexfuffeMxcpP1GYU0Epx5zo2WZWfjePbKO/E6uIBILGtRe0k33QmawyH6g7MlU4y5m
DI3hjfu5zTUsiCVX1Tvt3iZpP+hCekqhkeYC/r5fF7xp1hJMYX6+DBtvU5Com4s1vcessfjTJNvG
c8egUa651NWoA7ttsfRq4IsDr3+8O3Tc6p8zI0OBEwluMaboVk8hCx/2tt1XVRMCNY7AqYdUrrln
dPze2sLxWQCSQ071XUAuxsZaSsBcdtPhDyQc87aSWcvFa0dWvhndqwC56nx2Qd/tdZrl652WXO4V
+ySIeJ+qHjV07+eSX5wWdAcfozIZ77XhkCxBpPQTiDwJ8N8FegBGAny3SFLzNNy9bTFCubM5StSX
IhIEo1AT7299m0CCeH28BPgciaKtPT2qSqIP7JUEpZAwfz8PlLlZZd6jBygvlzD8LJidScraUF4N
qH0DcJ2p+6CIpmfjhKh7Xr1OTH528pQ817tiPK7D+QSc0FIVgjKrUB/UkISIInGQe68jHgwzu0B1
0PCaXB/P4dM9FQD7xH3i7zgHgTUIETPqFctm8D2ijVYZAHD7jjWuioSUD/m6b7+VN/ZLjOY6WS8O
oG6s3DiS4Zu5DilcTKM7gyLwQnfpoToG9vw5nbHXNBjehCsBpfFeg9r+S7+DpuSPFzCgsPzZToY6
YMv4D6wF/A6a4C5XQJxxsxeICUL+YkytXY36N/x2FAH7l8RBi4xxXfNN/Xmykm2ADRBDvWJAbfMl
v7QTLT0E37RjITC4V2N44h49e4AbMf+RqydWvHPYl9hZSmgMhk5c4FpDClUsvr54Denv5802XpVG
vC8+GtEjHXWWJVjxxvV1re+QLctuEjhl8APvUzLGs+dqwwngcDg+UGJTqJPTLsebI1satR43ecZ/
w+IFn0YqyGD61xReIc1PUGj6pVzH1VlDeZa3MfQK3G5KpHd3vxDtkg7Wl6sKoPrucRqIctdN4L/l
YUosDjUMMwuFt7o4fmPrmGRh+hvjnJWxoNbLuybzLXn1Y//UGBN6n62Yf8ZXQwsc9yZCIqRMEifw
NXDyRBy6rqbv7Ay+3Xl0pKQ8GODqfuL649LbY86nvvU67nNdyBe4dgI0LXwkAuSWutODj4Xr0dOk
LLyj3SnGLYGbv3uEofc+B1z4kX4y9xLxzTYwjB8GGqD+aP01PlN7qz0sw/RDjQt5EGkIHVG4Uwzk
OpM92cCVzwjjXSMyhsCvO6FkmEgK1KCuvocoqYQiKZa1jnp9/mpZCj8oYQeqrGdqMC0SBPdiWHgG
/jaVMi5HExgUl0CInGDw0GHaPRJ8P6NSt8zsb14FuBfotlPI7BPru5CKXpw56QyiX6i8vtt3owt4
MQBzIi4JIsqE/C623oJWzrf8B2eFOMzvdosz5SA6MNUApt15KRG4UU6dsKu/eMtAaSI76TXRnww9
S+YPxZmesSOdDxiCS8F6PRLZRjQxCKYBfoFgLYY7UjDaEPrpiFP53nDTOo5lZgR3XoYU/UD7VJEK
9Sm1bpFh2W8gK6HtjPuBoc/V07Sql6ER3RMIU7ygq9bVEIElmIhxradnlHzAxj8K/43O4Rs94V43
TtOzR6e77uKTRZplPcKHHRL0gzcwEXGTwiZVhPl9ZQxPdd6FoOEv1OBj9ssop/EXyU1NsmGRfDd9
giQ4UDECPMil+rUqoyc/1XIH1TbfeoblUYzAO4KFEiFBsWGrNlevJPQkS5kSfkJM8s6BeT1CTMPf
4RxcWB3HnWBaNS/F2lZDE/xCg1E/3fimdFbXI6GFNNUPKXY962Sp9P3YsJSo1eYqXFdHZYWsrrZF
oBvYWR3UUmxJ8FtisXWzNYXY53GCHpGdXYZcVqNHf56nslHE3OOYiamu4DzNvKWPJPjtCJwy4ycz
/PAE3WXcOswVAE4qMb4RaoMuSrYoT6pACmbCQXyldj2MY7s9p9ksfjPSZl+sHDUqJJbwgbmD9tXQ
j/KoWlFx9IWF/rrew3brRH1tSZOzB/6Nnv4pPwJTvus6/guLjO3tJa6yxyBv/iyRcSTOTekoOfVP
2GpCckQ3CmS/362qYzsijUxv5YDhJVPSjihZTyUq3t6DcjzoJigRMhdY0xZ3LFK32+4cCdqfYgiB
qbv3S0jpBsnHuxe+vpVpBt+QmG3SZxzbkQP7CFvUHCxSSnbMCE7JlLU/ppjdD2cu9aUNHxgu6lYF
cAr/vN2AcN+yuKLvg2Gb84cF7CCzQDpJVUowP1lylXIBQSpyg+mcl83TTkFi5Cp2RDEA/3d6EOE+
DVmglQK5hPXvOHpgslLGd3Va4FUcfXuyUhdCLBUVGOC97BYgRcp76QeasDeSwzgDoXIk8a1IXcqU
R+sr20p9icSvBsWRUUDCQxalgKxRj1PushZ89LTeVjLXxJPYle5tJrxrDM56b9id91Av4Q8CeWWo
5sAKdq7+rJPre093BmOkQni73Uttonw6ly+Ago+4wuuMoMUNWD/xWjCrS0YxPROQu0y6ZJaN6d4n
Jk/RxbDvbxwNWTpX/kONx/Qwmqm3g218pXgacVaSdW/Tras3lMSOYS72pHevZF2R4S+WWgQW6TnI
2FEc3XVVrUzxkrzf0A7onxFeD7QRi/Kekg/8Z05IXj0sVTupvb14hW1uOUSHZHpSj4CoHEDatUqX
1hwwH0in/uxnEWExnNd0Jb1k6CfpvgNG74oJxx0paDLA4oCQa5AKdd20VnKLpzfyUB7p8L+segEv
Y01u7zOWoDDYrxvDaNhQACLUbf+jhj/4fp71Wt6tPHezfUgDRBKo35mZATfEgMBRsFeiih4ZNmpQ
PWdSi/GU2vP6pN/A+bhWktDgJ/7fMHglUdnFGp8VcoyQTUvWvKtl3fcXRNzOYX99tDDdpPAKvRMM
xaN1rGraD2/kySd5eW+5tOuAWjF1Mcb2/iSubJqKdUGpTyXazOkg2YTPK43BHEWrk8TT+DJX/6H6
gJ0EnwVIoKiNy9yJ2kzI1cRsiWtDOeiQP3VlQaieiDioh7RhLM1IR9IIJzyFUWeVxMt+dFcgAuZ5
sF9rc5DIZvynM7Ghej0mSrURHvsPm1iYIf631j4ve37o9zrj12N7prVAlW2q2YIJwIUjTzolVFVS
PPnJdtsX99ziPewT9oSMRaohdsEAiXYd+aLfY8ZluluKz0Pn99qopsEp6U8kcmAVxhn1kSDWXKc3
CK83KmloIiKDPLYGxCGOBeJaIp1NlK21mcApWmr7+r1Oxvntc6t9qSgeEp31+nrxsgcPE76ixWu9
0oQELu3vlPPRc1vw6b5bVm+RWbJWhebTGfFzLK7j8wzf+Dck9Nb+zFFireHaFu6Z7A/UIFn3sbBc
ImrXp7XZIY9f+iG+IezimgHDXcQWv94rZPpU0d0cpapx5BC5FRZNZd0z9VxZk2ydh54Rv6pCg9fO
tRDtoq1lzG9blJiw2UlCBgX3TLXM0MiTsL2X3GjKU94RArA31FCCGJtjcwTtH07jE+ba5QAqLulP
Ch3Ab6dmknkj5Z8d0hn/EapJi/uGV7f2bkMh7Is7CEn0+wS9TDlgnWBq72rP5Avcyz9EROGQ1GB5
FF5npYiqOZytM7Bujw/44D8TA9bj6uvEwx8BOsb/Ne5P+JZFhk3FopyqNqxWJKWwTTtRzO/29Eec
X9poD1lnxzQCg58zmUAfHwDHl0Ei0K73WbLZXPQm56A6F9OzglnRykLbhAKkCswfD44nNr/inDs6
SQzhqd1crLunFWpJ07BxjmpUAUxmaLC2GUrB52J9yjq6LVvzgElIIS9yfp/T3RgKm0wz36pvb66w
JOIehyMwXsu5y16OmfoQzLApwGuYqGZIqh1bmAxDK4i34FwDHAR6AKiv0crmn2Q6AnA51mJlFcTX
YJC2ckFWDwXGsjb36fZSvAhs0YqpE+otVsRb2wXq1C9jGXn76Zer4asaKgkSoIycQSH2cQdOMS77
p2jvYO9YH2b4Ml5bvDhKg/0AkmMzQVE0sbUn6igQ1+3AF1b7ZtNs0ow4IQemU8P+zNpD7xwp9Hjo
KX+YN/wc6bonEJWYf3Bgxh0LGBhxSvdnyfP8hqyWLnj3JWpzl8YQnieUM7B3ZkSVYtEaIn6LbCVD
2i4jPrRTmqRtYa6S2cP5QFvK/k5q6m+jMQPLf9Dr75LGmexgcXe466bSkehLPQgJh15hS16a6VUn
ccvwUezhucZqBc7uM+1cYgLYva2xki3N0jTMuiVKhwYSIb9BuVUpdf1AOm2k/ODtiYRdx70S4B4r
KZdnCDnqKqqbTkwl4Q9j6ghZP9PeTD7v9XsPq6U9HGIzOKge/c9ypxalOkKXGPNOJvdYhx9TAqOV
7paa2tRBMtKf5+j/aAxgag3OuhbJLYzKxA5HLkgMR2xD9k/PJmrBM98N3CtI4w+5wDXEMOp9oa7E
t9Uxgy3HdSHsoyW0wIuyC86of1iTLiPOSXIA2PZuexyNvOT5AGNT53JFOP6w5DwaoVZ43+vd0pLE
W+UIhjMJt2V5u7Gneq/B+jpjnw9uhzkqBqThMc9SeoagvB8FbmYqfAudKVukxbP3pXSkTzP9mFYi
YXN/7uqhA6FeXfobdKo/7kl15JaMfy83xy2w0gANNCBYHt6T6AeM3bC86EbklU5hfvnUEkwgFObk
jNjKr/+HDAi/KTEvXn2RCb6bmU62TluX4rZmBq3H2L9jVFpfmxeuLRi+RM9g/QxNNlF+ZFCI/V0+
BVeI3iLdsVvqFMUI9ZG+uI/wiDazjyAUox+LTezke/FWNtH7Nqd+gyMi80j7tHAzsoHhW8h++iOt
gLpTHsTNC3aoRFSaV2HIUUinfp0NeqEZmYHLaoKbd4aRSNaisw5FZC2klOqM1OrQudV9zHK8n0Yr
OUEHAJ+JXcuz2WXckQopZ4KWAxalNDpglbibghmdowWhmP+13GJK51y7fMLgeBWw5aah+UZcD1We
jZAmPcp7jTAeF4mZ4IDu4LxjyjstgP0jZudh7wjRIs7Sac1rDplP6zgr6AQsI3M4aczAnxlWzJGq
zEX0MdDv+oSAQPFUGZofPkwCyQ5YbjondcFpo7IDeaLniBitWzdRaFY9kA2El2qRR9il4fw3jvmN
KOSLrLuR2odhUt6T7e0mX6SczTFrhq83iWowNK2MMxu43yidMTVqhe2V7mzyfTVXwnx+0I/CbKGU
NSYsiMR9O9kQZb1c+PMaEjvXddsvlIHXbkd9x0bHVVgWLMsvmvHI3iIAdeiDp/WFZQxQ70M5Ao51
vDLpfGkBmcMYcQ8/i5vQJGmOEmCYKeeA/bpKklcaRMlhtW3b+bChSHgLN7Bu1XE6FHN1yPIaBlmP
U29kaw0XDNGLdoei8lRiwHswzBG36LjxrUCDDOorF42JstXfcvQEtHtIsDK/YmSe7wsosKqEWvtb
HZCprFtAOcoecJ+wpPmDmEaKzfGZEnGiucHtFHpYcx7eMrzOwUUjXGDyE+G6yqeQdMZlVwh+1zdE
rp5ead/KTz41ClnOMZ058XdQaqkcgmOgCSUp8pYa2uq4fUXRjyiXwz7iT+Yz4YaDhBWA+7VrEg/e
U/UrvSa5CrX01Ucg+pV1WPYCIBvvYi2/r8M0CG/TdkTt3UmnE6uHk+Wz0m0qVrtXMxRlWuKYALMN
PjdgTmtbP4PMtPGxGBcgPzEzM6jE+nAUvgTUzNkHAUr6WiApLnERMxUfnO+t8xDGrKjtgpH105Qi
G238v0TGsiJwkfvf1PhduzLtNqekdj5bGYsyjylYtPMh7R8pZNV2/1cPw9CBUwp4duv0pwECdOVs
nUldrt/ZrbTU7suyQ/fuEhbLOqCJ5QoU6vQ7ruAI4nXogb4tE1H2XlcHN+OTHUxuZOtj/CQOITsx
XcFfCptIZ7T3JZHVtp9VEhLt4hsoasZXi0zFTJ66g74f94Yic4G8hsF6Awsxwahv5hUDhZozinvH
9U2wO8s3eusb4IXJTsVXvo3PhKaSJ45EaHR7YV/ixf7YNqv9KiJEwm4EYFXi/7c7STPl8dZ9LpGz
T41lJ9oa8UlF625Xhk3p9Qqh0h1aTIe/ICXYGCTAzb4f3QnWlzIJG3PBHdmgIdMG2GDetiZ5cYwi
BN8L6RMAqq+laLOfu0WDb0x8GY9xc0kQxNiQkRSqvBrZud/lnRU0T8p8i8YOIzI4PzkOtEdEFeIb
onMmxZ3LtpOBFpcgWKxHu3h1iCj6t70aF88E7jiJ8HX65OIgThBDG23IbSLpzpVHPS0+qkU3RMcT
Upr3+2NQJj2tGCc7SJRYU5ymQM7OY3FrtvMyuoXkdHJna4tzbcvJgsLb+rKdx55F4aksi6feNsX5
FnN/DouyNdvV049u4lHhOG1XRT74XapmZ9wEnpKBFO0HJP+iH2+FzmxENpXz4uOPnW0343tNDToV
loQtX96UTOerDp/Wcy5LXZCjzUX9vULwRrKiopmfC5PUFyHB5pbOA2r0DJTcNYoBL+RYydzGCwjl
1nCK5LfyOn98pFvaONgDN6O3KYcZAV3cD99j02ySkgMNJKbNdfB0HNo2h7F1GBOpeXT6AO2S0jo9
ZKPS1NPEJT9JYWQ4jqNo0eMZPgiaGb9nZIfoInUHYMTMDwZRfD+Mv8AQsnOgZbVVOCjUw8AskLUS
tagT0eH7rUAEEvReR1m3bRzLWFBSqDQXPZnz6cXlNIreG+20tuyge/2z+nbiWv1jP1pCm/rieF6X
CSZa01j7JLzE/dA/CPowKN4I7uF1eZoLZO7KOqEGwItfOLspHlPGkGCZ5EmddA+mxRytunVuluJX
ENxNbTiMy2RZ6x9VOyV5RhwcmZdX9A52QsmTIX3Pd31K9yv6AnKqen3PbHiUifV9WqpO1vSFcamY
0fOUGaTeABdqZHd/I4ges9k/i+ZR+SlTWrwUm81OdYUaM0lbEaycK+mdFjQrEZ8iVUDPEhM8Ko2p
dbwVmHF2KPovXhqV8s7tMYTL/f4gVmcz3DHQHfsUetdsIt1RHyoW3GHIbP1gUnbKjXRxoyb0UZeF
Sm6aD0nTE2YvXNdTF3h65yZ2tTd38jMjL2R1207PrOW1DIl9ftRr2aeFFlT0oX5Xisn0uwscisYt
2VxtcPtex7DfxkQg3CaC6oHJfS4NQRNyW/bZK+px6T6Cu1yTNhcqW6Yz8XCQ6TyWV/kWTevE+UNs
OIoiijg7YP02hX4s3D/ahrCaEX7cDov2+INha3NehXqqpto0nRXkmnyWnLPmCxyp4jqmrfjuTrqP
a+WceWLYVppmxlayOI8oqk5jeTw6+TtaFOx28S78uxwWF6BSTV4PvotfA0rjFpaEUl+iy8mdKxdK
2pV4u+g21cyLGsgIbxq3K7YzI++1oJwB3/c2iSb/Lr19PuCTLPxJjTO+IpjVdA3gQDakFIYE6skm
1FqVn1KiWCuFO24JzBKUAzwkFU3AE0xtFkbFfyArkE/3e4vyZZmiqgMJNaapNqKBuYpLke7tk27V
pf/jIVg0JKcNSZ3R7KLf9e7W4Yf4g/mD35rup/ENrcMRFuRpxlXy4r6rwfgf+5khEEBHMMbBic+C
gYjd8K5r3BcHKcIrdOvgyW4y035HOs1hu46uf6e7ONcXK277/vHhYZq4lgsOws0zV4ahpdHHSxp9
JANOnEUaPZKStCFh5K3KtQQTnBKojy970IANIJfPyrQABA19dICSp8RquvdJdanweS5m2IdpId8G
PV5yxHBM1OsANNY3r0uTMzlDISEYe6elA7uu8VLhi82u4pNQq6SKrhkuOIg5ySukTHPdKSmEXNNL
5wUnDWcZ031gWZ8fVztLPf3Ab4CZOqxteJGJiYP2tCsujb4V+zgGZu1e3HM4C5AUGAg12i2fboQ2
EvCfMBZn1+iQRyK6suh67BxGohnJHuG2AJ12kEkKSvohySyu1IKThENkSO2ud5TzUf3Qh2MXZJz1
odcCI1flxAeLrA8tj46oHw0ImNa7q4N6h5tP2aDKJPeWp2yKLruBnuqvSBZwn6C1T6VmxPPVasOa
3NMcgIyaZZgQh5qodQlqEs8Z1DO8aYvn8nr0rkfuwcZIpaKVS5Lny4EvRIdERRklOozgVu1+IErs
3iPemwmXVkwjCI3+ufVp5uw56fi0etDTpcJMjAvfO7GYSLqvu6k0zbxYCEVMSylODgeDxZ2xlWCs
PUiJS+nsTQR1MXkCgo3CuTj25/WLuk6RXgNP4kDCkIVW03yR0EcqARiN9gg5ocm0xcuq0z94OgA1
lMf3ymXUak6WlZqfaPH6EF8tV4j4JPKv6FIoTeFlRObpfbIItZEblrVqutFdDw51PhbD0xsdlU5s
ZG1p2vH7/Ju9s0i+E1eNE7NLFvsWa3+11YG6AiJlD436GPXhVLOlFS17uuhnoE5PUa41JNUerD+1
dvkOhUNXX3vJXGFXB8CZrd25vRCdKOBQtPSCWJYopl7+fMYLFQOVOvu9vN2+Xfi6hYz5mMrLqQwv
d7vdTJg52hQEVM98l/7JglGl1vBajcMTq1c0aAbu37G70SEGZEqwCxMqmjJuNXVLJE5Rej/gLdAx
KlHRrEasfhiC2cYoJlr7/Ukthjg1C8M7LXjJh84lgs/hhngQXaEpBthb3xhquC8faq2TmFN/mnPh
n20b0fv7yumlAAaEWfCrrgFgmHyqkVE8EQclOgGreGiptWEggnyhnOrwjCiGDnmdxcWy4e7JwFTL
3T92Z96yaJjRqAh2SfLX23QBhapBcuzTgEsBPUG66QfkcBjvmoR/mwIyKt4004NYnVuM6abqpZtT
nCmqAnQhNxTFgHBtBbwUK1siBrVgTOkARtOmWFGMeMDkRcQkOK8YFa5ArlxEWQdTZW+DIY9kf4AJ
nmG8+dsEO7uAGgXrrtjAJlGDvdcycQdJa3nYAkTpBBz0tuZZheHHXATLrE+1YJ4weKA0Y1OexSbu
uoSp4YOXw7ehQtqSO3Cs7/Nf7HOC5dMbvzAwRy7J8yraMsUqfpjdC9K2YJEQFyJBRofWGARR8esf
Yhhp05gHtvhztOhi8YWA0Bq4wvEci89CSKkg+2osudcAEdWxvdqeW5lmHEeAAhxqDAhTPZGV9uuI
Smgy19Ya9YJHEU/n2Y16wCLc7K/DQZFNdvwvlwxhCr3/WEycqMYylEYvkJmtEXhAANes5VpSpO0Z
9uQENUFJtxfqdnNnQFKjsxhQw1/EKbrrZ1jHshql1ZFB/1RcGuHJ9jWCUPo1QecAgUuftGHLSxvI
0VSC8+8cxrz4nKrhYj1EtwFo65Z3taa2t3UzCGCNkIAW6qsBgHwIIzLca4mfrTkNzhJbTMtpALj+
5BQw+e/SdSQuTPSHeGv4myQdEw3leymd30AMbogb8v6qaeBFwhordWQEHMnTpnu1x+GdIA/hw+5S
7H/yDzA+H55XWVIqfiEBhHUMEr4JnQDK4VuV+RVVaMFRCbvQNrIGsmCJtZOPxaPZztaF7tTVqMHA
vQNkYsGgfTdjQ/vQdIDjuT6SwqgfMiKtozzFGsYId9M5iUG5sxRCpKDqmdIzE6B6K2NkSV9OuHLE
i8Nb3eEQGK6oS/HBMmKEF+XrQZcsNfs6S8f/fGVbYkGib6PZjIL5+BsZezEMPYNX7Vp8m6NfyyRC
fUFYNX5Gv/q0dOynF8LzxwYv9a4VSW6nnR4ekV5ZfzJrrsq6rNgQRaIfqW9NE+JJlhXIAqCUeMcs
Ul8LOCsoSJgI6HzbTMWcjxBY2fE5wFqniz9MujpbsYfXRSlyGuObwvQL/GMSnaXNetGkovoo4mPO
0TTg2B6+UHRynJd+/kAWnaPIH7IW4HpUjELgRkhM6Zr1pBrymu0UEuHGAdJ2B6d/tVerBjIQA5KM
my9lM6pw7H/+WS4BPlSv4ttodUm6ntifmWNQd4qoe/gOQulJ8uryNlsIV9yI+6e0ERpvG1fWbQlO
xa7nXMgezRza2uAL2aK/l5qXybQN0acaXKRJPTBS3rpR5+Sa0FLuIMFZCUreZYXOGZ3YL28Ag6eN
USc8cQAXAOI3LUZQJoXnjbGfwyJS7GX3q7DhIlOJzevnLT372Hq3iCnZv06xskjFqxOPouqfEfOI
aXB+HoBEM7/h0OT1YOWJ2z1EhukofNpVjo0Ci4bxId8/GaXbmLllqjnp2oakQ/9bzhggjLhmmrG0
UPsU9clndUV5Wrs8Dn0h5OlmpTiXuPWfqFsJR2U3dLIW+HvPMs0iRIpsiuC79bLUj5Qe0ZFjMWfW
O0L5I87iLl1jnXqb7Ev2mF77OWm/Y40J61S/w+76uEZlL8vI19eNz4mHxTZmGJPoyFxS/iV2sZ9X
qYQeqrlUXhStkFQCDwIxENYvj8fbVx2nGTRtiSvHWJ5RReaTBrM86+Sn8ulW7WrICVDmoYkultSK
dGX1UwvixIyAhs9Mhf91xNFtHb97J2FX0BveM9P7fO9Wta8PHiZICX+npV6ft5A4zTcVg3Amf6B6
Gd9UtuNSHeDnhVG0UYPlWUzwlxxhdhTIMId9I5H6d+5uDOqDZPVDySY43Bu6BIdm9nUmSKM4cEgO
+KIx8lhTVkyDpgtH9x3YS5VP5aQM86ll8V7LZ76qEy/VRrsBMAzz6qyxieP6GE8kemLxo4dXEGb1
SQ8dJzq+exWwSvmyQx904Sw+67loUZSgsrTNdAbZtjuQ5oRYCKJAg7//pGfdSGyEiC71uoHS43BO
zOTwRg9OADxfCs6FCRra9nCCe7vgc+BIYwaHrVdd6dllinF+x5ka02hzpl3ivnYsYDSV4jv65rAp
WXbzgII5HZstNXC8HosSX1DHocIIMGsSqDEFjpOTc2d58h185GGAgLxf/2Y7eyXkyzKyVY7Hmq6e
tcONayE3k/dertCNxlaqc345G6MsFQnrcIosvZbS/JRnMHlPme69gQubiC7e6l9MJxPjXNxqppYK
3bf2RCQQkn3WjFSYljuWA3qvUVlAx5lfjAbkC8eCBW1Vh9htxp/hF5fzYQkHIwAANXJYUs7q9GvJ
BiMQOCCmyGJbHDXt8yCS4gElcpCaQMBQ1eLXp02Q88bMrqnbYn7eNkwSa0l1K+PspEr3TtPgL5Cn
UFH/ls5prYWCU3pQeQSLaBL5osqV4pEHmjVS8lyzg/hKLKzZHAu0MTbK8+6qhjbT8BUX+Vkc2HqJ
Qe//nAXBWkKSsqsc9H2+l0Z87qYfeunujOSrGXC5d6iCDoyh5Fds0F9IAqMOcvDurB9oVGFfSpna
N8YlaoFPM6CxmOwEpUZRMlvYGGKpaEzIWK4awmam+uC1mdui6E+ht1Nzmsh+d053aC6YUvSiH+dS
FTtD159dT8APYIgsmqfSCtkGDeQZSuVjXP+QRQIxC9Z027DUtNa8C1OW3YSyxPqIEgYvl6WvZW9S
LdSoTrHpmkI7P3JW8bFAxrcrYNnI5wV2DIdUBalLj6de7gmx8O9qw6Wq5CijiuYgXp/JBLS60AkE
wSel/XM59qkaCcDT2GV1o7S3r/1bnxmEcp+6cBub11T2r597IaBNNNzi9RlsLC+Bu9X4RK2tK4LC
d0bDTYAz5JMqK+FlezVJb+9l/6uRSu/UiVy4sPkdZQqmEMFVxWfGQMkrhiACTTgsOxP0kMNvRWKh
M9wAhDu7yIOico5KqzVIxfFJxX3S5NzJlnEnFlecnxWGXwuXYfS+JoojsNIr7jpMbdZqgPBRJHpx
AHXsixojMEAL456qJVJ1D8lwZrXt1vpVn4JevyycLrB/8Nhv6ttPyOAP7G5aBGiBInG1/cZPH01S
Q5/rRqExFUYz2H+5wCnlo8eCrJriMIosZj0P+GKA81pQUD66RXt8rNpxR7HKY5nCrsNRSleeFIQK
R9PzN4bC6+tS17tATqIdHp75ykjUJl4e8rEG1WRA64E3gBJkNfG5AOF8KR/OMQfYvKssuyXsfKZg
vjAKT548CunIb/mYB6XPsEBjOPf0Dls+a43+ZzDfCG7ofZLBjoO8AeDCgaA9OcGOhoEq7zAhLKI3
0c9uk4eCCbxdtjJT1EsEARtgdP4+hUjtq2xQX4mQbuprXw8QiS87JXdS2EMK74iT6cxIjpBBdc6T
919yNkiZdnSjIs0rsSahv2SYNt0Z+d2UXI/tCdphvIYWiJjD9WhzjHcmojm0/ibAiGshgo9ljan5
Mv7SP003pPhNiVZoF2hYpdoW0kCpdVJNXqlnndOSvJihu746XeshMZViwb//X62YTOSCG4ZRYbqD
eCQeyd6KVWu48kDOdiWMCddWnmZ8Nbin8Sh6Esk3eNYVVdLKrzLvEkrQH5N9v6FrnJKKLH6iLN2o
X5bewcO/9CaKuNO/9nS/b19c053ImSgiCsdOHq2ry3JFRgWvLV8Tt6v/01DEKFzUeMBYBaKF8fkb
gmPgYfAKXqVcznJacx2x1lv9D9HjHLhqtrdeloBGecuITYeJpUy9gcq0Dw7XmiB9VVIKy5V8clMP
Qpr4v8IYBlF+FGFSA+6LiMBZKKwEnH7s4cI1RogVPBx7AcBInkBaBTavZXcb7mNbjyQrCYD9N4H9
XzLcftBx5Pyv5+akL+BqztnwdGG89N3nTF18LGn3WAgcDc3HdGlEcepi4G6eFjS5pYrW/49rKsNJ
MY4pio9OBNlI5Byv3LI90RejbFAK/bp9Vg2X09LW/Ognd8HAn15nT6o8bE78PET0l7fRUJXfHR5n
91hnldCvAskyjVfEZfa4qr5AEWP9kmGQvhq224kvVPSP5yZuSl9ZFXsYG1SvszoMsZxaUtLrD6Gk
bns8vN0HdgoWzeSJGcym7D927Gxj6SGkjGWjQenFojAqGA91yeDbvKQ6uYZm6LhCdIKXZssXklfm
+jFTKXehq6CW1fLKiRAzhCdOu94ezQWYMh2Wk3ort7ehGONPK2HD3SeFdXCqDTH9ActflBMBdX74
XZtfUL9rE1eb8Wot9rkbvU1uUY9Da+BBd0diPz4wKwdOAAGwFH7QPA+8vHx2k+lCG5nOn0v+49a/
zZvLbHtCAhrCI6F9qnOoFKqlhjbv4vIhFwkuiYz3ABtz5Us/J9NeHOlaNsxzeEYKvZINqyo1jzR7
iDc+lHUt0ylt4FQN+mHUJ7+Jvyy+/I1PbUJwNbfA/YtHHuCBOg0eLVKODXRAvPz6L3OTwzAJpOjd
uCdj+vwQJ5BCOLdaf6H5IMy/r9ZVi+XpKZIn7mKSEw4ulW5dW9piCemDUUQo136O86epEqM0gzp7
BZh/nxN8S0ELisK1KOFdwsidQiMdmml2l9cwyVuTJ0FUUs3aJc5jWW6qMkvNjBlC28BvGmbrLKJf
y7ufNJLZfpJJvODk68NPSKqtckjb5C3eAnryTMgd+zbf+Wtb/okvnGf+ysik5gotpwJPVhHWYbLp
uW0+OtHpbVf72o5epkvuXBqKdTPaRPaijAbWjhjA6bSGnnvNiCebtfmySHzOMZgI/A2DqZ+seF4n
7wvF+En3FQS4pQGf8IbJp6FGBVXNQdNNJFhq0en9qlQob8FV1vxbXJSgSF3t2V0372RPKy0D42Db
rFCCtowK4FHHnGQBZJWwcxchqIpCq579y0C8KLYagEBF9/tCU/+zcb4yzBREeokIw80lroc0KoL5
EIGuSaoemzb4k5m0sRZeUy2SSbNPBFh827gzFraX1Y2OV4aXUsjGQEq0OC1RS2Oq2LCX0PBqNWcX
cB1lJmMugKE3n3dYA5TsOXoSPJw3w2yXab5B1mJgSDGbw9C1MEcniQErr7idHRxZj9Bnxg9/oUih
MsP+BbUzWslxdPlZYIj6Fzy+Ge/2VIgi51zHtPueOSOe5VWcrkWyBC+oYr3zOA1huhvil0v6iFH0
/C50169aVEHwanc+ljj3vN7uNMJ1FYVtIDtA4lCbhx5GRHLuhnrxdVHk4fWOndwiuwt2RBWNHzGx
By1zmgrr23cHvICTGsc0nCVVifgFFfthsdbTzzoDlO4xk9WQJVuwHRW13bOpJhTjMA00TcFCTWUm
kxLccTPzqMLcq3oiQDFzdzFH5yQ08hHo/RaGT8MlkBkoWbYfnMtbGcLo6uChdCb9lyiBgTCBnj9N
LLGrTbP42TQjf/eH5BISnIXXdqpBbFmIBEcS+ghHGGcV0Zcw1dEiUJR4CWXsVQ0fEWHAZqVGfyyf
U0fSLF5NoxkApq+K4u9qm5B/7dVy1qBieTQ4jutWgGoVNZDX/oX4LFbki9eYb3wKjL6m5BYuslta
DK206ss8FMDRIE6rmnFIrDKzlWwYlv0Z6+NQL33epCR+qi6De+p5i/Futwx6lc29xY0IDSaR/d+5
os6SSt5Nj0oytlEvny0rWUnFjGHGNrZgBoL4k8Hu2SHLChXF1VPhXY1pI6rVXM7cMC2i1pl8/Onj
F2f1kPTdjXyzkYmsjJAlJKiHV0fjvmZg0iiuoozzvSui/BB9RaAfIXlUxDV4iVW8vrGNtxlxvJwd
yReU+OjpqLNHqrU007BxiZc6OiK2HQir996biKjvKve1CydFWXYu6lEOadjjxHu5hA24ap2j9LrF
hTfzYwXdntCD8U9266Omwtqz75tH//77cDGnOjZXpMV7pQPqtz79/yqGJ+cVP9D93E4Ll4n8A/mC
PVEIlEsBxaROa7nuw3IpxMvmgHOL5u3uCkxunqyY8aQ3RwmlyIZTsyjWFXLDSOfZfGJsGR647aAi
sdHWOvOu4GzlLIP2Lo0GbbHAj85yXdvr9Hsm9hKsWLZ0iArVtdM1+q0bmxg0lDoLKysstbQxC6bX
88s2oPAoasPJJeeqtSbTCLdaa1z1m6sm4y7Jjuug7NgrZy/mxcx4rFFjsY1i3qS14GbM6dRpYdYf
Sa06VZdXnhs3yHYQeOBvy01nXISfgHN2FrL6hNLj/ol1npSjvdPT4AUlkcBd+GrCM/PNHeTP7NyE
PNdXn5vbM6x/WTJQQRW9c8tXvSip+PdahDpuRTjIZ6NldBLtHdb/sAlc5qTiH2g8AxipIZ28Ry+F
CPPgICagnz5ckxuYBMoaGWKEK/PdJqV5stTw7Jb1jSBZLnEVuUVQ2HF4qu+gCmETF0s6gTHK2IXQ
O+2Vk43IEKCvcMf5APj7Daqf4rIN9+RRApw5VE25bliPFNjqufLwSqWZmk/c0lMTNUkqqxft0iSE
b9BbERN4g+4yjPWeRc4cMOFEFR3yqlZGH+GuC6Vr13EhEfJDyKB8+VQKtnvZbXmG5l6co22Gp8s4
KDYSXsrxDxz6sO81nnZ/JW2h/id5vQdsGmD4YoimuhRbxKC6h4dxHU5ewd7XSW5io3b9/uP4ZOKx
DduVcbD7nXl95SPhoerPJ/Vqewt2qN4IpuEBThhitpJVttwOeTxAErPK1oc7niFtTrgsR/WwzQq6
Z5T3NdrRAfIYOmTfGQcjSzD6gDvFCpkn+SyhYSYEUXvU/dfIhh+mEjfs7ThgzmHezIyi+zWNhapm
rvN96shqLlCicHUKxyHrxMlF1ofGR2JCD+O6s67YaKrjP6gryBXsKBoNaD6JcXXMixoKkw4IOhyL
/aVkeBPd7h9xP3AEZQypncpDpG8ofDImzAuKSXtNWhdVqGH610LOZZ6j1RuQccjCoOECGAXdswDv
qc7/ACHPGGhGE+kWUhKhm23csvR7hJJibj3X0+3M59HS4QdU8HrLL8/qgS5Lh5t4Wz+ImQphseft
mUaxkcgJqnsm606x/AgP0BL6m7KxDXV8jw7Fbg3YgsUL874rUYMYYWSYwVkswCcfqZkQ40xeIV5f
bOAny+UixwY9L/YFBhG4XMuwtSGjioJ5Y2zSvZ2Jfl6sbcVmDwW03B8XEwxLM0wisv5/bt6W5gAK
I+weWU3tGUYg2jvybRMGVXhTTJ4Isjkbl88/7pUvBK1ZF75Wghpgg8VIX8Sx6C0hZka0ko88nEvn
M3FCAprqEJ2OTDJHzJfDDHX26OtBhRd3KFVoGJq7N8knnBaBrU79Iej8I3RxRaNjnhyGp5Q6PcbI
ZnQYKNJCYrH4529xM6mTUN/SDWwjkwHpM6hyixvTneHhnpcwZCrqJ61g4iZjlhqg0mG7a13r32UH
yMHtYL+Ch5d+qVYSuoNwBvDLEp4b9CF9cNubcjqkgCXVoCC4hGB8Klbo5skX7W8ULb9jHnTqVkgQ
JdCAgGFSDYbGCnlif0NslMh16h4WGKLSLAq+R2yGNVRFlvNVgEf8WVOU1L53+4yon3UHMRa7KqSP
MbNSNOc6StHr+gk7R7RCgNqJxYjr4d83Fai+UHrmq9JkK2SlzDJEEhL28SoPf7AsCXj5pxlknkPK
VNbuGM7vqtzlEbVblKDhXKQebENtFZuxHlmKG8OHBHTRmQe7441VlST7bdGSgjjqK5o+s8sXhC0j
4gud41VjEJSNwVMiFoyCSf4ocQxOHJivGdAHiOR4UdvhOpXazIclpHfMuNZ4m5xeeMbXldlVq26u
fGwgBhhMaW6uMniaHgI9UuOdz18SxTCmvWz7uRBAGIgydu+x8gdFTWft8ILy0YqHfh2i+tFKBmzj
WUZ8pFyKdxJA7jck2UWEz6udf4hZBp4C59ioFipadFymly9ShO9s3SC0CNdCONBX0MyV15C1urqJ
PmLm6ma6ZI4LPDq+oN/DIjSto6H6wFo3AD7UWiwDg9kpk8StAu+pLL9AoIfuroJbQB5KokO0y80e
Rkqm5X80k+xKIXcBvlGUkk0ZbFjJtIoWOP1dfR1mZUaKsUlPCu3NxZx6NzWhB4D+v6GZZpopfuxl
D7njwpu+JzjqChaW9HizBRiXmwzkUCtisFJsHNxKwl1ET76W7il1/+SDL4s/ZOpy2IQ2JO80dtCb
dis17mZyFqHnuxx0ZyDvGpBTwJE6k9IOQFwo3ovL+cNSppu3+ohvHowBlC7h5/6nNp3iCV5xMq4d
YALeVxPeu4WWWQW3r7dCnwpW7BSCUFz4ObL87f+UAO1TJ7+SZi+Rt1YuA09yXPkKSFOBgSYsVXZ9
1JyodNJkOtNGPVb9Bu/nCYNXs34JvltrA1VtzCQjR6+2sOeRcWobDe6JyVpkIftTDf+1ExOQBRin
faoLkCUnKVAUZYXbClUi+bC4ee984UQKi+IGAqL5nGUf8+ehmc3az5ntPmJ/Lff5MUWerSS4SJu0
VAvzzqM3NCaE0GKUZdOSAcSU5ZkA4k+5f8VMnSgQM+OJRken2yHACSiUH2v8O1Y6E1H/Jmna6MQH
q7KcGG1CpmOWt5kp7+jR2+6Odatw+d6N6ADptGjH8o0Y/0MTQLQDGpKnXEbgYZqQXrakiQAEtvxa
toyj1ePLRXorb/VR10nrTM5BJoAhhvypDA4JGJCoLgx+he5ugrfExKnzj+kWcycdvkvUASzasKJz
n+uYJs+Q5FYGJe6OJb8fcNoKISzU9Mv+RhrdEzVINZFyVqp8jxvAlBSP7C43pWONpzwBrd1Cc2Ni
Y1BIjDH4eZszuMSyFbPhACFIa8lmRGLQPNcD+qtyuv9qOGOrQarEOg1nYm3KfT2HOZxUX5sRZdBS
Pgfxxd+fJbXjxxG6+Upi5nVSzINa+kDVekYSYyvHw1106Agb2Yjns9yeXwVJ6DX4yoi/KeYBv9Jp
metp0Ec1zay69a4EGbuP2L2JPjPvw635of7HPbP9KwBWIVNCijiVAu4+8UZFeRgIuMVLNtauVX4N
MhUV3fdVhNc4JCFb/JS56IAx+6BrSe54tRVa+q677u6ur3VI2GYWPP0kMXBj+EOsA1QqjMtAmMcK
Yu1ildEekxtdsgxsZHZrWf80u/ZEL0uB4uTQP+93iGxr/lJxXU7z9m2zttxEfu4fa76t53NonE7i
1v5Y7NRMHrYRUjJXlu3Mo/uS1W969saVrt3h/pGOgmHp/FH7HlUs9MEWQNrP+rGG0elJ61L04diC
oIyQqjLhoe7/M3QxjqzCM7yUyf7OyVJL2J6rK9CgMApgP54Uo7AX34rjei1jXYPDfpmX1lIEECKy
GyCKLvi2YwBrK6ApGgoqm8oweIFV/giK4x05UTXYw/aElNDfXF6ui+17/CCugTI5qOqpvKtV5/SL
vcziThFUvbp18OLGzJ6Jv2Obxks09JOwyfhhPLUEJ0tAWVKMGf/bNdAXHQwtd7fqxQ7idF0hKC6u
4k+Z9iiIRwCdpREk6jppQ4w58TFRohBOadngvVig4prbYy6L3UChMBg5zvpKVDDJzaGGA+1aHwGB
hpE8DJrudk1eoQJZBvElqPFytL7uT/IaiqCgC0wHGokCPO4660MmWfVL2auTCTZ7gGpj+rcUjPqH
f+D4zapwVbXC/tupG/Vhn2n7l3FUt2E4MGqtMwBJE35XxHL5aKG6kCVzM5DUUMRODHMjuUWpudv/
ZbpfYR/XGJLrT9omIJd07YQPX7ldpyrVzmTK18M6qwu3aXCsDQZB2a78xQkLOOkO69oKJNT/SSRr
Ts+eJ1L3JF0Op5L+y+hEDaaIL+1UR8Pm7uOiK6Yd91MX+Jes1G8AMPueW9hQUbu2QSBCxeVUhrbA
JFg5389Rgsowg/ykMbEb+A/3CwPn1PyCKAXhNIPK4ZubYuZktwM5mRxQ4UYb024ocZ+kxqOHEiMl
bW8OG8S0JNsx5QLrqTOsR3KHLLsRDuBIARuH161FbSz83pDzZiKDqcZ3JsheYOhzWGpTmEwPOrGR
uRZSRt14LYNKe7gRFCBveCWa1GegbcF6apL1UZtCUgczQ4Ur4xzkWWwBAqBQV6JteigzlpfQLhB+
iMaJoV8a2pOYoppqnc4eb6ePwNgA1c5iYnJK3KdKrEWocKx9QUybR2yS9D5Na+6BFt/w5HqV2Gwu
gjJYhPgX1grOggimiZXuXPbBfiMsNelfms6D+Su2FClQ7G/uksz7EPLo3CI2GyWp0jKXHwMDe5PS
cVROw4naxqykp8kuQguuzcTEaPMiWrZIBn/TazwKFWQ99GoQ0+0PIvPNqWXy5U8BJrvHLnGlKQE5
14K/Rboj6I0nr6MFKmT0KsRd+VPpPTN+r8g5eT0FyPbMpgC2YuIwhb/cUW/IOlYUmfrGFJ8Y0rO7
B6Dp0Lq7wgUOxrs36+dwsfPvK+VH7UJsH0/FpJi1EySJYbcJr0PESGgLnYiNgBE+hm5w8hi8/cND
JvqkPkylttBnt7NvoHHVb6IET9JX0kVtz0ZOlyNOg6+jIzBpYhUJ0fBJN2zqRnROKtXCI/f13PAw
aCbNGMUIlKFQlsMpGOdga1xlqhh7sStMOUo7CwH/XvxXiDSq6HzQ9JPczFLb+yVUtj2J58awei1c
SQDcByvTGgp2oG6VqCdng4uwrp0ENBs/J2SPHmHwiywiPaQ6kX6mSmhuXnREeSzTbUfKtNvoB4C2
11XCvb3zQNViJWWYX97tNs3q3VNeFlBtlZAPmAagl4HM6uEEBNWlRhtXwnwb2YVENrow4EgKYF56
lADXyovvpvyWR19Bkc1E8aU8SAU7TRS7GDphoxoe5nywPeQiWPDodJftnnVLkYaGHtRdOR64bVF4
jaDx6lURFegCdBJa4mKC+eG5O8rxvrGi/1O2kV+d2jcBI72Lqbs4ZTf/ZHmPkUqumQDbH810mCF/
mYAb1a7sjYMruwPPc/IMiluhoUqtPWJvHRNyILTLi3nnmKsyrBB46ZSnxZoGw03rZ+xisd+7iWhm
mPtU5z+gw5o1Adi158C51yGuL4ptwSMrvXig6WcozzeoOgNRMnBInP19/UrzAJEIhovnmMpCudpc
7afqbYz0VTRSqMWJuVkc/i1htgFhlMDx805jXm5LUz5SQl7OZxg90YypIarf8lia66O9wLAZXp6a
qDTS5tZYtENpp2z9GvaAtWB7iUoDixT2OqxyDHHsEh8SMsSmh3XzPfQDfPZcgiRBP9Vm2ngwKwMW
QJNFUf/cJJwuwtd2FkzeZ0x2xAWvnuClbxjVaRsMmv2/G2MArRvT7Ei48B/tGM+ZxjL5q4ZCYNvZ
U5TiDUWDQM/5NxbzaH60b+NRX2iZHlqfeTfdO5Z6dzc0R1VpOK0kSc/RKafV9FWcEeW+Tve5Mt4Q
dicoOjjco+6s67kd62XYW1iMJxOYKNIj1Hvxkg6Rx58/HRiio2PHlAbI83CtGwTFgNxlz5DufYRn
lWl4w5TSgR6LBXJbfJN4Ea4C6cSyExCxVGFLWoNAgM8JS1gwnLRU9I+nXDZimH8XCRrTKGvwG5Oz
C4tO2bE9Pmvrb0u7B1h3OXPPaiiJXgasFiBT9mYdm1sL/PhZhx4l2a9eaShGB3PeNxDL4NPeoIW1
C824EPMNascwtIBgDi546sXV6vpBvMe7qb1Ox/HY5xV2PSJeJU7GsOJOGCkVGv0LziW6dcdi9GA4
TcxhFV98yaKwOWhGkYs1sz6MjFFMNAE5vGRLQE7Z8i+PhQR21UU/+wEDF4i+ssD4VU+8JlUPdcEu
yre4WZCPOW7IRzpfjlSNGMXjwE3iIe/ica27XAH1yefFLakIfRamUiicY+RbZ91Pf5WdE7k5pu0I
SUfo/IUrV5K0ka+TWbYYh1ug47x3jguIBL2zoLaoBwD9exzFYXw0BbXejkss9ia3ljVMZOps4Qko
u8Qhvad72BerHYcAla4YdL0wNzGohY8n272XPpwNkhBq3zomuObE8FOUzlQi+Szla+krFsE2/42n
z3CI+fhuLum/Qwal4pV5ysgWj8XF3iGb/4P046zZVattbU/BfQu9DKo7s7n7miIFMFyACCX0nIW1
Gg+pnWL0PbtDtJf46Y1m6+QBLQAsIEfGqFNYt0UhFlChfXza1lYNGnVfX4ADVSQoKPUzgg6wXi3S
BpD7s1N1DjbHuis2tNuoqql0PbcPOh8cH8QHhcwT0ekFXyCHHtk/D6xOrmtWbyzC6RVHkO3wIxsp
mpdk2pavzzt+a7InflJ36tjuk8oi3dN+aMWvLipOMzXHRQ8hIcRCwvtKw5P3471h5p3i71vChljV
wS5jWmvJeTXoDlLIG2KZsN0M4sQlW/XEPPopBRMmBb67lhUB1v60hMLVALR5oL+EiDz7DlshrO5c
CmCcdlE1dNa+JfAHvEsy1Rl+ErhkrQQfYIod+eBPmORpoL9VxXjz1y+C4SY3UJtjtfRV8Zk+ortm
Rx0sX/zcrdaJKYv/BqPzS5j6jZKSAFOMSbceonsJ6U5Qz+vnoTtiZZJmyDB2IdPdj0E9/PoXEu9J
Rpjs0CxF/20Q0Psxlz4n1M1apgpTl4x2P2c7tHfsw66POwRKfymmALV2uvqMlr44r0lDF527/OCD
37S7OMmi9vTUZ1cEK7nJghkU2uI11c6PVPZCyrUzAQ7dlYjhNy7oiPHgpVPNV/Sd7cVrfMdSztXp
2eCPBTOlqVzNYzn3R1zIrsRdpxzdHlxU5ySLhK4q2q5ipcm97hMVBOCKExaEqdLd4KXEN8v6hhDe
+uFqbac3jI1YBux9aRu2cfS8jv+9y+OU2eddpuH3+/zIfd2D1jJa8x4b+ni4XNZd8nKLPW1GDYoK
WS37Ynyoa43MB26oMMHYY0ClfMprIfKhrMqQcvXMRvlCiLMMYOvUUVz0HvlNuFNMThGpg9AvPCjz
k72lBA4V8/QwK3v44wLgiLtiqBviBizmCnioLZWE622LBHLa7Sxb2oEQynHpFiKfQ28K2EaQ54Yu
MjYeAUudKrzdl6Fd0iFl/WDv95X+VNAAgflHd3g8jmWIGaOugtY6E9+2h7ZXFO4TD9kt8oVbc/9s
Myr4r/Sq55K6AwgOXfG08O16ggoNRpJ4AEx1mq1ymQvsScJXJwl087WIoLp7crU8k9Yc7Fu513id
DwS57ZlBKSBIyPtGIJD5bpwppVkiOjEUG10WGruLtPtBYv2hcJeWt6lbDoj3EOXhprTyPdykQ135
JVfERBDDt8cJChjzP8iAgIkFztSnUuBH3fXkuHmINWjFcFr3X0krQhtzVMBdwGgwPK8AyPlHE3f2
wcaUDND6LTcNXYcAz4Il3ltfnNDD2sWpfyfgcsF312r15vsuxQUXN3cQC4huQo9bPluVFVdph4W9
ZgoymBQffqhaMyp86/DijW4srnEt/D9chzw+c4mupe9uNLA30S042t58MKhIuCCwgLfiquvacvGK
3YMhXk+5SQ2n6qb0MjBrXXyB8HEdv0w9a8b2f4OvD1xEa3Iv3X7eWSmIiZTgHjCjhA+NvqYDMTgY
+obRSLBjn67xGRxkc0Mg9FiUaHNtA2Z4tKUxQFBAo4WBseqF8ld06+/5/TTiQORztVmYmCbZ2M/B
n88RbPPt4ZWrGoTUQgdcADg0AcQGcmUHPHrdo651a9qyTAsq8eZY7gxGSkhWHkYUbI1hmJTZ7hJb
onHps64e9152FLTl/vHkIKkVibNSAjTcJUJRrqst1ElcAZMcF87c3akGQ1+fqj2F6hnbPDztWeMH
YwhqVpbGND8Gj+Xohqu4swPCcNdiGb45Smh4DX8TPZvhrpLDJHOfOJC0DacBGj1MaSZwSOB8HbJw
PMw7vHXvFDF5mSfEaHALd8M78VOyrDHCr/b64V1wlD+rqnCQT09zW6OAOt00MkRqMIm3q/4EAqxG
8tGlqNVFjcVqleH59aGO+u9+H90Tx+LH7mroKn7mGXBsOCvO4YzEY6YGx1hI2HSY0Ss7wDOF3G/m
yCoJi6NCnkjE3EnjKdkOTG7hPR8u7XyUnJ9DnJ+v20p0zQ8Z+9P9ceP6oLa0jCuSZj93QsVRT8IF
TAmYhLskbQRxYs4bqc+yDO27h/o1e3nXZCXDi0qPpTDWBypsOqNwhKOU72WvjolCk+ve8Fwk54/U
GIM15haRkqUkj+tRKwSES2sGi8Bmb4CiKhs9/gzpI//AoFC915J6SViuYcVk2Y3lQFYIAQljVdXv
SGSFoxER4JX7ZTk3PprEkyEz7GoMdl8gmi/nIz3Gfo1NmwelfqtI6u+qWeoFFJmoJziHCX3re6Ao
DaeEZetpoS1EFQRNnSFAg2sX0h49TdgHMawCqLuGpz2QN0WI6xlJTOLWKPO09co476BkqBBtsJbS
vyE5ugg/KaqY9L65WlRskcQdzKGDNyLWNBmmifiV2kG4OpSyYe+4NVFVzaCUS5Xk9UkFAW3vo+f2
ebe6HmpzSLtX3T6EZNLjJGl+TvKdzWp5GaXKFfinXFHqwwJJQkA/XmSTfs5CmVWab79UTYKBLkZ0
znSP931reu/THacGxO90U16JGtiePLmV9b8bwpezkVfKil/Ju53WTyRW0GppOzzY6AMa7QVCZzwt
6dAUXEasJrPcG0Wdet8HuPZoyWClRKAwEWlzkzdosCdF7KGm3eNJLwiPl271BcSylD+Q6SHtoAsc
9t4WkVZyD80H5m14pKA7xrblVIrA9DsBAGUY1XoxxfiJNz7O4wgYTbw3SM0Vbv8CaBuF8YIaKhOt
Kx9b7W8MMFH9cxeT+NuqEoBOXu/4qn8hcoSWfVdAiGjNxBN/qF5SyCME3UWViSvXUnQj//fVSL0B
XncPYKKDwc9y2ZTj0s3014E9EMlGaWTGZ+Jh+KRP/52lHLakX+XDUq3wn6JKeRjkdp9QMuHoK6I7
o0ERmBtjADUmTjiJSuVTabkO/r55msNQ7j2MehsqBERM6Fsmm5S+ePo2GeejpCHaBRG3GVR1vjpa
c/se7I6JLjZiQawP1E1VvR7wGu2PdEZ7DjQcDcJ0qz8Ra+xMjZWLgMp3PfjtdzUzoXlhuh6O4ty2
4V6meNOnGX7kDGUSrA2YXd3RAwiCggVyq2HEUcnarjMgIyVJb1r2O1LZtk0nQztaLJPc0B3KwVpc
PwPjzVW5wClaBX+vXrsGaWMgQNamaW0TFnTzruWmClbfOHEbHaj/3kOHjj6hC/xB6CzMPGrTDuRN
1/COXUurDzpDaBqzt7nT8ILpJeZb63gBkcFhCCjxBwQLTXIKfhpuda4wQpaykruYm1984TK7qe0r
h2984tB1whdAjdg+ln7IrwK31x1dSN4g/iJEBADdO3LCjKRHwMJ+rgOPf2kvLBf0g8cFbByCvs1Q
++kqs6ZpYHEuU7j1J7J+JGAcjzZF9ua6Vbjq+HQ6B7ZDPs3DkQpWtXkIAHR75NH2IQB4vwwo/Ra3
O/WBKGP6nmRtWeCfje5GH5xrnm3LnXDEkam170wyMXMDr3Qmc383X7OAg5Ij1hy8vbxrGSRdVgwj
b3kS4Zm8EvvzI28NGxm8GxDt99FTmWdD7mhBoKw1ztEqsajd4dbfAWAUz967aDjlYKLrhldlB8yF
9NSGzqE721HVgH2JCR4d9nruN6mKy4c4v/WbM3Yr2d2Bp6/6/6Z2khx2SHxzYt5ct6Aq8CBVc5c2
BpgErXkfKOs7M0l3ZrJWSjaTmToEbtPyEaq42bwoiNMWndPMIgt1F5aTMqN70Ap4HwdmDk+iMKYV
0cgXRXPkkiCQEkAkgmIJTjQDZMK/gS5Tkmvm7Tri+2CNhFnJUudZ3pgMHdY29BUj8Lvcbyk+yJtn
cZxrLuWSCDLejxsNjh/+Q2KgKH8U24VxWUyXF1TxKqBn21CsmAnJy2/Cs2LYyzLun+vnVBooqeql
1fmrlG6vXFM72ZVu6ZaXd82FNy8hHfpb+sCl8HeqI/imKRSAqk/KUFI8RAA6p4bur7AkUf1PI1A+
ZrJJ0wo7EovOFr+5DhdFZtRgnAnJgpVF01EebgbAeMDb1h6wTZcTWiaKii18RdMrn9BupU433VnI
Hatnc7zOPl/E0b8Z1CDZTf4IpxOv+lgAd4uvqhk8tvHreX+CyLOKV5BRQer1kQviXnxmF+MiYvNc
edOCC+FwHwTPyxKWyuTQga3W8mCvKR3JFYOuXfMaGN8MwJ3n6BsMT76dbH+h7ELZ26zDhdBmc+tg
OkHvwK+Sc1POksTbhp7vcMLsIs7IJd7fvpz8OaFo9Ehmrw/AVyUwhK0tqCX7JlASjh7EA+YAvpEL
JjfxWz4uy4PoEev0rP4keAMJ9ySlU+9vC98hF6MO81S60VSEbMAtioxs0IrDIrTGWgAoXAgH+4X4
SPkQwnbvAej7pO3HmHt0Idj1rTYYZkXwPod/l2bq5rJW+rrZbKIs+d0JxLBpbjzTtVav9fcXkbDv
LmCt7u+rP06nIkKv5vlzzmW1GMbP0YfbPQGVQQqfBY1a6M1UxUSLyzv2NxIRFxH3r7ukBG4VK7hw
jp/x4PkFSJ5wGm25Tm8cYpCnC9wUV4acWzvXnPGWTQXJF6OspdBDNkowANLdvdhjJv+YTLzRbM9t
uSeZTo6t/Edv/O2Kkyt7O9cXWPbm7mKmzr3H/DuYNMKT0qXH692PCrdJccj/5WUsyY/brOS+EQdL
pYQVJYGaFcHGDy4AuEJhjeHsFnoD0iOBZCvZUxZBJ+LwXYgzMTKGXUFBp67U0KqjKmnvO679EqHv
aAX/AswItVq03AtqAtutGw9HPUJx5We+jHhQwn0rh35dFgKNQaAXpbgFSg5xEQSyqD6dD2Q4kP8O
fTnR9mfQaQIZhzdT026yT6/e66UBPwfSoKRYbh/w3gLXImtC7sQG7TReP4D4oSLvN8OxzaJGlM0u
bmjMxq9/YdUL8lOM9E6KGGxh7LqBA+oaF6nimm8xNy8DbqP/OObeIzbEFb/3j2hZZA8A/2ylr4Ao
1ZrEnqdW+HsyEWbDoSNQocP7O5CxWxO1VM1lpoPsv0WulTj+Hxt9iJOXoPuTkBrNMAiI4WOZmO93
SH8qA2/FpwgycUzIk3QKvBIeWT2GIwyq9Es242NRwrq2QuhXYqkOiA6TqZzjulBBKgt4VLHEnC9q
K75+AZvjXa1XyoL3NH/RE4a+j3Pa8Ge+byIttlyIDoofbwLd95Dud2tfwpgPkDlfKfdVFBEEKVgA
DmakKJFWMPQLhPoS+fPCWpbsTxi8XmJJ/3+WrWwWEapR5iah+ech2CZfERf+xMMXad0NkyWsMBlH
7hendrLjVqj+VJXEVg5rTlEeo13NJ1IcZD302OYcy6PQNP/Ojkw9FGHHosiJhuTmDnMPNQkLtmSH
hZTHqcW4Z6ELe81c9c4kv6dcZ7+W9hawr7DARd/aqhXFhATHQRN+AShZwOls7nBm/pKB2WyQU89h
u9quNDw4wek5XzdHsLLXRsFp17WiXojQz7WfH/6BrSJypU5m6gdtDmz3DZN9zs62RoQ6uArcZt4E
K9cDBkz3dNMEvQIULv4ubf6VyytnwnAn50IsqS5W9wI28E7p49wP9cBJgJ1rgFdxMTfYiXV0185T
qy2XmlOdA6USfD7dNiv835dbSDKtWLuoZUO9aF0sCbAvZ+9AarEYlcIaMO/NVk8sc2uosr+fPFd7
VFk/P7mCDZ/u0l7QBHV/HogSPxrKZVbtVnA4ABy8dm5QxLuFGIjfM7MYxIctqVoL9ZXc1+Mk40JJ
gbOam2o+4M1pKa4yqhySxsjPcZSibJRfBw9y7+rGVSOy57ElDrRwuL8BKOmZjrLlPMZ7VIlFLRtH
70LyP85MXEw4kmpkGZ2vUUGVJeK+IAmyICcRqDUVu/SKkLrH4ET7xzjME3+nyetoLWXmh3uJP2ex
Sv7NO9Mmd3pv8BqqiJeo6+YBWWdnpw3q8z2DB4TQoNuamjdx6PqWeDA1OKEWFN1FCO2B4ufQi7Nb
3uVcI/oC0pbN7PTtFgzu4DLxnTyrMxJrkx+dAELfyKZPOM5IglQIbHbNNVeHtWbRkGxCthQpEVQ5
Y5Qjg2eCuvW6dfeB5xSGJo+5lfPryxOw55A0AsXFoGDQON1mPiZ4NM4sZQZD8ZC51BD/a14RSxBI
t2ahG73u46UMnGNT79YRBM392aGO5ez/Grj3ynqCmSIcqXRLVmd9+bX6laT5/+otnZ6NIhdHScef
/7dkwCRx0jXMkHY5vYhYkKKmvUmYpd8OSMWh2XUn4m53GUU1B8U4qY2nJ0+fUcQ1FtBxTfPgqF4k
7ocESKaOMYLMcB61s9VhWz6i0Lt0EjTDtSOZfsLydK8BbOhRJft8Ntd2xFRXcOJbSnQOoWeDzrpV
Mw+T/6AnA4RYo7uoJn33ILlcHeX2Lo1wLNg5hJ/M1VFwkgFfmjBJ5ZlzZreMVbNkEtaR4ynteuG4
cGZXMZeQTVCYVUdkEJfANV08fcMdx+8uRbsQGpNYj7p+9/B9UePm0zn4+xuDKonU/IXzyQXmp1QZ
TcPjSWoN+XPFwvRLNKRVKNW96Je+drIEoEDl2gJ7nGB9c/KnWqQc003nPIscbUXEw/W3r5s6QPHC
KMSsHYJb+HqlcAzwYPXzYoCJKSGxc9hPO0MyGYT2ksyWW0Clw4Qgjwa/TIGA8WNOkIzk4vRRs4dQ
umlJ9TgfUNrA8ycJDHJUCw/ti//s9/lv9YxKRPSjs5NRA64HdWCvHpVvpuhDU3FqtXpcOiNMP/Ds
o6Q08CXF8yYyGEim037q0SFWTPJfCPB2YOWKdaD6HW0aoMvK/eVLCBETInHXTo2eDf0sRxmvJ7ms
SOhnBeSJ15C8ERkSTfqhVfGLgeHGrou/5TW8rQlzx+710JD7iXpBIbZAV8vRTv+tLKbd559XwLSO
5vQNLdPa4Caxh4ADOPE2uDnED1kXFF+7nkorEta2jgdEHYBJA5B41LN+2DqL2EenQK55am5qQL2y
9wBbZsAAj0X8vnnqz5+mpnbyL+8jACpXSbPm/UAbipcJ1cg9tBOLsilxpVcpXKv0eEIbR21DdSRV
aXm0s6yHFFLPSJZcQ0evizGQAKL86rvnmdNbkw1zBzCQZyNdWAEQgAnZvXVHlghv3eBgahptsmkp
KYXVQUL+Wql5T43ZtRZQAvDzl5p4k8Lwk/dm9HdCmh2Jp5YR7NgZkUm5tvQpITNoqiVm4S0jJ3b9
hoN2RKL1d4/dgjJ/7KczYZyKjSkPd0//b4HNEk6wcvFG5nWsBMw6LLJfWPlcoSoBec+MYQl/6rgg
Bmznxx11DxtMcfMepVJxOY+MIvHpYAAuiFfv4OjK/arV4dDGdElgUKsseIS4FCv11xqtSVI9TXGy
dxupyC6/8DVUJK4KperJtrVrS8OXyewR7cMwncx0ucFtcG2LDrg0LdrcFTpFrwdpNgEV43f/BuVm
X7fcLjiNp9RTD0nN93ZiUmLGmSnVKOnWrbTUc4cgbCi50ZQGAlWZcW/UGleV0iPcJsOwglz7BtZI
F6jgDI9wF9nVz35SptBTw+vQLpZA/Z2KMybkahe+sw+kpsEvWznyd/+7wa7hhy6j849OPHUwD++y
I8BcWgTlEYfLM/kBCymGytFLai7XkT0G5ucwMLrvz5ANmqS35C7TV/TGBbLm6LdCRTq+lIU/7/ff
Qt67nYyURc4TIkacsT0/24bMu9SRs1qmAtxBDf2OC3dGZbUfObHCce+o8aYq7sBMeZP9GDOLRJo1
gCBaYWvWlbGNQ6mQcDcsl4asXNW+eURXx5C+b0BBRRZH6rlC7hsEdmkr7lYxFz9Iqr15szMJV9JM
X/eL0dGwk3okxrKsU5kYawnnmd1jQBnHjBUQJIdAztICE1Svl1GXvqMTmCtcezVizXqY2rrzZKvS
Ev9ME9fWBi8FKo5thQm+BT1qpFKF7uGLoeZ4YaT+RAjSsmfZB5K2pj8vaSR3iG4jk6xpOckMHjjT
wB2E/dbATsUUjnt3UxAUvPoKZdJKJ3A3DT+BtaczQ4ngLPvz4/x6wkbW07iORasJ/J0vZz/nKDAC
3yde0akiDGnCbwX4ANfQP9yz5ou8zz2oNj2DkKMgOohyjk8S5LRIb5xgZMCloJ2MGyP4a7pe5UnQ
NcTFO40bFD8Ew1G5iU931JPJz9yKUWxVOswTqx7r/R4DpUg/DaA6qDyeSLKaY2SCGCsDfd3pBTNU
ZtvS1eZR82uHNYUwcWAtlej1FDJQQ/O5/p6BNVV2F8lizAl9ZsQjy4rnFezSRaI77/lBtIdQhT/T
iL1nj1a/hXTgBfcgSsno6h/7e++mzDvvocrF2pkAXcFIBQha11edjM1PF9E2s+Au1NWX5/H97bLW
Hc6b3QgFJLTUJEm4f1aNWLllagklDb5fV5yLO1YjXrfG45srxdpTtYS/KCbgkBXSTHpxbYlDlkB5
QqjIn8Zad77M7lAJZPvQYk4TCaF08AXVc6hQz00DFOc7qx6AwSmJfw1rs5eh4Uvy0nQgTxDn/qK6
HVKf8WfZjDNtGfLUqkQTpPJHknpy0mfvnMBD2NiQcbavaS33fmQjN/6puB0G/JdkldNodZS1SKq7
fIOj/LiWP8O3KUUQqZv47dQtCmBLNLC/bZGhTUmKGfmObvtdgKmHrpbjm2vmuBdqfJUS2W9RZZu9
mftwdv7+0nboONMQXGI6e2rkYGpVQi4d1Yd72WiWQ3SJOtczXKICiVFkj3iuHnsMp6+zNicnFi4V
phM3mD2SaSNzDBQJo5G0lGczQuuePq87yRLdA4qMivrURUudPDLcqeV2O728jG7ZUcepBTgEnvQC
wU0vQM3zrWnfKGae9Zf+V0n84FTlcMZ7qWTFT+3cwLbS734si796QxgpC3TeYKKukirC+MilQ23l
/AUd9sscJeoei+817V9w47zQ4G+VDFoTOA4ARt14NS0k2TqjsuKKWpi0YbBhCkOxaxFPLKiolpJe
QO2KbNg3QODZDpwRNN0BO25xGF6J2VXXH+RaKKfb6jDztzd7up9gIxY2d7UmcOlewLfjuyKPGElg
eFlD94mGz7mBlYUbVYieQ6zkuqqmXVQge7nvIJJ2mXkq85ZSMeYZtokg5gXyg+TJzdQyBv/9arfb
6mlcS+njermy4hnyUdmqhF5dYXnPZdDw4Ooqe3FuT8R2jChb/q3xz19HinE35cFSCrqR+x4Hyw3P
lXs6H3RSXxbKQiCmMvnpk+GxiJkbUveY00fEcLorQHTWC4cUh3I44U0zxonrRGBMMnYlg/NCm57x
NKJZcX+qiPbKah2oxrpUrj0CvEBDwZwcFVkF1FjmjnJBTWuFjNn/dm7p1biUQ8IViTfVHd4Mz8XQ
MHL6mkWcHVsihQL5jVau53CBu3BifXykp7fvb4Nd6HAIKMPurjUqGlf9+Fi5H+ZNDUOfo2eB/BA/
65meV19IFPmndCCp60iCpx2FHedU7eUGQ9uUP3ZogzIiNeHlSpbG8FQrhraGr8DwdIfq463uyUp4
9l+9CEKmPaQS3VDddMUsG+g/TMgkxywMHrZGwfYP+5g7l+FOLyNyjQ9usLTx4jZ8PVslgKbwsJ2X
Fb8CGVd1v8jiUW3c2bZPjwrbpi8RxDt/ySES+DlR7OFQQmjL2XgC4fIeUD0XhVroMVtYEWKH24DE
0H+ugfrIqiW2tBItYq4epTRYGB7ELZCo6BFhHLRtzsemktUUe8JmInszjWDZyOrrmY/8zSDVSyPN
YgHeyBXdXPq0D2JUQlBMGGDvofIN8wC9uOJ6l3yOopEM6dT8G4G1n0Y+0GYxSoGJ/Bk5Ykzg++wH
dAiWX21WKnQCZW0/3h4ghBg4UaGMHp4vTx8Ira+lv94cuWmuNuWPPmhC+jM7zqmxYmwdbovSYN+H
DnOEZp9wdzVgt2f74Egt4Hw63XBAw6MQEaO8RvLp/UovKNK16SL+FuLs9ftteApuCfE52Hwk0ZHa
6stg3uG8oMesa7/nFxEcQ93u3+Q1pt7fvAzOe7gvLX8dmgrYxg3HD3/BQ+pjyqmbw4TZtvVQiKQi
1xJKTWFnx/PITQO7je1xzxCTKRZn5kJHzoMtsIKFigt2phJo6OVoO4XCha1y4gJ6WdGnzlsrZBMS
geRcYzp7ixW8BsEmcP0eo5+oXC7dIJO160c3Mh4ZXqwiwRit8TkCBx/dz77CEQKq324dF9h+wjc9
qPdJuQU95io56/bAvDodWdbNQgR4cm+7huTywUjGpc5IEGA5v2zEcuH0+nuno54rHB43kqvf94Ed
KDl/vOlHCPC3miAJJXN+jxXNhZwXLoAwAHDaplVIwDRAQFoccHnSg6SP8Fy8ZN0o508wVOiJD9aY
M5I9Oz7o4TtV62rCEfEl8UhqeYzGh4YOoOIiYz89LEqNXc+bPmeW2D7LmWxG3+Z12zYPj11E8gYW
Pkr/mdDj8b/UvGWshbb4B8yNLHBaPoaquBrLkxdwHObLflmdf4bsTPiqlDfbrnsTPD2SSV7L7O8e
nE3y8oS57/IpKGZgvWbyz73J9S0PUr62YOCSylgGFn44X532H/lb0g/TmF1+v7TADoeoZtgbU9D5
WxrI4cUMV6X6WiCVV9p9CVMkOLww5+tT+hyQSEo0h4T+nZDYp1DUV+dpmWib33oyYg89Sil8D4Sd
JR72UI6ETPHI/rxltjfxbqjn5jCy6SASBV42OpBWWWqprozl+A/+CKj6CwvHMAcF9te0cRjumC/e
8KXlLWghH3uApMv7XLq87xHXOhhKh1KTAu8Ng+F+/1h7Y/xIgzDnxM7WtGeSWsAT+aO5tJ6MLr4a
MqlJGq7KOPSzqy+L1xGimQImNH5YDh6IYe1bzNYmevnhE9kR7NjpEkvW32JgQSQTW44hgYThcB3h
wizhDUb2uVFPfsMXyVRCCF52dX0JOSFFNYP5r/B35cr1JlG8Zx0sc4bq4nc1ZyEuXHDow5PcK3sb
xd10M/RB53IQcChMwlXos1FEgAy7mySAYJpjrDOmT6cPVrOMLMcAdEUbE9gvI52KxoXC9bNyQ+4m
f8p1NCxYS9EXgAJYcBJ0O8d51q0LMGm4N0a7PA7XN1BSWm1s3i+UZqORnt2OyIlBEFEPIaXDhOB9
Pyv0iDlceDoXjPOqLTKf8vgLwVv4LEGSR2VuV2EXTD9d0rZdQfr5Y7j5aSJdmVd5a5O0uUXrRoz4
4fox4fu6U79ciQ2nZzbWiW2T7OAzR6M0luDjEsFSp7RDpvcki5DOay6Pd/OmeK/OxqXVqrnF/idF
Qe0B9dZYv3GMcC+fLQrHIh9DOxryZVtAjuIQ/9dUiUhdFUHuL0Dlu5M7lAq9IBKRMndpm/BQws/5
0kvdpI15pyhISZ33Co6f+OMuv8u5V5K61sHx8qky9LXSp0vdg65jyvyGr9DZEZwve0kZeeWNBhuR
V6lmBCBu+DPnYb3503lAwG9OZpSewv7sEpI9UYKki3/MFpvWyHvCzXgUNZ8zOTHg5ee0Y8EPERY1
Vi/5nkManCplBPEpg+Y71xtG/XG1GhLp8q3eHxeWB7nbvDRluuq7UTJEnfxmCTH+Rnwmt0Q/X6xN
iMe2xkHwdGVN/ep3U9GeRW/jf+6ER7iTj7yclex6qiN79lrBdl6bJcuo1foXdxZts1I1a/C3rq+c
sRR0EWnHzRklyIcu7KMZqaAZ7Jj4i7rBfXsPqo1SqOHXx40mExPtWAVFu6zqNlr03Ro7fuLieg+L
QVE/9s80/LhEe97688R70h/CXnWiQEtuMSFmY5P1oQevOKDYXletMmkXyKYerSkAKaIBlY7MUMuz
D8YH15yDvhq4I5MUD667j+T5n9U91HSv8vp8SMqSR8pp+yQlCu6jT5ExfqjzSfdGCvNayJ1+jDOF
uX1VZCCXyu7r5uQtI0o1XwXUjRnJKQjRTiQMxSCXSS6D5rCliyvDy/b/mNlbpwvG8SGlhLwVmcIY
0n330YYt28NCQWzMn7xvh4P5HKW21Mr3irSjeZNyaLlEb1RLn/xJxDiV5oaKhNiy1g4KUrhkarKY
wop0CtkIzoDcT2lWyVirHkcdDwxaavxFSZ4+G4RvefptGB3ULenKore2QXm25XXf6yxqW+oDmTr6
7Ekx2u9MAWMW8BS10xhh84Fkmo/T7XbvOKkXCs+myeT4TgJWUc+HlKOvzIP4JYGjFLmpbmcj8Idm
3s0zgyrg9cVoSh2hvnLasbtv45PcYs9pCe2xbGJ/u0lpKbjbGibHANhzFvqDt+RkX2yDVNJvhtsx
9GTtXhpCKtxo+T+T2Jgu2xyVe8A64gjpukEtBHkaroRsI+iczljBjrERZ1c3JOocS8iv434fdW00
LBXzr/VQvel4eyr6KhjQOu1yiFOAAxobQChHBIsehWgl1VUlhUabbbmwVRLZezLFxWa/DI7m6ljJ
mKomBlPpBb7hxS7CJtMe0sMJACM/SRg5NOTmPPVg5SxAvk++Dqf9nFws/F7WXbFn4zJJwCkRhcs8
v5qyyALyYpXcmrKh+TklRc/rfT771SX70ygZbC96G6cN5ySvPX8oje0xZBWqQojhyXgw5ECpo50b
uAhEWTCawN5F7eCkKpunHEewjZ8NH6zYrRpKnW2AVKwEagJENVN4A4+Zt7Y6oVhJxnFGDx12oGFu
S7ThHhp2mdgK0tQAN2Mqha+XPSLxoHhlQReTEMSCWFf2PE711dLT9/KjnskAkcEd+wpaxULbveqB
LcsN+bFDYLSN6MptVNLAc8t6klRQyazeLiNGCPLji0LjnlELL6tdCAIPoLGKo0q5Cik/eKs+G2RW
d9mwBAv18TEKFtPPW6wYy7oQM2ymUgE5v+ranKbL9mCErlt22YRjXjg3stoF3ZjtwUjR6wgGr3IZ
7Y7dU4H1J5gMK1znWlrjoFHmyTDI1B03if9tEALUWoOHstbng9lURvL30w021C4bi88KxYMDlz+p
O97d6iifV26XUX/bYEnjoMOtgdcHQUXDIXCusju0X8O3mYRUhjPL6xWLRtT2my/75uNPGKvdXILg
2xT2izdV/KY4U7hgdVNS/UOSiB6euhgnmBGLASb2LU5ioIbilTRBw/V7YymkdkG+j6JLDLXlq7Da
Dk1S3kWfrnOwiLSe1v8AX9ReShWWmwMB2ViJMaQpsOsnfjHuVgbF0e6LIhXcvRp2W2HX6pC0cQCI
HeqJqBIog1ztZ3m/uu1dX1LhDiFsP2e3NKKaBY14pHxHtclIDef4Wduc7jE67ShibaquO9BZAXMm
KDTaRBpVujODxOfbL1LpHKq1s+FuadqPlUK0p1S8odGpU/zMpYOsmTfUByODBIxBJKTDsI6tp54z
/QkOwWH9IQp0WH+masLT1N9011VHcw3PzGZwVDPeuhot0777K2jlPlQjyI8lEXAwGEWbwHD4ASx1
KCCG7cZ0Ley+kCMVYkKq/5DVGgpjmJDdi5UK+A9DSpmiCsTQxVH3Rh7JraH+ojVqUPk23ILbrhuP
6ZSD1lS8Ce2qLFg4c3sle7trNMprvFMLU7NINyvzyVes/+kQJWz6aXZXfykxke0dIoRHkU1Rmy8j
us1dHrE0ARtGSuRhItBNCr+v7/MuRfWDWYsAE3yyhW1SzNGoTEhHwv/NaDVtg6rwrhSC3ZYRPXGE
ZHUeISrBZ4tM1UfT+Rwlus1VhS5YjDKtu7ZCws9BfH+vIzyyjFU+EjEJDZOhlyr83LfPPqHYPUoE
mCI6v8KSbHtRnTIZ/ZVQ+FrLnIMVamlDxaBNFrDSoNKhSxwQTT5BIJiZNKhmN8VQueI+ucPCCqg6
H9bTa1jx+segYtx1oKOVMpSS3NQZMlh2nRoAA8P07oW9w/cktQhzMxTOfk0Mmoe1YhG6RD0vOnJr
eruMptg6Gm2e9A/8a4Q249Udu6WVumMhkpPjJIIU3t3Bi+L7XmQMFXRbxPTuwgHniSwhKCLyOUZX
VBNQK21yA+r+8pNH9ZjSPvhzYilVZVMszqQa6E4mje9HhIYk0bx+jHYHDqXbXrY5m3pGfIWWY73F
IqtxhRbP63ZXDNXzdH7Ad1G10gIgbjvA4hxCyyvVvZESyxZkDUyG2ssokTK09Du3l2OeAGdf5DPx
+PlazdoFDzdi91IOHuUzVnLGylp/lp5MRgP6PZjme7OAQkUbTBWEQFoDCMfoawq2NFQttGd/nzjm
XW5+EROYtXS9VrfRvhxCp4My/3mZY30FcMkMEmGQa0e7pMOI5AdQ9BtUBpmwbBzrPXPACGSQH2QK
ymY73TXntmoI4+jpwlRwhrPn5+/Sf8XRBD2xY/jQm6ub2lEBI6K2WAxvnPIh4FPDC/SjA2C3moTQ
zdB9XHLZYHFiRcIMoo7rcEcIIwTdNR8jGzb/4dpaJFXPIzAOH1Q8+TXyVQ1JJjjwuvCkswMuAGvO
IchAMAy/qtgEZrK8s4E6eUdKlSeh248OiQ5u19qNfjyZ0fImyQJ4GIS6WRrn4gDFk53QU4EZd5h7
syrrmTLMD/0meTZsz2FB/qysRhEocNOjuKjNH+9MrtwzOq9s0d8FBS3mQ1VEZSQ8Y9q50aAo5bV0
cx6sycrRiccH+h0nOfXhFWlpodsadGI1UCfJUbxPkhbW3AoBrK3zDmBIA5UX4IRBCqhyny3uDYFY
krXboro19e7JjnitsNdbyK7hbCYvRnSjjUk4gO/T6CeN1T5tAKS3NIh4fzlpXJV1VB8Sq5m+2gk5
VtNY2af5pRgitYg3AFqTVgJNqu/R2VQthQ7g6qOwID01ZLJaFw917vzuG7kCm+m2kz39XJu0QsxW
7bCg6rL7GG9dCoiQ5T9HIsi4C2WHbHCTa8kyJI52Q/qKAFl9ASZh0GBnnunlOOLBaTeZI1vuGdmH
F61nEPJw+1k5gy8lU7pZlQMa8aVplcqdYKp2fUr0j+n18FszuuVjCUzZc6T2MHZgO2KHNxrvlA/x
K1b7TmTgyHmra4k+8jVZwaflGv6tJf6hWO7u+DYJ/sWK8K9j3EsOLYZpGKGJkrR0pKpm8zXdkgBz
o38zkSXxhBbnX7ZWxH1Vk+oNFE1WUFt8uEGKOLHNciTlFgB27OO69wHBPVQJm/IvDz4qhgnJjdFk
YdF2VPbOYr07wo4gWQ94G04Rgaaf2XqxpweY1kX8zz+1ca/aP/bgBiOIWvppnD8LoHP98AOyzL6e
++FY4LYOOcm8KAJok4BUV0PEEYE8bXXAudHuEAMzSaTMNA3yAbNxAP4dFiQSorXfwIq/zTeUbxIA
QYwxGd3qk4PHCzbYlUQeDECdAYLGBSoWj8N6zIinITbDsNZKA7/enrWl4Mtn4cFHo47qbi1JVnpe
WAAWoUYnz5sYF04tbWyMTohChLGqpMBtbTyijSLitpYUGCijJcHO4sMKvYPP0D2+kj51fXUavOa9
MSbK5MxG0hmeNjtCXtwuTAI2m+9TZMdfh+wB3YlulOMG6E9Ijvu/YlT/F9rlQRMVuzPeQ9YcgiOI
fbiDb+lHg7M+db9TwAzOdrAh/tUSVQmX6jlQB20EZ0JHLI/hth6nPbKboWqgeU3ENbPWvmpecW/R
TJ3iOk6KWIYR0itNFIt4aQD2o+dulcuz6I1BMjiAA4Dg76qzQQ6i7TOKQoWchox6JwCCNQxJT1wk
e5AuwgkbjkSpvYv+K5CS+94RRpxvfxRmowPEGK2ADztUuoI4fl0ucXPOGXcK7txDESZIw+i6zeSk
Eznf9jZwOvrALPioHIWpxIbbouX+n9NHJKReiRD9RE2ar6vzVv2y8o0LIfOURmiOSiVYSzOWJ9QR
PHa96MqglrmW/SxIa9iDxZe5XXcFiyPxwQJa69uQJZ0USTeheWDEpIsuRewqIDWnfM24d0w1MXcB
YlMsEhSnlPj5OINqtcIj9TB7uxJuSALMHP8RFvcrWVVQqHHkApc7uD6byz5V7mVpYVwF6kzmPFHJ
u5bYBsAdf5SineHOpvHOoSoRfoc6S9dBdGF8YZrpqTHtdmtJzQyeVaDhY+AzhajxVNel87e06w8a
+LHPPFrARLswwsUFI9YsweRPF2QON7XaEJ6EQCF6gw3K2pUvIQquVq0lx0hjP36PthfKzdz5g4vg
XaBUvv9pEQyLQF+FuzFQ1wEH6Ukwh6YYo64yea2+1RI+49WK0HTV6/NEYi7+yV4R3Myyt3wvANwR
g3DPEt0ZRSBEy/80J4f3ZuVnbK7GGUcpHY+yXjCieT9yWZkRt0LedL0DgIeZis2a+20WV9pKtXK0
FEV3Ieinepfo07Bj8v1LQkYn1HgrzlQzNBVSMeg9PtEh6VqahVtkhJIk7BbBez5MnsD7ZpML3lZm
pHbitmXqvticEvxew5tjRBBDCmVycxjnM1kc/SZSy8w4+VLl1RSH/2o+5hrEkiYhLwp/rxl5x4/a
ACjPrcsRu8URZTcmB53YBMlhxy6RCgI6PVBtFuKAXuZ6mNIToUpIDwfvrS+QciFXcAL/It6i8sTf
nA62d0i3Ti6twvtjULk2qQi6O9ft5fxvA3xoZyb9L9oNHIXrKeOw8s7ORgLQrCXDCdXGdKkQjN+S
WJLqd3K8pwFnQaSUYE8puFHv1RCHhryJKCRvBYAUOTSO02bZ0sFvgAqkimXObyIbf00pmM2JtWAg
cwPtnmxTBR7GyL+HSav5PFLCV5vlljDbhAN1mpAXLYE9qjbAc5+VManXNtYwLj59iz36YxwlMqj8
2qeKtw1vUbz3Dxh9nrrEtPmGGAG6RP6gDScRVFnYQKKBlXjfh32zo06w/hN7Sa8XBfNJChEDV5Xm
v6IE0kdPRC1v56mh0nhQldkNTHwkujb3Nw8HOeOzKJnGN74Yu9ufPGbOnKV7csVZyXq7xL8HFUYp
tdmnO4w0rRKXvXgvlKbLmlpPvlPYk6i0wBaw5ERSBh3qq4muO2VHOMDHerjzioPDvAi12PP9pAV5
Hydu+ztwZToaky1lofgQIDfLg9dYvi5DQo5Ayi7zvDq0fPX//unsquWnvbcyWkqcrgTzmsR/5cgz
EwqiFVoBw1XHWJehOUFLa5uuMKCcYhVmJBEq6curZw79Dq58piJEnnWr+mKXJwJRc3WsDSBhDBxa
gvyhQQg+QQcfnxRWZKLBqASlYnSgNVRraQEzOM74wkvUQ+sQpd4tQzO5DFVpC5dG9YD+iY/IOxXX
MHZ+clHChI04cE4Pzdp3kn0qaCcdjt0jHl7WolbPBVVU1MQV+J8oBckc3sKB/L7TuvPiBoKfJ87n
+I8JnhZtSzPU87Za9WLGpwXi3+ypXk2ekAeSuTBSja90mZeiyffFAvIZiQvoXI5HE19d1jmg0Jln
Ar+z+K0mw/x2pOvSS6JalYwj60mv7NpdfSnAg0Z7B2plhZzlOBYEENmfIQpbt1r43CHphX8NXTOQ
/+zxqm3MKXZYyzSvAPsm88oa1mPSV5f2Us7bWY8Uq214A2h0phDi3lb4JM4/lao8hSbQ9v7HlvT/
5JcRMAefIS0rGXrw0VAR0bqayPHChh5fq0qNoh6pqIHLWFSjuaP/J6YQM4aoL/+JUWd9zGIrZxuw
aRY1DOeSUbHr64sm3iYKx9F2Ayc0UPjI9EuFRGkFsNrtXHPo4rIherr7CxVakW+9LCHSxuf0OLhG
upwpN1F6WQcjApwLPPFQkcQbc6tNeBQ1xPXnfzQnoF0ONc90RSWRi8DAex/YaM2f1fP15beG+5lb
RNiUyi6kETQ09BINa433usymTK/Gw/mNeD78pKLvIHQiyKXHxy7zxLFHpm7k7FWCK0nxwG6YRHii
LZ3XIr4QFZT8MKUsfVFS+k8/9VHyl7OsxreHmd7NUyXNHkLl9GGhUCSURYt43mpxKPG6Ohmb3TGt
FgpbRpxyx/tkpH+murSGzy5mw8zKoznoA3AsMnFBaxhH+VElgRRgjYCLTm3r+FsvNuKFguo3IzC+
cqEWoBIOqV0GxI5yn5a+DOqIlH5dnJJiszyQRrrrSa7IPl/Xbbg+hw12oRDq/GkbluKByXqn9qsp
Q24xV2339l6co0bNrLQIs/v/fXBY6QeGO9CtrX9s7Sj9u+Lasdkm0NL+3dWAOOscqaclyldhYyHr
bNPjB1OL6yJTzIGHVv6pFgmxDgm3poe3kQdz7nOMgfrqO93ldv8UsonLQrFS+B5WN7zLYbxTnuRB
lAtmJO7NpZgYDXH7XeOHgWOsxw6LE7EmJhB8vukmv4nyNG2ZbSxTS49b+UPmCWfx7S6MCWPFeRee
hWhQonX3Y1AEgoS7yx30Kxw70E0bJ0ahAwkcyivxvDPMZvKpvdRO8pcMmoUOpFBOilA/Iw8F6YZa
n1pQwWg3qElb0PM26lWtLONVBXTckwqY/TjPbo6/6Ut7gIuUUk9w+51Fkdy1Q6J038VagvenVOKD
SACrX5Cmmfqu0Y6iHySKa9+99zW9jbL+bnT2N8NTMcQsEqm32Cnk8jVAgdtm2dxWT9iK2HxuBDIo
uMckY4L3uYPlD82ggk3pUg4TR0JMH+qhpkCH6alaLbvFEwQMZbbK1OOf6fmv4xlU5pgvw0RClLV/
AUbet2PxMEM/5rdoUVunGHGIW4ie0Oct3apNW5U0FEvsG0eQnR87vuNi/m/IkitBU8Yt//iXI5Vt
efPoO3nnRQSZ3i/QiNNg08LvchSb6SkFbVAdVaTKw89auHz/niuDCTUIUSGc/AmsCQq5QWrW48RY
MbCTwAL9j7yb/UdgE5Xxl6Y3FmKcezwEnau0MBnfkfmXdL5ubX7WEDV42kB1rSwhWzNEj5usspuH
IxoopotD/3xRa+bN0NJDQzmAicJTUX6O3rI36tFal6o8UQ95YUWoSKpY4AxGYCSEH/fG26oFeJd0
R0j+DlF/mbxK4lZdWtoFNk3Sh9dN1IuC7Z9cq19yqyCchDk99WmI1eBlZ4KlUfNrbSQ30aDMvtAL
PhmOS85jmE2z0tCaT7wOL19NLSs4VjVied0doAvVMFuxDh3qFm5/Q1dH8n7jgYrL1QVFCoXHWCgD
1GA83udC7oR4C6vlIfFw15Do/X/+0aEFP+8En3ky8RySP2QYXFO6GSfy22cDrd2ThrzbS9NN7fa0
0+00zSkcU4KpXCqE7GSr1wsYLC69w+0YlZCnksvzy70PxhK7EoRvg+NBM/lR7YDCO89s1E+yAd0F
B07z4Q3GHsdx1eQxLnAOi7H6GbQlxsKB0Xu5zEbdAgf+fSRkiltQPg5/av+YS63/MGhQOhumYzmy
zpZTJf1njJD+mTfn9uDnDQPH2svzVS0jt/2m+dY2VhF6TSs5ne9wlNmWZD6h+ahukq8ZAQA79QMR
IozNg1SPQeSqGyNtOEmesiePFdiCAMf4aoyGQNRziuRAxqljQ4bGZKjgQ+657IcGyksQoP193QzO
sw8aUxrxs/Sy+SMs2of2s4hCv+Gs+2UeNtzz6jaJ35YZt1Vng2meH6FQVTWwBCwdFojN0pYzgNSe
oJH2xnNQ2Y+9+BPNYzGCRRCimtMgqlUP/Qo/MaqZQMyc1V+pzLPDE2TdOe1KdbHobLrpS96XjQBa
eJCa9+PA7PS/0W+xhcXZKZUVKTyK005LsMbEpxTPnSgDkiz85rbhLeKZVhyqCfFsHZjUMwsVI+Pd
LhDS0sY5VbhUvFV7KFyxJeo9M9r0c0kXf4hRh3skvz0VWtqOxbZBongZeGSm4fFuR9v/ymTL/hJH
IzkAQpKjVUYJ0UZQYoIB1kVkIK2epf3Sn4ZjYSmuADFR3R/VSNE2RZZL3auMuCHoG24VeEQ2vVCo
/TPCzyEApsownXw+ZD8NhR3Exa53BMNQVnB1y7Utn9FOG73HrSUVIDEZpE+U9M6Yd6ZzVDcCYluV
hAn8jrIkua7cGQGYw80cYO63IlPTXGdPm/qR8BdI1C3VqsH5Q4EBseWjQqzg/+LR36l75G23h1IX
X2gbk7Zv4+yCdgdcIPRqfGK5jeUTN17eEUmHsR0ye7zsIjiAhLabou8jFkw17H9TTFVrSvph6ss5
vpEvajX8DWzcXdRn2NIU/ldFrVNil06mafrpWKUbkDk3V864rTV8vnyiGOkrfJIN9UthwYPwsfVP
vUDN6abiUsgL74+6//k1mpL+ZwYE0CHcg/pKgAcf5WU5uR5aMSAi/vAvpXQoeUGwuQCGzJRK8Uay
4F5lQMi5j0vhJS9D0VjDTznK1XzSsgg5GHWAA3bUnS+4Lyqtrufvi6jL/x1Sub3aBhcarzUWORLf
RV8yQQBAvG4Wwx3QOhlj3oyigpQM6h1vNE7EajWI1D1t2GmXFEZAl0B5wkUvxboMp2iUB3sxJErX
4OLCndpWnvuBRBiiEIKgfPETqVM2jo6yWL15Iv40xSO5harxm7l4MwPr0jMPBohb6u/47+gsVuH5
pdR3aQHzXPR0T511MXQehlEu1DCZD4wFYvVrAqeqrTcxY9sK80sCwvWaHxjdqxZmGSziNfDMj3VO
ChElr3hWHEhgqs5MilsET2KuIT97kne5r6ND+i+ly1X8pTByqa78GAgjFdaJWhIwv4kCF/a9hDwb
GrrywbXxXgem1KPNV9wp+134ISztmeT2vFVfoi7wtRY0283THnLuQr5/WpF6dVKjfwSbQudAwZ/U
E1wbiEovHOcAmNdZ3kCKI2ElHt+VKpYHAElExl6xUidAcjhtwubq2hE7w/dNd38DZbTG3VSzjAxT
yKKLtnjZgeg4Iz2v9dvcRxxB4giqhpftDGDKzc5vmzKuKBvkZPCUWxSAnjfpVm1kG9l3U5ckOgKo
VEkoLOYwqJEwehEi7Iexdt90iAb6JzpR4xN0T/teDe1C8luaueqYHW7wsvUMr51QdAQFtVx59wnc
kX7yQOmf7Q7aZWnPJeig8GtIdZCfB+pYRM7oPBwT4cmmuTlliD6HYfwZrOWJAo6UCl5RDUrJb311
7k5XV70U+CHa0ugrx2lBJnT6HHTNxgBsRDxcLSvvhVEjFudtF+/FwS1uDBwFKux+rv+1lx2yUdJr
MlrCRoictvtoAXILokCF/bFkzsGFpzCg+23bx35xayffUaYTPXXwCyZ93jO7CwUrSLuV719Zq3hS
59eJaI5LJfM86bsE6rZWByUTtkCd2yn54nJw/sFgqKhRX5ALWR8RUPiAO8I+FmWgHhLMPMzMhYsY
4i8JC9vFGEHcrAfIBpOOwfrHVT4wJ9fbUcQXsrS1hbhjF7Zyv0xWX9ycfRvQSgShFW+r6EW1bjO4
A+oLSfwgNxLGV4ouoJQ81ZYgJ522obRutJO1IvUVVItozhtsSeboH/65IxxkyT+7m98d5/B/C6BE
RU3cxvbyFW5ZpdwcYh40W418B63hBzZwWV/VswH8bUzyQNrSYNzkcZ8X9vgD7UyCJOXqINUxEPMz
CT1ANizgYYxUN1kiwK399+NhHwQbjmdymCcgMZxVUd2G51LP2dArlRZD3N+xxJO/LP4VoUVE2+2f
A0yZnyOzm/FVuugdRh68okz2Ztb+CB0kXEo2gzIsALX7biMClHvVwCz2MUaJiIWCr16tIc4TcedF
c+NypPT7QkgSyrr0SmOkmpoxtZAAOcQTvtL1boDD++hI6S8AQNHcXksWjmJkDayF4w7MQXjQv3SN
1uROR8j1hGbby2Cqciru56O/PE8FiW+E70vsUV14OzxgP7OfqvoekW1BslYrWruYn85evcu9NiCK
9qdqCVURBJ+QvNverCOuHdU2NVAju6YsZRqvIufKsjOdlVnPszlv2C8MipdI9lRk3AihLbcsksuw
QUzIszCvpO4Uq3zVpr9AMWqAeSGoWdEXjBD0rhoFRYml6+yzVcfbo9aSgZYQiz+BDCQVZ2/CpK38
m1VV3qIPyBFjoSTs9u8aO+ujHwrcsqR+fgMnVErGKkqcoJ921UpTYDfDKYreF3MeotvPaorar85z
FpS17ASJ4YswBYWse3iR5SGrqKPLYYVpZDAbtW2Oq0dGGi7Na3u0WDajcBG+2Hhm33OjHeKs0pLR
ev3DWlBsay1lxuqFHnIAAkaDnE6is7qnW8RK0IAoKRO7YgFbWoHgKOGc8x3IinZfh0t52Lr0dS8t
nRpBX4NSeA+OqKVsKexMcRzR4rlX1In8Ym1VRz6zndxS/IWBhM5Nm2pHIQyDH9XAwCeDtgMyxXOH
PEMlHWPerS0KcmvmytZaK7RYfGCVQm3nwkvcUZsccTEGXIy5SXwlbvyHphkgNOb4V9QsR7283Obe
Q//G5R3k4tVN9bTKzC7Ip/W/MBtKDGTv2xTagcEZhPz49xUIJ32sAxDLfjhSSUjpUxDKbzn6dfWC
QJB1/gCva1r8DdEZoh4nKIlHp651c2QGlbs9CWaE6XrzEpc1Z/osyQSvPU8pVrX6L1Yg0PN5k7uH
cT5e2ga0F3BCHSh+ONnsexS1r2uzYRrNBKPtYZ/xsjacqFRXQkcm47APXHChg0c/AJZN8EMLTBtw
YhhcssCZ10K+3yn6ZT/+T8F/ny8sFOCHGyGLpA4YfG+ld/2yh9By+Vb/hkC0xQDlV3LKI+SyNSu2
C0/i9mDahmozXK6kByi0ggJmyXe1w5gGoyydvyMiNhv5vAEx0nldjRMIQ/Xg7uBgOptlWADoRjj1
ryDnZNBdVWmP0URK0p5zrBWajNtKURRS8h+iaNSoSZfb6y53mc3xZoMF1HoZBVSlwCGNBc5ci5y4
sxacX6bhjtJIk3M63bbpZtlHz3BGf7g4dH6T9yOlfGSsRNSFOQJQXeHELiAQhpufB3OjsqcoRer9
dSnnFPJM6QjN9dbs4q4uf443kX1MmhkPjnl+SkAoOxTjX/lrwI6p3xy8L1CQN8g8iD+QYkc5KQZ8
1YGugyJGwXib1RPOCh8WXzF0R0uTmqPGEdMHBJN88va3F+4MOPuh8Ww0XxwKR6JXhjvIAPBhHieZ
aXhjgPuQbYSXZDQAEVkvCqFK/WtEoQSwi5k+/yG7ks2T38Rj4elg4qbhsW+7GovEoB8eCxu0WIYd
Cizmj+F4SoxjtdPbLMDHiJejZJyBhA+vDsehC/ZIa5rzSPJYKliwGfM3jYUYeGhsoR9Ef/MnyIqS
BuT6CVJGQZgCbhAyVf+xQ/OlCXKPAJjhe+oMbXd9+3v8c8zC8eQLAAn0HLZe3zikhnLPEz5Jj/36
vwTpe9cyzNx5Mvcvyx2AQ6p1DKTPzOwjXFy1KER8Fd6HxKs53VpF6mnEVYI2gBiDIXfPkpDLg6T9
cL/mJWnfAY/hkyG3VPHuDbLp54CRd1J0CKI736/U7ZBhpnO5Utw57aD9kJzxNrLZFjbmI5vrfYMD
pXwc/Ize8X4N63LAeXhC5GPqt6EqeNP4fJGhaodPVxeReojAJdZ0vjtWu8BPBuoVmJF+sji/vmP/
udFdFRr1Umrm7W6DbdqD0oaTepXhXrDYcj2yARVkoUgaR3qwGozK3WaamslKtssTZHe6JVHskBtg
N4sjVIpJoZZia8WUo4QKaHoZl+rcV/Jef5vx/PQsGnmEQpJlfPMawxKmxzyBUFRQ7ytACak0YTw/
v+gLVWe0tYhjViPTZp1tdE8ko1WKR4qP7etn+8EeqrYK8rvMMW+sZv5BFNBafeIBnS8xhZLnC6jx
VJ6kjw/U+sp+Llc79vHzbX5zt7bAwWniJha6sioFUwqSnmeTkEyvsqlmxceN7XdPIuTCgVPtNfwH
QAOreUtT3CpTZUYRQSQoM6wW4d6RopZl5nLIXYgGqzu5Jb9B8c/GVw1vRJj5z+RiClmm0MoGbrv6
UVN3vEHwEruySYMJE6s74m2bUPYVvptcdbELPA2Q98botowaIuaJXRgQBFJPbxkAvhNhsPdsfr6z
4AmdxpzczYXuwlrH+lItM86esr8DyL0ALTKXd7KWSNz6SfEdZo49fLualNEmT5m0mTIRWypKpwaH
XwUHBt4PB64o9fC1zrRln0omLi+6BtRLVN51vW/UFNGRM296zpVPzJsu0Akb2qSVH0PGT8qdXef0
DsF+HlIgK2qCEXzWShyPYaJCX1Jf/BmvwUreE+P5SodtjvBe13RnZkug3wANWKOuqHf2b8eijpF5
mkKlk/pKUBfSbUrK5hZvjSJlSnz1fXOpVEYTk/ZyJSnFcQM+OXaXh1cWMf1i9fFSZMon+yUoleRp
VMn9faYLQ26+T/MMQ5GGbFTkmzJJQOc1gmBeSKCY8wn1GtAKpKGGzayhf/4sOrgDrK+5Wk79Vexm
eqjWDhnddsXV5YCbGxV6fQsl+JKVQ6CAI3IrlaLx9EXn4YHbWmwg2FOTq/Gi6IN0kmm7CbkiAcV1
Y0Qv6o4CxEeCAQMv+u+K5GaKBWCtk813tII/VB/PQDIlmkk31X3pqNJLKm6ccc+gEQuapTLnmiUs
kvHnAtM4z4R9YOym+qeTqAnnGZIOs7A2SH5cJJ1xbe78FP+uzR+z6lEcS+5lWZ7boug1Z3/tRgi+
abTEo6iRyy9xDqAvlsqe4ebT3mXOfx/bjxB00Cm2ddbL+2L4xHQP0K5oqorfgW138+cA18o6l41T
CqsvHvRlFzeQ8e2dZ2vJjmBViNxH/CMCdyjtlc5ho1KZmDBp6eZAzII2CZUhXu/tJgyjPtpPhBI1
Ba//dizBkyO1MvgAH15IjwcN/kNbsLR1XYUyVkhbmeYPRUGxqlYs9HG0phFARg4lyuZEJjbg6UvF
aNzu8E9Rgl2KxKjuXJNnaLt5L9NZCUKTqa24U9JIkjKpwnSgPzDVhHvuK4Q68wzvf6vOZYVW/NCk
YqR0Otyk35woRf6tNhphPtsNqf9tF6BdKxVOHCAuP8+LuZ3tcNC863AJDH+U7+yJjHHdXKC9GAKc
z9RbQjow+yj3ec++b+tS58ihwGzwnhEUjLlbqvC329UOxt1bYbbwmRkirjfLGee+LQh//obC3N+0
rEtftZm9m8i/tD+yAnkDkcdOeO36h3FiLBREwUl94Yl7NWZW5DN7nkFP05n3OTubWFjpN0XZctsS
sPQFOaFEl/YrPIyZVlqCV8UQOZY86skCU1ROoKXrl5m5Nx28t02mZGnC3FbqioiWXJeQ7/xOggPo
NXAu82laDJVGKa5CJzS9/CUBPzvaCZoSSfrAid22J1iSS0dtbd/+FsS9s0ECQN1q0Ie2iF3bbkof
bV7EIxbW0AOUdJTqRrJrod0ONeKBqblclo2EjkgxlvvPU/YqfAYj29teliT5NMLcEbz63OIz+ZHB
llKIAc5OF3jbOk0PBl9brw0EGaw9nLfmncq9O8FrPnvkbT5/Z4gfTRlRESblzlpVMJmzzrM/TIp+
QM+pM4NTCqxR4uFiLnLwRNnoTIMW7uXYH+bwFGL4JNdl8pfF+OcOr1keMjoTi+tuoaP1t85EYrr9
hcSxk72qJxRXDjglOf+29YDWc2g0ZsVCFbaAcyNuw2oVjAhSGivrvArwfLGMuaZdNgIi/E050BGf
5nlHWMpg2gJa8vVFkiUOUu1a1fjfLfIeichibSC8vNwQq1Lc46XfVt3wfPSuUNATLjyMgEgFi5bH
8bkhhY6CCPRQj8PfEfN6GD4+XSgLn7QC8ACV3QHDPnknkqQQagGxiQ6B9pkYdAcXzUKMWbBLdcu1
6PWmS1V8BwyydXop3jgON5OoXaD1UnSrtsEUWQIkLOY71cpOjUXnUysenw+53h0ENOm6tvqO6Ctn
UIdEyZZ7YI4EuDPMvZzdKHZbXgm4dg10horku+FTzcq735Cv+pmE7dj2RiTq7yjueMsbEJqalC1P
rz8uylwUTpgcdBInkQl7eX4WMEk82/JJroAqn01nXnpY3llGhf9gdlHidrVSunP6JquC/eZrXW3Y
lUIo27lMAqsLTzgF8ZO3A+qj6w3bzpFwXUkWMmXe3u2NesE/A8Wt0dQY39BDeK5buDuxTgtIxb6q
NaLOankObFbQKedz3Vgg2AGu337ZCajDfojIcMck4tB6e7MWVev1XHnujdQfPFJSEtU4iIlCEPFf
xByFb6tMqWbuVrN4tju5bw8kn8sR0hxUdihxHLCEzg75b6VXVSg/yH8RuI/IQ/WrfNosIIM6QG6q
hro1WjinEMAfqc2rvZNcDAdQv2hSt2QD16AKh80WhvaswAbKpTPPtys9Ihdn7YKgVM82cxFwQuxg
7EnZtcXd1EoEkjkgElGEpXjfcVOVD+FWi1f67MrtosAgS1aBQmMvF1n1yquQhP1jf7PZzoDQEPZu
ylFIzwKBuc8CZ4n88N5npBn2Xt4KUQDI/TdiIQG9+8B8OaU1Iu0Nkw2f8d8uTSd7LmMrcHO+K0Dt
l5uDl8/QmWhvG7kvX3JSziXE86blaQg5NnCFWOeevr2FieIn9RPNAHFPhgaMLBGYKVFCp0c7MfvK
9tvQsfRVBk0V+Km100UCmtQqndMkFCfFeLDRH0ZDK6MHYCQrqbeFaDfbLF/pyf8AEguCgvLzLOoi
aQVN8Td8Ao3rZgP1jyoXo0Y93q3J5OSMLpeWvOSBdULM8Y7d+9EZGetyCuzOptdgqa2s349ALzUf
W7tnPV5HSWipiCRE4fRqMusJwpTHFI4Y4l4gFKO6xPrDmkBfvLxbZTa9fUApc0fixzstXM1B/IYL
zhGN2+7L4ZkOZtVIOG/4waKiX1fia9msMwepHj2hsXq/qzNIf8jALrn6vP0Lh4NZreHVWxkkVVJg
ji6fuf8YV696PmaXJCjEmA6XBUhJSNe2IH8W22XvBUcYFo93kynKePfvb+JqKlEOAiZ/SGm2avoq
dS5JffTWXvctdy4ZFuPv4T+MByB2Sh3JeEtPcSGHHJbRCwBOez2MjbJYKBy+6TbszPoCNd5kRK4e
NVYAFkVU8l6/10uzYa352rZaPFqtsVBrVQ4w2hKJFnfJGQsibZLBl+AgKaYXVLkSE9GEr7EMGwKP
PNv8C6apfXgOsUi2zFgJ4Vob3BMs/EPYwCgyLoFD27xf35BH7W2RNIYvKAg1J3tf2ypxwY6qdBuF
7jVURni+4pn8LJyFa2ZZa6EIYebB96ObWSwDZ3vjqS3ukXFrc/9jbho5TpQgE3O7V6pj3mJWJGNC
o9pAkFvIp/5K6MroPIQpnltt1ql41w9/0ghXhlHoGh1pKtxpR7KX6WRbmEvDrV3cZ/O6C68m0iXA
epLTTfRB6lJgVL84Kieha8BuUVoCABA+UK94bpnt+fOkWCwOK0kub43mn5e39q2fbbeYnT6fp+WO
x1UbwA4DaI77PmtUWlGXvkbj/OuGfgVCd5/WyQaC2unI4FlPAILeBaCOADbHJeEkeptSeayfnHkd
G2NdE77ydrB+ZdHFe2OPojGhqzI/hj2D/gvOx7pmUykb9m8aITt7vgTYpJyabLEN69A2sSBAD8Cu
9IvAAE69yADqMiUdEp4014y0KYOFj3T/lw778Ha2E3JaQC9pyzGLDhuTwhiwIfzvP6X0NQg2FubI
HpQALLUIL8FG95QO+nINwHj09S/2O8GCAEDPfUNiDhwfKnbicOTelazOGcgaElk4YtwZUUzLOBt/
y4i9Gz/5dFuV7dlUH8qTYUT1fX21W5H3kYxmIPezZPhvjflibgjSpyUvu7Txl9JDpw4sxVlvzlTI
ghSL6K/waYi2OVhDakIbN+otltoL2c75Votkr6T325qb6FXktPp6MNFiPkuHzDoc7cFxIIc+ma5N
4Ucg2Z/Uxn3XeR2XYanfyvLjiHuqwIuqw+5aZpWNSIWGNH4NJgeIExVDPH9fOXfjWVqgdNZ7oFCv
3lwjRJQ3ts0szrNaQYBqtFPhWwWuwNtBMc9X3oMoKscciKTzOeECs+U6HVuwBRhYKUe5a1ICf5w6
akY9lKbvRV0K4TL+8MR3BXUP/iXR2NOnQzRlS4YrtIeSDSp1ca8A4H+OklYuMmRmVbtCwF+DG2iq
XSNvjcOUDGd53gYQSbeb8zgjMuobKxnCpHAFs3nEVv9SbxvF5KapeVPwQLYV/dGdcce6vd2/OZIP
C0lv4Ny3unHz2wtLhyzdVZxi0UKX4yli/ov4Q/s1BppmS2womGRFyV6p0ZaaCvncbtMkXUWP+o1L
+h0s+fs+EFfKrT33I7e0LPcDDB1q2574719MF7dhihN9/juYEiFdxKfSEYWGhP78pCvy9qyXEv2r
Pvn+ZyzeUf77TmClKcltT0wWwwrcCYMEjA4tKXMTt8azQfc8j8D4+IFVuINhT3LTa5e0qjmYL1Y4
jqyELSpKkPgPPj1/sowduxj6LFb3HzHCBLp5Kt/CRQSE61F0tvAaRShS3wX1pHKygrZ70AhzJ3qQ
9dxev5E13BkTon8RJDbMD97vsHZ+4/IGZccFyOwyf6bq30WB6taF11Zz6zAoAwXMBipNtceqgbFW
+OSiV62a0+EIJ51gbTbq0a+tN/HAXH7pz/bcQ5tjYWet1fSaCh9q6GyCyG0OjGLEhM4zLxs0R431
AfmV0HoScvic3u6eY+gFI2jOxSDMaEEOdjbODcLQ52x4mzY62OSlmlLfQxUbh714W5bbjd+vWSHl
WNlwHHx3jApmqrlnk6zVzJlMmgl+ie2lyNw/ePsPsWOuqu49K3lZYSF44nlgPTRoyuOkVYemxKRE
M0qGSulila9UecryFsBJ7sTEOiAbU92p9AOoblhb/gzTkm9yMTVy4Ucr6Y2jAg1uon/2TFaZEsAS
Qr3Yx6GsHkU03B0bLeHvEyG6tGwggaLiMBY3J5fpuXsJ82Gfk+YnDMv4gGuCulpznYM4FQWrtWS5
bpu6P2IBxMZZc5bLS5x+695spWuiXfSCkuGbwvAKjUM1VEQAyPOxkGxr28MF6KNMYRUbo81rUhg5
XZwlWyHhgfTPduHdCBnSTAhCStIe7gVsNFGH3UjafGzqeLwe74BmaY8sTGUZnnIbOwNvH/9o9HGR
H7eMnbEHJWgqffPRFKbJC7lkzuLG0JYWAnQmGqsAgSZi+zk4JPuqhyBCC0qMJR0pLONYhBnS7/rR
AbFxCuejXcVqPUkXfMi+BV9tj2R7gKRsqFTUt5d6Z2l2XLrcDgqLO3G0/8//c/pOZpkhNCR3YGWi
E20OBTCufRtgSy5EAn9B8aak9YhtfaN6nNxUYNZR9/7vOGpjwVrn0unWmByZJNOkp61JgYSrzI9E
2BVOBJKXvo8kYo6MIOo34fYyGWiwgkC86FSNU29UEwFMCuNzky3aN7dPY34ACqWZ8XeFZqov9tnR
6uhaQuuU5mDtnxjMaOxpU4slZw6+OmmmB5hvgSH4CqWHxKrU47ezonErpqfwZhcBybTUuEvVId9s
yEEghYYu32O5DGacUob/gAkinacQrzMEMBzu2Y1ugCXKMkNlVFVV//Crs1drAwQuj1iMT6UHPyGW
ugUez7zVw+3oZQLs5BWE/0roHjMPGyivp1s1pxhWTLgEJKNabrUSGi+5935s7DgvL3IU92X7o4GA
bcfI85niAb0GaLsdkwP3cyu7iLwg6/rSnCZGHQ6SohX+lAG8VO3NRYH8E8AOsP+NXXkrlkxuZVvD
GlqF4pS4a6sfmrDbvmIh8URwSGFMIfoAJDr4xroNVMjFoX+jNorVKEH9mBajOaG8uhW7YoxQooml
Q8qdDmxdr+jU+5TeeJcCfZne1ZnrdyxLnjevJJVZoW95zmBbPAKgmkQoUy0axa9GQ/hi399ZAT+H
UyAQZFO0JdCLkuBi9ulTWarcp8DRdfRoIyoBofuaKQIQJQGz4eoKiJnWkGkqpXsMcTuuuVWpKaix
JePChfp7SPmYBqdUANUsZGbCVYAcFjXi1r+K8EqvoHz19Bimppt3ua+UIOAhVPBUUSMhS1UE95dx
oP/YkCgUf6tIH6XgWGIagY7xqraTa9DUX8JuJB9NJh4y9ggqyx+mV5oybUsgwihbcnhrrj4IX2V0
yVH/09xZMspUdrkL/2f4zMEZkdRBbpfQ7NzPA6mb2MZlbF4wys7U/2fUJjEC+Zb3fxnFSnaoXjZI
10c9eDCYkIotN8ZFIHOM6X9LpIjk/eTzT8TPsBHn/0Sy9cIpwU5IMQNHpOyIE3SdTqOJgXLlnhWt
OLQ+9rhp7sDqke1MjJGWEX48msmlaZK4uJctzHODIBITFNOg0Gkqwzo74T2aT9JfjyXzUFHD8odS
IWl3oiTXeSTaeuZ+x2VPUg6LOAUoycsorSJ9Kx+70ssmo2mEtHp5v3MwCmaXdiV11bSuotyJE0P3
HQczYibA3J09d7vs4YagXTKlRwKqWRa5foCTCoN/eFCcHUbBRnnRAjGo64fOoY/XpsCCKzXRsJDK
v6Tf4D8XbYcRyFQCeC1IrS6R25AJ4tAoTSuO/n8y9b37YWhRJPayPbcDBtEgsCyi//CZqmVSYelh
A5Ycc/5cfkDvXCDTIxCCnJaw+K5in08Gu8x2RedQuGck2k6UUrwzQqZo16jfMSa1RKrCzMlobCgK
NMNBNKsD7X76J0L1M8RFEnePT+lW90EpMmDk/ET6Xyol/gJssolA3E53ap8RSwgSpKcptSVK52t2
dSo6/n1WtYXr7lfB0XFtWoh4dGiecIcuMzUbqk0q+d9W8Sry5nvb6JcU5aN4OWNl29GhUc0m/sh/
Z1jtz/T0xHiuDdPtpb4VPY0ewDzTXzFAqodVMEOgtVgqfkS9Irb3erQm3CK90BC0Wz3KNeA+Lswk
qWZ2rnvyOEAmRDD/zweQEsjIspru+/Q2fG8061uGSa/g/jmXBZpiciWrsGLalLRKE5vGLGf9g35i
4351UtV6guOYJKWc4AAxk9l2eXKtjyOYElTQW12gQjh5OZrGRgPPDAXKojpg2ateu0SUYq2LJXRX
YB78dQRNc7wuLXMGkNfmNriwy94oulSxarMtY3aIkEuZ2EapEwidSPC9OQZfwPKY61aGW4wv90XP
uRQbocLjXkXn+5RqBYa1L4ycWi+zCVDm0IWD4g+30USgn2IiGFy5S0pchNH4c+j9JQJbJ+PfisKM
kDpbI3X/Z36ABSgXIZR2VbgxfxBTrEDu+nXjz0/8qH2uNURqye8h6c2cW68SocuxzqfzUM0z34YC
j6VWdktCc5cSdvUEFjraUnck3+mQDdD8EsxBBSm+RjXqMS/woLbhMhw93Mcy+j2Ed8AknFw1yZjh
YmsbLa0pb8IALquNA3T9r/XltMxuFHkbr6bpjKzNFBclMtMx3E6fStOh2oAnvxLFMZOq7VVKBPWB
wz72kYckKyNbc3u1LvJDMnMi2qi+CUN9FrVxksWTF8xQHiqOGG4UxWkjNjQOsrW0nasE435Yws0H
n0dmNnmME8XvbJdHGMhwaG9dcWBtcbjjNrSFiKwuvDcA4elhRwugDRfTB+NpzFzsvVxq7ZX/2vHH
hZsNa4q1phb4m6oZLtRDQAloaF9Ycvu2t6rAUDSFutMIb8bFNMeCjpKev7NiQnmuJhRrEE1DQkld
LHLEPb60qCJw/hX0krT6kJoOcr9c7c8ZwbGrMbnbingtNeCjmYwgqUW2htAbfmnHYSxaFn9V7tR+
vlrlZqmcUp4Un/HxYJ/rxEC30eIS/1SmjgA7cwbK2pjgQOPWUelsublq7xkto2aGfCR/uvGVrAvR
Rts7xwZ5X42Qnfx3RAYyQe49owMN3cYEH2S4YxJHHdaw06yaCth+liRP9kp67oPtt0577mp0WhKd
cl5y7vxvIzgxV0xO0T1uGkkql8QYxRlxZM6TtK2onMlIBYr/sbYAn6K8ujCWHuKuIW5KVQp0qfD6
g3cX1owNyXUHkZW3atTDbgV+2Xel7RqqSbTt6iU6Bbw0dYJHHfUsIkEWvOGF/3TasTYM/zifOtiJ
YpZuWgMAiJw1EGKUb0IHL9RrCPJi1p/Zw5I5CjrAwSkJnFcu6pWw3eLX7d62ufKWVCCa4v0iccSB
D/sX/cUXe4Y2SYV9RxweRyMCSAk1aiQQg5Beb3bRGb3s0ujbzxfIqxfBDHhJskz8j166oO5yWVPd
ZmNoMA6FyesQUGuk+SPhh4fIl5MvsjWYr74p+2FZg9oNVc2/Dkxx8DmLCunRjdg610wRBYwvob5u
pvnU1MgEELM9aoK7HPRzYDnsHxxxTuJqoXDzO5Ds1oYIGxsF6uXvQQ8Kr0hn7v4qS8OkBKdDzi+e
aDMHP0R4xmIgJQ01nFUnzIGYnZlHKhl9YBFzrI8hKaDzG21MXoZ2fbGrbfZiC7TnhF9dq+TNji8N
WLBudPdqmDkhi6DHzekVy4HbDB9EW+djhwYazPW0yEUlz05C8iqIPMspDQ7cXW/sSAjZhQpUo0ey
ZW2wHERsmIW58dL1f0VZl/KEPOTRXYrD6kEpa56lw1ik0+stw9XO4oD9xG5FTxDVhdXQ0g/DgzyV
90mZ1XJJc8WMEJUBcbLDed1TuTT7T3WfJK/sSizcTxlJ8S8Hq5p63gkZ+IoL4S+deLvxg6ymMKHa
Khs3CX3odxkIbyiFSsbzcLPLeauoz14Dm48Rl69KRMYvyX+dQC/+L9HACV8qBoRQGE21ZID7uT4c
Rs110N85GwJX4/KtI32wmakXD7doh6IunjtGTY0dbCMQx1oY6Wb/5tkHuoZdllW6Dyk5O0m8pyG2
7UpPF0Ny1lqbUOAYL95OlnJgLjJKBJGAlRk0FA6mwG2ZDQQyF/rS/NvAVwCNcVYC+sx9PjUoa/tC
YnNWwF29aXghIxprfmJYwF/si34PjkV/jU6rHzJRjtetPfKiwh3QZxNFrZzdgnvOc+4xfQs9+Nq5
rw7U2i1Z+pAgpQRLXl794jy6tkd/2CJVmQz6EDmOHC3ULDTWs+pu0bkjvjA3SXXfFR9bw8mEO+b6
qmCZnjC47CQp0NDzJ6PTf/gJbBrRgIPFaOuATEV+cuo8Uc+ujtbpE1ZPSm2IpD+qc+irS86ipU2z
ckrWiQUvguCERm6Vko4QX7svoUrD+Zz5oecCDn8nX2iYXhEj85JoerzSzmoiKi/4mDzKGsJHGZk0
qYcV4jH79qGl2cAlqX5CXnMmnkXueSun95jDYRE27MAXbcd24nhEkagXvCXXbQ9KBIsE89VPplto
Q2PsSKqj4MMaWdno9gfoMgpBKhezQ6PffM56c41IIwmpj+JnkSwPRicFAIjp8qfMXMA7Losa14qJ
13baDi1xYuxOt2jch2pzhCp92zj10ruFWcg/O0gQ3TN+ryWFMCY1E0vrxlv2zpz3/6ioiMFKbMuO
jo+HnI1TeX5J5D7356XUHD3T4E29hnAMob7uem1WOUxg+1OhsJH8Y7vOy4r/iTyjyNHvVbQ7XXdI
xI9ws39IFd83UBFt/yfjq5yPFXqKz1vvczyj5LIfhlJ0NsYeEjRWApT+im0pXS8CnjTUsemZg21i
sBrJ8tKz1VZOd8DSKASwz3GqZe/7OvwKH5RfBW9k+30LUc2RRqLEkwEAwNy5JfaM9psgq5mnPPCW
jj4eVEIUanFzXKAOCL0Os5wKWzCNiRokEPRu2DG9n+MG2Vy7+bpI6IY9WbQ0cEb8JqRbtrtBBUgm
fcYpU0QWSAJ/4QR46Oqd4YNIdZjjmGb3hWL3qpRfViJnFf8BVJfv5fepbvQNNPR5IcFdQKxH9XmT
xVmSvNCxFpQoVCC66MuHBMRduFWrOfNXeZhtby0iopXQfM8iK+3Xi5nCi6DORAYyYGcuSmp6I5f0
DjYla64rNSgqx55EqdPR2MQPc8TaygaJO18Kagu0Z6mJSvRLP/GxSnvdAoJLIDz4yKhHVsDsn8Rn
E1nXLwSXVU7AwzzvS8HpOft4FBIU9lUbl+qg7+VObRxGzoYJ3txiDiewiw3sb0oHB5ppTjPx2DR4
yoosjzmM4iUR0WubaA+ImoHzzjmigQ8GYuVCdlBN4orckF1MVr48cXAuUPEanNgICxvlmYXX5Kpp
kULM4UZeL6WhI6hvX4q77o+rPq5QaQpuUQGv1UYGT3y/XkFlDEdxgk5rsJ4n1MXw5k6Z/sxBZv9r
JJZmft3WFxIkDlQyZq6HYMnYmxm51O8XBJzxYKgqfemxOqt8EmYlCi+cBovCRnrQAkTeU3wneq6m
vDjNNxKlRquLUnra5MNaoI53WxJrq0g1j/ZZLPbzAW7DrMZWqYbNQOkyuiC6NIi6IVm1IZAjNz0u
0LtSyNqxFJtskHLAX9ibBFHhL8q6IE8heAWGpwIBOZx2whGq1YTARbiOeBmuLF2+vgF0sztexCri
ufUJHd1R0Z7l8RGpXZcfOwngigpPTG9IuRacBD1VGGc3nMKWzMI2VfHqx9OHWc52qAWNWzPA01Q4
xWFv2VTdP++g7cnC49+qSvk/Gg+qH3OY0RZ/rfu1XwLDaPCwCbChzJ6wd3xJuZ2wSWtkvpbZXqQS
mokvZA+Z18JI+kS/u17a/mnbYZJ7ozw6v+wOND8fIIiEnZj2fPk3IG3apDbraB1qQE1pcGYipCvw
7nmeTzrwXLRaL6CSI2HV9xPN28tPPZRAxVcBtiFQqqkmPEeDzqaNczrr3kvdRsoP7x4aZEeDbCaP
GC+iIS8Tu1t7sM9rXgXMyYAy63baSFXG+XT1zRfgaF3ykPyWb8NKtWZPgwtK4XemMviq8688fP+6
56Tr0fuGFbxPK6OBfIXBKvrcaMVcvJJ3EL2KxbCuG3xyey2CHNOgIDyMyPWFd6FXcvDSSnj8mHFv
7wf2VuvxtQSUOavGteIYc5101KSix+Jb008E57JNQjN0zw+bamGehYc5RfIH7DyGXOqwpjBpjZ9E
bxTzu60elRh4xpIjvQiOwnsmh6rjNqQ7HMbdFFbd8PuDh3kaFJqQTu31JdNTeMIU3ALO2WRkMZHc
mlWMrCVvE7mWFByinkKHegy1Va1PDM8i2RttBU7jnu6sWuZCiJtbTzTMhqRLXl7xq7sDjnlP37gc
scHj0i84Efypexxiqn7SEkmTT5KGxyJ+DW9MQEeADqfSdh0Vv+LvBJx7eUmoBFf0/hnVuiJD+KFx
XSs+L8s5lpAQUvb42EahnImZ23MjyXMFRs8xKTRQoEnuhG0VJhK/4lI5uzBq6VKWUhE3FEPh51DG
KhxdBcACYDA3O/zyVVEx8aSDz8UpMU2GyjO+xRtA6r61VngRsQJD2nnX2WVPPnr1FOJtOdY3GcDT
70E/S5opiLP075FhO3wcn0Yj8XvWh1ZC5oPddbPMKox18HuTnrwxFmxQ1k5E9cJPjFszFLBOo8dG
EUTpru7DGbTj1XctGRejFAOXKfJCde3yqPdC4dz1eX8XBPE1WcRycrs56PvS2XtHMYJiGxpeJ1MG
D4AlRKwQs44MXVsEXeAqdx4+9Rb25AzlTkymD3AZtCyFzkQIgETLY9b+svE97/fQXsTVNB+SadYp
pwq4Z7+nTS+/AUKfwfmFv826IMhVkuuxLNvrOyyw83q7aGScgBJpDZLizIZdae3h1awJCDLHnr0+
NSPrt+CJSreqJxkp7D3cZYNnYmkDHlyqclk0EGmojKGyskwztl1oQ4WXIsy3mjWrXV1TPksPAvNH
r2XwQwa6RfSPPkBrsOylk1lsoBFPpVUTDyCvLJt8v1ea9Z1sS3PvhKXx/MiLEu1EiEyngiB2AN4d
HuyvQ5TjChqLjn8zJ3dTsacbDVa2htdWgnBN3LaOOAYjJyYlJzjRgohJYu3blyoA02K82lJMoo9l
G5MPwMAFV9exS/zo7Quwl8UKmV2tQC/y3YiEI2p9Zz+GyGQ+AQTfxuB9I4eGPQ+X4jcMpZLVBZTP
b5o9rfU0WqFEkG29wfKrCpVLCCzUoXQiBXxQ9VfCjruflmUFcUPwwrfpqdRI83LCRCmEuK4LzI0G
lHlQeB7jmvSj4cWBshhL1teboQzg+OFwHte8uZs3cAw8tgouExlyy+aU8DbZygn4h5uAqSiS4JaQ
QtF8nkTMkcWWa73RB8trMsQRzhsedSnmmEtUyNih7F2eV4f3xxl/p/R9jfpwNQvMz2sMD5KStRXM
MwbN6On6lNy5ky4KZiLGrxFh3CG6xN9VvKYDJFaOZ4OgRO3useCjeOE7crlh0SE/UurMUiVlutmY
Pg4t8YTnDP/lTWD7sZT2zgIX+6HtUG1lRNS1RVDPrkPwR4F0NThQ4ee8K2j37UjyqXBvFvHlq2B4
UrcuXoTvUNb986MCsGrIjRDrl5PtOFH08i/sz6fBkzSDnc7b+LhFF7XN4SovzLVYHFQkqkj0ilZk
QoqkOfOiGFv9zMuRx6BjndcR3u8ISfMx02i1dn8HtHtHwRDWGrtCOBJp5znoTqVRa6Mm9NNeAobm
HzqmOyj3Jb1yLjZDlHYz4y2Z7W7T5zswsq2niJhLBOZ3SmVbv6O2CJ0Iz+0QPcmRWweYYQaY4dw8
KSg8gnko8ics8VGPRr8x3nTNBkEGzH8qTaTBPa7HmMsFFZkqJD5qsuFv4VXdixFcIRlfm/vKL12T
oaj8LU3jThP3rwUeikcod70V9JgaqckgSwzTXvJ4ZcFFr0QBZukEP7KzqYQXrJV9M0JZacrA+rHk
nV2DdLIZDmVRJmgy0bJpGF+eHXB/UBxtHhhc4yA8gQhwPGeq5wmQvrUkY0KmFeXHAekbzgC3GX2u
QA/+ekfRMHTVm23vjJXFPvyYejNicYgGZFDO6hhSoO5cUAkNU9dNmtySZOJRgUREGL4D7MsWpLsq
ny4EUjIvCRA+sK9JZkKnFtN9hWvmI7Njik/RSzNktSLgdefx9vuhxqospw8E8VyHTWkXbiamxotO
bsUiR8iUydLlH1doaVpnrCHY6+CHhdRR8kLuxagAaxq5FGEiTxs34IoipN1QT4pq0GRSeRKhqj/q
/lFe7t9ljvRqbGg7uY3Dc5Nke89oo3kZPVvtGbWKmQiygbaUxPlwSs+4pFM9WymI4ez+ZbAnDkn6
AJnHw9iyMjSQerqbCSK8DTqUvnPP/JZUzCCi7wc/fnpP/BX08XKvPraX/6zO0HU53o9kMLPH5VFw
wi2Yj0si3f5jzFYNk9tRvNZmlfSUGdXAlLuWh0oIxLqDLOjiFrfWEk8FuvYLW0EYZeSpW0GMlgpy
35yNCDnVBOuxYbLSsbafwwzXJHEP56ETYOIJw54X1mOHprlI1ZLr6kjbFaFCVfEFQr+AWfq5rUYG
Ysw4ohdXv9w8dGBTDRsQ2/aXBqcWdsIYlvOIZFhQGGZrltH0El8tk1l9yIxG6c96dJf18dn0CnhW
3UTTEzCeP4Yz/W5O80efH11N1c9HNi/96pe7qtXhYz5tOrF0ep/tGmCJ/TzpFSjT96ZmkJN7ecFe
t+VYN3L2qmyNpLg40t1eJNibcaBfaWpHUGKEu7bVSPq5B3MtQCD07190rSn+YrxCpvxmQOm+l2Fc
8fMTCgzPUX9bz1F6IQoPSynmudPq83xwjmVKDWEWd57gUrS8/jocFmFVOHWUj1k86sEMKT5UDMjl
n4Y3vbQCWLiSW+G0kVHxO6i0z+qMQy3QB7Zrh7B1BjcUDQghsKaQAvoR/nyaPD0/AvUOYBMK9auA
WhCUhOJ+LldwKxTmCNJVS9MmDekP7ykFwr4wewhHZ3EHo5P8Ca7iHiDA+FoAYI7Eg2m0rW9X6uos
8nYoZCyMDQnZ3JiDRHDSuMMUwLJxqHz0WTDSzqhVcUiYhm4wV+zVXjIMlPkamHlHmgAP6G9IQg2G
/BGbnBcIEBayQOQOviocVMJNLq+4TQQvCM9PyMc5tec26qOu0ndSn3FwaUOAaE8/vLGwXHV2Iaxw
k327HlWxQ3I2mBItP+y2k+i9YEGMYVVBFMBS5R4wVpCyrSpGExp5DaIiKriVlarvHq6EqikKFPRH
p3vQktp5gy9JJgb3KOsHcWxMtOv4u2aRvzFjVZiY0GYRtgEcA2P6XioJTkE1mYtR/2sZiFGgv89F
XwbyHbsw/ibe+C9GIHare9GQFW1a49CwjuikybWUPCy825E7RdZDnk7aSYCjoEce5sATKwyPdJAj
N4S+bsM/8/SZ+hxbEWV/Y30pE+3L77T919o/BpHw09qvcWOaoWQ272WtBQIn/Q0gKxo8pjDlz5i1
PBEGyXT53MkLaqbMf/g4gHpQOEr6aY4uOHkeZXiqu/t4JPOYf9Wv5AjKEBSglKOHyGvlPT6KzTp0
B6hFLEBbORF2HIY5ne3S5Blnr0brvIeAHcbTGJqovRWRDRcMWURPtBDSQKRtaMY9m3rcyygIhiD+
tXwLopln0wXkFBHqa73bvm7AilIIjEE0nhgm7NZ9apZ/Y+iS2qfNSKqFzUjLHpthw3CqSBHaG8fd
FNwhQor+fK/oQeUwR5eIHf66S2aX4WUEbajKEi26ONS3k41Utjbol0lsd3YuFnyrpRgWzNcbuQ0g
Rcx4QGqOohUYUj2bDiH94QojLOUKN6gCJ/0XQXK/ShNXTb7qvnywDWhUh6vtvtP1kvyk3Uw1pFvy
WOmbca2itk2NMeYtVWUw+cigotrKjpSbFZHbR0NnpUIGN1IgUL7C3+3GZ/6R8P0SH7PEPmB552wY
zp4sGNua3roGuQ7uBMU7VtGmcPI/q7LQxXU5gLdyMe2EZlEPktMQ+IUHVuGA44ZrCzjX1eoYa3sd
bgLmTqQ0r21FcSx8PAKykVqCbdhfdoI0L5Trhyc7WIF8Nm9k5YdPstR0Lf+aj0ArUJbGv1x9uBZy
cRvLC2e13KNod8ktGvIe4SVpeNCPlY3FIYUFl7lfIOuhbgKGjJxbnx0AUS7Q5ecf/4B4rEgMSoxY
5Hz2/8Ik3ZghiDW0fwyiQGi5Iqeb2vyMhhhdBgKlqMoN7G09/z6JL4NcCCsHAPEe8WVGiDHoNDQb
WOvXLVYXa/1mACJCHELaRShmYgsOWD07wipenVYP3r/MG7pNFfg8e7vAlk/o1nHgVifHzebNn3IL
USDMAXRA7iQtqzK7psE6koDfZtCSdzTtgKpa8u2hVHkisYpvUx4XemQzE7Z0SAxobL7L+qc/GTXW
T3PJhbu7bF+prOdo14k+7qS7P6ffVNSKwwjjcjHm9RGpliGAFAizrWPVUaYIP7vBaulGLhBZmeEb
4mKY09lWOQUFs8eWA5wPvYmXMSrKPh/ojhNQ1KiDhEQoNGv59GDD/95wU4EFoIVd6TtAVOBj4Nm8
oe8Ma5RSQe9H+ZwWRa8Vu7WzwK1Y5SrnrqHnx0GOWFv6cLI+3RHtrITIdX3Uzn47jCdYu9UBZBse
azaJDORzvcj1keFC30F6Qx6CBR3EGA5yPhM1HgH6cQH9zAG1UJMK5prl1JH9aaT/bSULrbXH+zJ+
nCHVOeEPzBcrLSOzbV3S4KtMd4m3rJB7+bvC8FCPCYsdWMwoGGB4NoFIPaC4h7Ecr18nGZnB6YMV
dBMJpyXUAEIEsRTDOAVB4nwxXvTkc8KI6MTzUjkL5o89fDsJ84FBhrHLZFOWd6x/Gv1+FiHSlVn5
GFVOsR0RVv8yUKi0641XId9Jrd+7grbgZ1y1K994VEGdOEX589CowqUXIOQFJr++YM8AFCP3GCUa
Qfy+eIdOpFtu9vLn+qi94Iu4zufhKCpBSZWGYwlMjvVf3y+rDmwofEEPUNifHKP/yjjt0i0BsnLN
SC9FIzkMc3ZsU1Gk/nvk6WKMBxdGFaAESoZlw/fJFpDv3Vif7cO/kN+7wXAck911W/nmDsotkFTh
Ij0pfjbkmVuY8S20xppeOI6dcSSEBCmKlwGN5c1FAvCnB+42P1lKV2241E661ghyBKHReaWspYkn
NXQnZ4X7CfVn+SUuJ+HuPyTjYRIJXLzzgIDhGv1laBY1qrZJNNBfigV4lmJGkCFASloTMLDrBvpl
6G41rHEJR3agPnnPJWzjQ68GRJ+DnjF9T5oCdDTRYDYls7jP/3ovFZgzxBJcQvkRubaPAiF7I+KK
EgKuRLsZgqm5BhgJpDd2nt1PNPYxoYRAKQTUDcpUQGI8v18ZYPEUVh5cPwX8x1olEqhinsrzFx1v
sozNMz78xerOoCzTk2peYL+GHJlJh9p1OA8oVRu2z08H0y6kuIIaM3BUFUmjEMM/50dGy2x5FiO2
UZUC6l/PGlClmdj9AiHMRkqsg+llPTye5R6D875wUlnbxAevOoze6QtCdDdaxoqsCfyM1Q0n5D0h
14SEN92wzBZUZLeYTK3eedoMdiUjgttKzkH3flj0nTOD9QR7CU6ty+XCBLseBRkTul3neFvdwkPJ
iF+2aVRf/HuAqWliujO4qJOeMcIi0iwQN993kDECJ+YDraJrvLA3krHPR90Xd8/JANVZ9YR2GZkB
AQpoIeSpbHIzgfMJu1Cg5fsPfcrieuE637Mm0yGH6s6D9JJfLPmFUfkhrezRLjcLUiyLjjXSWxlo
NO5Ysg9eW3fmdsa5xxiNUkk87syFpL81nh6iIwWtcBRGgiYzptNxJHlyXOpEdk54TiT/O8aBgxgV
eVj5CzlthbY7/BGhNKLJ2Pj+eyRm71YWKjEpXtJ2RhLjOMgz9jeNC0CJbPnj/xR42E9OUm8OSDwu
ooP7+rZvtXFll2ohiS+A69MGA2+3efGJZeEm1VeGbC8YNunxX4rHHI/5JOw6KWnOC6hE7wHWNfWd
W1hodw+JBSwJWaTREDwUTU3rLgKRi84GeIS1uHN1Of/pEPU+Oxn1VBUiCj3ND25wSLzr2hfCjmeo
NvfH8Y31zflCH5SqqTOTuuCN++5t6yl4m4oEFvWagTC8pRE8yEtP7romhN6mhwCo6RLSxcci8UBz
Pa9P5t8Y/OZ4CDze1BOv9UpBa6CBz+71ymAoyOxk70ngLpg03saMH3NF3/sf8tyWZf/fPJgswmrg
4TeO9ylgo1taECiPVcHzeYJdJdQZ5TrKTGSU5ah3gRuwcWVbq1LeSRMK2RpJV8COlVWfziPgOGtK
xT7WaVPd4JONS1ll9FlG6YtwHrjM1zMTQyFTl/QUiWkBFT+mLBNCUKtMPP1og/GL/qrZLDOyHcWt
6nK7E83ZhgcT95TNGBnWZgvDgT/7na2a8x87EWZ/jIkc8Z8npRBTkLcQKLksR2T7H74Kuh+/596D
FJ96NNondnceUG2gBPKdD11JN4bgvDlGMksBb6ESiK0+G2rERJB8OCpumjtV1Fl+qsOVmaFroTjI
xn7I8oJFuQdCdQfuN0AHOo502P9RWuhiVAXU5CUjYIHp6J0TuKHM5FxEKKHEMsOeIBauAUe4/XSH
erIQBVQ91Ncj7ygYYYeb+jmoRJKX9BFbvWOgEVEQJU/lwuN1twCVUpmO+/bQ+mSzcYiwlgld3UHt
lHeh/34rDs8OydnzIF59u6jA+B+KXuVuez8H2LnrD0iIdLt6FC+tcdoWzBqgX+V3CfCWHqKJL1P9
slraFIqOU3D3R3GG93Q70plAecm5EDQ6t3TmOnPPnWzYFybS8ZR5v6YVaP2t2uSDYOrLVw+b9AJ6
NdnVl8L6RhwC04oOwfoa9f1kGv0EJpYqch37H4fUj2sdpayUOhlvHbJw6A0iDlw3ENBvbRhulClx
PKfwivBLsxiubwlfF7983RGRGWBqPffDqHe6xcXWRd+V1SMWf9jwCKt/UEDviE0h9KOF4ReFodR6
2yopVReST+r1AoAwfOW1bV2LtAWmcTvyTGbqtYX2CJ+5d+Phcupy0LbB7jZ//DgV4x0lQtwMySjP
H+lZFXO/Dh7LOJJ3GwHO3WXZT5NTKR5Sl0dxfmugI2f7rPvrpyI4nfK+JzZmeisu86TtTBHtGLbj
JmNQtcvZfagWnzYgxbEmViDgC8Ht/P6sBtGXluVV+PcIX50BrvgSDx5GmeOiCnJDtW3D4S6eRBBJ
t8dhe3Aiq8Tsgz50tKGAd2aDF3Dm/AosPg7Ma6hO4z240T/SeNqy/37VO8nqHsw6YGwqKOrAJzGC
pQp7FwxPCWIXxbU08CsSuLPWbuLEd78LE4fwUSETTWxtkczKVreaVl1TliFvTOsFZx2VM5Y1gPM6
iybqSbbQunMBiHJryo4cLFkVivm3SC37l6307l7aTA4zo55tPuCntY/bDePGOGjySywxOdybxJj6
dlXYsYeWVk6RfjVSnGKaj54J6p5nRvxA+ZyKsbOlq5xEMiny+wz4y/k5kKy5uBRaaAnJ2sSkwk6F
YUghgB6ImyHXUK47zTeNnhfEBc+Q3iD8MaAMMKijiznbnsRmIPfWkFEAF+WgwC9+r2EoM79dXRI9
hglbOANwu8scDNeVb+45zNvNw/2mYTQk4df8pdYOyxXA34cAae8ZDqAichg01rBsZsff5VFWVsEl
6bdooxrYZ+yIhdjUiaEak48ICY6C+bulCrY2TVxtT5ek3ddmaLEdzaYVZDfV4mG1E9vp08ZeJK1t
+d/Ij6E2kL+vX/DbviOK16yLeKJ/sL9uNvJo42ihrUnd3vvYqg7S6zSvqfinRQYeqcQlXPIJob9G
iVxcrBY6T40F1QQYJ3+fEPBxZUKtnDPIY9oN6eyUXDQGFwD00Bp5Xr4ROG4pkp4W1NDJdGTOqyfO
NBaNQCiTgH0B5DM+fQGav9ZvlJze0DqIIHrFw322Rks9cF4Q/WZg1tlLqc3SpWtsgZ+w34o3EGMz
lb8sxb8ikTaNlbG19FHd3gQ59Kb3VtngwH9gjtYiGMW5QIBfRxNSDD1BoDOilvECqHWm+QTVrr6H
0d539W9+1NvbskAG7bVVIgmu8fK31RpCXLtlB0zO6+N/Id85hVsyWEejG5C56vgOY4S4TkHQByrG
s3s8wcjB/wNkxnCAX+K/cGNAChyDiVyxP/HZVQRqRQSmMf7N9eD//KHws2Wci/MtgTqEAePx4tut
MDUGeX9ImbHAc7YsW5oxNLq8p0UuDPr3a1oK3ya7Wm7KNV6mvREb7juHd8Gt3AX7ByXV15kXGFOI
Cbu3Ol4pLu3tK+AOvZJJVpPh46Ui8iDKsKTxvqsqtN4mIIps0AV9VXWrY1v7j54Cb3IvR50fhsgC
ZSDDnIegGtdXLgNxrX9wZkbJ05KF7HTR6VMHb+1W0i4NAIU6eS9DY87LZP1gLXkDInzBpusb4plN
QVzYS7jg6NXg3P/0FTacVCCC+xOH3gB8EbDvirIJQpayP/cO26JqB+k5Z8OfH3jQ4bogiVlX0z6d
5Ac1fNwrzZi1e8zycWmG/36PjS+d4F1a77nCYrUf9mVUhZieLS7ZU91ZdXPEaLXYsDk7mMyacn6K
mzROEqhCMZfbAzcnpc5vQFTXgx7B9gl2f7JMVY+jIuxCPJY9UYpRDbdIqDxk9pD5kr+ELb3wSaxC
uJefgu+Sfi+8sb0A9Wpfrgj2pWymOWhGAXWa5/9RwNYGIoB/GclTB9gl9CtLf8bhu17CZZ/cMRJQ
w946DAnnYVP3IblKu4RKLu4sN5EB09nDy6QBTEWp/n+mJbshRAbLMwnwJSJHIwVopkGeduAFr4pk
o0jWRZWT+pMDxTRgJ65nYWWROBUWXShSXkY9ouVkpc1Z6ruscjjKmo24ZfIXrFoQ9df8GgztU5sZ
M7ggoLZLMg7tTDHZjnk/KSOqAni8GkoNXkclqzK4Tu4dYh0LGu6YPZ1pA5FBZPIAF8poozUakW/N
5VcJdCt2sqvZ35sCsT7i0ujO8eEu/Zy9y/mNp7YKdvpfrrd04tG6mWOVy+onrQhX5QHfp9cZapaz
ilTpLI2qabQBcKOzhZAjnjKXzycFO9J5eDVxVxgFMsfgYamgwKrzJyIPB9QxEq2ApLjZgpfM8x64
ta4ZDO+OPKePa+b3X9Zi100AOLHAgZPm2+/0vUJJksuih6Z2dAElALpfFe4pNih+4CaH64JeWo3s
qFgpecO0e0aSF2PJXXht0lgXS2V5DURTNxe0ShprrIAGdHWAP24QTCIfyfTvlLhVlyvTA4+sdwum
BKCpoLOARyYS/bevzJ7zXbFsDB8KmYA8PXzaxqUIYRoc3hlOyij8oJY77gDnJWPw45vneg0ftJOx
s2rmRnWUWeI6udRcH6EatxilcyqV/PGQXAP4e5/Ahi/tENiLfJgOZenOLm94zoljLnnGyjfYp6aY
p7tSsLV4a88hSeLTpIWJeRvP6B76HSnRMOOtJRU6rXJk3TQ3MwwWALt3D1RlUYXuX1vX+a8RxVLf
s8QM6MghLPLY/x+OgaWDNzgTFYaXeKH3JfJbSlc4vTRccwDUQfnXpceickzTckbSZHTJttuLfvYd
2Ntv6tNSeHZb8OhFN/oCvjvPwKeS/jAzwOozMZYMsQ29WgQzr7yiuCfMScPnApElNIoOt1cV8KQO
n4808btupdaYyhG7rwUAVjKPgkIuIe9GyT1yNMfNclE1RCTKYVJdolkCVRcjzn+HF/yyTz/MuyD+
wQj94JmMQyFAZdXU49UY+C9ZleAXRe3jqV4p0+G2hI69NpyjJ4RAjaScjnbD1OXRftCb3MJbBavl
surmlkPlH2nl9A8sEG2syOEvz2RyPdDTbZWF9Ry5HQxtKcQMiKjvC+jVQksnKetpJHkngDA1n4y1
lEjSX5bvr1AVLUzho0pjZ3/jxmuNYiQjzkYdw19BOeEJPqck0/qa7CYt4xFDjeev0gxKfCxv/YiK
eZa1X1Zj8xL+WAZrL8B5f/40RmSz6eA4v3wN/BhvkEd/fI1ZlO/Q5e6NT3iCfBZUyTEcLlpnxmJr
HK25ifFNz/BaOd6TsYyjVCWp9AKB2GRJsxb+CdbGrBeMMPH7EMpflG8/LRowoM5zSvaAhRWeCUpq
pqbunxDAtNr4X1J14ynHlHhjaP7OrR/EZy6jnzjMXLxwnoA8xoEd5a8r5O30ijBKCQfyorPR9KtE
d1+BrZWFCfiM7TLeMkaTiM3j0SOypMxA6o0XCh0dMcWlGcHYImFqp0ptQ6KeMoynbR2otuiMB7Js
aiXoDjfatVMHb62I15SP2lmswotp2SRE+tglBtmBELVvsbsoDCmtB/qlimwOeO4V/ryafykBcPk4
9ToHJJRTGH96Ycuwg/QbrNtXV4cV9uY03WtWFUBmWm6wV3IX2HPrJvLCLnmyNaG+r+ggyYyVdhBT
rA59NMmeVV9zd7eV8vUHlyhrmX/wZeBoQWVXVSC7f7RblQxVe9nPEVXlOqXMWFIor7AUFpgoOwX5
b6I9oKA6FgDwf5evmKboAOyN0ODxZC1J2WsHU2b8kTn4bfcTLofwwHVHFpRUMKe8/JiyZ0t7aCrs
dFMgGHJPEDnIMHbUgZ4MlRBj9XX47d20OlUM/umVtIiobM+Ij2w4Bmh2bZK84MRrLGSZ9+MOCY8B
zOKmjN2f+ycNirdGnkYDNKjQ5EvjMc60w6V7cB+TJ+2v+kgG7i4Qjd8dSn1HJNVp+RQhOJAP1wWK
XIwBlkMzCGc4cqtbH07985huQNWgalMozKfljgI3bfs6UgkFsVZLrlqQ2sUCNBiV/PQocmN+egX2
NzFQ5rE/BPJZy6VdsuZjeVOhHHTeaWIdp5Slp2AJjewwUrWdBEfu/nOqbKC74Tg4rVVGn2kvG+O/
Qr7Ei7PCKFeAdGKNeeRYJbxUtbW14TtJeg5s3+jQRgrzTVQ4cZIZfpIKyy5uHW3zxb4ncVZ1hafY
qUdnpf+rh66EGu8EbsKOfd0fZEQf31iF1ouTnnn0uyrUj9KHr2Oazzg6hLQdQjZDsYD58APMdO89
NVi8FT1+jdm3uPb2EGEwhziM1d5VuYQTMjPLHBjPUrwnmdI2D1h1aJyezkQJ87wqEYgKOGpYTrXS
zpwevLiMsrDkLdvd7+uZSK7CacqrbqdVzzbwfIbG8R9vdcPQt7PIOhO96yMZ5S3nX8orMKrJbjKQ
MCxqlm8eRWN5YsG7oI/GorRjOyeHdv1SA61V7dvC9fxcB4l9sGXtk3QHre+qpYRMr05b+5ymdJxe
En6ailPAXOrRGFGUJKWjfCLNjqy8z8U1UHg5tJITBd6cPid2uCTSQlO5Y6KfCDRYuEyHDMGfrsTO
vIRWLoZzvAHLDlPIRh8H4W+teDr6OpVzokcc5MX5Hwrte8aVsJhBDwxngNzbWCUe1PEe7GTSupdn
b+f1qeUI0utCShqw6jXUCAPeUed0MDXHdUmZvtNjLUDCpQ2o1ZKcalVO5DZcdlgLg7BoO4Y8eudZ
6kYkaw+O84OCLq3nlKg5wK1ZbP0HiNZSnQKl2F2XD3zEOl9f5wsKGaEEUyhlPHe2uDRwmI1CrJmo
ab/Ln85vMj3fLOwxjUWmlxuxEhdzX3gjWN2P/LrLsvMlfkDlIFOOqTzjXeMpR1mX+SBjKzZiTaCS
epyZQ2WKNncSlHzraMnDXj8mKTWHXdQqHOKINInglUCC77T102WwRv2bbWVjYwVYp57mVyCQd0gY
+J1JsDrYK3mBwpDYWf/N3yL7TuX7jkd8CkKbA0r93ySAbsniKkZ+K3JChPYkg4aVGk9vPWeuWIXt
rOp/OCi8uDhiIQ7zDmvEGF7IPp00XsiID5kIfxcKK4TYDBWZ2BcifFD+ePYtNiFTZSnMrS7IxLAk
lKqxuwqAvVPCL9CuJKhi5Al2D8ghoaXlrbtup3f2qRHGm6n7og8KTw58r/TpPQSg9NxM60bnwO7r
l/XfLv5xXvxhbPD1+ntEAYMlNt0pFUSH3h+qxQpmag5L9u0YrD0XkujzKXQNHMbIIm4YVAdgjVk2
J3vSkhjox0mf23AxtKLnT0kDprJPZ6ICQy6OW7XL3PjPl4F62escRMgr3t1jQe74FylBdohE8qEH
TxgDm7D1Fi5MxYXoNNS1jE+aJk1EWOmNtevdaVUvixy1+TeIhs3jW+A3Wse9uloOe3WnDqplToRB
99rCGrlrRHqZQ5T3CVT77C+5ZVxMGfxv3DCVVD00vid9nt7Lys+oy+A96yfOi3FkU05Phy7hMckk
thG6niYg6R7L4M+qngduL8F7dv7XYnjNC2i7J49e1X/88qKpyEn8jwEI0h6FMhZm5+PyzyrhJums
G7vWmLqkKjGZi2iMw6UIdPSHwqCQnpxQ2jjKD2U7v66aftWB1ly5oqVoK8dTDuSCUD07k6/5WDSS
NjaEkhl3iVOB/PDEd1cZof1Hyfcjce4xNhMxjvmiSfdWrKz9o34cSZZXSlzNyIXG2vm5NW6akbXr
8kPcZouiMXS4oiO2LccpA+/ea3AWKsqFyfqQ+I4BiH6lVOcPdAvk5l1LQJc2xWngpSu1AN+7n1qv
i+1PthRT0dLvjrHN8/zUAjMPvNvSnfsjraGW9E5fC/dBbDhVjDrsESccgz6gOAMe3/VwKWPEpWXr
cw9bfgpmcA4/gjEQwSpOJIX8Ihsmerr3sM+BWfkGQS8spTjIR2TaWNw7smzQ7dwmVtW6eq/jIJYc
tTTVVg87M/AsHb1X/AuwFohWIFhPfsofRnNNWIhsHtwzCO860XhYEUWFr3uLKQXNH10w3rffUDHt
I975LMKiTDLK2ubT6GAfpnG2ni254LryZIOktRmdEzeXaqorrBcWPbt68LUh7qrbJF41Z5XNJno5
Bywu3xt16uo8Gmwb7BkC+RM9x2ue5BzVwB/rruym4jEtVmgtE3NjH+ukVknEfHimcquMOrP0i13S
11f7JoWaY+dv3WNqhWd2nEeDOaS1sHaIV3EuQ8Ug0BgCqJFjxyKfIX6UWXGomLiwakVpIln33LvJ
BdCH0e/iQyNqSPaikWHp8htXwU8XRRY3ToSvYJ/kv75HcwHyUjnqMkvfjA2oLES6Ru9rg9gzOQXU
53XNpnNq32FDEkjhCv6U6XL7+BurQCdiYfRYmE9WQnbnIpMDfZ0A6UflgpvEpRi4xNUuVmhXXaDw
zDl8sV+byDV/IR0VAg5Jz6cz+tDNFj9d0bsUcdKRYcjXr5nwd5/8F8VRrpybtwgjSC50o3bbPUz5
tqTKxMR1+/JZ8VKCSC+ISf7ES1S84Mq90BwccORgjSoWP01LmNR8qw/IH5Sitb4JSFZuYLxUzywa
pwpwsibdaM0D36XNr1G6NSs2IKd0QMo7pz2Mo3CxHw4LwBkaJs4pmpPr7bJESlrZ4V/auBr5+5Ly
mcXb06BbwmQPR+MysFly7TnMC2atuB56IbipEu75gYb38JQk/E8YPHZQgpN2pih7mKxXWVZimDzW
2Ptlc5s0rXXyXKi1M54c2uOFgodu8tJl2qgu3VrCukooBGnrg8viNwj6OgQg41SoDtwy/zz9fdqp
z+BWhTFJ2Oh96RuVh3nNQ+Zdm/FpN3mtf0AJ2U7ESrgMWYW6seWFtLfQE6aMGJisnERkXpoH11mb
+JY/kNglwfYQUFr5x2js8FZU8Opcoxmc/gBdf5ePf7Ux5wA+JmXnZXHyiKuLH/HYQRdIQ1m1/0KQ
uU/NQc3bO1q9ZeT+Y4iHH4lNt/xtxMDhvg4KSb8NkBS6CFtEQ9HjJqJI5akmD6pQu6x7ww6oDpXe
3qXn9R27hA6EzXChCTHd47ZPvptcu0AwOF6cN/COMRqviVW6bu6tbZoNvdMsagAyUPNjIa7PJpb8
PhlcMM+JbOEPUPnBP8kLLWg9V3+9q5cgkx/UDZFhVzOd2LUxPmDuDOlqNsjzmewZWIIlTNLc0ius
OOtoMGqlQeccy4NJXyU2H0uu3V9fMUBf3t4vEVW4NxU6d7uXpKMMMWF4trzs01a1yGJXw6WOSuv8
Vzk2IbwCfzWMLrEpkY3TnSqhh6vrY936VDzfrCCLQCVRYRiPB7MEMN+HuxFWefHojlsCF8V7TqOF
vYBEE8YXwuIoDUvoIGhufbtadNyaUwPu3lLoc9223JJ4fro9aQbe7/jY673Sv/FMO08nZnQ/lX2F
6W+jm6RnaD33hXJ1tk03FflfVA/CvE7R8vbkPa2JWsl6PwpeThsYyHH+4b4R0cKl48zspCPlGgay
WM04r7X21l+JTM7KodKEQBeMjSbM9nrP0yuTfEKKdOOBIASh0sC9f1tgd9oC4vOA74Nua0fM4VD7
NG9RLzNuhItsGgJ0IxoRnDILGGeiyi2n1IRwgAT8uTvE9L8ZGxF4zW5dhgIrmFGVhH8QrP4Egtuu
ZtSCisXjmyU1GzjZevjlGAJBsKWIjmeX0PgfKatROX4DU5bIdkud1p2ax/iYIcQCztoP7/7Uhzb/
Qb3e9joydrv/Y5mKipenNUpvsy2050j3+uEsszycswIkKcDNKu1Qoqhg6hZ5ct5Z7RkST1l1CCUl
XS9IFVJwBbVMF7FzdS4mpf6M+XmgAjtjRn66ohMWT2cBcHG0/033xMPRIH5gk6P7eVZ+iuvEmHqz
gNIOFse45YexGZWRJwUvsQ5m7nmRLnJG9KsfDImQGbJDe5/MF85XO0XBp6L1rJTIVEET23gy4SvB
K+GtOTSlr48vI1WJT4e8cC6u9U2Mv2fOhBzdMWj2v06rAO8ho9BWPBEY+/oDk0iFdJlwS9FbHqGF
ebf2L+VmY5G6HH3sraKBv8P09UtORC79XcNjZWm4XkGoSQQx/TFlk2wZE0rzyPV5blh8T6MnRC2a
XG9iSEzT8rFaknTBnHaaPyMbX+D5vmjXRw8OLFsZrVSltaP75XVwaJgl3vRNqFpXarI4yJdTIDKM
wjzz2kAWcTzCi8YHEZ5caZQnkcbT88qY8NYBfSWTKZEYEV7D9G0SdKzhHuz8zy5t94YSQdnNC1Uz
oojKiFtGnny5uHkx0dy7pHYE8Otf5GweL1h0P68VfAnvAhoad0z87ILXFzxhuLk54PmaYlgP9bcF
DOe1rOkz0c12Dp3jnOQI3JIJnb7EDT1fK91tCkccKGMFgVgKnoBj4lcpdPcWub5zwzmYGTntdyNF
nA+68FcXr67g20swDPsaf2B6e+QfOIq6oSzq098lMCyFqiVLWKy/l6OP8w/e0GUr0Hz5R7HwFgPS
qKNlrJgqC9QMc0xJxC+tLRXKrLUjVLT0suAXIEBPGgqAja0MieA1pJ5/xHsOrBZwtSlGK3BW3TjE
XWf4q27ygsX4O8HEeRgPl+SSbzKnBzJeEWYN29+qqcFZYTmJU96g8K/jI22K8vk31O3FuHJj8H0C
Jv3XciS71+BNiaZ6BJPlPv2v1DmzKBFl0rAprD1YYTMn7v1gqqRIgbpIRvAvDux7cwhRiHqwEEI4
6ALDbWDUzMXYyDJWM6sgRE/94FKoqFsINMv17Mxh7D8Jda0G2ZsK9g0y1OwjdM6vsHhWdyzR1OiW
F7fgPnvFdPTglsL7C6xOAMegfKX1KIFOV+O1qEVa1uE07hC2AnWbqUQZcL6//m5yFhCAXFnpb8Z5
lRddSpsNcujwXAgAXjjL9zKz84SaDwZ2GFz7PrroqmIwbNlJZfy+fYSb1N45vlFOPvkmK8qt2Lr3
JV7vzksDD04WEJWt5EZN1TDJ5wfAv0XEC2vIeZZcQU6UueSBTPOGszdTsepXH1ibnemeKvRxXXV1
ZyUXyILF6WZUZUzOU8rpK3a7Jug0RNQQcDb6v3GEwcG7DJiqhkeA2Oc7wQ2RJYYlnO6U9c5RIMUb
N+32XBz5j2OhR7SDgZU3Zx5RZoL2vbDaySVzSVjKekCeeGBqvSsBfuzUxWHiy+jVyYSMCGIzz+ox
qV+vmtbYnJ/F2cfTXM7jx0iA1x37lSz0wX3vdtNNtZaWOrEo+xxGyzBXl/THNPeewqb3n7HDzAqg
Cm5zf3WiF0VeraPjSJxjq2jSKONfgVeWG9KdOsipxzZWUtLuVZ353JMCgL7+vrS141AbcTqeD20f
apvFxFAWQog6NInbFcHwOcXLN+C6Syqicops+uBgR/TPiSSupE/UBxFAsOGQPyeac1IIW9ZcWaSr
FTb7nuhjgP3E8fPvHOE9Sko0Q1Tu1ssig0dbJ6nLrwTgOYRz8gsMBUBFS/+HU7SQXBnD26LtTJhS
D2hilB2N6YsYpRfqK790Ugj4cilBGv0wKoN0sAf1Kq52zixH7IrEsc8K28bKyvb58G9Ckckf7eU4
qUHcsk3nWFzoDMwel9eXkEz3tTG1A1cCSTdhO0ibUWdynX82XeGNWCyeBnnGZjUwwZgj85gNwGka
ErAiKFN+P/uZeEAIwcBzrA++tSf6ey466GEW2qndCRqkSN2R2FbQnZpKHx+LMofEy0PxRZw5ls01
dlNW3CaNQnTtoCtvgiEQ/qcp9qrVgvHKuRgKmDw2E5hdSoFEscczW+6BIXBoSc8Xpp6LXtsiBFxK
IzkHd6jHHXswnF4L7P7ytFkcPPBjIuRWlxn072v15zEGfSH5R4914apopHqz/IU3X4zeDFmCmewF
ib3spLymD0ZtkZlUxcrmIISsgYrTjMwELkJ9KVWSkYUUJsUQsDYhTK0L9HJFJdNmm4UxlgpYqUfv
fxJpK+eJ81xwiVA63MRhENavdVfdi2ifdWKsXohZhVpZOA/V30UwIOtAk/upAcKYMwA7iX+3PjTv
td8PUhleqmRiqwd7UxbzhPLjRXZjNEm5d+4V4f209mYvXoTcBWbnt0IqyI76CY6fgm4c2KJjnIJ2
UKarh8DqYQF7Hq93JX/hi8nDTx723uM4PIPzpMGCg5Z0VOS3P462s0/mWZ0pZ4o7r3lloFe/VtvW
ApiPRqEy3A3KMLNLRhoNXjMAQLrQkexzAU8MlQHZ168cW3/c7VnGDuQbFx+x/GUe5YiBGjBzjXlu
j/X/MyOA0ithaEOqz5BGPCelx29eqHDdAICqAdHwr73ld+Csi6dF91tSPRbFaJl4c102UuWFOwNv
SJADYB9/7KB5YCOVyvHoTtDkV40ESEQwhuSn6oLBvxpI/C+4bJmuqiDnfPS2oUm56WPuwfJS6czB
DXcuQXBQ5WebVgJFYP+qyj2kihwpv8Ilo6m52wswd/Qg1h9HZ0tgn75vFxMJKGrVFoq5rjNe8RkP
U9ND2GAsvsm0MRnNMXmwKxKAj1G8IK7vgb56nX06MvD6xQffmOS2yhPxC3eEt80608Cy8GUclVSy
1WZ38+1zKakTgQ5wftPx3DsRJ69uufAsmdqR/Z7VQaBBbYeybn7qvtqRp2l19pwIw2fyxjZwjX1f
A0jESlnr2TwG682pazBtOJbj3s3KNYCKc/BZNmJILx2V3o88E+h2QaFeDXI5dMZLr7/Nop5HM8s0
tdQ+FBaqSOA/1TuUN34cHqppUGM5YB27mTckBRWfmECXruBXNnpcl9P4Z3I10NNG2fTptNscPNTa
emRJ/uurckwPJyAuDnUgr8A9c5wKS99PmmmZQX1mSDsCF8qFKEbX878Ts04+S8/jKfc/6NoFjbky
hsg+bFindDyX4BE2JBLzr876PRR5OFysSrZL6GonOlyPPjo1/wmJ4RjRF/om3q0QLc2YLkINRx1T
sI2FMV6Hs3VTfBhEQDUzrUJLNeOUHd0IE9VBrb298A0ByntCxcV+bV0JxfUShN8aUFufKf7lZDp2
VGc/D2GG78etn8JDSI8rBZkG5VGBzMyvdQV/gBREUWyS3tKmRl2y/1TclUPcrWLDIlL2wyz+prXR
XaL4PMfpQsXR1vYROha8jQXg6NJbsPjdWQEGf189Wk6A7ufg2PPoQp+yyt9uTEjbB5BMYFDyqXH0
MdbjtVLoewZlqucU69xaFDqlyA/MaRRhFu/RK+k/kDACZRKGVCxhLA0A0LgWC/WBvNh4riX9g8HV
OVoZe80dt8h9+h2u28PGLYo9AgwHHcuCDEIkoS3Y4nP9IcGdoEqowXOL61A2DD9f9fUHoQHVfBUm
aDXbmuEXZQ5jbAnb5hM3KKxWpjKu7B6vxanYyvQEjQa1oQCgCrfHENnDHnchVPM7SCo5ItMjUntV
SOoeuJkqsmI6xYbBgqpdarOO+nX0K4iXW1U/5u4yhnt7pdIpfKux/gKmOYJkQW0z8qZNsycN3Mf8
YlyyraPrPf35wW7FW5gUiVCipzTUNlGxkzT9VrS5Elj/U5vFEWIUjJ6SMCLahUaHGpPKby+FpfBi
qwskyykAaYDF62O5MQFDs8mKcBJEc1SirZ1CqWoX8rs8yuFTkJv7R/2d0eKGbgNBbq5LMIl4CSzF
3BsEWgWsKlZdtTjHtW2+rguHm4q+Hos4djs7NdIKgqeKYKka9jx7ZOaf8F8bF6UCchDrKvb5GPQ7
0j7RsS5QQ/6gfDLlcObOaamMBbrjpqic5WlaJUO9C50iRpuQDHwlQseVy+zT2QGl0v3P/X5k3TG5
OGAR3bk8h6tIJ5Fzm82tDT6XS6HLDCZRrKzSgJg2B82EH8W5TXfvA2q8ZW3ssaqsvEfsT8jB4ZqB
0imggL+02OTpkKv00ksiuohKEf4rKarWiFRGzDgwGGmu54UCIFtIvioBViT4bkSFtFPEyb9Ehyt/
Bdwqqfjxej936Q6WVzn2j05ecEmi+OEYlDVMU2xPG45PLdN7Av46Kt2jaKRAHMhfoKyNE2pe3UsB
qYmHekkSKXoHZJvl8JOUrZKN6d+JawrTOX3YwKCxZM7Tz9F3FwspoqnWPBpfj4recKLs9vvVrrIA
HnizmtuNDr0DVR0k1Tu7PIqAvEBXUIVJ2jEkRTd7ulWWrJWWC6i7/dCr6E39AFy5JIbR2OuuCEZA
e57l1VyYSm4YOZFss8+FIcR9QGG/ptSR3nsxfQTxH+9nyRqEwE1TztxczXPv8vnzTUn/8QfK2s8Y
EDJ4XrdgzBVLCf8OFu9LEvqVOxLoHP/78PCKRfh5QlYYJ5f+1DrtZZR53Cb4nmtyIm+WQUJiT5Tm
qBRTZjO0jpi+D+W0Na77iSUUETuA2maPEdiitRK58G0vWTfLp7KzgxTjE/zjS2WuxQCaDQJuKvsV
vTbHNTfiWYXx/XDZHT8mwocKVEcbmYZWAVNwEubWEAUQWbhncGvMtGNzVAlvdDH3go7CD8QOzuYC
fLdEtMstLmjDtcyNuXF0ZPjbkBwX015bXkl+ZOwNRONmM9ox8IMppqxZOunUMuQatze+3aHNFH5i
tb+Xl2653Q5/r6+nqT/ipc8gPXbjXLkRWeW1plIIBabjPnWRRNPPL9Nt9iX4N/iuc8jcMa69n7Gs
Bmkp6cttaxnxlpAVk4lIlOJrV5jns8aczG2dZyKK22HbJjNAP6//jShL6ooE+VZ8kxn7K3h1eaW9
q/hWPFkbRjLD20i8J6F6qhsj8dn4S3NAr5+cr1ZzV/Dwzfrq419IQj+MN050wzBcsegv1M241kS9
H3ZAhUkNLLoykMLEMMxTUXa9OmP6MJojTk8L9mNFotKif3nEKMFNKuY9ohTKT61ZM2bHLxYe/kCu
MqfHFBgJTi5b0uULDz92hqI15MAcgmsPtTBxptDUKqSfUlMoxvyqs271QxHo2ANT/oBrZH4FPC9W
TEIufp7l+RdlPlDSo/pD5j4XUGnVF/wykrX2K8XQNIM0N146JBqyEu3LzRq4mkrhG1C5N+/sHFOZ
Xw5qNV5dLbKsLsBd5QEynzvo0ZzDDU1w4TYc4xUKY1VdzqJi8QVNK0bW/k7TNViRbBfikT8quIpn
QHIgYx31gkhfuAjB61odcwjx1LHOJVXAE+/DSPRzNa1LhGdChdjjkSuccGHbfbdExHU1EyNCpxyp
UzTgTYCE+DgibnMsVCzSGrsWj4uqcnDPjNNQUq+MPYAz5d2aDqQFCqcDxRxx/KkewQVbWk5tP5fi
0QYPafOL4Pv+N24xQHr9CCh6rsZmPgx28Y2f+bYV1FB8NH8f5AS8nbYKcTwBLG8P9lszwYw+tUsD
8i4M2Opk3JRpx6qZ1bzfk2eeM/x2sOBmd85e8p00yPKlK+GFEnb19wONN0wRoeFlvihR1oA3FTjD
j5vf9fXmA9fkSETq5vvdmm3NBD19jQ447Vyry8lLXiMoa3KVPZaxHdZXfxKO0qAEkUG0FGp9VK/p
iC3lQKnymjgjpqwBdeY5wX+YDV6JvKrsIRJfqJr3IOL4wcKKOyEGV4uvIgdDOZgJKWoOmxDGJhqU
XHjV7Hh/S9zOUjiTTLMMBU4NbIqk/BrGgfCtBjJjNg868sv9fBAwtHKa28TXPQBD8OTVrjtwX2U7
SRFBdWxVcucedF9Sr5vgyQM79VKdehTvv1ZkFbQP+RNL4zypvhSMawYZFppjRxq16h7OMLvx7hmb
Q+3o9uHVQMC3ry6B7Gh+srNttpJftjeu8OU5onIWFZgjoEO4qe8Pujb5HM9hRvMJjjcAZN4lbfrT
766+2VpC53CicyjGx0NHbV/q39idHykSBvKR0asBXVZnIdamRkXpUWzmTQBPyaTQ6D4yntEtZ0nc
LolPu/EpmekI/UrV9tbSbJqaE6+sJzunhrgItLe4ZqQEeXRkb8jsScuIO7bhlggWKvAfUE1L1815
fzK2P9sEMaPaOJYxheNqrufS/hyrzPKFyRewkb4R+JxjBbXk2Bj8IzYqX5AwaLuM2dQTnuE0KJtC
+1zyzt4msRzk18oSX6tlhj8QOu7MOqFh8leZvZv0jJtPiYsYcxwdYHZgHMwX00rXkfpqZzZ6q3eh
N9c3PLwH28apYhZNLS8oS3Ss6rSP2m9/sSlj87+urXi6OagqP+nFDxrtD8NsLZsqd8yGG76zWYqp
X2gbWu+M47IYBOUGs5hfb9GsPqAWRvaDZ1tlT2iwv/37dxBjgrTndmq0tSyQ2G/zAaTZ+44y5Nj/
mSyXPRBENCyBxD1tM7AjNdKCemUi8tV27/2cB/tkA9dVOo7hrlbSXsd4XYRlQdsc1Ew0BPTldPfT
CKm51/yuemUTEsxfGOe1jJAUAKYxlEIDeS3XTcsF+E2MjHDe235udWvjolOVHu6S10sxN8HcqiZP
LCP5VHatt8nE/1Q659BX5W/9YNBJAlCv4LIYlLGN24b1jHqiaFJ2uG47p0sG98ONqXVuY/JVQc4m
6edh6lP7ACY8duLlqyHJoDhns0eC6GsOnG/kfGq8oGmFB1ZladvderokyVjLUTmzsqp9bhofcJdW
4YPnqjHpIEYcy/wd+gphJXBuQphv11qbhJKK2lBqt61EQz6RPJwwC4Vp3NQFJc9dyj8dEJ2Z9tlK
v+/snEKmYo+AS+lSwdpjdASID7cje3f9yY/Q2J8Xo2wFmY257KdBIKdE+/6RAVPEtbsuCnb1Ok+z
voc050Ef9kFqDGcpDtsOGrzzS6oZE03RetTe1Orb9RscGaEzw9xdO2ZtJaS5olxnpfcMdOzcbqfM
55NhBaLfgo7PuAhILVy1TvBP2A0GUYGpzm5lrJn1+yJpjM2przcLAYVBHRv9xHSud8SIUzZdGWU4
aQhxmyI3SNF4w+owWZJIbMrtViLIqPK7BAYU7YxDIeEIOGEFMvGHCM7LsYgUfFYP/ulX1TML8Sxj
GD5Jno68G7p9TmkVaB6BBManLnTc6NELhafYa9wk0/+upyTxD2FXGxR8WFddid0LPrYwprrJto7J
nVc2iK1IMhL5Q8dZjX0eAM+iwQ0YP317R0phAr2k9Vg8NG4koIv1IYoZehBYgPJG32BLY6sOcRvb
HTmXjkHUjqHEvB20TNpNK3NtJWQmhsa5c3qhjT6DIYPeuTQX2UWgupR+LyL908ujXanDTaKWgjGJ
+j9mMaKopyOFbJG2IOH4f5SoTusRLIIPIbG7CuQfrfJUxXL4z5Za4LE33GCl/yWiPpkqGe3A3qGK
Cl5UkFLFaDDDYgIS11lAAJeGBnouH93LFA51XxcIy7W4pmghVf1GANgaXJCne/80bsZSJkKxxWuj
hO/jTgLXIb2gTBLgfyhV7wdw6SbbDCKPNJXDcQWSbzncLUFs9za8dZu/008NHlIeeMz5VCwoaW2i
gt9aJoO3Y9J5fe4+mBg5xUpmx2p/GJDY3lDUE6mrcXB8+8I9M0tNITxtsgltLGKvLiOFcw2+m4iW
S2I+9OvM7sVAslaL7AqM16IH4a6bPjz4aZpm6rHNu6TfHoZNMnFvsXVK3/bXTAlhDmeD84jxux5w
wKYQMz94cZRP6V/R8+PQkarWsNw3IfLFTWW0qTwSDu2ykYd8HtcYV9FHKcwlCrRMH7lhOsN/2YeR
REHZwurPIepLPi09B7soIadzdbSJ5PSupfD9/fBmQCdV8rJ+ztaDIhtBdg8I/gVvalZCXEy8d5/W
bcfEVAIkiaiH9Bo1zB9rPyhko+ZEDSISsxB645ldclmfpHWPhaglo3pPvK/Y1KXcgPtSwjRCgYOe
nhSt54F1fGTSwW22erZae7HXN+3evRi75gp/Stb2NijCx70eoirSIlRNS40LBnVi8BzyjU/TXkAn
R9MswLbgPSuZ6m9IkV/+DSZhZpwD9NaSVuBjPmQk39JipKiyRgBBB2LocCISgM/eHgQ016HQ0Pni
eFDsPTVGCo+8EarH3dwunV6l0Ms2moAwQTN+ovHcAd3XcqPHYkFbB7XSG0e+X67L3lDLwRsQMzFp
96A+/ouYSaplFKjlCZMRecLROHPpb8GA6ZHe2ZD7IjRsHq5xv6Kus5N66xckQpZlPKgfFpgZe+pA
cb9ZXXrO/zxRSHu48qbmhwqNOe/cymDA+34mQbAEtr6LrTzDrEIWPoFozO3CHLsfVgUtdMDnxWDN
OOeVBofDUhjo0T8f2DiUPzLSjGBySuBjK37ouBVmAWae7+sEKa5eTfzjMZ/eNjpxlvSvNktpywAZ
L9DhyYpTiOQL0yF1rkM5irK4Y0fyyDGcdoddFZkr7GdIUHHBCDt4zhNWPKxERTPBskqqWTFYB6uv
ZBNrpYaCwpmVJTBXoypNHJIZgnjLxl4qcvAH+sIFtWAbzpv0gshvdp0j7PtTNozk2DhJERjL2UVX
4/22epDE+hW6CTMATfkRyyGCRscyq5yBmlEj1BCafchhjvqZtfMPUHrDB4kbMs7q8w4fqu8zWWIG
ac2gbXiVrItUbcd7Sg9Al9aicZZfkrJLgZTttx1ZuiOK3OmMmQnrL+QA2MQrj0s3E2YpicaEuIQW
uFcAqsOSniu5lnIRgQiqd8lfYj8fN8ZvcB62rGL17rGAADgirQxUUBAK1DcCMcNNrJezCgTKhjYU
wwCiUgL9/Q4+DNAMPkYZeIgk5MyavFz8mThPOmyMp1R9A3jEtpxTFN/T5HTGnFD3rGqGVPHxiJ+q
E6Yt3cGSdw5zWWLzna+IdI+RT7O4sEoHDT48e/AYz4eiqtVlT4edwih5aw2b6CAdpVi/OqkZkrwT
GUzCgjLZVTx16Y6my6D2Qo4Oc+3SYGbiC+yK44G43NTXEwhay9BmQwVAdz2vF1H8+WTc2UiOnP5g
hiyeXn0fUEhly5EGZNEnwJW+5SlKFbwiVYGRGtCKwsjHsVNxi9aabzVbGKIa9QUt8r1hsMQfMt5Q
d4yn0VsUVeG7jhF2LF94Aq50yutYEAYjDfiJfLJEMF19woU8jVkyWb3KdGh2oCA/l0868MafFVUC
KHZlsKbNq1XEuebfZICUXcKE1yUzKjgrx1aexo8M5u0motQCLne4ytBuV7Ne4zAbtOgHsrZER11R
JnjfDePm2T0EO/KMZz4fsxv8HAllgm0n9PsQV/39pr6dadM/v4FGbjsB4q7gwa8br1O4oJugR1wh
/SwaZI5+k5rxy6dN3UxD+MITyeu0kRlD+NBv0E5gtfZLvmdfHcSi+N1pvHgtH6YKvGK+22uKRb0u
zB9C4O+bq2XTAzXHuU3gXnhOU2lAJQz++CkPCHq72oiSmbm/laoEzbbp6BQ2ej0kiR1mduAwwZTc
OWjGkXtFYnOSloTGJXr0vVnelFJciRT91U2+wF+n1f6BThgMQHnzxMyoimxGhpYnta8WjzowO3CX
lKH8xumOoDbvi+vcy94T2r5tZKyxeaHPzr842NDRJUVlqU0mlh5gik9o2qP9hjmOEI3rMNnf/NB+
dp4IdQwR9YfUpkkKCMiqcBLWs1W56VR0rErfirCAoSkQSgClXXUya1mQdr4UW1ZFnU5rO+X0xcej
FW+VXshImay0rIybgusMV5cu0+PTdcurUxsitWJXpESI1t9BPz5bfOV+iLzrW6xGRQ1MpIbD/D0j
p45/7Pb1GP+JtbEtgJhO6vvaAJs2XQZX9NP8xgbmMoENy/3xCkFYdXPDTyXF9LwjDWdDUUn3b/fR
thKXESTUraBVp2JQJTZlVx2tFCB/2UUX5EqjC9MMjeb0aq3dTLUmYUvbD5FE9kiiozdXBdmfteXh
uGxuAsvfZhizJpy3MdUrJyVBNwmxMyNP/+0THznnklxlOtfiHl16Ar2TyZgpVRm3X05JsaVr2ilj
B099eUMU+3Tu1Y/dIBcB7H0p7Ezw3UojdvktWZmp9Xn7xWzgCMH0NKSIeh2dUxUd2l1UUXp+fnFk
l2qNAUzBp8+Bu6fUO7vOqmNCKHwZ8aYbImywtHnzrvJ9S5jQWJmbymRvca5XozkrAg6QFib3Ogy3
XtMN5pxN7LwkrdgvgGNFpnlfxGgpcqbdFL7pDhT/mVQ6pgeir1iV6RV34PrLLpjo8B6nBLoJ+n1b
gJIQ9o4UHF9rDMbdugpvpv/1e0UoifOaqxmsrnOOGxKYKTkoINke6BsPnnjhLQ2L9f6taeh1mHFZ
vFZMKsWa40yQJN+2WmCaeL16m+MuDb/gPwh6cMJkVqUdxceqvIt7QLjtuH0ncvQ0ZVGLODCr33HR
uUYBjgPj3y0z+gCJE2oKSkJkPpaEtQdjk47DXJiyBN7FWqsxvqQr5QiYxOBJiW4nH9mNUvDxsjC+
cQJ6ocf1WX5GlCwoLHb0K5bO1gb97KeXHdNDXNa/ZkcXEtQp5z4o1Uf8TxbFTgRDWCl/OaccLKok
ABAT+atFK4ln3/xivziNuY0LseCcj+mKv0Zf15J66MegyiVUkgW0UyauKPo8MrEJaUfjNAyZNJGJ
ZCKg3vA17bw0Qk8q7yfFdZGuymdBnqSIMCZPbR3P4ypXkYLSs8YzzF1CJrruTkhu/7ffKomGqq1f
RNuXblOxtsPnl2Z4Ke6L/O+4WgczcrfJqIYh3ilqhFDxefFSahvb07Jgt62KfX69pwSEw/SBxHz0
3bknlzWRu0zRiepAc76nblJfTHDMuQKQJxLcQ7Ikg/jJACaHoLStCFidtfPCMLbrzwqM22Lnf8Dc
PAOkRBoIP4uXSsGfh0wbHRAxJdGfEzdhBaAp25STqp2jx6+wiB5lOelSRK5DnTsG58vg5CCKI4TH
mqVixORMwG8xSLERRWCW8LrclJfgjRlq40l23wlxWc2sVRnF7K0MI4Rev1hnSxaNNYto73Ka8iar
AaAUZGAPJ153Y9lWpe89sxxUFGf3FhQeWwLHWQgGImkfOCNdUUzptX9W5SSt2sN6/dh7jn30WlNB
yzg55pbqn9qQzyXhf1hBaDm+1KYi+obAD0KgiiZJhue1DDxvoappTBT45ujvwELDaMx95fSnWXN0
itWtvcKd1dn0PGspJwhHVoc+Uq0WDP4OXAVO+L4qV4LWtG8FU7FWELSYZA++U5zbOWZvsqIipNPm
0AggzbLcvO4xFy55+FqFyAvh0ehylHD3TOWvL6ngnxUdmrnJCoYkNEIBUgv0LqW0GEO1FNPk0zu4
4jEhwT53Pfrow0EnYQ2VOjWlKjTFAAbTn2DYagTJWurLL10E/qcXnSUve7XNShmtO7s3XepcGu9F
Kt8ykVAEj6DL1VepsyOQLChr1yIgSHoIOhdQvCKRZycRZlCYoI4FPXBuz85WnFENnb+SAYJBwdYY
Tx4pqH58veY+r6KF9F0iyWgw7YifwGt/24edu6KnMDtM1cu14yfypiA8kWUtzoLOkHD2Y/u8P6YX
XFEd14JKvZTDV9NY0+zNhH6mIS+O5YnfD1fagxWYi45ZndcJjGhWmWhjfFVDjFqTiYp/Vjm5L9Ve
1iQaORB6JL79BgvHEYxSdFFIvVESrGYv7NtKkMLssUM0oZMVwBn3mfwVJkn0ztlMG16l+0ELGm9e
/mZBWRWriziAl9SpY8nNO9RlrZbmkdfWdB6URTRHsS/eIrSQF01jMUZCk1JMyhbH+TwAwRepnOvR
/cyWydfTniz8tVOEEJ04to7c7XhMFTcVKF1refONrjpUl3jRTL+VwBq+pZKnVufGemf5ObMnS1AP
2UvJ+Ad6OHeZn8wQDxBQzneY2Kdb8vWgI4FDEODLbanTKlUBHDS+witY3fbEYuGQWMpT5gmjXZpC
TpSFUab93FDz731yrPFp+gIC8NkHFk5MmydJy2giCPegEvfPdXwyRFIx4cvCWbks/zI8UGfGc6W5
0a5iGcldiDB1AT6Gf6xyvW9BaYB9f/cUYW9jXYlUDLYKDgxkm6EN/XvP2ZZ3IVbHDjynrvi2MIsp
eqbfC8Hzc9g00fTjhL5PUua43fG12jDd4UdrO4gr0XWL1+qLfqiHRoWdUsiNIo292ku9gh/MarKQ
iv5D8TfnQQA9gZvDzCPn3AC7NqYMePGi3SoWmMvXXiETmVFTPrWk0TPOWn6sCMO6qjX0cfS1JTp7
ootmTQbjvNPngbRXbwoieel11fKrKHHZaOlweKw6Jj0kXNmyQmr0mFtPCMJfZ23KYiLFi72U8IPj
Mm6Tx9UYErEd8mKOD7prpA1dokzZlyaS3xwvgbNsv3F1m1JsDXCeVaCdIsil4BIHd01/WCbXIEMy
/ttJJ1wCYGGjoWyGTKm2/UzXpb3Sx+mfy+R1EIJGOsCCawVM0BhcdpheosCJMIVRWl/jY1Id1q3n
RqsCV2IJbqNR2noPeD0Grx7ZC3U2RlcgZIVLDTTVKBtuPUgtD8bsPXnmyKya2sPHEVfoQPpeuf/J
D7Lxi9ehwCCiHIo0+JJEe9bAKsGIvlkF+Xv5BHQp1gMoIKs8TCgEuCEs6HVCyCWAykEITx167lnG
0FwLqaa3pWFE0Up3KozVpF19wBBDuxPSk6s8/eY51u3A+8/7wErW860u8WRPD3+0WGZyYn2oyRnQ
Kq4ISpQDVIq4aNCn75W/Ig+Y3c/gnXTTV9i2BAqxet/U6+Tb///iqxauWNPh1+FtpdZeyn53VIaz
4FttXVUBKpEof0oOxDDs1HE6l6CMMZnbsRzfA9Bi9iP6ENsMkbVNAQHJ4jTHCqIkfrOyKXONCgXK
y+gmUXHitOLYcQRgneKyYN7u7YKYu2zdqbj8EiC/xz8Gizp0WvgL9xPACT8w1tsJfcI9iy7z9JnG
bQEQcnu79Yc5G4zqjKYzUf+KXLymgtrN0+lL0HDcJjBjVGxeJAe/QYtsBwL2vEnHeF+jCyX70U/N
eNcI55ksLHk5vrfo+5CgP0mH9mLaBVJfsrUTqx0IjhIIFA2QworjhmZ97URzE5agSHYjY7ulfGMp
h8OpI8Xivi4GATztB2Q8hBzDNHI1o8zG+uLsiDx0JXoxFkN7f3cdWAiBXbOlejaA7yrVUNspGUnj
S7l85QYvD+yxwWCEUp2r6zVjmLvoh51HcRuoGorFoDlwUqSDcSKi/4z/9TAMWgCDdz4Uarv6rB9H
ZqqASEyxAN4f6GCvQSmKlJMDoTZNNCdp2NmXF2sfV/e33qjskF48bUmwPuk1Aism2nczuIeZmdFw
Iyqkyks+mYUCZurovqcDE/wxgfL5sm5dCXc+IgQrAkZ4Ocl7gVp1eO3Qkb9MLVyxm1I8ZbFbNIk+
5qXkG8oJgfj/c22L0eKH61RAFDnYGCssPv+DYmqSZ9ASePbx9GnDah+IUa1GLLYSGjOXDuZrdUj1
23X6LGD3z573SjnBiXZwMDxeFhp11KM4nVaTjpniYtLVFnvCta5eMruZRM1cTqw14syRyzk4RozK
6e97YiqfOiEEaxaT63+M5uRi9/eHI3+4xoQnXpoGT+2BLX2Nx7MCExRtgjOn6eUxAx7WluzRNOpW
5569NiYKRC0eLWUkXKKadYZeUkPKH08Frlph7s+G284QtQpkzeSqztPNkDmmSXPZB12X40lQHNgk
Tb5OXflURbUx4M9C2FSWSbtIgx1LhqY4NZNenpP4h6+w1vPUNCSMCUDH1BEVVZPuOfMJDENcZnVG
n2wliR68QlT0yxxTvHGRpcXhu8HwHXfvjBWuRoBO6IctOcmg0mEviBAqG+oJ7aAhx5iX4gT0jTED
gDmbdLukjApXQ0EmTHU1AgTszLT2ANMdo3I/UqMUBSuAkbYwzLunHjKYxbdIqujM9KrxUy6rP9qX
vGbcqKCi6G7xgtrnDgcBf4q7uiBvu3ee7SnKNU8o3ofXT1UeLq1w8EfL7TUdG/5VifxpqiI5XtzY
Td+yB5EHyVV2QZw1/DA0pxO+RN4dBlN3eY1wLUNygt0hs3oT3ALg8CXiI+T8jlxiW9jYoFclGiFK
s1ipyooQo6aPnphXh309B/UexWfVEVd9zuW8u6toIg+AbpigTmRKpzhM7LP2bTAnlrvZsvm3Qj2N
ppiurr4W38+waS1z2PoRe1XXBcmvt8vtIPRv9t3MFcik2q87dsiAlFjLIMWQTpvOhkurP38lI6Dx
2djzJNqIBV0b3xEcWjn4MPyDvWWkWawHGx0Wht2Jsl+zaDJM8BU6iImwRwF7RgDEibg7v6yXIFMR
iR62Y0bCf/zxF+yw+VqBmzj5y5WnDO+S2osS9nJkKR4x8yHlP6ynOf3wfFvSCXD4ktx5pn7rWLui
jyhEzFo0uV0dx0ps+1a1tCiYGW6s+U5hCbhZvOi/MwQTmSlUQLAYgpQxT4VYPA5UOI0Jxm4N/Riz
vnBXqgs7zckBhQuB32GRU9GnKl6qB9tIZDFVjZ5yF7+EX3C9ct02bVtW3fnjKg5IYQ5/oKjfl3Oj
1rTsVd4QhQcWm+g2WVS8MkD5MQXAECq89ZY9QVyc4r0g2Y33rIEOGwjFNUhSV1GEYOJoEJQm5bci
ynEWwxpNF0K2RSp4cpiLz3ApYCPKZ2hCHlzYNk+z788FSCh0tY9KvC4eXqVCcPIW3wzQHg9ED+qu
YhHzkGnAIAwqHmPtcfJH/oNDUoQkfzjkBWs+LDYms7SJI7oL565jfcI215LMfgyIFA9J1Y29uM5r
OWQHWBWusTYwTG9Oe4t2W/JwBZ3mRQtLdDCNK/m2yDwu+dyxSDg9pNlHP7QeRNHh8Ti/CbzvilBP
jdjjn/Pxr+lLZqtR0zTqZva7XdDaNRqoof6/SyXQbjyHePFiQEdEv78ZM+s0FHOdVz95OG4R0XYe
2AS96QS1D+6P3IQ5nR93xcLzJr2u4RIskewIQ8/hrDmnMMQ09X4NXB72h9IwcbjS2pK0zHP37X6W
K3bHWR4gW41C/y5HW5mplB6jt5bMimjaQXhippodfEao7/cFQpwEeGcSaoZobGRTzfGebhMZ+cwy
uu4o69Mf8mo5AD7tRoa2ar6gNiu7WiTZlKv3lN4Ot1jh8xEadhS4780YYCd+57/GoD+8AlOi4r5f
QnmT+JDJbbGkQo66htG5cEYAB8X031zYF8gSHs7F/bglBR9bK2VeLUnpzX6qQfcN7smeJrqGZT1r
Up6fTtnetadi6qTLPooW9yM3byvImNtI2acmP7Dti8ftoZroRkfoNFzP0rgEmr0OVjO/3wajedap
UXk0RaNDRCVpAdvhplGkIKfYN5Ikm2KbvV4HLmIhzoX0tQXah/VLt5cA0L4WHpSFvkG8M/EBzeh4
+TGBqp4ZvhRF2p/t4n/M/cFiUoc3pIsu3sO0wIjQfRjwEtTnaXe06xnD14Ex/Du0HBCWH6Vv1jUk
823xIDu14T5F49DKWKdG4f9on+Ag19h+YeqsaeeJfdO8oghpJvGzWr8xEUk9IiJaI0LqLYxD+IFh
UmxILT01L7ScUKLF52OR3aGZ+W5U3zh1bPukQZJ3XNtWPaQgW0UFfajyWbUN3kcUikSUjDORH17J
KNl2vS42mG492DB4Z4rOkWywzHQZxh0CZKzgbijwCsCYqaX0GncRhnc0v9u+eG1oD+NsabzUdREG
6ot54U9Xj1x8prIrs1vxYd32NO2gYYaGFhgR6ZtLPE704dkkqeFpjEJ5eWYZTq3ObSl8cL3L6qyy
X3b1kEQ0BHdEwfTPrz6o4pMbBuVhfuIuuPk0LaXKSjCREQaou4Jw3iuh7HkflD16JHefdxHzB/0X
Uj5dwAtJKcyuZOmNHdyGsoHV4ZN4CmonsR2/BlhMzajO+VM3NmU2huM6fBa2bA6vX5fdQPRqbkqO
NZ26HfByCflAEAiEa+rAyA3k0EkEnyERmKVIa/J8+zGYGpul5QbODgH3FwzbqMsxN4HIZ18yXqS9
OTfLY6IjSix7w2eTXA2QQwkod2bhx0rkPUZZANSM0fTzP3TZx0+JbdDuABLc3GkolL0wBC9jmqXy
q+I8tS0Esx2fKKuewgk5rLE9ed8d/I4aepVgKcPqLdRou4xWFURmK2RZ2KVbo/9RteaFTiy9ze6l
QNJLO6owWi5f5oG9Ff7bj72EXhL3IaU93C7KDPHX0v3a6F87A6yLzAUOZjV85qKXZZO66bHutykx
1JL1V8Ih8Gid3H2JAdvXrHaUsuZwc1ouA/USBd9VXRKtfNcyi0udiMYeYL5ncQDd7WWxk9chk6Py
1s3YhtRpg/bkLvHIJebDPLSKYqV2joH268JKnkd1DCrgQfQImlpXYVfdpggJd8yxxREm20Sw7Q7M
AarqdLY1LMDVfXYG/npKKKzAezQwBoJ9EV9KKKCX1e7CssrdvHW2RKzPSpfNnv/cUhMibkL2VG3O
kWQYCrmajcJjkvNM0Y2IteBXhMsIc0K8+0PcC8nUqFr5oUECpUNpA/t1H8kgccKpTCjmcnbVGQ5H
+yu3r9LHQbTvxgIGr7mNXxl/pSkq2D0K8fRliztiW/lqxwa93GME01y+eMCznRMCfrVR80+EGKBS
hHgwTFJVaA/vZ1LEh3bq8lFJboWzyEDKVqS40cNU4JT+njiqrrJSsy8R5etgF4T+uxLcnXME/tyG
RmCbKGDZR1dbV976AU+BkbvZsurhQZE8cMSr+CuzlKASwSXqpdMAuSLiLCsUkziOqgdSQW63pi8+
OLidMRYZURU1l8QsWIVb9QqaHkZtFRf+ckB0MbVYnDuuIoJXlb1ykAXWdatLQRS9SyT3sRqCjOU3
D92cYJFbg3F08MwYT2QAdl5z7AMJgjCUk3Ut8y9HCIhcvNr3jqTgJ7cG0WudfqaRNXHUaOCS84xC
gL7SDLB7oCYmnYH8hosQ1K119rtQ1vpXgUbvKC+Hy+QEdYokaPqUMnLyQIkyW+x+HTt8oioDFe9e
iYSC7JsMwhoSv81t8xIwNuHFpZoxvgk5CVL7eoTuEYzmK2t3SvEHdyb3R50IHAsTdiFmz0hL9UXn
zynmGrMVUUSZGH2eDXhnwCi2ouqjs+VdHTCXSSVdspVzZ/klSEVZuzYwIpAjJJ6tceDU0YXvIZ3Q
5sJBilCECAPlmsCUfQtlgWwqb3bFriaThagHeRJIHv8zZ12JbLpTCr4klD//xZHfaEa2g4fe5c3X
UA1M/uPVovxt+WGh04hjzwkviCYNOdS0SR7vsU/VHz8b/1VRnqxrjlJinQ/4Vc0iXOP3C00J/VQt
iCDTrmybgbHw5BJRQGrlWrmkYNgWZrqvaPICyCBxUmr6CvaFkv9rG2mGT3ZjYDQAof3kPVSrZs/a
rAfGp7BvleRUjXnGb9YuILBY5zfuteoZK7rtfVFE82KWBw71PDOdSmDhsHp8uDFViuNgW8YPfWBY
J5V/TxVwsI2/0VvwkDNvX3MarEK6psMw2zDuReHEwhqKezZIQ5BYTgJPZJdRIte74SZvcCJbezMk
H81o1c0VB5siPmaQGMKujeG7hBtXqO//4aYiNI0nrM4yg6wckT64D6HT6CDEVDc/TrphrZ0+zMzc
RaPi3mOmG3HRnrV0JM45uIDhHoN62Vnou7R7GoCiY3lMsMyqqbzAgOd5VOGYAIdzbU80FmyHds2b
1tECpE0BES2Dhg82AeHfeun6mCdPMf6seu/g63vI5laRwbRJHgTwdhuXrpcagnUEnTVFmdyF9zbG
upi36BySH69eildlwYmCugWt6hHQC1g3v/a/MakgEqUJBlESdyE6hiGlz0yxhjwBteNzPYDu6lr+
o/59QxRnZ+SubjqR9fTjf99XzeZX5KdnvQdYzKgTXwEiNe1GP7rlkV3XL1KCoZHPNA7YsqTPOGbD
mVmjo7Mi+ZccTKLJIR5bwlFeU2W/PriDsMMmDBOOHC5HRHuexFXBHbkt7Rqg4Xp1XPnppBgW5o0Q
dR7tD9VGFZ6vfeflg9aUk31onYtpnIhqgkPJlbhyqLKyKMiyv6gwOXSOCYAY9jgNgTi4e7sDdy/i
ytHDrVZSONH0Sa1VIIDfhwG0BpJ/dZF5kZp+sTotrOkjp66Cb66dSpjbUh+2pIvQqNxrL2mgTXXd
mb8L/hqQ1sUKAQERmL6vh3SYujdr01gsWrHY4Dh39EoZNxr5Codkouo7oYQ4i69X17jRi9JOCn8A
mYVupqy261YJmEhgTtmwVGhttv2oUBZJe3Rpko5uM/QmpbYr/jtS2sFVHJSDSalN9fZiMrsPImeL
UN6VT7gp6eWddqozRw/icv5UJFzqfeycxy3FQXioWJWylG00t3/7J7sxq9m+KiAcEqVzh6H85VBE
HNjXp01b0HNsoWVAshvy8/IXbF0y++RcduYIPI3hUr41cOpKzXJN9Z0oQ4gvVxJvuLyDj4TPfKrc
+ZTkIS5XumZSk+vdg24rm4R8fll+5+SJSh3oXczljVECC0e5gyMLIvRYetjtPpd1AwOW+kwMF8cf
YO3WR2s99gTiWa0lcivPaciHVh1DHLm5QY9RYjcXzk0ke5aacsEKF0Ug1Dba+OIYrf36MDK5MJuT
yG+oH/hS0i61TjUcirlsgL3CXDMImqkxUd0v59F7Igp9Shl36oEQLFLKiYVFI0nJrbbVFJJal/ti
NjqMxkCsYxF3O1rAdjy1nG1eEvcsVzA1fnwU/7vwUKUFlm4Cbb/sz0KbFkcpiNM1uMfibaoQ2Uk8
sK3RGmwveuZ1+xlfZy9D2UsqDZtr6DD648GZFN+PghEkjkASaKpvGK47q3/gRvkVse839V3D6r3B
2t9A9tjgfrYCBaUzRsnp3LtqJ7jKgDlBpeZOWjDWExTA5QTS/6lGhKbnADOPcyCob6QLLbwU1TxN
xQqmN9YNcJElbnfWpHeCU+npzgk0T0zrQJGTPWgBA6X+yB9/x41b74WI3DqfugGxaLAQeGEb5dIM
a9gW4HVKZ6ZiuPgXUS4CCkwzalhjZQgh0i5ldGjl69Jy7v9xokuOiHCds/g2RGNCZ+2JUoBJzv+r
cDsZBqNXNM3ZH8mZKK0EvtU72WrCZ2SXfZAcXmlMlysY4fC7v3YWqmQWCsU7FM0T8SVnRAm1tIC9
bI8Gv5IZU7QGxtM6KcI9XSHOgD+11P8H5aSNJ58qsWkJoHAA4FAJy/c4v28mt8jD6QrhYS669sN7
EkBCvqOnqOhyJEYDwXly7dIk4oDtudALl4HXxleku+7cNHc3SOMgDa2/mCOiWaPjv4J9ktdFSuAz
3V1/bav5/97QAv7Gs/RarvgxQAND5c9CUgNN+aQwlI4WwLfOwzRC+oF/7/9M3J+NsiCOkjdvoDW8
7AYQW5t3V0nZCPSL0J+grZlsh9AINOqJUFLMCrd1IIFt9ms6s4BOL1SFKMcjbtOJOJuUD/vUPzF+
ZiYmah+4QH3zdh9ws/LDBSGIyk9bX+1Hn2oJ76hGkP0iYVWJVgxpjJnOmYjhvLzY7s/rL6Sd2bo5
FpZl8KRiM6/p9VVhXTfIB6vYBjJJzl493SZJGn+gTVYHwB1U463unm3UE57QLNru+1nHXxPhmC5R
Oqu5vwcCsDNxTseH66eKtP5WyyYFpPVtBi4WzLMhui7NKobnaCT3RcuUfZ+mDAFh+a0OeB54YzPJ
QafshB9AaZZiohweQNUxCizVHhkgorzWwjH+cYzO8Y4aTrCnI/LYTQ+/S9eyUcypqh9mo9mKXLH8
A60k/JVLiuVnVvu9qkmYCrYr5mR0M6jr2RRJOkR7/NrkMqF/8LBdpZzjREjFwCD4aZQAJW3MZxFH
FaX5gj/9ZwPyFB5fmZ0kBdnFHk8QzFt/8pzlyLZAs8vFof66yzBicc5O15XAjSXDNys3VxEJTWT7
lGpqQbf8Hu8vosfrSA17hfc61aW0/JfHIlXOBXXzgvJqf1t9MCTH7cBK37uF+7tMULuDnIRSQwso
WriuGYbXOQr4wfHW+Oad7i5llawis6QaRzvRosQiYeohdXWRO8aY4cNgYjy8EflnwCm9nOSA8r49
ZNtfQnnq0MdalEO9eBcpCliuG9TS0SEutI+J9IA4cGiZDEsBmS+QcRASSfAdABTxgN/pcnUqeApV
yh15N1cERqUn2nZDaXSwNvNsgAu4jHTruYehm54Nl3KLdTU0YiMquTxINhY4Rb3JohBKUM6urgZU
qXPQheOMtyBzNshg4MoLSq4N+vskdZ0mLaUobsFwTeuHQdT8RzVJOoDHoit+LxefIrw974SGAcwq
PFUt6C9/mhyFuitOa73nattj2Ro9JoMeqwUeQ76kNCT96Gm3/TWUdYqqO6mrP2vIGjOumanFY/Yd
M7MDKmdwwqF40logt4NtgZcuLU6wOH/u87IhfXrW6r1aSAIVE+7b9PW4rWpDoCF4e5oTlTBRBnne
FGS2iQn/riVe1u2YcYW/S7b8KSq/kreNo4ugHy/V9TXKHyETEPMAAgGS5gTkX1oMSifkVUQr7jhU
WGUh5kWwt7HA1qEu0EvP+KYClEK38tjtMS21mSDB5z/PHpGPim/l2u/to30IIDrKFnnn87QcshL5
3eAzQTH86kUrU2KUP08t7GPDwK6ob7vDcdtT132HRgy+a90C/lXeRbwege3fg7w4hah6I1881feE
0/l13D4bCmqxIFn2Nm6jDdHxCXmFRiCsgZSconrzq7nvCUWAyLpv2+ZE3GNXd6IRinttdHac33z4
6yvXaumB+i9VhTCvVlpN2nYjcIsZVg+9WIzjsh7jrEmpW3xjDU788bdyWicvZk8zsxb0pt06aKqp
KpyNPOgIsgjOCajAtCoUEWw1N59gVSXIt7Iw0AnfStBvKwf2UdrZukXKNYhmEQ4WOmKNSY4jz1iG
qxUQep6aC1I7oNwXO85OvcSXtwKCBix84MYKIWQfwUYxuiJ8eek+TlZZwI2NKtuPM2MJ6cWbV/SZ
Ms8zqFipQGl278/UyasIiojA+j04yxkGx8Qj2d1JYvw6+b3z0w6jcVLlbDMibPowtzqaGXAFv5tR
afP+3T7Gc35HbF9lCORtv8+yBfgxIvqzAeJZSsovHuJaU3ItxtyaKcrLHYIjdiaQOUDqe1j49FJr
MDdPz21sjE4zxGcQf5lG5iKUPilcify/HQij14wUdDZi2JT5kF0Ymi9xf5rEyKsEqogVCDyPX1r3
bvT1BafQtDUjCcfDleAvOPMIsM40eYfGyJufqj7HC7w2/Y0uCC4foBzx9DVovx8z4kHAK8A1gL9E
3Ml41IBDCDtvz2GxfVF5YPdbvoItyRjSf60iFVC9cBgtwnlLJxjDledYqluFbuvdFQr5XshNZS5s
LwcJp0zcP+1DUgyZXtQO6bnjGiNIpWnZEaywVrWHinvkbyzXRQpDvVqzcMMr97eY+1LgBLgXHPjo
XF+1w0tCtLN3JTPP2CuArSasFnXSHc5zRNLQJH50MMI7+odH0idRXg8bUHdqzDE4MjrAuyagACoZ
h8kUvl8v3Rd4T3N92nfCA+qIpC9coaCWnXpJYpNjgrj6pO4AZFHpZegnUg0X0mnyjXmDmSv/wSW8
DiVGuF9eEyoV4Rreggo554iBOG8AC/+0aAhegniZMqGdcDTRwqQK5kJOJPXoQfMQ5/b/dxosrFm8
6xnRneWjfghoXQhbS41+H7ivnIrsrxVEVnxh7HCmhWDNfGFm2c1n9sHt2gYprjSCqMCUk05K99BT
gZtcN3RylcTx/RDMnw6HT3YkHgg5JAWCWwmqb0WXZyYrWliV5oRS0Z5+rPLvvwryTfbKgYyw5bI2
k3bTNvmZC/F7T1neLdpVDNHVZaAS+/3JMbUF4cdeDiULExJRLk7NsbvUccGjEBpO1/D+8s6gaH3j
6+hdrUW721L15VYhxONjA/kPNrcWDFjtzeaz2qQZ00KSckrVJx5tlDdeQcXYWc+N1yZhw/NRrcib
CaY2NOyYr42+gJgwfg/HSTyiasWJk576QQH++Pb4ynDIOPzmWjVPXK72WcqqsDUDDXZ/6XI1RF/W
7gdVZ1WGmGBwScAL2N5YOC3xFg/RPnfnJT+UtkrD0KnUIPgsEHf8BNhb85XA1Eg/M7Q6w58vvel6
tvFkHrawBe0zQMvLOj0V/jzO3B8QW82V4LVSOJptxCzZQiB9amYJQkwINfLbq1EQJlM/7kHVhDYe
MnhUeNamVCxiva5WKauOrQpI80axNHJXr6/omqWuiIcXcd+fx4cm/oO/5997frR9EifnaqCsj1Nh
Q64iOkP14AU0Jc2mhT9FA4g/xXGQQ33ZIWyosilqRWgpqW6yfb8XmuObz3O2eKVcDPCIGS3Q9Ze1
dhitXbIO4a2L5csFMYNODfeTwsfzg80gs/4VPBWRSxYXwR+CB9A6xBJ5a7Odecwn+PJnY/YXeLKk
MaV0c1Zpb/xBYadp4rJhiU0y2eyOJ727O9hjcOWkdU4QY5AeB5/mX3sRHrB53F6qXRjAYIIrPWqO
cfOhK+lfzHarPJtnVU45zz+os1P7FxRgfOEisimoXfxbfgiWibEMDj/X6jG81dhuDt2cOdnbDahI
QjNILs9XaeV7TlyZ5s8zXvd1kn5/0hU1xfn8ig8jiJxwGJzcXR/FjHlmkOyOiea3nso7hCGKIiXO
BQlzdtsWQInnhKzMClnFSMDgRlpO5euMZS56dtmnrgrMY40oRYfEEBltqb+CJaSPzpKU9qLpJffN
wqpSriF/brntjFn1mcJrXJ//dl+B7EIlimUlrC6jY5FePEUkvXzyu9FP43F5faSR4L6yomsq552O
Th2SNgZKh6Qb+NQy11+UEnFaYGUC6MzaBuqTwuSlKv4ZMGElUslWFw+sgNudZQ2P2dOwI7KI69K2
pGZcInFY+KuaOrRSsujuhRT2Y2fwDOze74pIV9t3qiVPwucUp2CRJMaKCKS9NtVdV2BpgkfiwM08
MtjioBSvHMldcgLiVvqkQnBcnvTnwcI0uTSHCkv0dW0B7FSlXuSMFcgfdsKqtC5Pj95AWL6E//tH
hDofFpAxjd572hf/BtPOKj1vcXW7xzUouVEcFGVZ6nWPZ6LY3CewggtMcBBnQGmCIXv7DXpU7cUW
G7/w+4aXuwADcWTqRUkehKwk7hEWmOBN9fCE80n2Iec04TQdW1UkutGuV6okWTvy7IZb9R8UqLlN
PID9ONUUsutqeiOmljHw8wLp/vkYjUiM025HARWs8c5MG2MaBUOWc1txpsfm4Ypo/53q+gz89+tQ
HMMKVxHYU3TZAQMqeD1MQk7mMAUbpTVcG30yfWyyu+T+dZFx+mCu3olDlGJOmV6hXNT99U0yhf7G
yA0LePvVbHvwHpoN1MnPcPVw2YrTshbPTOQjg3D7C1TTWies4ZR+MOh+GnAKgrCQ7ZZj7sUgIN9k
4hnFk3Rzl5FkA9A5K9EbFrrTEr/g4EswLSQyXdnpby2WAZ4zdZkfU/bbeP10Kfb5AN42UbdXpZaI
IAdcOPXnEiK6+Q1iIKM3P1Q8PkRnoyDh0zO7P5qv7+yiy8QQcGryOuF7jQH72FH/oR6AhJGQecxZ
CfL4KY6eLWMbdqxqlysaGYfjFXNv9ZMAb2Mk3bvAoo2fhFkMIUsZ2zLSyhBwlNUNbCbzrI8+5CqN
sq2olbaKvhzz29xHgKQ10mXm6l9/wWF87sMqYpeQW22Ja3C/jo2vVdp73Hjlu6saVYlM7zABTLuV
hejcCzXlrJbCthJiBrluWG/izg9qzkPcb/YJwSk6XOBysjNbe81yLnWTLSsGeL9/kHhni6qr7jeP
dW/Xp8vMAMBXBsNozFMsrjHWnRi5JoEXOCvUYC9Wk2QGjDPp77veiiINi88o8l+H3lElqvha2Tl+
qkkqhXp6QBZ8S5KG0+4hqDe4rNKeX9NHhP+mYvYbKfei9HNfqFI4S9WDbPCosyomwKRj2OXHHrla
Rk7KT5w2EDftlJsUyUUHDRkDDqbVUWNa0xUlG2+Om8Z+SBWBiL4hfGxsEr0Nt++So+RBYTa5k8FT
+5723pmreAljt6gXsMDsLXXblZiJmfzc//1zqQ/ASzpc7QvbwJq7BJuSgeSGNOQIK1EuL3lealBV
WJJ8ElOfGTQp3k3pzKTD+99ZikbVCu+MQeZmSvqg3eT7z0IXY1a7YDUyhS2ThmCpbjv7T1ct6qfb
Miuc79+l2a+UDikkN+N2J+ZmSBJ8CX/vhcDVufTbRcGElJs3kc9VVm3FUJ2tmvBltmaKkLYkbDLQ
gAGQHrKEektaWfvgHvUml46Eha6QuonvRAem0r6jkqoNC5pea3rNYnDIGW09lRBg4GxcDVprTIGX
3aRhPJXIHm+BNENWjp3AqVudMmPei9dPMLvr+atnRlmmwyPyy1pO2UdSqnOIushFtu8V4Wb30vSh
jIkKYgESM8acWpw37q99lCg06EzmKm3qnt7JVfmP2lzt4L+lREsacE+jX8YYRmxnPK1GIz8KRBT3
1FvaLYg7w3tm5l1MdazABZ6iK8EQH7JyJCzwDr81g3FiSSF5Xzp2Kht3Zf0wr4egxI8Pt4LGiAZC
3q5SJlFUJA/ZIsnMDiOV621UXw/sDFbhPsRyHOjSYLGyCzgGzbJeEVNQWMc4vqI1tY6IRAh5nUVb
uVI0ls7DCk99mTgHHz9p/DsCH1NiFpewpe1Zt9UYIU5xX6+44Dc0QDc3xDqIIRMjbG7eEz1p+QXe
ILjcbB9AbcADZnw+s9kOOR/4fIzCUvxsXL5cpLYm+aJ/gEmD+dsdSw22SQg4M9jAXCdgQMCbLRJc
K+MvvlOM0R6j2sYqLcMbTMFEgNALwx+wYhvg4x3Cnw4sU017kJdVJGYDtlWxXqK6KAKnglXgW7QQ
G1qSdQYBg7ogVPaoRWOYmRuG8ISYgBNpG0IiJtZSG9V5BolC8+QWYP31j5tnhOnWgtQ50D8f+YJU
C3ku4+Ba0N4Ilg2W8T5PvcSdSCgGoQm1qzt9VR9byairgKECAeV7YScpaBzHbIzxB0IFvB5PMDwl
Qe+buMSAk4NQaq80wOopi+gpWvUy4ceLhZqvlOzUQPV0dzTXbH3cccglEyVImYSdrYiLqO+T8ILa
xLjIJF3DgyBuRzR3OALkkh2xIWFwGEm4hRgZ6LDYRySt2CABcQSVoZL+qH5glOUxNey7b/ApUXRL
0e88AHyaNPjGQKvTb0SpjM70Jszss1cI3OH1XkadTzATu6l7DiDmBbV9BptmWV53SyWeYDRJ4HaV
xZ+P1WTuXiwVQeR9l9STTuFh2f304Ny8g48tRazdZ9WYSGELCMz5adXqhcXcWtEe3dPh8AwQC4ue
DyJjdQJJiRr9cZIO4LeRZUMi1GYeMk9xkQWLYq9sL+lf3KoxCVT9wSNfdcoV7BUr8NuPAGePQDAZ
zfOUmc9mvrEErV6JKzMQzXIV87NYgDkNEhrnQN4LS9KoI8oGT4Z/LlXFnns7GTwLe2buuJ9qrrP7
Rb+vxDvjgpaubOFgc52mXIwHRaqDI2MkKmDwndYqwpCpnqwkSNixretcG3QgmQrVgr9cj+0p1XD3
OzfZbRITQKKsOrdcXzlZqTpxS/kr3YCjbA3lkbBu5YRvZ9u/7QELD8//9V0fbmL1j/279/bSWtnL
bD3L1YjHztNBkSQv2hX7IMozJS7M7H3BIWfrhoHFnehoPdGre9zJF8KeBiO3dO4CEfqvDal6B7Jq
ipAD9wcHqRLHpKYiX/xFzoY8tceJ0sFCIg9MDQP0P+f+3a2eYoK2Vv97mU5azWq3qmZxg3T7oiAI
R0Eqx6xOcLISCEg1wtUsshTaMUxv5JPJ8BUTiPSHPd27OsvQBL+1edRBkaP88j+tcLrUVnMpfBxq
5+yJeqn2K1oiXCF0R7hoB9uzCTPUXjmrRDXCOEqQfibxlyxBZaeXqae2gshTWiNIOb7b1fuhJJny
VnIoGh0lTga7BIVm5e+OVdRUQcBPv3z5deaMpWcnUDGtltzf7fWudONQk1QvZypCOC/HREmJYIKV
/93gJ9gFhP0+qX7bPNzvTFRwv6+VyNjNEzQs2/HKMHco3U+am42bTaQdBWWimFe79fRhKTYwRh+C
NBWXy1GJcFGFdTxW4RKmM9Mar4hQ3L8syFBifGSxFDobJspCqTIkaHdVxJR3fciX9P0vrKtaqvcu
XerGF0gi+7dAszSs1yh+8ym/Taga+rzP/HQCnWvuGI6eaUNMuS8S5X7+9VX/NFmsRII7+3dBnYdS
r226BgPlA43+RPNJUl9Nvb61dhMvXI0U0pYLn2/YLd+kiM7ydAwFoRm4wsVyMyOTz9Cmz0UFkxB0
T1CV18r2pjRnhb4fs7njEoKsMYZUkau6V4VxlsoY4zKRs/+ukpank93ckAk3qo1yyhxg7J5pFfXE
PyM/sjcivLwizL3qyTAWJAfTap2JPpt4sBotgeYck9wOW/QO/K1mvdV1tIUQwjESSTVhnP63VR/G
XSlR3uqlgceCSNxJtQj0BvSwAtI9egN10GZ+PhD4UwbFsahRdJKXEfr3J0H3vk4M4vtY4kMOiOUZ
xCfocmHFTLvSeJdUj5VPBXcMDX5WNH2B2a7qbS95K+6vpnPCXeU4HjJwuQrR3TuWoaFdW9nKkvu0
cWxR9chaQVHlGwB/c9BrG7wx4Z7dBpVCs0eZagNdVoPRnlCuTs89fFysUZCLdtH09WB9YOM9Gymd
C8eFkClsF2ZAXoHLTxcmMEVSSWufQrEICgrFfHz+lsz9TsfiKlNNlNCnr6lJdaWlsqgj743V1yv/
UGhlel8G8PS6tM1BlwoF5E21rQRI38tSwVbrDqDa1UH/My3aOTkyB57yxuECfVrP0S53rPKfX/xt
OZCS6JNFrteHm1CX6IZioxmn8AJ5vxSm1eHFIyPd1vyMUNZxua8WToRQYmVjM7KJmb546g8tr3Fm
QZ6NS+6MxPo6rCqQRgGheweIl+a3j8kIwCFaubEu2jcO1WdyMPyXKaqkAHFzGAvu6ciaCzEw40zI
OPTWFlZedzLEZhhA2K7R2y2UmAJdBexqDQbLbBxxIOyUglHBIHGBsdrjFBXLuAx6LmFM8HMXdjm6
ReyXsO5HsaFx2ocyvN+mvh0EBxOSMZHENAh50H2o2w3XjLKwGSvGhAhPs/H1/lu0YY2GXSLB/C7o
bGusbFDf5UPQP/JcFnkk+iuU82KaGWypYfqP4hYvr3BhR17ggkoBS2cusCN809S/OrI/TgXVKYgP
7bGsH7piR3yQffSFdcK0Wdfi9Tr/7cRXLegi9y1XtfR1jG94t9LH65XdgdelekNq4t8uWL8crzIT
i0IEWHStGiWnaMg4/IXtoZ1c+z8waH8np3bZQDrDD6A8GUBqCpuP6+w28m6nP47SOqYfUrqwTMv+
fCURh1TGXWLEoPFBPpr1XtsPRwCvRslruTR18YqmbrahMqWqVo0FKNnQYwnyuLFvsMhcnd98li9L
/EZpAabSBvtkEKTAF6Oe3tqXBG2oNd70OpuLsi05hoXLy+VSwxPKpa+7vKa3W0+f2TZfiD4AMWSp
9HpwouvCy/JaLnzga0Twvw4McvuMFG+Vu0DXGhiVmeIK05JVW4SdIGyV5pqJWK8Q+WiFtMF6wd+m
6oRP8zdJru5vslGQdpOkKkqi7Dru7m/V/IKndP9fs/fPEKh5fXyYo+m1wwy+ISF4Xs4kjb8BINGY
Vt9lrcvnK3KnTbM3b0+fpDiPSJurHFzI4jfkOixxnA8QcgjrMhNc2Ago2tPsWtBocRjbzSiTvSjz
F7al/0370qodtOxqTJsKvYaHqSA8meLDHW/HxGZJB0lEDFVZtiO7iesH9Hz2jXGtX+SSSmMxd2IY
zq/k5kXbgF8uBdvBqKfTS7d+sQ/Q2A7NjKwt/IlY2QgmJutzZ6ngR/1kXWaG8THp7fythBAMwF/o
vaYmXjlmvdQbqYlTUJ+HGFUzleiPnkBc/M6wUryBk1DD/M4wVHn+S7vZxtMhktdd4tUiBqPXT/P3
ATTpYRR1ZJzeh31jKdXK2Lzw07aqGsmHZ0lb++USK8xZzRePTP92NzawQhWCMdHsej9nHhy7UqKC
dastwvOo1ovBnDGCNuxZAKygbmtEVxzuIfiYxOWJ2StV7h2LGIa9hbNnsDIs848IJOy4M5C6U5VL
Tr3gffXV/i9yJYkFWkxXbIiStW2rSBGHNzOz6n7drswo+rIf7WFaeV2U/qn8ImsQCVlSX+trf/SR
hgOnl2LDeq3AdvnQOoNiF/HR4t03h0SQ6iFopdIA1bitT/fMZYfEXeRh7GnJpYNNf+qoeinFMYsn
S1UDRk+XArZ87ZNrRR8idh/0pmh08dt7WvUilBKpWH8gHzY6981lnjKvuf7LNkYrn9oBsidZ8MlW
CIXh0Px0XB+k6ZbeJZKNLER6NoQFtK4h0S7ei44CQ7au73s8YGQnVbtKpMBozDjzVBUT7jn35aPn
0n+esYHacw4bvwppC/IrxFMADEcOVP8hMBfc+38545PYGb6NtcN8UHDToL4qOur+p3IB6ae+VDap
TC0j295KKYlSmPnI0c0TO4+g6NUl3h+YhutnAIhz8CNkL3tGW+fmZfBxQnoGrvgbd9lD2l4ZfR2I
3g4KArBxWnmBUm/0BlV/D+Zj3FiGph68SO5p3WT0bEQhI3Q5iI3g0+BzS0JRQbwJ/MEKtstyeags
zCPcdy4JiTMP8ihh6l1WmgNk5Syy69bJRPu/ZzcTHCqjz+RFzpwyC3sEbKKgZoamu3U9JJ/MF2bR
25q7JANqHmQdCGzarlmm9Zvb6g/YD3j+i0Yx4LniV3L0B8G6ugKnIi0sHbBcTQoQSZe5b48vH8/0
Qp9DCF6D5Y3UtEejRKD12cJwbXw6GmqHnP0RkFjgYJ+B2GD6FhG8qK82olDbSEUvCcr4OffZ0xxa
QLRIr3k2Do/YwpLW3k0Fnj61OPXM1ZzE6u7bMD8Yd33NeYDlfs+d3Fr08KqUEr8NRJz4eMxYI1qx
ysLQMHf+UOmM5NOy16SQx44BenpQm/XVN3Nmlso7R7MsQmgP+9gYeluCzZg2DGzM3/FMLVj2ekbo
I2jQGmnTSj6mqCFCgTU8kUw/3SkFNUiAf9vFviyR+hsUTH+xu0j0aU0PWUzGmCq/vESFz8KQucEL
od3X0dWe6cG4AJfCE5OFjjt68ryUBjaURVcSlgdgh0+vqaZG8TgOAWB02w+vkdi8Fk74aPeSt8uH
o8GWbRhPwfBy3Qshc3OhLr4B+22Cxi2R/sSvuAT52haHdSahaK2EsWHbiLZRUtZIUeu2jtOJdaLN
sFLFDjJBa21CRN3KbKiJ0SZTBSx0CcwX9TkSis8v5UJL74skvJPQs5WXCpavUEsEpyPjqnRJfLua
J1N4afXwhWjyV/DfBw8z9UCBHioWgDU2LcAImPkRQ6Cy6bPETA2ovHHDPtABevZjRY3tlhTUA35K
drezXCl3uJ4jg8jQK9BKni4H6ho93G5vGzH6RkqFD53gNuXmTh88C5bPqDcOle+1o/0MKa2Ho2cR
5xx5upUyWIExbwpQaph5xFYGCnuXmorvClZdKH1vhk2bXTl4NO8vJvZzgf1sANUnA7x+J9w4zSo3
yXwclof+gMGfCXgIGZrvhwNVbTc37haJESsMDhmrtYm7NRYACy/P7R7p87LL6VTgi3TqgkLK9kzf
PyBQ40blV1bjOgKu1Bc6n2uxdXNFni7Chr09BK8qJhF37bniRihTy+kCVJaoZoSunBplnxxwtewg
6/Xp4q8YtLU/It0ddTmhWZYiTAsVSQLprFzNmnThS31E5ErRhGGmYLtoUU77I0PNuGv0ZuLmt5rZ
RRU8TFTEjnAM7JfoyCP616NjwGyYrEBYTcIFwpyR8lW1WeF18Vd4HrL9jimA3vkXHpJB63o9AKos
TOuSvUUP+MApeE+wihWhkrCZ6vLJL0/5vCfzEH16NDAskz+KH3o3byPZeMt5Gy3ow/0dnXvNEKMI
5UjQYKKmak9rIDH9xNl19W61QDQ/e+mOiKmToE7ADHCFE0IuP5rGhgcwqf+Qt2estJDe62g+MkG/
NSuMYr7eof1ok900Da4oqebmmHY810DgjUKqY1QlhJnon6NTOg3+cnqYFykbaUJE/ghEkKlT24El
IM5nYjcDavdaCYlYcKnvEh0bjC6yry9KqDqjUOLqLO/IdJrOreS170pzvDfVA0bpZXmwjHiuzSU6
AG/o6TXM9HONAfUyEtJ45XNkq9DsKSNA/mE43R9UuQUerkPoWVkwUwa9vYoMYNZJ+UNDD8V+OBeT
WgWvLpNXIhit8E8IUyyCqRv85ynN8lgIPcbaAF0FHN/nicUpoEQMT1SFW/PcMGcHAYyMvSp/QRHO
brw680fMvzJDDKb9i8pujAZU5uCGceP4quP9tlCChtSngjW7em3ovJOlbiNLbL/NQYa1MFAgau2H
WhjL8AZuMqcjX/UG8U8QV0r/u6J8nkxYk6FYzFFEj/JsiM3IGSanoluGehMoKs7Ng50kHWC/9OnB
iKkAG/CpUgkovYYdE9r9HWrMshnd0HV7TCBr51Rw0osMI5S0QFg9HEU1FG12eJhOSCRcgcy/+Yn0
4wEuP6ttaeWFBYpBvgFBDoqFRnBjGz6bvmCDOGPgFPoi7XettUJ6PryhRyQ6zRTx70p4gp+xi1YC
n3kjtzaUQNNqbjr5VNbKuL5mXq3I223wfq17/thvPsremq9xxNH7PZAn1wBwnEPEf3nORMDwPKxq
AL+rrC/lpk/XISMcmEY2zGs424Yc/LIuOWPBOgj9qeET6sdCDifFGGizkVL3GpJ9F+EUaolJUksA
vphIOlxj3ybqETqlrjSQMuprSJZp4XxaoNPhmEYsL7Eh+m8WAvgVumGPhvVMEG0zJKVatUsli62U
3kj7aqRTYM1rFM2msGOQT8BdhODjXtn/1aGMmwaBCXL+26y5qMBVOpBcNwn8K0bjbJgZXfa4yDGg
5PLOGoq0lVVBwy+BPF4Pfqql+VGsD8RB6b648DVvcqxtHvvk+ZzigItpxVVLriDkk+P80BYCNkyT
mm6qHYMC74DlyidKqQ7Ub4Zh70OoQyyWwqpd4ri5orsYbLy1KbKkDeFPfy3yyb5POrJ2sUSLHE6X
LHV/jBWUDHm7ODLNhOV6LTnvXdGyjeZxprYKnYQnnHNCokFcN8N2vAu6+/zqfrTLw2SBFEHI7eLg
fB5uGeYZYxWz/d/JO4vl3PLKdZNDFfeLk2Cb0iRLvX/Wd4br5oEEosW1+8TFE4iwp49r7j4YOv5y
OJs7AndqQCHYXQXxTyAlNvOxFKjWdb6FSOyTY2qbQ6m0UfgQjlQO0LJW55cs1MhExX/tecNgvTx/
Tz3GFA+uBa/2FPRu3HCcK+P1sB6RnlLbo8/KiKGDP8dTUjpQt9KGVdhsTWzsA8RREgBzfETKyl78
439vGfFQJ5uaqTiJcM4SKQI/1wF5qrzQtxM6sxjyYVa/CbBpRkX1SgRUHYn+DUdH6sLqwLHsklWL
5JsG8IPPmBYIEixIlEud3mxftjs/azaAv5DEvSAWm1xesf6ukPheq24uSaGKcPdbPlBwRnqt0sRJ
wQv0h4/zNFuKQXihkdEW76Ie3awleJECDEK+QnPDrQOIrNTwxtOk/tff3VGuXsd9UMElTW9CEu/I
KWGBWj1C9+JMdXwXz7rf6soy0/Mge3Zb/CwzK0kvXqiuNrNV3VnlGeO6/0mATksnqzyG42zvWg10
oTNtsQ8EmIy72HNKP8YJXEid92rFLztranLnI8lW1EpnHaLrolEqvcMmWwhruVhu0kZiARHl3LgY
PA8fnyrocEtwTFbbhh+bLdIazF3jQPxfuXGFhmT88H31yNJMCVCDlh4KNCGkOkzjC5PnGHTTGhzx
xjZj9QayHJig5zD4o2czIzYrZvzSz8tJCWXfuzOMTWH4Q3pjX33s7WqHEt4cEGVBO5DCrf0VoO2p
/okTw9zZhvBKA7ArSprZGTC6gaEHZW0ihxjaAfB1QgZzGvLhqDvMsxtkQXSC2aC1UC2hdj4SRcME
xGZxllNapYXAfZ9dH7W+SrEHmrSrfic8H4Rsavrz9QiBS0P9jXiHx3ymbiCmBXq6C2pbpRUZ2RyT
f9RIvijrRE8Wzj3goKVEgj7yM3hX+o6BqCHeLjfLghL4S7JyeIQcRj/IV6dwOu3bShzJSav2NHD8
vOkHv5L2bN7lcpb5TtNU2cjZ770H5q98b0kQ39rliSxOuXZES9dXdNDccJjmPDyMLCMbiWGsHhAY
LV5r4eOlnUZ32mBRTzVLZYz89IujjWmNlS7tCJFncJf57AcrrDfjIHyB6DwzazAYdd/dFqq97Z+n
F3KeTYaoIZJ1cHVInavcytBHQ0sA74Whl0IBGq3YUxL0bazIP6ijfOkhPVT8dzWToApuqUGctg/t
Dpf5vtD2oCBujOfKtEx44s8trlWvgt3Ypem/NmS2BMflTNSi+zJP7ZrPzxZyK7rqFCli9jC4XUnu
9fCbxsMA4cHlKCaanFQufRUv4+KoQ8v51dFuKF2BXeS/QgOlGbsW/SU9DXMv7ZGERhdFH0/2Yx/I
k0XSfnMrPSZStpcd9wkGtgaNFMQZVlHx5qfvR1hwoKnYVq2SMSgVt29n6DvZhMIRXreY4o7LBQDA
DPOdzpj9uUdxKWfqFa9/quyBNYNLdmqN4lL/7Iya+iieTh2bppJiryn+O+bPabsfOVMCy8Ca7mTF
4J7xSG2gzkMlq8/m3ScfL6PlELc2PLoEn0FMBGk7kpbbIvcn4k0GkRejBWTD2iIMoc0i0Jg1jgmW
TtpTrlE18m1e+AVOAWJkuhllzNmSHGhWnDrKPhM6U+cW6DnzCRsv71S0ywKkdmRjMn+CSoB0Phd7
PHOHwkVxD8ZhYnpjUKngEdgK+sg/thUmTbkRXwR61S0JZ+h+SxjS4qfVLpWgeFmeJFxxcogV6Q+o
lH+BqnHJAYYIu50CaiJr74M3gpEej5+Q2x4i1zpi+6Tph8DTwigr3s2SfiDa7k9ZGdA9daqMGyuy
Cfsb1mAJrgbEdBheAaBy+p2sFiBVzS01QqLcJC2/OxewYBuodUXNJAYbQc9ZPb9YubRjfBCDvUkD
pwNwNFz4S/lilttZdXOav4JMm/P6DqNv7rwaT/Eavj3cYnohXdjJVC7jaHVgLjYs0pS9e2zncQ6T
WURf18i23O6MX7ZuA0oBybgzSeUHWVieXo/KJ7qJLX9+eHI/RIkgDFN03lV6VmtV6KFWyXC8xjE9
AizqE62Gbg9ee/CFb/3YtErauDKjLmpTal27eMxLHamOPDgSszZiX/Tg29UTmKUhDnlhO0KVyVhd
yYzTiNKFi4ZRTTSbq9h4BDUKaJenq7lkYcwFYC+NW0CYblfFMtc76hY13lUMxPgDFShJL6llKAiE
IZr5+nPVW/VMZgV2ajdFDjCoYdv+C6xYbc8ZPd124GlUqVKWHZj4irP4JvBbwbPzY3VMFA0Icmpb
gyYpq+/zLpdiHO6q37H111KrQt0RfOj/wT/NN2vdIHGq2JNrPLVVYyItri60LCtNPsYF9NF4+6dZ
SZ0RV4UibVZCJa3IQO63f3j1nVXb8GZMPtpvhHeoyQsh4A5ZDHd4DuThGjt0HLmOFkkMQ8r325lK
Rtm1+YwfZEVj7tOS9XUxbBm1ycuBhtTQNXi4YJLegn60siTyGkd1Mnz6w5xGq4NYyC5ty2BpN7Sl
jAkzbW+Fm0pzkODJYPbu4HuD4ckrhh48wNLIZoDMtgNaeQktG6RX1m+ZcQXRKqLtFIB5ibi8EMh+
29ysf1SymJv6RG3M4cQvVU3QNDMnffd88lnJesS+Khchqs7EDX8Gokg8YWYuHIPN/d70zZ92YxbT
XW6EYGwvDyCWsxSiGjjAWkF6ZJ2Z8ReHR4QtCtVZPtdGydJirNLDjH34w6jBHxIpPWqGbIgQU7AA
AKi3eLFBcjgqL/4MpTSVTV5GFHE47TLHq6dqEVjJnGTj5o8mxzNFmqP3SUMFUdTAeL8Ri8icYJ8n
F4nURCSfbfdg378EzQWV+y1T6ZDYcLgJ8rAoDi4uJyPHqMCmHmidSuSc/yHGL+GzaXAVNHWgCMHm
nMPAQHrj2UytwYYhVrbQm3gUwYlR63Xi0hVp6cjdAkSF3dslqKPX31sQdUSV32OxjRHi5wiQfAxP
nXA7/HGgtO5Pdw+frswh0dHj3cq4sINAbPLP9wtQnSan85pthJI7JS9rOmrV6ZU1EV4hhItzcBIb
kXEACl5KscrjZXA63nq7LOtowYhQ+Tm1b8tkWKn2kr9luGPYedImUYSl9u6pBmbN0nEhhP3jPTBF
rspB39rFTrnP3SbBeKYdo52krIwONFo/bWS/kobjSdGDDzfRiMco5AGns343VwJwFM63NPjFD3E0
oikmqCBRTXBz6fsgvb6q2z2p36ChyIlcjMU4afzs2QirnTvKmsL5xj7VGYJsReoyGGvU2hhj9WsE
O4zmTb63DMiigBbrVZ0Nl88cKoGFRyRU+WDwRSIvLKC0z0yb4Ac7W3adNQ4UhmJhnHUzhLWRvP1v
Oy8qhbGESVR04ZjXp77SIqzzF6yRF9gHi92T6yVUp1X9swtvTauMumQzioacCtcRaHnBk647Nm3o
RWuxV8a5ZfqcYAtGRnzK/OBsf6zj70JhYBA5BdIpBJOfMjhTJS7MKJFmwa8nGwqtUr2Ubt48Pm/g
a3scH2mgvi5CJmgi9KOrsG8UHQiRYmFzp1OeV+bEtAuOy2bI1FkUnhwa+/cIoR0sZlfSw+OI+MPd
yIQj6XyM3EfJ1znoNoQb9jpWFx/KQfB9n9SqMOqXhiuPz8SGlKPZB99begiabEkdblYzE1qpms3e
1yfbh9Fb+flpjBdcZWsu1Evl6c9ct6wYV90BdVhrFtakacInE2U9XZ85xen6wbYXSP1mteSsmNsE
lgVCqbQFKI6Hfw0r6UQpl1esJeB6t2lvRZPtdE++wRLm/l2dijZ+y7jGJKFBYr8kK0kWAYCcuAk7
TpPEJU1lHSXWtx9lHgTomnwTiTe89SIlff3v2U56ZLu3RjIiG2vrM22TWw2cMQUfo5F1V8CemwNb
epjLVtlFt579sHsfCEqSV39oATXFDW0bI/4Pjs0p0Jlfm7nMnsivCSqFksvjUe7vDcswt1/Nf6u5
+zCgK0VM5GGAgXjbqhyLMbyGql8jtKlhSvoH8gSj+VwjwafxbCw64a6aqq/0mkt4BFLf5hBh+5xT
P/Cyn+ZM24P3FkseCSfu9HNm1wxKOlZTceZlAxd/SkKCKldf9+RYf/BZkKFTXXxLLgsjoyaByP66
855Tj8Hr2HNP/zpKpH1ELkfAkkp9pEmRK/Bmq4J65XB3iNlkcuLfEUNbGkuFBQd0fGQS545OHWVD
bYjG7hh1IwqhTEtrlGTEy9ovt9+D5IaqJXqPUMSHIqvuGRvaqwTIYnwv4R7lXUpflg3xOVfCQfjf
S4CSHA8tmkK+I72bz9AJzcOLrZ63NWx9uLve/g/CjLaiDzzBjXlcLc6wyw9rahBZeyQhVUuwvXyV
g+90fGPdsecpWyHOc9I8PpWEvGYWLYQh4LAkUYhoan+kRfr/Rxe9XSuUCtS3FvD1WzloxRFLM81C
WFdM7mMLbZtX28WwqOGBBpFYKic8kEI//9S8xR3z2DYcyu4Wj4AI2KEXHJ9s1AlycFCOdAH4Kbkc
WVIBKwYaV7dqVbn6xvvX6wxwcTYsNuXyDX2QUMThWzboNxgKS9ixh8rgegJviN+Lvq6u7XevWehS
wacDBl9dzQ4IdiCGaJvEl3f8uh7xtcrZRrgXjOkjcL9ayQyMyBSwEHWhe0D9pEXP60m1Ys4/stEV
U4UP+b+i0lBEH/aiNYNNZLH5v/ErLyJEswIYQP/bYCRa28UeptNfVgvZ3ZgQ0/jf5BhFaquoPHOF
67ewCjK0pToD6aFpRP5gGC7D5HhJJL140WCXO0oyAirY7R9Izg0reb7hXwwLwecvY3Jkh3i2Zsnu
GeTi/HCYlgofPL+/wib9zIB45YjqO9FsUokBcDGoNnKVXVfK/seNN8kQGd5IMSQPhO+zTpQxn838
sZ8KY3lppBoONY6vqYnBsgT8Taz8Ibo4pDCFiWJbAJhGhDIJfIPpKVE5cUKAqgxCsS9YKzBx9Y+g
+xVaqiZ67FnzP3e6zNza7eMNFWn8lrArXFwqwwM6l6wrgGIqRshvhXZ16hyvMFQwL0AnZng/ryjR
NDawpScnVglgoHpq/VhUIvy8K/qHRb9qfJIOdSHP8YtKrT9oga/a4MLExSABdgSZ6Kjho5rKQO2t
jcS++Uaj75oUQ3VRF39ApLj/T0gCAt1kLtj5GrQIUG9U9Vr1qMr3vTQWrUC2dYH/aL+OJQTSGCTV
x2cBqa2rtPZoEXZ6YPp6bD01BIKsau41MzTb0PvOlE+uE9EnBpfxwgxThoNG5krydlzA56NYq/pE
Upp7tUwHsUirk3XbHrcrAcaa+VNOUw9NFpg+V5EWULP4eRJmtSygLV5hmTqA7K9zTqlM84u19T/s
t7KZR+SsvgRBjNY9IKT6A+fqspgMIaNuXKUg9UW+MpgaHbg4b78prJiwNSF+3yReuzckVeCcGe01
2vbPFy0qwVUUu0gnj78kGH+fMn/PLu08ggNE3FLQFb8nrAUfZx6eEJX+9ZrulFUFFOJr+pODs+rN
f9hMVgUVGDpYEBfuqWQ6LRDgkly0n0lyQAnVWDggZ0uhfP4OAu3fAUikFc0h6Ggga0oz8RCor4wT
Vpavwfw4kBiigEWrDFMYC4V0qBOog8w1BzwWsuTeZslKSPtruQHk4tK1N734Pq9hhQ3TGtB41wtz
t7vZPYXZcbY7JQUvLCNB+YOR9+Uu43I4Y07mSA6o5Cd7ac9+lwjt+8Vxipb3aqNQUVkA693WyWGw
HWChhpTvzLqNVLgMyXIDTuGQF5yQH+t7MgA351n4gO45U4QNBGwk2bCvScRbpPOZMAK4BjPNHF/I
J4sKTAu9ieO2f/fuTUGtttwyzTqQw/22E7Hcw8nt8SwsYUyqThpe275Nc/Z15JhTnHeAukWszMrK
J4jaHvyfq85kqQeLzLus0loQmxnCD4+w/eGcooiZy53dy9vsfbnwjSiJ3pYnmn3ObR4tUUUxe8F9
rL1vPrcTVNbgKps+70dgzicWZAyfMuQIucp4sJ8xV3YJBVKD+Nw9XECOaGQMZmAfuRR3au9NSHbu
4BlOeWexWD5XQvACYt0bSEWE2ZGG1oiWU1BwCF0IsZ3WkPRWAIEj0T9pa+1Y5mzmXRhSsj9tDSjS
TryOeZ7+hoWh6EToFZgqKVEReino7L5xW6MP5gr2B8IucP553c1pRxOkiQ8HyNpsIDBK7wYe1fF0
8z10MP1rE1LUbd8Z6hrvNk5tHbAN7BZ8uCcEu5fzj5shcwYGkdHvDDEeEKSNu/X1QgMjhpOftXMJ
s3f2KbBsElCS3bE0N0qRxsebU0Qj42OB/5rgUzXHHufH+iQvEXdZESOPY7KlvBoWv3d/dSkjvlke
9aBZlIDYWUDLsR5tZNbfbfYPb3S9g6lxwe/W4IkW+DOEKb3meQb1ah7A4C/Sxv1gEz8NgGJeRBh8
i63ORHDlfv1lZc3qIKx5M51ZwF9gS2e+Iz2qknJBt+tN7cOTED+V6b8JuTvVw6y4PMQ+nJWByjYg
jSmcIOLnj5qOhS5eLZUXgoFr3VwZiaNJZY35riTspa74dLSzWhhu/iMDZCbExncJL/1RYLxW6uhI
iKof6inHIyOmLK4IhLW5YinGIpSbnh0kPY23gw1x5Tfqiyveu2DS8WjeBCUuW3rZ8jrLd+auKiHs
GC3iXy6t+GRmzBRdR78M6NHyDthj2EKA+2EpKKu8hXUcGXvmKREmSlEIL30sNthd1ul4UwTXVF6g
8wAhWhumRvEaFyPaPKOGhNcKvOGfz1kKWK7ZMjxjbxqeTwnUmsSWeAMh92NQQ6tXlK0VYKrnQBWx
RHYBjv20oNbWGE2AqbqBpqirKWvHFIu077XdVP0D7BmWeLKlUeUDXJMUwOROBQf4HRLwYXZsfvgL
Uyfv3P9mo4S/YlU0ahGxI8Frqb1Yv6Dlsj0Xj2nzPQtTkCknTRjf0o8WcKVRMQUzqMvRz2qyG0oJ
BFu8r2N4tgXQtBZvK+3VE6pCDYH92g9t3CnGdN3lSQmYrQDefncZoCQDH5PXD9sgq3qQyCrZv5yH
MxCR6hvb4gYWjj+LVy4hpeD2OMPrnTAhfJJXfgkpdrfPB05Cs+Xk+f8vjcsY5JRT1+PRnrrbYCKj
INCoUUisSpW7jjo/C7w4uUOJAOy6o+PThhAC42Eh7/xUXjPhW7nyfkEQWCHBLK/AlObBW15+jmX6
R5MmONe6e5+5Oo8rhLnKglBj1ILMNlwCOk9JZ9VR9gKPmIs+p0s9VaK1HbzCP+LNDXCCnkDTo7uM
ePI/0wMPxA8FtSYkHFI8LG2c82N0UysqQIPQTzF3bmghUQYB06GWvxhQxSHGtHf4WTXE/N0sXxl+
JgnDkdJy/JM5TuzBKt5eb0U08B+rBA6yjqY0uoBHDgzee7qILNi/jWYuFNkKwB0ec9JBvc2oE7XY
tcPFmQ/cNtA9qcHr+eskN3VyMB0dNr/PVvlHvVdEEOXjWu2eles836lrn4YiaoN67uTQ3PJpHBbL
CoSWY6CN9UTiheuR7BtipFIRTHjRzp6DZdhFO+pAYNgqNBavBwTZ/ueRljTO7ErHaAolJtRMgVwW
B/fMAmdmdwJV1ESWPk3vITJh/LlochMawrUsI87ROxFLbXa0+LOitOZ+QZjPejoBNxIJtidvzKDG
ORhqt3upxmbr0wUB3hruEOf0hRiSuaqULp4zPae9QKs1Fe8u3cYhRHy5zF4KwCLzlblF3nZ2LchI
gAH/47a6n2wfGz5sJlydv+ZG1xj39IAT+D4G1SmlkQr9td+GtBqZus5o+hbb7htsMcvQyIOg+oMF
/r8ZtzVtlfo7n0o70kmXrNLQ7KzuTI4MrilYYjddDptKbMd4biibJh9k5V1cmmQGs5mBJ+Xy6y3B
UbHNCT960RC/YPtCTai9ZMamuKDIsrLF4yesOtYYP9M/aUHlOO1p4aPfQ4Ru/auFBpO5ggRIwp4n
SLBAcsrXdvcF7IahodH0S697+pi9l8ICHk+eaq8nVE7Y1kd1h81HalV8Jee2vcfT6tuQ7oDDFkhC
xvKDsr1wAGvnnwY0Ht+ax8jyn67dxLUHOdNwESfI3EhOSGJLo189tVFQQMK9A2JwRNg32oqjzHvU
bUOpTspYYWkP9mwhi+AoQ+cqZ46af2HJZg9J+Phs94RZ5TPdl6bwW2ZPvuoBVeZDz6vFgXTP9LgV
yDWni34S8krTCRWcli+9plWjd9ZeBD+umxCHPQbfvTZLHXKRi1oU4oXMX2bkDzab48OXp6stfIy0
+NcTGoHcRInQZn1YPYldGKCywYN0P+jQHRQtOBqvKUYJyo8iOHUEPf3ANrs0FUEKMfTr4iCdGzf/
QSDL3Wf+1yhHSPZp5SFmLYIBZHO7gfcB3eCewB233XdZdSxjxcIay+3qW+ddU2xeNKMqnVXCvW8E
Y4q4QT4Av8eu8mKNpCMUotXdTn5zoMv24qgUTlS1iODByZvdRqbt4hGx1Upp4+omvv/bD0iBvvvK
Q9kyucOp8w+h2t6XXcY0DbNaGxhDb/RlrApwnPWAMD6vgmTqPUz41eoqbqA7QYt9pHdQBUpE/V4W
agDrqfH5IuuC4jBEup/WXq9q6a2DJ2fwTusByKXFY7R3CrS03ncIKBGUCiBez/X0BC+SFxqg+8d6
E/W7tQ7N4/WBfZ7urPULkehCtZIJnPraUG9zqXCw5ncaKpZ/M1rwHJoXNva8DIm/3RaZD08dcbFo
ckiAlx9oCGrfXNa79ac/OTwTLD6AvTM7BktYQVjE11R516THev6AnuUR9tPJPLXA4tFcuqG6CK5G
n420nDbmJ57W2SaQsxbEM3We2vXQaydJXZXygShPJPKT/k0MNZIV+QAZvOaPXfTkfuTM4ggkTIT3
rdVV0Z2d6H3xLh52Fvi/1j/Xgf7NyKXc45rWYfDSdN2v/6rBs47FUKgNzy1vF3dLibHy2BmywEv7
ko9ROcxSf0d+m3fuySzogOCZ0xdkMG5KLkujd8PbnI1FgoSTbfAFRWUO4wUZWjwz8iKxJGbcS48z
JcVPenGOkHBcpdWp6+BLkp0tY6WhJZIVzizySExF9KZphxyc33IknWasnXJDKjVsFTXgdy0JWUVk
uN4eK+JVWtbDKjW4O648Zmr9yisoxdwhekOqrxhVilICttNHfwWegrZD7hYambf8NYq4AroOJjPM
vZ4jgto+Xrtb9HUF1v5d9TKfKivEqCYFG6JprQqp0E2Hl0rCW/6NYs4IpVNrK0Bq+tlL1TNjmyUl
Hi1NVVle/UysoOjFCtJfur38D3+rFJmly8wW8pq3dAukK9I3AhOM1o6LtYSzCKYMvacHDkpfumnh
z2ejO6EPcFvvs34hRCPoPR4+Bc0XjtOa0Q34RYvhIWRMU1iscXvfwxYZTIiKhZXK0C1LffYLb3t8
4GESc/vQhIcxF8i+bIswaP1iIqDbWW0GCpaTov4QKVHodhYS35fhCgl4bU1How3vNEwQD5d4KPSk
UcZQvHPi5AwY5bzXPoZazSh+r/j1jIRImEauHY3l83Z3lacDUr92s9H3s4peK+mdSNjGFW34Upra
f+cWWCZP+oAv2VrVvsYIb+2jzIY5hoYLlHCoyz8NPkqJQTW70NFFXtQd9fJiloYeepjTokNn/1yz
iXw7mnSnwBVqa3CxAuPNwgxqMvGrtShjZx5fSACDhJp1d9wLDZzwsaQkBXFzTNE8C/m/qfdzPiFS
1UgPEHEPH7AZQLqOtUTtlrGo/xJAjmi/ku/xCYn9k2pq8+ZMWbp5BQMV2riNKyZm1I0/lEWitG1N
dw8Lh/Qplzc0D3Dfayu/IBWMIkllPayGfTaoPcfsz6F8T0dxX1fWL3PcDgeu/onHlD5oHZp2OvYG
Y7au4VsUduSbEvYKIkOmXePyZMLmE9d7RTqnoMAFiJHN1ssAl7fnGsz6OHtpt1ydAlaq3+JwSg5W
DcXPHvgtWrkyGsDbNkFntaZrM6tEKebK/euhfGrqbrtWWgVSXZ6pSURS8kp4KusL6b1eA1ex2FpU
RRqq1mMy3Oo+tKCb5K/KFNG5MA4fU0HP3/3qrF3OHytwrYVlKBkTEivt1GrODy/0XA9lis21fg+C
vfG+JE3ER1U4btTfJGWFsRH9wYMQJtBeqH0WnH3om3JwNXxK1aKpM+2wYNRFw8ii99J4iDHJQ+BP
5UWQtnxlFBajrZ+Bz1wmvr2MZc9Ro124819JpHcJPOCJVijsbUFb38lRxpXrIbDN8SqtjZdccArX
5rtBEzs2oexIZ69cheCYVoqrvtd06qj1UWsKrdCjyVx3k2HRxnmmnT52sxmouSWAbdIOiKL02lLM
N2BrPPcszW+dba4UKIrBoRC5KFAWwg1R9lw6GAYpTlTjQH+QuwUFyJWZT1H0wewohSGa6uA6DRKT
vjlNpTExu0iWK+E+R0nt+Zvpu+LQlUJdziBo3ldWvGACBc2phF8ZTMJAgZzm9dzPYCx9NMAwsO3m
eJEJzuJefQeWVU9lIRcpoTvYmPpQxYKfXZt7Ea50Yj6GYE4XAXC4At+BBAZr09x4W5CgfX6YvEYp
UhisisVRtT06CYRZvBRIr8Nz0DFKpwE8wj8dKtmrIi2wuEBFq7Xix2PUda+FxCuF4f9nseuIptaC
xXU+mDx+he2h1RAGfWe1eiXG5wIeERi8claskAIUywCohhQ1OPIFqxGMsOpI+4n2f3ucXNiUh8CG
Ytt4Z1p2Eg03gdDCWEvC1ViCkk3n+SnfKxxC5T4QiepLbkkFd60abEUuFmjXrGm0iUHRWU3i5ofm
Tgcoyk7G3Wqp+h9GIeKNKv9ZiSUwXp5tj2P1xhfFPzxsrSpvlgMuwcvydZeZvfq1HQ9ocFb4ksyd
SPwrQS+gCr3NdpWHTBumyBXt8nsvHW9Xcr4Fv1f22p/JL8guSBRZtOVdbWflkqq1eiY9KhRycb3k
+BHGMj/ot0k8YBVcOMRLBImoB/bLMCWr1YfFzOc5k/cIRSTT1GtZ0YhdVaNSS7rqeX25Hccg5VpC
yK/GVYK1BFoYV1qRuFGrayRb2ic0jPWCTo8bDKmc8hvxGqDsRn134HZGgb+Bf1TqO8t9K4fq61W4
47b3affmqpIeuYn8Ldi6AQU7vW4ofsIkK5dXa0jZl5iByVYYsQPqoiz3rr6f41/s7E+9e4aoe2K8
IOE0zjcJfglMF0GWOD3yv++tEtrKMgeOmDUPVhzKeozpfgDJMJhW63/wEmSGRnqIUakhEDtHnN6w
ifjpcxWXQKWWubAboAWOkqvc1jbzLuxim2qRqqumQMQAJQxLFe7f/UuG2Aui1PlNP6zGqA9KEQk6
x19NMQdiBZRfNzVUF2scWfz9Wcppim29SyiMS2Kn4JnoC9qcwEfbxrmPuuMHP/jYWq9aUMMIPpiA
8tXRVeRYgE0zkG1Xsg+H4OVs585XihL3l7JhmJ+BrfrMLN+zVNquQx/49O4ShWkBzlEXmSDguyVD
M3qsPxBI9ANfpEBp5/nhKCe+S/ltchas8dfdHuGKQQiiYdtQDJ6JMKdpdzFyrplZW/bEZkT/CfCg
TOrkjewzJfxHCMGTmU8dnG+NJg2D/gSHhwlwM/FwJuFYIZTAgzZ57jq2vpJhmynP9BWYQvm+t6Ui
kgFFV1MDZoupYR2e9VtDk8F9QOgTSPEgH8s3ke8AU8x+A112HNdZvn/2yT5FLb3hbqxsyTKrBYz6
wQ5/h66OLfDp8VmWyzEUddq7IzcWVyauZ8wcH0r7ElMqejMyab/l0+gD6bb555NBdTOQ67veoP26
LKAvlnNGMRVcz0EaoIeEEqbCwqHcAKPxrJbviqxK+QK+lo0sFSlbaxa+4ojRjAi7jgw1h6vDgKv0
i3u89Wd+OaUenW0n/kHk3d4zPCxmGqFTaNuWEdynpjpqcJQG4CdsvBTBizf/OwOuSSpK3BduQ+o8
ZHfL3ORMaMhefbDyNNyRt/AUPYelAJ+up+R+yc4Az8NbdX4We0bULzqfV5VX5S7rRP0QZfL2Qwtx
UriMXKcmwcylt8TA9a1iL/nlEAeURdx3xQhcXNd01RiU5bYJM4jiItMBX/oGpkkTed8Wrn1Vt5LL
vR9Q7QjumdhEF4sX9jZseOVoOLOmv1KertN66Jx+N1suHB51vJXMWKt4EUevruKt02ZzlgCEj++5
GapXFEDAZq9Z+JtTi8IRVa4VeMAKjp7eQM6VlER7KTe3h2WALaG3akuIGOL4cDCYEc4iGFVSIQEN
RItDjKopnyRGJW7vc2mb4Uhpy5/6zK1FZBBrPVvljgHTqoUKOWMn/Iok+elLkSYh2RyUJXxSjfIB
DPwZD7zHeoffnYMGpLaXxCLU0NCUfspOFYD1u7swbu6PY0E1VzPmPq7nVCV62cGx1ia4mvdJGAko
v4G290ewROs8rgqGkGFgLw8YX6DzloV60uy2srNqGUu0NUxRP3Dz5xC89CByMaZg7WUZ6IrUYWb2
yLsJx8YXB3yFv+LVwVwLlHHUhXwfzoFdAgRmh9yTynVe7kodp5TyHVaacGZZbH3KMxAdhG5EwN82
ZLY5KsXEywki7s3KjIfAbG+qvo0IvC9yrrWNju8HKquKFjWBnycQQKNwilXLhqkk0ybLoUumWHUb
rq3ZNNPzQtQekUUq/kR6o/ua+keE/i/690n7a4WJHgtik6x4Tur/X1teFTYK06T8nLoXKDTa2Djm
2VUxcttYexHE4VIO8y62+FkgSDJPefI/YKbKuZ7+Ko+fNtNBzGJ9+q2sbzm9wbhLV+zvKADwNSNC
9OaTdf7ChGZUok0TRug/r6hmSAp5SZlKZxFX9L4wB8PC/Y1NJW4L9HChJvJnEHq758Jxzuu9VXMC
dAcUbpzjYNtJhBARAYuPmsvQYIePRi0SBFd3pMhVxYPfLiYBj8u0WWZmyqUgR3uNfpDsvJ4Wg7xl
ertW7s0/8oP+IwxyUEkKW/ai1nzttAORvfZ7DYSW8kQlO9Les6VzFjOGB3iIp2slVx5sm9cyPy16
6lUZahUQckgfpAhRfMZDOaX+HPxZO1rahZobAQBmuaf7BGL0AcrXLBodVt5Gwp7w2mNdH6huqekS
MEk6SuGBUKBP6NHkLI3AMqlbhB6iF6WegBRdHwXG1x+a8MaT/T5nkANnHciQnxq4aBpa8B8BDEwY
lBhOZLCFGNuDnu5i/WU8KBuRTPFB7F3grEbExei9qplBxSQeQqMDsZKU1C2ij4PaEQHo2vXFSwYt
W37jvFkv3UWnM1LzxADigf4RlEOAp4gWxjtcR0kFMLoyaRGWJsGm6Cbfg2f0xwAH9QZ06ljR8uCq
tVJDcf9vjuEdyhKjfH1pWBklsJq6kSws3K4/1KR8y74NJcQRwZtwEro1YSv0datF0GgkLA4qY3Yl
b5uY/FP7ect5w9CelrfrIjTYijUO6q+exGEgPc59Bud5o25Okohd/gMrIK2qyjlh6dSAzIhJiHwO
pg8moTVQibUeNB69kjMhr6BvfBFWDO10ObZ0c6T/gIlM2ymsXATU9YyZ3/VIc2QP2x5h61cmfu9M
RaKFTrP+NGCATuDlsTkwx/X0IlzJ9Tkf8mrdUod3VJOcj17wH1+FmE1BdNci5FLiL7faILKINzKd
VuRZ/2nToO3BLucZtfbmznd6Ouzdwb/GeDrc6/2OMPyeIBQbGMMKb1BRdsWaIj8W8dT2w81v6Z3E
2u6q7jVCArmwOi3c+BNREeAZXqUS/xCWeMXCtj0jJJLS5WKCn1giuMmcY3tRcSjXKcyVzVQvUiRQ
d1sNjDplbfVBdTUVoaDUqGeoGoUPXUqTbNLDW0VW8lsuBE6FbN9jrJbLnhUFUXuZxBevyLuWZuhB
U1ndEpG0pD9ri/R6br88G6ZJu2d9BMK3IO/g1FcgtPA+aYuHIiqBwfHNMlUQ90lbttSGRllQXLf5
yeKeLs8ce1elwi3vO1FAHlH4J73CN+Qble5WQtd5t2XvgVSmUPn8AB9fynXVshJFK0V1M1LNrUGk
u3rXi6rK+Zs6oma2kop0GCOkMrnWo5usoXu6hNAjWfpVizBpPwz/JMQFBK5U9esOlUbZtjMquX2s
bTqJPapcTh403V8nHe3vL2Ccc5kJYmxr3BqsqBj2MDPZaBmbAzdRUmu3oXuFP8FMm1lvbNqhVq70
stwSnYW74l1okIh+gJrLgqswNA3be7s194w5l38RGjzlaFpW/Yf4iVAQzL0cb09VO7/VzC34YGTg
Pt0EWKWFMi9XrheYDT4OebMyyYzfH+tdaIkiEWxkw6qaUoqMR5Mu6fP/W8YLMAGufOaZf7eJip8u
ndo1+Tm0E5O1qN1t5Piy1KnFMgdQUjLsEhHY8aVZz93HKTaTejDLIVZgVLke34IVwcAXrNylOarI
Dp0J7pcsOWhPUGE4aH6N4qo2uUiU8Aq7DpIs6U7/kD/I3j87x+znJF4CWkt6z77wj21cuahlAAvd
MVgDlKTNy1fBXFo7rUuy0ilCQgIpe891AmcjARM59sc615QP7fful4Vnjyj19mKT6ABjpasX9FQY
y+r5CwRugTPFokYo7NxTIjxNBR+3ArukPHnUMDNKWLNlHezobvyhnut/nQGNwVrR3hHFfdnYOOz5
fXSP78y0NxM0gZSqv2RjQJqtyKmf2l9BqObzk1UMhu9bl5t56HOSOoaZdt//aXc6o5witU1V+Ybn
37zXZ7xwYT1EfwbwjdVmjDObQ6Q2ZhaFrjJFWWP+8p9Xbw/y2Ym62lI+oCZcuUztociiMD7jB8yi
7B5cDblkPYpM9kDPXSrjrHaF85LQR3LcpksvVAitxxKUNwtH4FzCV8nVaDohzjf/WOHT+zTeiuxU
T05JVhfnqG2+sRFRC7q7vDwf0hyGJFQ/bPa/hb1L5XhyBNhQniB1EIHC0EaQfxG9J4KDNru5UqC/
s7ANRiMqWT09mVEvGf1TaqtXEH6IyeXKuErVyfphV9QS9m9HkGIriE6QWO7x5BHDY4VGQeSST8Vn
BfWWICeiImPEPNztCiuR4WMEPf6FOAXSqsvK0x26O3GBxdsZhYz28AbZ4aUqxnJMk4jaJk6WS5/L
B6QLty8X6I6f5NdtSKHslR0id2ZEbuYD2jcQz6NsiUp4qqM3L314PuU95j8rJEA3e9/Vl+eOtDYd
YUW+6GxoGXbacWv3CP5c9PzLrLiS+Ggpwmccq3eZJ2A1Xu372MRRlVbI4s3OOgsK/09Qct9Ci0Jw
iNi83dxwQAaN0k4vRG3Igt9uutdcK90N6zFZ1S+P5hL5PGFbErCeMoS/PCD67hVdUl7/DxVukyDw
TEW6iVCvgcLxKul49ra41rt5fwEFQ2XxrzGMisPfz4DDbFi+X5fhr63FoLRgg+0FBBrNuqUDhRxf
tPr2kGzh7JX10ga7BHyg3CgMRmvPvl6qRk1iWmaSVnprjaHhn4qSISZ8Za/r+v0FREfPl+tY8lXT
cH0NvytqGVhergTBdDxVwQoI3tP4zP9nM/XUMnUFhfjO2wMnRDBTcTCpxre5zIrccokNu5ZW2Ksy
q27s5WM1/s9fYd6N54ATgbdePohxZ4XjsBe3me6nHGz1DtnKEazW9E1DcGtiFdkEgs5l4JqEX9GK
J5vk8mEu1/T9EyRF9PGbqjhjNCfgYlUkgciRR18F3oee8YUxacqyY90QoEcBZEL7FAaJx9A9Jt1r
Iq5AmnvYQ3YgYjHxW62IomYUl5aDSI4gIL+B6Ndq0VPQDYPG0wRghqywIqgXPCj9Qt8OvsTgW0m5
/1gAnkC97u/tHTwL+2DbBZzaValb9xRsXTgyCxGk3JiXFJOI7gXAefhdP7rKyhu5srEVs9Hp7Ibq
fNWtwfU4S9SpVd1Wt/SGbF41krErpUau702kQAZai4BZAlYyp6AcTFYpmXyAn2KR13rzCwQOpJup
9NZWiibYMcWZB1+r3SKJzgtebkN13wsXdd23DQ/IovyeM4hkkCitfJw8J3+SsxSAAWa8fChx6DyL
Zui9JLc4MD6RsM0sbdiOIVLRi7nudAvuJqUnmP1fjLFwRVmKrLNWncBJaIXWo8eUAtKQdMciWpD+
uVuEMI2lOSSaSfoRQNvjdqAUAMUsKOBCGoWkRjZikaFQUCVjO5alSMLco4YFqxcdDfZ2NtiwgR3n
7ZusUtFYKV2pcRqgDDwena9xsyFWq7iZN25chDS73DeptgbMYwNgdadbIpAeUm8wD8nJT84NO76U
hBcq4MuXmrWlCNuF6XjHUT0zpXwjNwdSrCP9TnWBpy/wFEn+upIejx97JAMYccTxUe+FtGUcTGxn
0FrSLRSZPJyqkr48+it3i55lzW0QfplIDJuOr3Qj0mPPVWbwHebe/EO+rqcuqeGPmW6z1/bYS1dL
cEEUHp+wUEGcR5QWfP5Mg4lsiZI/F2k+144O90+oOGPUdgib6CcVYYv4/yd+AwROs05PruhBSisb
BVpzEkiyT1TpaiQSEh0QYgienki0wi7Nwx+Wur+JfyYIoOPyX4AqEwwvQDvpafvHvh+MHNqN3Rer
JZwNsZazECF8hJVxodciQd0VrYDGcwvuctnkJrL3ieEyWMnhxPZgNGYiAfP3Dbcf5FLx5QzHTmkb
Kmwgk2mymEaqK5LbJzn8dGeKMeuJOAPL3idGCXjUVGwiGSB5xz9TX9s4qva1sMnfO6BEQ/v/IC05
93LMsIyW8Sum7Y9YrnLtFKjsitZe5VMrSdxfVljgo41cQCvbtqO21l4Of5yy5MKogkURdXazO6mD
ys83Ljoli1QdMQJi0Gy5G53nS+hvPrPj/kLqgbCC41TE0ObSunlVFIo2R8zhfsDXcFTTxFAAMmFg
QA98EwbdlNvxEv93ESmJNu8PYK+zQblKnLZIO6vvqArHe84iS05mvwWomePPcntXxBlocfCLwbRG
CaUTUWAknOnHihm4T3qbr8Ftt2l+rsAa6FxtGyMCMSWhDAszK/DJSe9Bmzov+k+z1qBYktnfBIXq
u9ZevOLi8WmpwlLlFBhy3tY/9RshZiz0FOagU8TKwJEB2OgXEysPOB9IJ9KLQdqVGqDhEqJYbavY
LA0EmKhzPZyV4nqVZZml1xMJQIcJgUgjQIjR+bQTuut+t3VXchQJMYSfegbXk/QYdYUNzMOUKUkk
KAl2YzD8wEh0M3e2JAe2sXL10v1PjQxy8OO6LETRvCPLjH6Z9wWolZ846WTyy/NlRPHFnrD2VAIK
yXX9MIUYzMNSagkxgYEj9xjMk7BTwON0wLvezEsM+aqH80E3dxPVUClOt4YA8gN20Z34sErpyAl0
ZZnY0M11T7FUZloDhOp9IijKtnxnDqJywWO2j9+rNzWoopAkoNG3vqCzaBjcGmNSzCJsQlWGmUOs
njKrtsXb/FjVI6ePbPzsabBtJQGfUkND03p55a+AGMqCga5oVpETenZSh2DqNAMk4qpPHkoUNbJ/
u/UYk5qbxNbP4K3gQDQ/KVeo8j2Y5kfLMEKmeF8XNpRjioAPSWSu21KWV5nStW8bn1VDZLSax1R7
giAmjNSeUa6lquZz1RjX67cMs9oKQzIcrVI/GQaseQFL/r0gXBei5+IL0K+L1BfZnzEuAZnEOu7h
xEzG/e04+UI5uwNUwVvDQkQilywIO6R2nJoc0aBNHlKO9ynpaJzAyH0D6/7bKP53XnvCouGEWvFs
Vq7eqKKYlj3Y2IrLFSq1xlf+1VGOP2XOAdkDYMxbOXPBD9ipALRJRsed389J+jK+9R8FR0g7IlJD
LU0Nu1enifB8fDyupDm7cC5VPyIWE1Y0ntcyrNSXdFeJK2U0oHhhejqNfAvMB0+qnXjEIpHKmKu7
axvZosSQS/PGD4lrqUWrZMSwoA/Ge3Hak0FgFjccHy++OUxYHKnO0Q9MpuZAcHY6+G8SJRxiv/ci
QNGYIRCEaJGVAq7UqBAlL7+pZZqEzl6ifyDLKiaietufcRcuiMIEYAjndO+9vrGzBQ7LNmYa++ME
6ah2RfUu/eMUjpJNkrGXowiuJ6SQxuWk7e9Cos8JCkaP9QvuSHOU+tF0wtjMEuHswYZT0+B5BpHz
RVzYts0SR0HkKE5l6uu3NIwos/KaDFzjooJQXK7yYFnG6Q71bA3QsjPSast4HouwzfJGG/aVGrZp
8txoGT3r0xAETNZf61AEykPio/kechwMqlvpfbxnudUsfSnDHjbVX0T6nToaQmfZAAbOIrPy4Ate
Kgtvhm4o0pqz4HN4dJgkmIzJM/zDgGc1385KW/j2NHxQUEUeNyJ3rzJUdxwYJbugk/akJnpa1Rop
lAr+OqUyk87AR/aKeuwkGdi2sRV4YUdg4v0vQSNWWMhZdP2y3IBeyhM4VzD1mNIsuUoOxZ4UuN2r
q3LkTqf7Nhsps/zBktAk7MD6rh7TL6CrsIxwQKN1r3CdwmSZ/D2r69OtMiZ9RDXUZcIkIukontVF
8DG0fAdOq4spUhE/w3GhwLY9RhnRMlVvKagOAq6LuJ3cbYzBH2aD0EPGZ7pAKZzi1iBndn5yfj0S
IinGEtiibbq7CzRPOJSgagQyErGhrl22dMY5gpNH7w/elc+UWdnApI3LP5ngb6Pzao1B7WHrwrSd
4G/aOAXTt0YJLsddc2hQmONfZA2rRUIBLI7CH+zP46FO+pDQfybJFD68D00D5QCfGL6voWz6nQqw
ZHKh7PjaLgSfmhchl+PJeKfUh7agppbORefRS/85Ov70Lz2XMzuUaGC/IZl5C3tzUnZwyn6rLvFt
zNbBI2A8uiiHAeIwwUBBsZRhw/Voz8g5MojF+DqQXk0GF8mx3BYGhIO2/iffgLh/hGcCbkQPdjJy
g6Z8AZkb7n48QX43BkcCBhJElzZ1sUsnb8JM8eGwCyMjZbLtS3DZAaOljh8MSU4vM6jgJdDOI8nD
eY2XtagCVVdy7y2QltepBHgFP1Tf+frI+0BEF5G0G4vq3AjEYJyydmmKZQ3Ot2KtsTM4Nrb07m2u
jq3zQbwNP+u6pufcyOodmg9XpvfQPwNfPHMpgBWH7zqmYKtIfv3zQQz281dBPMR6RVWhxQgyeA+g
sUxPnTsevGGT2IA3i5TBBUGovyv4qCAYW7omEkOrbvrmDaE5TDEb2cquYoUXxeLLbArQqr8dpnBQ
XLg6g/5ZRiOC5LVTlugy5DWZGL7Kdw1y6ezbHxbKC3VosAYiFDZqtLoG84lSmN5LDXAVBvWMVSwR
i7o6MkpKfj2YBnf0CooEbvwP6uKl6Njx716GrZpnQUaIUL/lXcOw7+CXPsn1oULlvyjTPkND/OF3
tJG5pKsSUzIy/2sAYOE4xQQ3L6IrA8+TFB/ldfdCk1uL0ox3RO5BnsWzw8e06jTxMSkJQaBaDrvS
OseNJJEFPJz3T418HI6agR3gytxiu6XzVo+nv9foFUQCg5o5rh58Hmhj+9aM61WS3Py7fybizN15
YFJuYUEL2KLcMyW9JgggrdwbehbiqVoUCVnwT5OhY9peeLjAWaiqka34k3+qr1U8q06tskJTv8EJ
V6eg/9RxViqOCs/OQ9XIvHiUY3ffTBM2tEYcnTNjJXZcqrLj+cniwAam5QtxozTLwe2HkKDcgKu8
FYmzhJKwIJY+b2zJUYyVD26G02mGaBpKmJM+Rg82Zc+tvOc1gTDVA1zWfnPhO7Nd8LTJaYk4K3AE
EfWiXYTxXed2ckU/JqOUGvH6GK09Yhe1SgoXDwCVBY/hT5BDyjwqH+TETjOQxqtE6XulzHkTYHAT
mvzZv5+sq0DikCpu2kvqFZsxfvJkOsJAJH/7eJfksf2Tv6a6zjvtd041xt0egAeM4J+6HLo+9IK8
IdDz7iE+H3g8UxHw4M4hVlrvUTS2bTwP1JUtRceKd6G1u4/9RxCTEdmhnkPgcDemzn1s1p/HTL8v
aKDhGMThlaTeSdIzMhv21vqd6uNvctOZHBHiwenTYJj41fvpT6kHisquQ8GMb+6XiZyxTQrpqUGf
0jGRj82n8Geh8DCxnywkR4nJRIEMsBZiBw4Lmn0zL13zWStKSVQiiZkSCe2Kcr/buVPTS//2y8LO
dsos8duyegsS7TentSaXnQv8rU7C8Fh39sohJkQiRyzSNiAT7lZ2BoGO0tPxLb9IOXUu+4GxRuvy
0nxx+JdMf+r8Ow+IRwRWgxaacYiXTvabrKq494g3CPs/TrqNrfwjpPPTHxouCj4dWXI1cyxo+8Mi
y6NdrlGbWemMp+F3A8zxGFEioPXa4Ll0f0xLqpNgYp+mq5CtYhrh4wx7+Ah+4S4tCNIXptXMjQ1W
4HxTN1OC1fzG4hoycrazZd3ZGOJkkYwUEPDAO5AyMMibOH6tjka3myDYvix+l0MwHhCsqjTdxo/x
RpGMjEoqwl8g1dPrWswj+aaptR1OIPc8B7cfoiIJdyUllzur10WQwRWwxqtuJNUSuQzHm3BuwRnG
hgtXM3+faM/ZOxzTnErgAGYlcp/vYmgjhzaKHDoYgF6dNUMgTa4+ocJO685OJiIyPtKw06RwFwT0
SPlCjjbl2QnwcZLtr5d+vc1lOKLe5UaDmNt82GN645h1hEDufFwWYWN44ytdUJq0/3Su0GMDRDXN
GzQDSYCKlZ8lekaDl6D/lX5VqMnJYZZp6/vTPQPVnQE08+Am/xo5XadQmafAdOMm5IVYkRlZTd0F
K+mC55Ym+EgzPoeDZt+9ZyTpT81Qm956s1he5QC49eklZUD2uOhqj+1/SLtBhWg3Fh9dRKJ4ziHO
iZRrkZbjlmPi26oCx4OGebgOqEhc6TXDLIabxoebgggnn/hRpSQ3Jc9QXWTytZi9MwL+WugBMldh
BzzRWz1reCXcNEAGqU8iqX92XB4hspErJkqOGHYve7jDAVw4cy8xVwtTdUCqiPSXKk2AvjZJMdk7
Y65HmvTqk7YZ4s6wc7pV4eYTOh6g27CBDwQkg1yO7rX0nV9abhFCLcv4EZ+nCmS41oyZxoZh01JM
pgFP41pcJX+qqnj1rDAJGXM+WP98budiO1mx+OejTHcfwKqzl9r674c7RID0YXzwuZs6Sus0sFhZ
f3QgQQCI2lLhmDT995J7E6j4rR6/bXiL2eYH4uRdXXeITKo6R5209e3q/QZHMpoF+fJx9VFxN+J1
9AdERoG3nRca2g+4wBhnvWC5lpeD7GOuY3GLB8NI2VRnyUoMISPcB8NSeB8EshvCtvZHfoHXwqHR
dNEfsZ61dyWLxw7LJ2nsY6atqOWmhspN45lU4JSSAb4aN38EheWbKfw3YhRG57v7awiKRoITJp0N
B/fpM7Ked3sTGwl9CKfgMTe57DuQS/urqlkjGpUH6AOYvRPp0+l1i+x5G0cZHPCg5R/ibTqduV6L
bop+LJQJPMxi9FfrYDVItvfr8XiIW/fYTf1kJTgFi4tMGdqd6+ImgG6CDlg0rRA682IgkCQkyJ0P
mHdXi/m8mRRXKIffp58G8MXpj+x7EOoxYESyi9aNRYeDqO6WWx8SsVizhli6OgkeMxcW+QexnV/5
nr6Y146SZoFER7GBRFtm35oY392iHe5pYUxbrT+6IWuMXuwB93uNj5x2j8rE8/C/MVrPVcSMhmn0
22gn1iwoqkn/TArxk7zF0Ysez9w/iPLsbQwmKWjNy8cL9PUVIbcZggWaf6I5Z/3nd61s84k7QC6e
IfgvCy1CVbt8Sid0L90pdizq1NS/CYR5R3CA1iUkxP3ivqj/yAmOElSNjd4GnchkalcD6SzDmQT1
97ReDb/hfEj3yislpucVdwQi3wY15FeWh6Nfb5cVaEUiOnbn2AFyA/g1zt0A3qR0oZIywKdl44TB
DUx0U8LaGCL8ucEvYYIMaL1Xs6dHNRStxWiMpfKhIm11YQjo5i/OC/X0wzTC+Z5uONsx6FBCifux
N9dm33b0ZXd2/t/gyddjafWGO3/13eTpx0zD7bKwRNEjh3d421OGL0w/3ywZzvqE7zliY4gLobck
DfC87IZrCmwi1qynlFXDgyI8QW3Zn0fxizBFJq+7n/NA5h56KERoakuPg3OKcEqix1NMyx8+usIY
tatrelYhmkS7LJBrknArpn3aGlZ/pfS6L4W5lgvKf3mEHFiPobD/V7+yKAL3hVUT+G41m7D8ZkdX
MZQYxmaoSQQD36Q/ZktR4khP07OL0/cpu3VQ2aNhbTcb3lY6Hh1m3DFVoHp4URv2nFua5GBLqMPg
b0779wgqfdZgtt3/+EfAdPFJ8cTzi0WFXh0Zl0cpxXh4H47tDcFBsGOyIlmuHQcn4OkySETLIslL
sslynaB7YtEwzc0SY4p7KXkc0Ga0OctyrS4Ass5QtWLlehd2faygicAKmmIS/5QHlc1CC6hl9oBI
YVD+Tzq2mGQ5UYa3wtmPzVG+MzipbywohRifC9eLeakAqrzbcKLh8TxQKi3UCMCIZk/spNnpxUti
uaTZ3imnGUynwScvx+KmM2VDvfqJVNBaN1Lsaoj2oSrhij5GE0K7rHtJ5Rm90nemNu6ulRzj57KC
iwBcdWyKXUskc8Dylc1fboyQ1wSqUWA9CoeklO/rN5uQx4AGGJHwowxxvxZ2CRCwhw9y/vfY6eaQ
FyM32Ugan8iXsi2VW6VELAAUWImdgdshX1sfIRXV3roOjZTTse+wKY+TTC08cHrIdFk+Mpjluz5z
vOKWlXs2jd36J3m9mwe8fB25cNYqf8S1jVKs5zRDADQb61/5ZWhoqDVCK18WetdUGdqn4pNRxx+3
9DnrlF4QlwLMTn3oXscxr+KR8/YYV7jP2DZnro7xx+u5/UooP1FuYFrtZ0ySJuCbQ4ZMKWDhnjLJ
1fJvexhuKGmL33zTEKqPGvA1PspbVBzivCjJNQtg4eMF/1AceJn5Mc6I5jda/USWCF4jpat6jwo2
2M4nVQ8xKGlQ45AzwfLlhEGo5gmNEoqAmB9G9izoRaip9vfwogV6gOVHGRxjuGFoswFlPuWKjnCt
mMnbTrzPAPmCoihW3TRNFv7BFqMYvPEiOu04dN9qpyWEAX7yftKtSAQLjQ0det4K2DHQQ17RjRwg
KLV/1fu2x3rKwdJX2LWs0KF6LDpl4Tkhyd1Ys8DR0MCLMhAsvcIGbHjFNccQGHddYb6EGsEboZGf
8a0Oxyek5ydt17wVrYRCxdXrr0nLgG/25Q94a3Kw/W/T2L4i9wNluQFGDocp6n9V9kdaVvCSxk6S
5FCyEGkt+qUHsQTIYYH35bv4aqFvhvly2ZQ+t/LjqmlNhAQ4tcBbskoOnF9wj4N94gZumzrIT9GQ
PjvTlkCaDZosF4fvTqGVUXJpSlgHyg3IwnQtgcFHCD7B9ffBhzE69U+6uIkRk3w6r+ro+GQZ9qpV
KZDmkfphPGhJDlSDOhUbvKQMgahc1+NHZn2ocAGwYAQTDkESxbUfBveF4Urp5/DlRav3xxTCgaZD
VSA6Q7uV3m8qeUsDuo8X4ICsbARCIWEbYERKfhZH5seJEQrYOnb5sGHM6A7NicJEkoYqUV121a82
tK9Rrf5JH8zMNmfKbxoqenjR0Vnuw0vgtTKACjHN9FDTSGd9wxqOjKzfLljjkiNMF7C/Hq3+ITc7
wQyjvbrk+mh73YCUpXu7UxWdJ1a5JvXbjm1H26jpFF0qVP9l6F0nBiaF6snV+ToT18EuPBaH+YMT
Nf7viJHl6bMMu6OflXnBfbSzdU9oj8lm7UEImv4RDAwEgdxSU/3EJdc3Ymvb4qVdF0l3EDZmtxo/
z6IF0YlGzJYRo88t4hj+LOz77p+rdMiRgdchyC7IZYHVxuL6/DU7XMa71Yq+7WWkFA8FfydeQjpM
mxd2981/G0vtR0bQvWpj7OH7Hzlzg/AWWVl8JuzgbPd35CKf88J4HlDzGX9/fzIxtXfVKpy+DiG2
J3O9BV5a0Nwn5qpfdECWZ6t6gXjgjRxbTr2a/whKB0cDbWz7r/8u9HX1qaPjFT/U3CUMQ5WyoJwR
f4HHs206y1K64+KldfulydwaY7Y1ldVnWVTiqNemluSWbmFiRbZ2m+kLhLPV7wVIDTLLiC/dzglX
FZb2Q5YkD3gmPkGyFpgiBWEVpaB0sBQwikmNiejyazaYMpQeUl1B3Gtcr3vhEUyhnedZfdiBlCyW
HZx+jk5+l7DwEC1GdHqrYwPvIVWlG9Ed2052VjOOAmlicJJPId/aTK17YxfI3SVM+sinAuLHQPls
nyTB1m/PHwhZ20SbDkqsEQAcI8BzmocuIbtm2KKp6z+WMvd/fERw+rnUHYvnbUVo2QQZEkZsn7A9
qniVwoWfeQ6DumAEKAiTEMCAh69ybCega59bJSVNDNxsPnbzocWbW2XnTle24JO7MYBd7atDMD7l
F5oTiKApEVeDXVaytUpJu9ITz9vitBd5h9QEGtDnx7DRnkQifjwzUOMoXz7GPcPaZO4a9ZqOhCQi
3vy4i6yhYfmCuFx78q10DB3i61w/WfgzQcy/Vlh/9IWrSguhTGeDb6V73/3Et7akPhV/GImdoOae
VUhgnXOEfIFnd7A2WMRFljhCMtGrBkhOJC7kXac0MiFY0+F2L1sdF6OeOk2I43Dsbc1Z8LUzQAHx
MoJEJmZYZ+XZOlg9L4yoxmJ3WKjvvWnSjYB9A8ETPTyLfqw0DZwNcAvPHAS/8pGoSROSL/oieA0e
gyvk2s+xrOnTAjOdvdlt14wy5IHVet7JBhV8VV4MDlJ0XFsvuKtD+DJ7JdjbMlrIMhxhsESD0axj
LZxP544Wu/215ogg49Z/mppq9FYv+1Ie68WEQh3p4Gw8epAbs/4/T1wSSzacNPcwbKeKcNg2B/jf
qK+pHFm1+94HZmXwFPxJfb7vxgEPM+YDJb4mDlj+i2pYh20bPP8r4MM3IQEtFm8XrlnPzypc/h8B
y6iqo6zCI8H8OGnTq+FrMKauQgN2wrSZPup8eGLth0oQmh2o4KbkQWv9+vjPduf4z5svtF/zcEZV
CZIGZTq8bYzZx3ybKImMb8AJdEtrS9opiCPQIeC05N20HVNhgUzZf9oeoDgDQJ3iTxtVgsagremq
YsGV+YZp7TkcwqvrXUGSAvfGqxvBSgvy205vWnNIo5nZBPu1K3mCfl5PvlrnVVH0hiunH1u11SPu
cvDjdzdsBgkExlQ2KOWaUwOmXr9Luzq7V7iUEz346VGF8QsJYn7cULkARmqVH648Sl94NZer3h0l
HcBHTSPW+sTDiaHSux9n1rlMYUNqBhEzarnWilbCCHzzhzxymk9yn5K8prxjP+9O0tQH3/vRexxG
hDdSJvbbGHG4WVGy7JtlApNG1UUWMLH8rgebjYt3Oss098ZS1RLAJLki/iE4wKni+MChnk8TTzvW
AjxuEogbWgBUBdBlNUlEt0WAkNynPQ6YNzQR3E9YAMGzR6cEADLyndZ3959JZs0Z5g+jJRm3zFY8
QblWfowncEdAeh25tAzI6phfTwggYR/UaZ+/Le1LRf56ITc4b/jtKkPqtkBLxIqreriwmNjvoLLq
kFPca9dKV0nYukNne41vqTKNzq2KvH2rZ+vvfs5epbgpfhHzeS0/ZmAMQkdPfeeEDn8/4bxvZ4Rx
EC6rYg0RcM5f4xyV/Cl3fNjAiNv4mphmPAWQLapXA9pdN4kmv/gd0T+jazNoZljF1wO526AHXpJD
4NivLVfcnZ7oa5D2DO3D4ZhtKFC/c85/1iYTDd2bqJUoc4mPFa26qGyIE70pHLHK4FkdBewZZLsL
JSJHyi6+DDjYGaGZs+j8agoD7c7hpIodPp4HjdBqnR1MGg9lQpKWYqxgQD6GSm7JiEFqrTkdkcbu
lAh9GFnpI8GNZejmdrkYvI0EAl44ecSATL6tZNGNphZqswh+77fb9RW7d3GaZ5p1SmfxKkT0marL
d9k/FE1eFfcwBNLhjY60Fprr+qA4OtkNUN5BC+DVoT5VJQLpfyTEwNIYTO8OtAXJFUKtGpGwFYK/
9Mzof/qHaVoVSzudnyiNy5F3BQtPMSkoYjLq3i1wYX5dVmIfI/neIenFaNxOIcnC7O5VUgCXnv62
hAyrRpcNOliz6Qm+2tSAxZpWjc8IuQtC0NtkEkRGUemwsDGhOuzfE+pV/V2w4oplMPA8klUuXsrT
CQ4bOr9FuhaK47Ga3Q6gHytJYTDHUeLZ8TU6iQ4GDMFt/tWzzBgkCQ9hliTC/cvVDZNxae8Qe/Vg
UDpmq+1ttt+tK+vhpvxh3lLc5jI4rlglbWGytibs8A0MMyHZ7MrmnU8Fz88FTQjZepEqhez7gDTr
PjWcsryBPY0OE6Gz88gWAUnyxtKzpay+AeV5MLM2SNk2VXaIZ7qpjXGucpLo5dYKNipxDshx25Ky
+hDX0n7+HhQtae8HrnZNXJ4Vc0zJuw2bs+jCRjrRfkzMfk5f5ZeQCipUBtTgFgIVpeFQE8XYY9ti
8Jk8QD/kB+BQOh85k0HILffUlmeXzUDKC9kTKg0UmailjSWYXJujmXoDSZA10pAmdJ6L55iDQVif
JZAPS7pl4air/HT9rWa5waJIUTyHfoEK4uut92H/azhBzJt91Ea6ygXfsftqXUtSVcsbBEUT+Uk7
KmcPMSCdc1cjA4rmRiT1n79nEsE4xswf4v0B0ofVglzwMcnO7n6eSvKY4MtU7uDHGDsqvOs6k4O5
4dct8NfGZRsUUhl4Q9uacf8xuD54kMbmXvOwoV7Lg/Z7/u7MCkyvgkFL0qmPjZFLqTCnHC0aGPxT
iCUcCKDSttGOXdrZ0lVGOTdCPxBvdEd0UmTbvCkXBdqX/mkAEcv4PX7t8fg7X+q1fw2rKLj2g0Xh
Mk+otvshA0OSl0w6gob1yiXjnVuwX8oSG4ZKBfmxuQXPPyu7kj6ew3yQHiZP9BYUv5IaOxy2AUvv
+NHFoJFfNo3bqIfaupnPJGLD+ZkSfgHz06LqhI9hUwmwmErZVmEYaCpljspTtO4PVgOHJH8jktRW
9NfdOUHbCaLag7VZe29prQC79T/lbWlI8lqSwSj9T6bYrWj1rW+t2QCJbQ5tla/sEPzdrq6D9yy7
tXji49wcy7jxc4alDY7kbAbdRhK88y8S6+eJk7ijK219Ev2le4bWMF3o5oUvDLc/E3FuhRAuUaJ6
R8g/6BbYE8RucL/GP1pbTGDNcYryiQxowrTEhcr6dyccDv1FRkSFGz/Mp0QA51tjAXXxGrDFRakt
dAfsawUtVeLEeLdaPrfsQ2lXyi/IsPfAE5QIPAX8AOdjMXcYAwaSa0H/ZdqutBK+GKWfpr3ZPIGG
4+0B6RL4lhbOjkKsRdeS9DgUR1tBuD+pkLBSGoHN/HUOk1iMxVPYf42D2wUKRGt8IwpzO8fCuYF7
p0EoJ0E/HKyEPtpCAgmzTP4fQ0aKzA5/eJiBl/WLDVSPtuB72zbt0Hz1eeWbckQZOsljf2HfM/Lz
yymnXtVNFoyoeFgHpH1lRfKC5XiY70xlfqN7RSH88c8uynwd6lguMfyhE1cp5qDWQATgpaBiqE59
Uo6KCzv1+/gUenM9U3jQUFpsv2dYxFk5ovq79tovnKYqDu+KIBSjL8h3oAKu1zD6FiKqEue84XgD
H8MJXA1gvXQ4F97cLG8a/55mNilr2nPcRkCOXE2G9lEHGYciPsmZIC/dw8vViQu+kvj+N5c0ZtHY
R82Wo7EnD4Yfb9KPy/+liMr+s2oBNrdd4WuBvYdvx+3vhlsmjDstGPfTo5GynWBcnJNE/qChSc7W
3LGyRK8wZX1S+dGYa4MO8SO/QIpAd6HY9rYD7DIOfJR1LmheYh/iP438RZCyuW70d8PWFhCVgoNA
VGPjxnpIaPIhzm2Xy/G5D290WtAYq0MdEPgd1voMI+SX85aayoS1wRfvCcN+n3dGN6QN8EL8qLaH
IsK3JLP20DfA9P5feWahtTHPBWGnHR963/Ibk0xpQdRLDMH0L8QcxqAq8rn8SWgjZbz2Fc2ttGhy
bcX6MImleNK8c7rfeIcJuH96bFM+U2r5T/cx/hc7Qcf0oRY4ndzFa/fRJ2873hCJJF/V4AoFFyGe
AP8efoDfXG8BTZn2MKZNkvCZUe+Y8/wuM45Uh0/tfjNoK7XeDzkCNdqS53/oisT1jmsCTMPHODni
BI7ervO/BuEDF1Zu582IGvNuo2sjLMWG3EUXNsYFpEu2MJxeLXsHwD66F/scBwxxjLZ3IpyKbWAy
vxz3Cb+iExcn4EqYLqqfePchl2Z4zhVTb9MHzN/CjZQNHnzF0fQijp7xawJzS/PlPtWntn7hf6HV
MCCTAWw+XzZgKLfWI1VaoGXq4OCVlxCQ5tz7X2AJyfu98AbXvl6R3VP+qLDjwGYNTOd6dJ/x8hHm
EIR3KdAsPqUiYenBKbbRnLdsu2OCgB6RTTWv2WgzeAamGNxsgAsbMmDdIH3j7MISckffcYR4ECpf
EsPKKY/K6rTSpeZ0/SyPhDxRH9y49DKmjoOnqjPKdY4OuHsVdeICnhjFrLnLlj79QhiX20U6yb9V
W1dth8SmXyNRucKjgWdCL5zCg1MDb4XsS2KxBzY+GZv7Oik2dYQ0YAykt5jCMiO95m8kP5eAT6wi
/r4xZ+IFD0y62egvkuERlRssapJhd56VEs1WVdPAMEnIbScY+Z0sIN+Zoo6kpIwmIoMDz5qxkoRL
nE1i1xtwP0y213LXGXLgv8Rkp0p1imrbRlnBGo1ciALB6eVJ3DmY5UOvJe9mj3ceW7TPxCIx6Kto
Pqr3ElAjirRKu38RL17WnFwE1ulUjLduF7uii8fd6mYwUjTr1UaKxlFWegb+UXqyUm/OiInOhate
5Wv5HK2zTHUYpj+gsskIAp1v6k40h0sTPxwwD9yOdYS+0mV/FiOmGCyOOX1b+VtSc0E42EIyyXp5
STs8GfIQ36hcLdrP/70PBne/TKO9/7BP74o9niOx+ZPNcy4hGngWObiqCmPYX4nqWLWpW6bIEzQj
dhEDu54TshlmVBJOq/MGzTlb8OYiYr70ctk5rvWmjsOJautyG9H3/xb+CNWTucPDjcSdoM4efftb
6sbvfxPwIvgSelCGnOOMJ/3tfuU24q/qFHRaX6blUyoZFqOL4AlxFDjcMdvX/9viFPkrETiMYzLM
Lwzc3WZZvxsXhb5tBrXZ/lUc6WPFy0T6J/An0GJpVax7VzJWinsNpcd1EHyz3xOxbQeCIThbYTir
nQ9sW7GGAi5mwexvG34UDwgUGzes3oLN1luvrmxwpfC2Mo1TNcky25aN63Msa5Xqxn5fwycfkLdZ
yJv/MzDbCpBMT9t6SL7DBPBV+N9fNtbsde7DtWjuOyqaQWAlGkPMlhZMct3elLaApcv2V8y0Pi0W
katpkhSFngHGkb4EvjVtHf/ZVV4fU9rF2rGoYP4Ry1VtK3GVrWGeDmQ8vDvAxvBtR2u6FwQdWcHw
4BbuRnjWmLpZ072zbwb3C2bfThpI5uQPgzMIZmq8ZT0AavfraYovn7wJq4k/1egpwUnDaWYpsIqK
zgo+f9JwI6fHWMp0lLYjtHVQ9WzdIloA4EuqgmIRU4QEyzwQdTEfdPkg0mI3nwYUCU3CXMaK+Lh1
b6EU2OpA7mjapFKhy7wb4ZKsI+XDCiqeY/Q4KVXLeHepebhEqIVFjKnL3YIbzLnAMJoKhKCY5Z8t
gAjFTrQX6UZhNCfU7viAlKnrJ5ohdUF2rn71N2tLyWR/NxIqZ5CMOL6LsTHFfhZffK/aFkGeY/Qm
HEiV202DdpH2z+02PPXivlh9WGZIe409GObDVc7nCAgg//b1bPUxQsfDAFt16NzH6LYmd2J8bzDJ
apXmMaYxc8VOmRGYunrazHgQWXisKBnbsdOYIcnKz9PpcmAQz1aE8e5hgf5eJS73X4EkL58d2Hvn
Jg6eHdI7Rd1OVecMqFyobf5xB3kr4guheLbW483D6MPFDH74XhG2yJlpgqqaJpeu5KAw+1SPi9bc
/1g1AE3NbooQpeeG8d9y4EsZyJ+gtyy1jsiLXSzY71EcphFdC635FmP7iSOiv3FlTWfp6ICSBSP/
ZbVshX3NOsy5LEEGKInJuCzpgTtwg4xWQZ/8j77DfE3XqMEASSiEo55vbdpplIisa5u2zu8CZb9y
4oQR9YYVM6CdoSyDniIJLWgzo3Aj1Ytup0mZ0w1v1QaOwdW2GlHqpesDxvdQiqyJJTkIZeTYVplq
WtpDfh91CExWrBbu1a/VCgbBcwVhJtQLLdGcnnEpz8+ZU5G+pazNmh+gzy+LPpXlNSUjB8rwDprL
eF+p0Sg6gxRP/RE0PC5O0/6FiaatcJF7LPEXV+9r9LED8vYPOv2l4yeyF+C+My1Vmv7e08UdWKRp
9E4EtzCJ6f9ZxLpCtXQauA6RynyOlGx0j2s8X/NvyGttn4p3ozLhviGcNzYgp+uXK5I9rcpG0Lhw
87ZZnbbEWTSiLEKsbZ2xr0PcIBiTMMd6bxvS0GCCO/1DaP6KjxjA9otcVZ/h5JeliWG168OHHwX7
TObQvHUJ2m/BHlI7UPzHXTXyT2O7JBtbK2dKEnD4/c2Bs6Mb9faqnLGu3YDBFwt8o0rqnP9cAIG2
hOu88TOhwrZ+hTsPcLU6OmOpbFCvS07cVwbeTKkrXsHWEf6jbeV/PyXWWjrMWK7aavslezxLgk9I
1D1jH+lPGvUr87u7N6I2mhDYlYYHUMwzkz0CD8AXLrQdQnRTHddRZFimRHNytu2p0riGvQnUiysq
4tXQE8Leeqe8m3ta70TXC/RIcYyxWKJ5rUtictmGDtzN8FVCb9IHWjDKLZ4zW7m0t1ooGdpTPXl0
4Fx97nDe+pVC788J0P0NgDKlwAzLc1N8x5EHTFnk2gA5P+93VDRddU9tNDIwuycCEFhsNQEtxodR
fnHxOu6sOUNda+PN5C1Vl03oRDx5kC/JRGv6EWjlHnUkN5nSy1pxmUTLsjCBCScUBI6xiEWwgFDR
UxEeO/qhbiEkSY+Cky3rl/8YNlHnzvBPSKj5X0K9NlPALtZ1JV7FqFz+LbaCIGe9jTKAGVP6xENj
XJke4WvPSo+XqlgUoSQegBAt8YWM3Em6CyAx+im6XsoHDYHUuk/Yzz0M4Ud4jEdf1utHO/0FXgrc
VPfmHApeMfEmJD9xVFka15JDfhyMiEJdI+6hDpTsZBIT3dMYUMjUe33Gq9gDxJgrQUxyE39IIcv5
Yc+ZWf6kgjGncD4/YQGIzQFGzDHt5Pbg3yWlPzt7qA9e5oyZGF/wrowKRaZzIUGC01AvKc1VcTxw
h5mo6VjWlgTzdZr7suQ3p+msxWyQCtWiG5KL2EmB5OzkIiz5A86A5IB4Mve9xYxJ/q39kf91XA3d
vnoTI0D33FdxO4c2xzEZpZlJpOr9hUlCoIiFe/9WvzARY2rvmv0FuOP78UrCReg4UOZ9NINo29Rk
FggCTbCQ2I/+wGig7hP3mRnMIA4IvqSX1HUwTPDwu7g5+O7Wnl/xeFyBRDHKog9a1//KeR7Uel9N
j79aeexcqirpYij6oXimHvbjR8iw6NOHcOD2YeNULXwFs2t+t5L5KKe4ZmwAYKKBr90wLUzvXXOx
jamxKITixCIt3E06hKUgzBkP3EYZ65HcMYSn8fZvL2lo+HDosWefWoAtERD1M2X4S43J65n/jU5B
vn+P5ILNpEbg4x5ixQdfAGYOxCq6RorUYKYxTR6NcapmYcWpClizqz0nic7ZzZJKKvnzkJ61utYI
VWi8WNY1Y11+gKz5JrC42bF8mmk6hKKwX0j101r9qfymOSaJjfcUrkLXGWtwLO1FOoFF6W3/6tcN
h+ly0eHUAxvPpv8Uei5rKSyhCeGodky13B5KSoCtobhphm7/miyaAnyoFzzj4edRd1+dbI3WLbkq
jvzRV3BZEgFBTIuF+WzXWXO4Mry9wW/OH0sE5Po1/zsHk1B9EZTtFV5frDxpg7KXobsrpoCS+8nl
WxnR7CL/SSzFQZ9iAlo+4pkwwjk+/j+jUuEMCisODTZMkfq7hdD4aCi+xwrlRBGX1ItuH3LboJmg
I3cIHXqu1w7JZ7pF0t3olWyJCd7xX3Qz6Nu5JRYKbAsl9hgyG7nlMmMb8QkRgjnT5lHGyb1u8lkB
WlvU5RCSb0vCXC5N5s94P9CqIeuxhwaXIsmD5MnpSr4K3RhcI5nTxQSMzLoO+lJMj8w+QAL0rxbz
KU3rx1BU2nZ8qJ+jPuMIcd5QcBsY1jmWSRIB780k5vGkwS4tm82YgekUDwkWEXBpfGBfdGODNw7/
qZ1N4ka1wW+5tYWwZi7v9aSshKyuTocfciQ4Rzi7JFNYmFZ0XZs751hYlOroci8Lmv7j4lnAQH0Z
OqPCCtQDV3iPf037JI/laI0KaR25y1hnDxqbtmlhsWxX7HCXu4zDJKrbcZW6xUNh11eeNwbdzCJM
VW3tNC8rfioAKnXeaJXoPATg7KAMrwapn+MoP3xlH+KztYioglofqH2RmdXeSXx6Xr5PcWEMuQeD
U+oRM3S9ziHU2qA+bexTIwp7enoQRqGH7VGSw3uOQbUKq4Thl09IrmVit7e8kwK9whXMFKzY0Jp8
cD6Xt431thgL/59gc8PhY+zaqIe7/GWpFcSgZvv3AXmMG5IM2534SuThB0vOzSBVfBHdezYHAxxx
uwG0IIm1ijLziXXvbMlBJR4iqBdvr9OBmXwEHVXe7Zz1OE9qRi9zrfjOhPf/fRBQS6EObU8SWvps
e/ZC6DnXR8MYf3ZaRPkbQmwmtmRpo63bRt1l3QRpiEZphMNOrVBROtvYYSsBAFj/BqvwuN9Itgc5
pc+FUV70aUpa7VJkKCqaLK8woEb7aFJ/8frgjDRADGAUWrt9Aor8FUuzNFWDoUe2TD2tQJxlD9es
UncZ9QH2DXbyMsYAdtcvqZnZGdwwR6M61kMRrK2PsXEwjgLD6dtH/TtAwDH1g09ypjpKK8bINHpZ
O6dWALPQb4UhkTXWDNe8PhZV2o9H0Rx1Mxl7KQ2N2Qlyl/ugTS0eq5Lm+rJOXVRYt+kKSzTYQurE
zjZo93n93bwwR8ydPMPtf1fz1ISrefhFEq0T/h357fMVmWRcCJ8DiiEDCLGdaF7PM2jf1ItfGSaS
d6IWpNVjN4UaHj6cjMsKj/PgTk58AgfF3QLewSsHF494LX+1Okh4dUVo4636zgbAn3nipNxtQ8qW
+a7Ci+DH9CpKK6r+WEsmr0C7I5DUY4gcC21hZWMmt/2sq3JiJwki+OUQfgju6XkcEGCk0gwcz6UR
NRMzW5K5PAa5RQ5Esw//Jt4pg9gxDZ5IrB/kVhI9pdsgAIohKecJPD/LsOzF+5ga7CH7iY5shuW6
lCJh6GFq+1SnUPe7AwG09Xycr7hTc+S7Sj0f98RfUgOrPnt+Tb9yb5Pr6Vy9yUHuqPN0QU1I1/Dt
6z5ztAvT3eWRfS2IyF+y5I7VWpWWzASphO0uwUqJz9KJSMpYEw0/KQm95eVh86VLtSiDMwU2YkFE
TQwIBv3j92JOtNtxg8fSYYXE7fr6qxQzLe0PyegdK00oeDhvYjibSaa1tYEP1e0XXEzvjtxmTunU
OdyzjadZJ0TPjdPy1S11GYrqBgew4gblmD4jRfUFzRtsVFUSkMHVeNxnw0cAY1pmzYhf3a0N79Sl
KUTbsHS1ecKJzDiOVAabHGwhMNJxrHhSfCeJ9IxTrLKIFXVNvkB579xBlm/Qxh2LkFTnekbskzRP
DMxsG1K9knFe4W1JMG375DAzjyTeo2gdfFqrMVJ+VfpMK1+NfrgZBmOAlCxZh+qm61qqza777eoj
4F6ycmmjIkuLomYUHv1aBjtP5Zj5Q0+ETnomrPz1sf08YzRDujLejzn+C6kEmfqcPZpAvDbH8inz
tykDaAH8qOuztnIHNYnkWrT0KRTQJmTosKViFmOlwnV8i63nX5qv+3dA3whoYLq5U5SURW9P74+e
Q3U/lJJk4pdf61I0ii1vNnH2rCUzenhKPxEUJAqVZi2Hf0pAugeaRoH9BGXoMhf5tzGdJytgyAOI
1NhEzi2+d9bVHy6/BE8pJb4T5ivPYHxy0xrpjijsYZmtuZxYubvOqV3LzaCQY4y8iOdd5mP0oUif
AnR6KqyB7hzOkZkJF8MUSEMe9WaClUmdV8cKTZ+h64rBYimveKcWWTcirRhmO86YhHmWYPejD/56
r4cFhiDrlu5Aocrtks3psAu8SixZpfbuFqotBBtkZsFM6xzV2UDTnLMSLKDw337YSx8cdBmRhd0s
Zuwdnv7S3OeJcciNL4dtBvWORUHhbF2InGUWCdO/ia0gEIoJo/T9RQOpvLl646t1LxGAb9vzQmtW
Z+PN4O1LC153xvBWF1GVvRkCOhuXyzE3BrcHmbuyMkvEBd7dvojIxGvGGLdtQ7eYJai2baEMiPyW
dt1iHso5jf//1skhZ/Pao+EypCakumP8sErGYX4iCCvWVAdJzOL22bRuZpIph4UqYU1dRXEU8+U1
mqyMAqyDUV69ZKjGphOqTvbb9Gy+dYk/u8lB2+4Ak9B/netT6rUC3SnM7uzs3TRbSPq184PcoL6m
zyPSo/dzKBU1Je9/YuG+c9D8cZwVpyeBlyIkZTRlbKX3w3/4+4N2Cku9Z+KGwxNQhN9qzg8CBGrk
SNQCUneJ6JequRyTHEp8p+vyCGz4sikAm3Lq6MikGOa4LUK0fOvAUmtBDaSHoGH+vCY5zp+tkMP5
krdHIJSFLfA+BUvG+rItXLc55WBFRIbpLJC/05L8MUlfaE/2NaJnlQt77lV9axqLXrR0r2M/5QRE
NtPp/+Xbv96Is03XG82AkpwyHom8Shrbm2V1MrkXb0Njexf86YeghFPXmp8AtW3Ajts54NutYEeM
q6X7yaQAjpMW0IpHbmd8jYvE7t9JCrVwq4a7nFiMoDD0cLN3XyGsVurye+VuYZWAwEJ1PTk+BsU3
0kqymcKcIYuDSmEXHnXyApdOxf4qaLx5+90SEaz4H+i0fnndUiYWB3PSv76sKKD3gU9fpKWbkmT7
7fXKnDxQykqRr8vbfC0YSmJGC3Qede+aPNhPlToOhXFxw9ProjabeVpVuyVL8Fm9ElUvVIY2WiEe
LI8J2Zysu9bX9IYnncDx0NtZklT6X9jBPS2VCK7FCK/OV85j0x+JyG3mq0itUgeMCAa32chyTKt9
Aj0qKzXNgf6ZSMgKHQgWd5a6kkvZvUrIIx5/NXyJn/9IByWNUmWQgKKMOBsbXDCUAvXiAFjdFXBi
2nbuFhOkY4eOZZAkccVNeuCNMo9o9SfcfrbpyyWqIoy+B+rLQa80wS0kDAPBKozSXvGdmmyHaL8G
V9U8azgv+Bdn34bjnGenoFCGxulEPqTjujSdrZhMoGvEPSR8Z+ios2Sc3wcWYZwmjKRzA8DG+gYI
fRttHpSE6EyHWlUUrwyREornA2kSTZXv0M3Q5KeKGw3q5L+Sw3LZUwxWBnrzFELSbxrzyXuGBs8/
ojYYBD1jfDtZ2o7dcxPHWjt83/rxnoA+nzYyovKUczU0yAhkCZAqKDEkO/Xf7bFTK2curvTOneaR
21mzfMRXEZ7qff7xuKxH+Kh6/kaKQFj5fGMgtYPS2kgShLkxqmUA3TRk0apVmgrEY/rvOOZwhQ7P
Eywv6luif8jqWvghlhltyhXldXnwu32+Xui7IILdcR/IJlhjiw6X6lms0vb4+dh/evSn3YS6qHJf
x8uq2/8g0jNMlPBvZlDS+r+HfH+kW3srQ954RE/EAQdgPitW0YC/1ixd7qnnTJArgcKdusi+dRKC
Bs9SVRdT+dG+lg/jThqwIfwW/vloUBdLvo4huM74ozVyHGcTcAR9pJfM/NNl9/qT99YhxI1IcRxT
+fU0Py2zW8uK9E+R6QrtMbP+L+spLZrSdAaD8hV/H3cNIQJuqZbvbtckabi+GBNJEx6pN56Wckqy
8AOR2qGI/R2p5gcE3L5LFnrD91qIEHOFbrs3Q0MZxMmqF+V8l7wWBe82yAyKnGJjF2fuL2/S9cEN
cjqnE/ajzRdn55iCc1BH3mz8f7vDvlFmYjJ8bJ+8lVKtpCt7bzv/WOALCa4fbNGyPMG8f13Nj1fA
NPlamwWHGEEP30tNVaPDr3hvaiPUV/8iLvbvavt+iPNaKxZOWZ2Q6jHzwjfhL4XRG68+BNGAgNXd
/NG1rTTxZGpTZEQHcAj6m8htvXz3B+g/OtXVb7k0IMCK4j0lDfOziYxhTqkMWp4eD06o8XLw4Pt1
jUkBSKZK4tXBqZSqp5/5tqNK0R2zUzJoBmUUT45pC1cPpwZfTo6gdK1ZXB7FFGwlWZCtbXzc14RD
pvPZf2ZEGqyyUrtUYF7IzrJTJwQGNhue1vhFcApkVgHzWmSibTDB8iK89B2v9G5ewZvgyeW56bvp
PAFuqSIpui9PA5Gazlx6NOOzI322s5/4pwRB45goVDh4wwvN/FO6RvOcGemRgNP6pxQxsnbc/4if
9OGTEHtGXdoHx5LDEI87ej3Sgq7gA7rYKlhFwP825kaMwQJJVqmT953mevHUL+4bi8/zV1of6/wA
rb4/tyyWREkoCHe8L3QF0wJCohWINW+/Qyqqvmw0sDtMUwC4XmbkhxUq1GYxaK0rmkHuufajnxwy
T9RBeBGqCWnbAE6+Trml9CZtcKoYJq0Knsr/y4U7VTjHLpqH7ZKWa/WsUlSqbpLNGLCwPvWW78qn
Jl0TDyBVPb9jgkJtFWR609QpWGG/Zz9wfPrcfxpX0xwWt7xfOcey02grQgKG76l+RvLUjkYSbqjl
W3fycUUQxD3ackL5zpxiL1lTgZKxg9SUlPUjlSpfVvwj3GfOeL/ZbxVusvB5UGYJpc7h3zJzTFUh
xG4SxxXPQqgPZc5+oROug35QicrVFOwjUbqd5Eb1HTmQ04SOdscgLvbnjjWtUpoT2O/RFH9wolaG
MkNovEUreNOiTvW2ey5JX/xhPJF41QlH9wcAB49QE0q/YJWe/XH9F1+FrIfT7WcKSMGIs9aMQRIQ
K+I7GLVfDrNusPSwE/eYazwWzcW/wKU09wcYNRykiJRSwxg5ZVTJR1o3Itf7R0trbH6TfuxgZNVz
e8GN0p07M4kshrKH9SaqVKVRepxJ24ZnA/FNZoC3vheFEvsDEJ14+W8up4LeiMvL/QssUQtNNtqZ
EKmwG0oxcYtJUhO3ibVET8q19RjxkbET8dVbXjabsu9dJo7VUIiwmpONwQm9Pi7q7l8GEVRl0hzE
8TFdhRXA/iyE488pbq94awdLqDQpenhznIiXfWjgBgAqXoxyEOi+LkjsJxu4DmI36BIAb2xoVDol
UFiNrnCyxnvyrGEajvZGZxmJnMJscxBuyyXuzNtHA8hExE22k92emvq+rE+ZTltgVc6vQSvVJohZ
+6oZFWXQDxobIgMfMPucB3Mjx5GqFG0F4QwCUnXvTMu6HEEtZIBR6daY7sK1WYFs7gcASNvRqQnW
rZWKsJ0v9Tf5GUoVjFbT/sKVcX7SQKlWsb4tqDiUlRjp7OJUSTglItKVP637Iaq0Ew6w1bBn0zl9
zYG6AnrM/W7mo9d5QTLjPfaofvqMjmtbjMzQsQkyS+yh/IY0cZcL+0AzoYIisnDn760tuuwDT5/6
Umw3OAs7ToUkgvgx2A4VeiWua5Ga0/rY9TFUPzQiel58anL9FkPtoN+Btt23Sg2Km18d2S2qiMTE
f8pFMbphQI7Krh6iHTp+xNg5VGU5rf/6OiKsQqQH3qXDUd4V5uNUHvGxfwvUfyEHmnyDEEMC8iou
KjaCWHHXCWUqw88GJNFlUFJ4zHrLqtFgVJjxc9gontP+Uv//zLijz5+XuPic1kwQeSiLualMURrC
zdzWCotZoQ8lwE1FunNvxbA5ss2yo0iBlR+IDw7JegCZov8TA9KStxxUt5hn87Gwjia0w87gGXGh
+5UrjYDwaQWFJiIMbSakgJ8AYXYJlXYllr3mMYWHTS6wWn0ItzOTABAg8+jkkB5Erm1FzzTG1TiL
w4xHLdrGE9dbV45DY1SuUGPZMjaZ+W2lE2VBK5xw8fiitIuXSf9sYfvxRgMlRlEGLPCYyM5G10Av
WaoTJJk4954E2LpEESEq6gvjWD2K3Rllya7o35eLWa6HQoTRTOGoFLlfs1/74BI5nEH3aD2j1/7z
RUjhnHWKzLaM5339O+fd7YPUowjYKq0b9ALtURt3n/pxDAP7O24ZBaOh6W9I+zeH8HgCsfhs4YqH
KW8NwfdhSU+CE5TZZKoSqomFbyT6gva80GKKlvcSmx7/PuH06coTKv8nPaftrAY98Lgs48kz/1O9
ZOCOWTQsb59ITdea0WHrDW3YaDKISQCOaIaqpZnYbLkzu1fe4r8TkSA3G6CHEoiJ5l2VeNx95DUd
iO75LQwIuLMym7/17W5r8MXvRIAEGMN6YXoxOHHPjCX20lNZKfpJNeKvnDMTFzdCgwG5y4dlUdqq
XMjFL/ovdEWvAKqfAQicuIUz5eJIMrDz4eH/Tpgan0PtXp4+avfKawgQHdZGf5rIWSTrmSItTpA5
SA9IOIAD+vs+ViuXPl8CRqlaUqQWJnjhyc5+Li6U3O4Jh6wFeUUd8CcYeko4uopumYxVSj7D3zEt
daZJSZqbHZOXN+gWC9y6LIUXcMkiE/csby9PDyy/KsAb8td3N9qVqMwTJY3RMhZebxM4b4rIQEve
WDYr4DJQtmdvPfXNlyfyk0R3booeKPkIlkfMnrvtqx0fqDR3P1pOIUO7sPfQTRGq9mVquirz/pRZ
lIKNn0fKy9utmYPHMvnsmRx+c3tocJ30WFCvB1hH46LqmIphpOSg+CqaTOqdAUnBL9XAGOuO1ITg
nyAQDR4pyCz2V12EAEmtDhAHWLe5UxXgFSUnWa2Mfy8ckcL5FhaTVF83F0hxdYanD6hdr8JixwNs
x8pYUPVfiqw1mHuXZi5JIAxrVqcnHUnSdVl+VpSQQypwkgdQ1Z8QBYGzPB9ijPgJCzNAfXqnnjG7
02Gl7YNA9AbvAebSRWS3AgBwQvtQOpObJm1IP+mgIyguWylyGi+AwrssSPhp+MZT8q/VeWblLj6w
j/8NEez8T94+tT0HweoS1oid29BAZuWnwB3fcdFIdqupqPNCdGV+J1870nHKWXQNdu2GkkwUGfdp
gSq1FvyV05T81I/ywStnUxMH+uGc4L+l2ViAA1dJaSLp4gFjPlDY3Cfh16CdNg+TxGZSfg2/xXEU
Dde6IUITLyNzgKlOcUV6LUgpKC2A2JNObsO3B4Zdxu+W5g5Gy5/g6N7S9KCN0L5nZ1HVABXAU3RP
vYzmBUnWuL5pDZDJgF1VybPesSflqhd+99m5aQ7zO5JQGNLY9oHh/HbjZOAVboQ+tR9x8FKRrRmq
cQJMQK1QUui3LVMdUkptu5pN/lbLbItht2L9Bb1hHfx5v0FHu97lXTkQItDwMOmQaoPpDi+R7aot
kj9kc29sfP8x7aRH/a8/0OW/2BFBjA3W9zxHyFVSH+Y3D7J1Qa/VUij87XzLJw1DAOTHbdRefz6l
sb6IQuYO5BOaoYXvyXU+2ycHDLkED6kzVwraK/Gebvf14nM32EyayoF+FeUUfHxI+CsDuyQKDhAK
S/bPlKbpOdrxrkqr8A0HrQnGNp1KQ8p1P7kBLSBxvSUZLPEaZKW4sgONMdtbVan76izbPgGc7+Ok
pjyTSdpxSGrhQo7lrl668jxMS53JCL77TZ3p6dzQkktjDo/suuPSbOehoqoQ66OjU9Qbjb1yU67m
z7df5cIsETlhqgJAA6bOUt3eS3lyA40Etp+LsDPAOlVs2MAGqo+46qEn+EUnIkvY5dIhQo8mIaWa
k/6HKkpKAaml1d/fJHp7jXojCLRdVv4LGVzdPbucBA/t9D2Y1llrpuUlg28WGwc8hse8bbfVR4sC
k4d6bhj3Ca4SGQeAi4nrdNnu9b+U2aor5TWZthXXBlB6GAL1Oxt5jC7twq1tjB1pdQXqDy1pq8n2
4gIwn110lUvoWL/JhKfXhE5Vipogp3wJqE61sybPse8iwW03A184oPuUGkwZCGNM8cNH3I/oQAZu
6uq4tuxEvmkDqDV5QBvzIWmzVMRnn8E8bFUPYvJwPRjBn41WmVtzWbu6e/DxBfMf81D89Uh7MnKV
i/DMjyMFP7JVO73NzEYG6l4kMBnaFWdoibJHakElkD80axuK6HyPwsumDfaGVkQcynPiREGbD9Vh
ZUX6MNju4OTvJAa2/cYbeQw1hOeonf7pbGZ2rR+u9iU/gk312IIl/1JmxBYueJFH8yzuEsyJ4Mqn
eRQHrajMTMyWCYxRFWNJjDrhygMSLii33A3B9vv3foq5TQPk7weRl1fzz37lIrpD3T+nspipC8Nn
f8gpiBnoGuX/hZKWkmrJTqjHyTVCWP/HFEKiaMzGNpbPGwLC7LCUjI2+65wqtap1TleLXJ0d5bSr
d4sv70s4KuOertAINSgrGDMDEqHoVQEsR3YaiQRCDQP3jG5v6BOZovu++J/VN3lVSUmcHODMZi9M
14AoWjObS5lPIe6oGIOsVKew3m4n02yLxHEx8waQ7qIhhHcitC7jywIOIRFJO/whKzIwq1+Tv8he
JU/WfQ3gmlrRRVeekxrOBDM7RWQpHy3uGEqLLYaHk52/h0QMuok1svUc75cOIzL8/ug2DfvEWoLn
hhPU4pBmpzDxOAjytkn3BckOuRgJtl0rSmh2Wq4GSFE=
`protect end_protected
