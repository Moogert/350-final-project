-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RprZjXkGXQK8jgU2qeWZjSQjXHJyUXnbR2gRQNECMiENm59NUCM5WWSrPcEWjH41kO8uMTf3qli1
ECo0ZAxhtn+QsKoGPSI9cTjz4+fnHtm88HRmWMYHDc7ka1nPxrlGCgZuJrQ2NTKEKt63gft9jnJh
WzudcZrx4x1b56qszK1uJCVZw+LBq97R9vj0q7kyat/d9ufiSAObll3qoc3HDEsbrGcIIFsToQKP
w7MUR9idY2sjiSlFqndT1LF332td/ftuzkx2TN8/4IMt9LujpnjDFhJnBhV72o0KWSUflnyOYS+B
BRM093QTbAzGBx+l7rpisFpEr/0Q3T6JUBZNMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5312)
`protect data_block
LqlyyY1HYKnll17uxpCN9hg3R96FVIRMb2vj7QEb9HDwAsJES47+3h+Oxm8NhnT6EwUgh1sxdFqZ
qaygwARSd5EEphyYAySJB5J/koZIhk+8DQDBTVzfUe2KJpQ5kwat+5jCYkfPkVJxie2V6ZOj6EF0
yGfv3I1Nf7o5zJn5y+DKFKki5uxC5Jb+KFMfzX0QJIdpfLkpWhP01fCe7X4SwsG2KTuF4Q6WC/pm
F5SjKppcjqSk6XeV7HGwZmj7qsTXZ3B9bmGCT5ZBVjxXQSFmYze1qcEMyA61/KmCX+pg6lE+B8wH
qEbXcKSMtwlMga78EYFtdBsVKUnLNfiUePcxR0ARhYtRdSLqLMm0W9CxtwukPnjB0aXU08OQSJaM
O3PkoSCNuCJNfUzyn7eR3wMpgBjbRFneb9c23boRNJZalYKqkd/vzIarEXytCQA2HgDTiwttmii8
C4itVYQj0gKNzpjEwM65csim0XNXZPZxDLRYOnmNNA97yMY3tcSZS/wkmVVD9332ZRsDyRqP9j9N
o1xewB+GattI39iBZTzhFXtvfX5j3OzYHID5RsmzqYbvNpl1VNKnUZuQWsK1cfIdxf/jO7zygsRA
kVc9UbB3KonsYCiBOO6cmilyNny82xypjttGdVYvHp3usD5ZeQL9VOpU9hSDNmKkurHrIQK2TgsX
IFvfzpv8BVGPvvk8mcqo+IH/Y4QCC61SUKDmOwfm14aHSwFvVPEHXKgBTrRkgOCFNzcW/iDR1KlL
8V5SBpcpIaOL2PsvZkc0e7Iqa9JymEb36eOE0WfUgNc4DAs0Ex3OudK1DpvmJz4jvXwKrbBqpogs
e86oYh/fqxg9xfWFn7dTTrfKeOD4eut+dVeBYAJgQ1TxrOyd82UxqJrntjTGbYb7ezySHPwVKznu
fmq7CXyAxxqB4ppdjsQuqQlsOA7qHhu6oxbD0vNjWs71GbZ9E9JjUdLBNhz0NBM5mpQXjwO2T7mg
A1qBGaJlMn6VLPwh48tpq6+rd558A4YgMirGsOeeUFArNnQdBIwdFa34yBJdghogGoAm0/6B4ZkD
4OaF0mUG4HU/U5pJJJBv/Id8gFGmdZd4lBjS5g7qt5rVdNqSTDbMYO1dxV2AVJuOKZB3ogk8qTJt
b+OSrdXsUvX3z9WK+cy+Pr6zm10vL0Jkweesojm7kmyVNGYSRHKE13qiUAmi+BLoUakqLp/RTi5A
XTI5xirMboZ8HJla+/PQcP1NXfNm/fXdaYg5DgAOXd0krrR9244+CD8DXMgt50YqotThCRA5r2HL
l0BqWtSUl9E1TcpszoMwgH9j1xMQrI81cHnYfzfyJZTK3CxYXujM4k2U82g8N50QyQs+wLOV3zZe
qQVF7iULE7kpmgGLp+yfADulAVznvor5215FobyEURtLAltGLg1wI48BoyuzZ65tJpXpz1Q0Cls8
PCXEGRZHpjdFIZuO44NGrP38DIC08hWhLDSN31Q+zaeOibSuMlwiE0T5PKVBLs7GR2OdMzA9zpDj
huFz66jaVeaPpvYG+onLwcot00g8lBGa2sCBdP9jHZ+FBqbIYNZD3xY/IxglUU82oKwsk24wvLAA
mKweUAICCwH4dRQuQneYtTh7FG6aP/yzuel/GGuWol4vy/FXnL+Z5EpR9uG6unUMfrZE56Mli1X0
anb8pZ7jul8e/eYWixffT3SYgZOTAtDspgUvsZm7R/9uRD60ckx0LIARqe4NQudaX9x4nSQ3D7JW
z41yPlRBgyykh589JOhxoQTNrRLrGzzR2M3+YzBddWtAOgkPDkmgpUpXpdxHD1SoJ19GdRWA056C
Ypx3o9s17VAQgweHmb5b2l+GoSheu28N/sUxVRPUGUrE8v11KkwvlbIrcOeJE+opqqj2sBSA6W48
7LjOlVSAqu5Ke6xeWmlbprwkm1FtrdAVjT/Ct2dYTJ6QDRT1biEJpxpqYouPgm269MatzimxSXNJ
0u3EwdgxIBmF3JTLpxugRmXrGBxAIr+Tc6+cKzDfmAJ582q3sg/2RDdPL1wXEE3KV7K3N1wvIgWX
rGKcmKMN2I9TGKcVFb8A/S8xPIkzy9iUVpRfsLm5EXYIOFbZi35C7e9g9l7u8ls+44wC6xJ9x76C
M1aOi/lMXHUF+NT9BlY2Z5/gmpedHN7Oye2C8aONCGrr9DAE0iydWSAAb/hSzdJhB2pXyTB/Sh/M
+w/22djyCxR9GKcWLS15wzk+/2MoiOPFMtR+4aY6rvKCo3LCjuN7BaFSGQFWWqclv5nWx//G7tUn
Zr+l0E/ZS05puTj5RHI09kThDEKdE2AkOUOiWyrN547fUzX7h3ccRjtCE4N7B8Wao7uEUB25OGWv
Jg+rTOmx9fsmdtUd65XKF7AWhAA5IXEg4XQNWDUkT0TVC4gCmftXe+1buAsvLipVNYXjWRYd/OyG
eKF56Tug+Ix6DHlOXy36BkXwZ6b7YnwC7xdz8fatUDJf833YTjyQCu3t6QgsJi8YzZafTb8StxpG
kn5oADJt7BJu5O0x5woIoj8tzpjUlFJXGbPLbqYWUjvZJZebNJ9ZRTrl8wsVdwMuPr68kIWc02SZ
DG4AuuzZTzT4gbBQHH2nt7ydlX2jZODttWljL8EZRBkFyd5EjlKW3i3LZhYPQBvrLpWuXGeGKtgC
JLpdVTTGfQOmBV3DED/Bz4mPzWvo4rQIY6bppJvOcGY4x+iHO/BpOYe9z3cBsPq/tjphIE3shukM
QeP8P8SOK8ountki9E/5ohJ4NSlUdAHsRMggpZq/8D5iPf4IAX5WhxfqRyef58+fHkM4s/Ta/xpW
n9sVlnDM979IpFbru+YCnNHFqsxp+FwNKdYBdkX8VEtByN4uXPzpLW3Wdba1U+auFiGNh+E4XZzU
gaGY2Xk0eYq30yNQ87peVTXOBzk8fzzoP1cW4t5QbYk7AU5aGSl8sMCJyCzb9oAKQPKtpdMgyGo2
gpvFgq0RRv8fnBD3jsP/UHDO/yiC2fM8/lTqhl0P7lUCT5TNArgcjO7ZOqHme5njvZzLfb/ZTIGM
/3VqqcmXMzNEMN40aOhCVN0UvfELrjShzku/6cCAxWlt2wzxcbanpVIzjORU35oKGWFGXzbkaVFo
R/hSjwibh4P6uLhqbVHu7BJgECs7wmN3GpaVxbaX6QTsScOgcwkjacinlJ+cjWgRxcgeJCiveJp3
P1ClEJYCEx3Slno9sg09kLcVcyk77+Z2UkyP73EYyrR8itmQBD16B70DEFoFbGr6FKcpJI5YTcBx
DgtiUlDGUNXyfx4uTnp/RxZTggqfW86IUBUMOLHE8Lxv2h22uMOFqIhNt44alvJb2Z6pnb4pu66r
IoqsYus7RKoZzhvrAF6IPYOJrb1E5wlzfligSjwZJamhYJwySxCcff59tjCd8BQnRxoQBGtFkSCq
wKDFnWbrMO3/QCMAtYl84aH9pROLH+tddfm8M26x5WWMANm6xTe6DGiaYqH5fAfCAvhvqYyWyTY/
d6wLeyoKcdluUKpnzmvURfwYOMQ/Au1YhDCOLBfXElSLxGprlGFE1rlPiuCYzh05plCSsgiiD6L3
BfUscaae/x1MpVgFmmkR1bUz1Jz+Z6fEnWRvfIv2gdx99jWkfvi/wxBEVdZ5Bqc8uMdpnWzMQgYO
NQ8dhbnww5okccTsnDeHC3GfH0Al5g1janjYEBX7EY30OrZEUEGU5mcJ2dUb+Up1i+83bVgDfyku
7wzQKv0tcLxH3lSY03LHoftpcdCgWx9edoDfJewVN9+yhdkztc6wWb2zF/Nb1js2YMNZZyfzZFfM
kUgjq4RFQolAFr5XXsN/PYKY83TM4dIPoXde5acXJOUPQ+XYXYA+DhxZLopaNryUZYvGhXTYFSoh
42mnfjTtRJZbF+i/gU8/Qdnj1C1eMqmvb/ew+MnNdGb3hSQVwvBmh9fKY2aEMEnc7Dbd2pELpO+1
p2A7UVBHoL5v0iiNfZ8HFB9AeggNcW6fSxe7YGFrVZsAul9eXaCRtPWhGdF2ReVg3sa3gHQLrlYz
V4KIrjaBrqYYhonOia84b3Z/GUOUOHHncKJMLJqQKrgfgiqA+HIVgUEmBc0g/llMGTdK7FWVRgMK
1CPDOIiv3C9DF7wobT48eGy+bpfoxGW+FFoP9LSXIZydilWbESsnI7VJwzxuhZy4ims2CCwz15I9
vtzmpH56RQzkSq09ZKDaz1XSpWYATdimNQMHWLlt0Ai2jrUCbM9eHlhLix+gE3StsyhTBjycpaV+
FMTKSX1NTfCWV/aZIw4x4L2bMBKlLecUqzpBCQuZRGXDwbF/fLcRSeBhFPegs4AneMX9rhpFX1Od
TpnRwuFM9or8M16zg3zvkYWk3RzvzeuDMyDEwhvzE+j6FUQRfmEDQtrnVraWExsO0IXvtAY7ekm2
QYd80BQSA5siX3og/RHWrdcV9RauibGzCEA2u7KP5pzzxJBNgwXDCVIc5eVpr/kdTVUF2MeIMHE+
Gne2Kg8SSDujg0x8jRqaSjtRKC3WzbyGL/HB24NrO6RYVrkNa1uySYTJWLxLqIHLb29kZCzmNvlX
6fG0yxVgt0Yha8tQ/x2xGnjl8aw6hR0DLyZxf+5lbeRkxclX4t1UKF6S+J/AT7fHt/oFNw5Gj4x0
CnCzbSDKBN1zFPg2REJ4n2Xp4/hgznHoJjl19ekXMh+w62ayaKKqjMnIKTzZwHBXBbLxbR5lMwll
/T5548DjrQoxv16JIqLhKZDJQpDq8b5q66WMcFpG/t/8kv+MuwRsOKEsUIGzAbeSLozNksdr2mnj
Lrv2/4bgNvzTvN0pQXHEsX8NOuBkQBFmF8ki/78a8E17XymeG5W+DZJCAGZ4IDz8SJTx3+sRtmXB
AXrQSluo7QCSVJbKyRVqWwuogaQLqtXOVJbwdBDVQO5hvGZWGY7ARgpKPbMrF41lkDJuGNjNXsyM
Bw/Bn8aSjymjwKDxfdswwnlvWBXIepfzbdaqzOGiTxe5IM4yUoNhVEJwyE8Cym6Vc1AVAggSfI1V
9R4TZcGSpknpLC9T4UzQdOuq97q5tVAKhEEtnq49ilfW/60NUgdjtfPtIL2YRigGuwH7m2yRFGEf
nttBIRnFulln42HJm+Mk1w/2ULjflPk0t5kKYB9Bc0PO7vTTDiYBRmjHfxz2PMuPy6FEahjs2pDn
rKH9HXWCkf0WG24MGkbXusOs8HokHtLS24mtXIRsL28iqKS0M9hi+RhQOmwmp1OyG5GueZUGTrBD
K0T+L0frwVqxUij0/+g2chIhK4EVcSx3gvkOLCVlzmieRxDAd6HiCXrpW1Xdw6n2/fZnyRcGV4VY
c5JOWlQZPeIwXTFXQV+Jzn6ZDcmF5LYgfioaIlXxpPP9XoJyPOQpfyfRY07203XHkgifjj7Vhcuy
eYEdgCingIlnkBgAYK7a4sVtVHFPjn6Pba1kjWr5hD2WxheSejD2QMAha33eJq8+OA1EAAKJ5rlT
LTc2L+sh8scJ0akFuVHWCkY4Jb7gNVhj5nKBrTjiXdMOh6ZSB2XpjTeRG9OvsDiaJ7i6QrPocVpi
PXNka3xazEfJWub/Sshvvybu/M3bJWBFWMkr23GOabboMO3uLFXE54o6mGEJisG0KNJ/JBw77x6s
rQKVJ6XnXxgEBgPluJkt6+i8ZZCB2cU41IscYpRT+LiYns6o2ZV1IUJD/MZQ2kpr4TzexCW3NY3u
HhbM82/xfnCbQ9YrnJh1T7Ka9u7nDDXbUm7a2nWpxjJ17lbwo9HgTFo/PiVhTfWF7bb1bkVt0ndW
hxgCsGFFZRInixjrBecI/D4lYT6luU/ROG7rxCGy+Mj4rI7aaISRSf7tk4T9SK9M9kcQmCUpv0jZ
WcdypwfvJDNn1o04NrShHQD3/Zr7Ge8B5CGIZ0DuZBYDTzpA3sB5sKBFaGiKPGUyaVtiqqnU5oRZ
V01GWLk12TteSnKgSxW7AKsweQZ6j1EZ2jpgfE2ezrJiGo6zNpHiW/t0BElAh1ccXRUgosw2h/s4
VG9SqMdlXPtL/Ue5sBjMGvnXrpkW7RiyPnHXT6j1Hy+DCjQ+gmUeibknIDtuLoKdiBj4SYUgwhFW
j630umSHGSKLmln87woMil9V7RdDpKAh6vga6UL/8ua8ojLSB93PCRNW6AXKdNwjvy3A6+WEREp6
rPBBUu8y/c10BA2v7n7zdnl6B1I+dNkUzE2mLfzuBj8FpWtlTs6ae5OQDWd0VCHzZ/EE9cUnO2nj
9kFN8yMNHNYg6wujeoqIFS0bYDNogyY6ALJFQtkryL9jm8j9lCgXSGXA3HGZYMVk8Lgda6AVHgME
X+pLMINT0nwu4ICMrPGxrLkYotQROrR/0Xt/fNjDXLPkaY9pAqe0d9bKpzBLBuwA4n0wWeWzhgrb
FmxuOhTck17Qn9r3osvfQTwyb1rhpc7FtqYa7nn5qRSu3re1qReXFQihXJSZXdQar5knJ/rrUp5a
gaypRWIYuMO3bSoSpEXavTRUWrUSqvx93sSXFF94y5hwjzaDsynEmoQkoocrwTGfpDQ/CBScRkFL
L4mItLE5zhTgNFwtstHhsQUTqTztfvqHutZ6KEIZdQb/uP/WCuYESXP9YL285KFX++5yqWdbVLUw
Ah+Xa8gvNkJhxzTGJVBb7v5Ict97mOI13IDZ+OD/ps4qdXA5034A4khy1nvCCfUeDuGsRETbBGnU
oYZZDXE7fRdhik7+io63P5b5E98TDeP/jPCkn2yd8yj+2E4o5qkQ+N3+XXCLfZFIaLj2pUdpEQr6
g3EPwdyPNaHi4TIFn1GbnWeD36fvgW5W69wmt/lCh30dAg+6E6/muITFVBPKSjS8zXCVCohp9Jw0
ePU8Fx3gl1ugqBCmGO3yL/ZpmOWlI+yNnt+bphB7VmOoMSRHCEQMCf4uabE1eqOvFgaOST1rRjHo
u7b5mISE3ayrL4l+dYXUuz+rT5n66TZqlqQ/pHazoLOUJbDAd6uC3sp3RXkCOIdo1Va/Ka+b8Ydz
Clm1HYhD2iBlaPuWfHzy8ziO+KwlXNU8KsBNPA+d8RHKF2xu/Kg9Duzh9kQvRVYu6IIYV0zkJOCC
6faq9bIOznFBVi0=
`protect end_protected
