-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zsDcYXHk7vmCFRU+79qU64x8iUEbz8N80ujgy8DpOyWKYAUrUOjUQYexqPryIZnek6biaciRem/V
xd8SDP8Rlr1B+bDy4mDicfq/hiG3OS45Aw9hyuQgwSBz5SUDay/Cij9fAXQwsUETSg5L6FIM8WLj
OxDjsmWR2wVX1XZ5urJ8wc94CBSMa4uyQXflareftdpyyDD5FBfxrPOO8bbUTPsf4oIFcx0oT1B2
CxFDThy8eMPzu7dhg+5pbNBwsLQrugrsizmvLQXV7m6heZ2u45XwJAehIAg/clw0QQBDbAF5Hw+c
iMUy89YlXc6Ln4Lo9dusAYVrpUZPURlDoiid7Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
NNl/daYL0P/sNx/yjHhu15bS+XJJQqEy7EGfnjvHCf6TUaK5xl1y/JEvwSqTd6liH1W1k1Vvu9qB
ZWlzrVPn3qnu5V7Q0mGbWEmw+LisjIb4NiY5e1JLj+UMy2DDhvgtaDRir0p7s47tgmaq1LEtMj4V
SHAPR16UfztkuuOoaFnRfTAUQnia8hjGZyUj9DlDgJlgF4vpS8btA0NGCgJTRXRRU6o32DRu+e33
rl5MChpMmh6Yq5SO1dJgNXMwob5sD+GJD+onJdnTvoVjo1SithoKT+RFtHko3e1GnA9emlFKybJM
jBO6O/nP+yMHvTUPsIsrBdepfn2mpLdL+cmfRZPZxprE+6GOwJ6+2b9NT4ST4AfOaLZM3MgCE4Qo
jNmkPJB+IstC5ktsC892y3WroyqZ3W78ZqRAk4BD+b8Vi4qGbRKmfLkdzzaBU8aNWYnG+I5Y1wH8
ne3UtE+x7YFYOEkCc+vgxIiBy6AWpDsFT0RSPyRa6/syRJY19Vs6INfYRkVk5fgGpD1yIKaBjbBP
bRcV7nPasx+mbp0em3t8VloNSt9TsrSB9VuLEJqE6ruse6Wd+llVRKSdz66VqVo+60MEFUabNnGF
+G/RcCKVcEQ6kbho7g4Vw8EYcic1aagePNJjTVZHLyRXAKWuKiWxACVUdJt2PUFPLl5StZaZuK0U
f+WHj7u7Q6SnYR30DtArxRFSL4riaF7lVdl49MEa6kpg1xfDpAift1Rh4SJNmBMDP7AfT4RLH/nU
rtT9c38hOTId6lm690532XBjzO7TC6MJKqy6k2fCBAzbw75UMIUkoyCYaX3rDfv0C7Zmx3Zi/rJs
9H+1dnqwEaXvPh718loKHY8qjndX6IX/2st1SAa5RAc2Xgv0IBQlHU9JywyzPfVT1tmzyJRzoSF5
QVWuWaFjt9HV40AS7/f1ouYl3ACNtohMYP7IIuglGixm1RayqFiXjXivgM+OKNpcmheWKadd1ZYV
iRMHWVgy30/C27Ek6fAAQL8utH53T2BiF0n2xND8NZrcovzol9G+I7kBI8/f7qa7fR59je2By53y
j551gSlYiDKpaC4aGDT1Px9JS412Ly5J8LOsrgURkRi43SsxCH+mLaWlv7B/f1pc+3iv5y4wBrI+
olFm4zBVaD3ZlE0+NH8XikZKX6td9KOd6JwHEqCK42jwC498b1yJpyvXfc40NC43vpflfV2OoyJI
CAfuLoKLk/89goiDMhgnjAJgZmFvy4GUhFE/6t/V9bD4++Xm7fehJRqJd3/4e0uWDEMBbDjpzrPq
yEXTtibGeOdoQNpNjR7HQ3CFK3ZEpy/Z9T4HfsCmbNb8fQ+jpSar36gWvPgxZYMPZoDztYGu5pfc
CKMiVQVz0xhR9XoY5wCqG4RMhdwcBfORjmR/esCugqRXkGJymihiFjg9+ZQPDX3yjzqjwi41plXs
q/umWkLwcmOdPMLVbUb+eKfcH94rAMgR/NyNx9QqmBXQuWVdRyu9u8QWaKFHLrlzsHKSH36bfp4k
PnSJEpy1krEBKq+W53+8JbI5Dko5VWRJ8W1iLo92dNJFa5DUopbNcVaw394GrJFjzbkP/ApcDbIz
Ga9sr2B+AYr21KfscwRbfa5q/xjNZpFdxo1nWuDKsN12GtvmW0xtwOHdy7EE4YvjHAI7hXeu5dBF
+70h8QLABuDNn+qiZIKc+fVPOcsKNAT3qcy3QiYHt706EiJGd1yR/4RYpqN3dycRkKVZZSoY0BsJ
JwabIa7L9dpPbNTOjDa1VMFbw7o6vtHzkNt9ZSqzfzKhAi3vyvJh/Mqwe+Q9r5DNIK2Sb4Pt4sxy
X5TeWNwRzdZ9JQi9P6T8O39LTiXpcBw2/WpDuHZgxzldCqkHp1YYT4em7NqmFSbMEy/0VzQs/7CB
CbsXJkWMdwDHMYGs6UveyQFhT8w7vvIazgzCpzexehd+YXkUooqthSNrrdDp4hl3fprSiCbJTn0G
3h9NY9BxgpQn80buftiCs4tI383cqoRn+DsCZHHXOMLZlpX9N5x+Ddgmf/uSyltqL8HtzxUZkcrq
/uz2CjWkQ0wqy35Fs9Fl8bERHKiwrRvlFbo7HHSzoqMViNMfxI+iPMV5pIzsU6R2saQt2zBEKJ65
XnCQSAUeXxuv5pBPOubmVEgFlwt3BLJTkWFVTkkh0exfi4YHhwp6w58ZDtRlEimKUWUlTf8MTWCA
NQmSJEAJrC/HVq0KKwHKAbxkrVa2A/v8Wuffk5VybHoLRbwQWjGoj0TKm2qv1CkIdfnc/njubOdx
pQ1igpakKtqWRqpYLQZxMxldsDC4YhCj5mnJD09iB96kZmsW02Qhi0Z09CSKpbuPGy18qmvv6ZUE
rBcah82mJIMhwKRSYbDG8ApVc5/l2JI+SG6iNfxMQH6f3mi+8jmZ7bf5SQHj4L+r5oqoFUTjZyxU
ZOV9WX0Z4pSoD8vqDcRgSB6KkEAK25p91uhYO5g5w3Pa+qJ8zG1L83u3TWCoUazFrI61NB1PatWp
zxi0Gq7A3xoA3VRpcC6V7v5XSzvfq6lkk3fIbx2ywtQhAKjj6d8FvG+818w7krGYmFk9ewzXoHfK
MIEM3CS/xo/wSirarFu9vaMcZljEwqozZB59CLCECnr8rYP6pchRrpWr02CjzF/KJDZ8lgcsZMUk
F3PUa68uH2cfx5NO41Q5kQTlZah5kLZxyoMc0n/ucLblOggadVAULJQ9+NMWoyCexOvQLBZOObY/
Bse1MTxBgBorTdaKmBdChkNBm4U1zKf+BH4L99S57T4xWGAhRCET2xEWvljsyZJmBnRoX+6mNieQ
IxKiXycGzZRmiFwij5FRvERi5Wt/sgodLaPUfCgAuPWbSyR1PtK2znUlZg0cK2dx03Q5Vb9Yznib
AclKdj6LpdaCfzsu8J5Acz5DBaXX7soRIJnDtDrfd33mlL1MXU6iuRGgBOaLEWluADXjALnzSg12
fkage0vTD87+dP7WUIH3rpaCXIJK+5mbXyrYzTZQDSjv50ZWVhzd/ba5F0zPp5H7vzR/13yaTx3U
feK2AxLn129DuOPvgpFjlut9OqIBOdu116pkx1QPeU07HRqzRaHuiqJnlQDZeMKn8nHZTrD0wWsY
G2n3MdzYdEHrGRO1H+j6JIKZ5DWb1uTxNeEErZfwn5Gjr2GoPXJXzmp0KhbERJppFo8nymmBeY1v
dvftxuVP3J3Q+pz357FO9MwAtEdKm73bvnpShpvBDPW4NHs4n+cdIvbUHPErtsYFLF39CM1VuC9k
YvD5WLIQX8abxpFmoFLbIDFmaCKtuVz1pRjovjazYDJm0q/gKObOBsI4GrGcR1bZv/sl2ZGCmkGb
oQ4np/2OQ9GsbscrL5oTlNBBEjx1RqyUNKUjgPefrXElA2PhrQS26GUYSkPH+9Jju0w7DhkfSohb
ayOmhwQROdxNQEhJ+uJp6mRVr2J8gzNfww35iI+MTdcrFANOmTRA1C/8M8QEA5f//3Va4vRRBpqL
lOexjaBB7A3lBQxtkG3ULp4b98jDSLhAsPpZTnSkGZGLNaq/I0QLSc//DMwDs3MbKKZsmQL9fXfB
lLHZR1V6TN06W12lClJwnXrrQqq6YHn+yYMy8KBRR8jUaLDDdNstGC9sdXqD7H9PVYUcpGoUDCsV
7LMO6CLZuZ3CloAoD1TE1a4DyhkSDaZ0JfbdIz/vlrFdXayEdCAxBhN8nSE4C6DRxhr6MTB+7CAE
0lNJGZaPYxxtxafh9RbPZ4q5MTZWVEzJ0V6OTx1rw4WdU9ZtyI4Yshig49LNfHooWZUvhilU+9Oh
+vuei70PQc1WQgWB0Cw8m57Fs5jltXXTvf95ZPtILnqnWrDWx7SDnRUpIC+z86oyk8I5s24M/p6d
KsLnTiiLQqgFVVFCo8vGRoYInTi3Lv/QM38EBI1ikdnNGbZuKJhBP+Hvt22udEmel+ye/UHv2To3
z2chELrYcoaG/mhUSIJw36rB9Q3QbPGbDEB/jkd4nB6DLaVMVC5o7zAiGl5K/fd3vAk+mHKt5n+5
Tpw6FgaHqEE0RoE+vcUTRoFylUe01RPJp1YGdFrFg77h33I30GJJuZ6MQeRYdsguitAuy3OE2gwC
hOgoclYpYsDZ/9+OeVrlGi5c7plsFClnzbf2qATUXdbOJlEo45utJTZgYvCDbFi5URaf3treFHMq
cFQm9Z6AjFbjqqrSCoGoZJPg6VPayRp+2z0lN9EPE6+GXqmQSQncbz2vWhpcR2gOmrB3k66vs9XO
zbhG2rCAMlwRUmzqMF4utVRy0JsCw1HdeLivRnlk7ukvaybfR2JaTpwaU4jTw4iJM161BOnUf5Ji
6RAJY/kSkFlIK4Cbd7hM4QTNPsTYe8TY5BXlGog9x5lmZTCgzm0w149HS+tQd15E/uIHvGmwt8Ic
nNtJ7axzDQZcsC0cYgeN3m1BR+J8qJTaxg/ocu2tT5W4V99mxkvMOOlgMKd776vU2tASO9iZdPyi
lA3zTYqSMn98lAagEzIA2CbU6avtScqSgxKl76A76gD7+amKp7OfQYVEZZpOXzBJN5hhBtYsZfUg
dkc1bPg5F7MiWJMz5oUcR4QUxtLHwZtoaxOH8H0AALYCd1tVriv3YIoP99hrQ1dL2k63iO+Qb1kl
rzgb2oOeD6r0WZYFAyi3EsKI36k2hY/ccYvAWXDCeqbsXS+SE5NDcVqK/Ym4ZQ5grFkP7p6dmfjO
jYusAbg+T7Mb3eOJq+8T/wgAihpRrvUkjVES1d9FpqjCxe0gcqzpfRj1Osdc48eLd95OlV2Sugb4
YFKoYq0eOkViNsipcSVtaeXKg266YvX828c9s0rZcK/DhB2T1DOqB7LyBiz4ckLdiaONtQIlOs2y
sdsikinCmkUA+0ZR5nqboKUdMXYfJh8lTT9HTocRsgw96J1C6ulw8/hu2OGrJoIAQOOyl7HXdXGm
cpof2zXyOh7X+urNfR1JFgQtf8IKDLJG9SAk8f8J32YtBSvxsrN5bHMyH1+3bYW3QkULDoFx3sWj
HdDBUI9EJHFbhDhyGtBYBFU7vDiW0523/xMB9BsOh0RSZfZk5KkUsm+iHIa21mX4Q+2momLImEP9
IHd91OuQQYaEvsTsB0sSKASeKtYMujXZASKELK+8n17j6yz69JFTI5k5nZ1k+l5uSoiV8QAHnZE+
VZ4TqHnQgwOEqjVvK2j2ic1YPCZdHmG3S1EG/QDrUDfF0k/siXHVRFSpX0rlRHqjnuFC/w3JBZM/
nJw7CHM2zmveGWEUlCeIwd1oD/fqDFnn46ax7dDLdL/emosOZ62oJNWMsAbNPgb0F/03oyiNO5Gs
tcxRy752uY9RgYsUmaQxQ02lCsJabRoONA2mfI0k4FYXz6gkp/+IvVvx+TJmEMy7RfTbJiGkVaeZ
/n0m+Gtpnaf9+5cN2poEkibfh9g9Svd/oHW3qm83LzkATqg7SPhQb0J5hNkYBwHhtibn9ZMtAm4r
bP8xo2XwwaM7bBFZl3WJmAmYly2P0Pn4du/EcpEjHrjUeQF47Br5db/fH12OoTMFIWd4sx7dRKCr
GoBJNtnHJydQz2CCKjtm+et07xk7o9M0HkNKW1q/3OmasyFPQyZga+261YhjsNE+rk+OPZ1XJeSv
nbUfQzX1xgyJxxSUWG6leNFrEudrn2QSX8iaKquJJ3HscOPRlh+UmKnptzZN9o5Hiniqh3V8Ije8
NLfg5ReNLxbYVJxXIrB+b2hGTKu7ZscjFYj9AFRWY1vdJM07lkHOnzSxuyhPQJrrRbxKP5WEnybb
VY9+ZQ5zVubYd7LIPHPla6vx8Vgu+EosMhKJ2rjXS8nl/IDDd9m6vBi2Z+mp1G6YVx6gdxynKD1/
zCvMiNUUzUP/vUcoK9H5AwYik7OHsQDRaVwDCiEHk+OTSiNVNYvDPjTTRodzomESDFruOqLH5CmC
eUlalNMEIX416IibT7LpXSvHLn/OaD8RtHCZHfwto2MuADeKClqniNu+/yojQxxhWurhHx6C9PfE
uuYv7q3vPMu5cYBkcTvI7fcwfknG+K7STfa6p7UoPuepOYaqtOUMO94Ij2CsGYH39c+Y3Qjd1Ko1
5JFoTa9B3x9VlFkUQEbCZBbZNDj4ZUbetRAtkXNvimVVf9uDrTOII566IWs5SNLKNCSM+Jkp9KGi
3IZBEs0rdIbiBX8h15LYflyCf4cdhK0Kf7Vd1MP5YFopLIxc7v83o1jLKNu3N/GLegvjTNxx15la
jqZDD1EbJ9K6rPgTXbEGOvUnBqpaYoUDWQ60Oqx/fuDsyCUOpcuQEFE1tW7RYfaEJnOkFiA69PNV
fRJ35/s8S/QnOuEpiUV73lQ0ai00aS+UrydZO76LUYvW8qwTphNTAUld2ryEXCMLdly5ZR223MWn
ysXDriThbBOfjw1rwisTGfdq07Ew8Nl+YWPP2KT4jdKo2QYmys7QTca9w0OnxDhf61Y2xUF6WykR
ZK8BTCjrbBXbcUpNucFRCH+JdRzOy55d04dldhtZYrgG/oO+hPV2+uaSovXQ9ge9ubKC4CYqYS44
yNVAjsqudXWtuo4eR733zdyzygXG56J/NNuIgo8A0pUCviZTOYCgc4HX1G5wWk9izGlLMQu30e9A
TGy+nIChem/uaPvfqtHDtDivjeHh06N7bUPwAviXxqjoeFXa4l/oD4shc84tE4+wcAQqY+Ov3x5z
t4R2Dk2KGHlKRoRA2wzWD66qhkOA1uIHW61AvksKvXwOsV6+RpQDjGRvkI2KeLehpErXL8mmtLZ4
Bvj1HKpIGKnh3rlfLCEDMljYnqeaFAlqJYtCiopIyc/cE7FdQX/xT5Qs36q7pqcv3rVFlnn3DcM3
p3YX38sI1pSxwqaW5XSyDwQlIx1+G4j4pphCEJE+1IMgJaArTTfpIt6zkHgSEcZ0Rb8M2bA79Ol/
5xVlCUGfcPU4uraPNLzmzgWobdyEdNyw7jZw040uKFrYqRk0QCnj1ZYSZkJ2OVdSHk5xMLr9tk1v
yPSYTe80UIqu3SE8kdWMZXIqm+Wze2oWieOLxpGdvhYf31uXzRJ7JFHR7zPXc+snX9TZsk7LLPIl
1Dzn8FawOxFYOz4ZcyBNBo6URCcn2uAaPtu6m/g67cDkItyeVO1xwL1ZtRhwGIHhYWu9fETwXEGO
NNsXpGV20QPI5KCws2KY0GhG0AobLve1krCnAlOf74oVjSv77ZFXxQaVxTbJ5KejK9gwZUOO4o0B
/tYDSLnH/JHbej32/hGO/2Ub/ALYxmfgQ/VLNqtEfAxiD00LBgMbr7n45ftL2NeX5oyJEp74oNu5
nzhZaS9U9JzjjA4ZluLsCJ2kvvkY55gLlmiPVSD3aEyvm8lYNjdZUTNLa1uQE4WgJ4iJ5ts6F/hD
0ArZRqwXp8125n0ilkKXSekSf+aCQ7rQGL0SxShFE4P3TNlA1ptKD+toNux+o1tdP1YYI0QF7nc/
zcXpOwc7sBiTBah2w6TZA/Il+FRE36J0Y1LQ+rv0gA790LgNkLNJC1HxQSpeQI+zqaXZE+IHYuSE
5qOeMKnYnQL9qsNAoMRw2ZaTLjKiGxGT/1Fvwz7I5ieWU3yM2zuIj5rhZht3Y3xJAm7Yx6C0e+fv
tAeyNPe+Yum6TrtFkhrnAqPzBip2V4aKMg3YFVD6xicvp3lhcxlbnosqdledKOOYCXiAXA9YN8q5
5sL4Nj7YPW9RVyM2b9IBVGszYl0hBUeA/NHKqYM6dxq1ADLmByCbcciktEfUTAtzy5/LQiuXExzE
EZJl+iPpSTKEyCGGxZRTE9rKPb8n9TcnSJdIzPGovKvF0UyisD7il9mc2/oyJ6xJY7wJtgCCOAtK
4i4xLACGFAYbWTQ4i1jzaf+xSyUAcQS1/p+oGAXBN1k8umDpv+OeBe+P0ZzB+jonz0beG2sb62XN
E8EWoFRTuu4j8p0okyNYR3LLKDoaCjlzEZ77eo0MyH9RxFP1+YH27o39JkkqscKYUG2OUdChYLyC
HuNaMs1QBsYFGSTnNejShw1gQLTh26OfwW3kaVbST6cjDq5kGgM8vVPZZaBjSHO3aK1934JK8yjC
mks/10S7DYxqDr9aQ9TEe5rRJolw23w9WczwXNMyeoof0wgzRlXeDHhOhgYo+PE/YWeToVSyjwGA
6w9/7z4ARqDOZNx8jQ9mTxkBsi0uHDiUidqOC7vtCTnI66zB7zxma2gTSpax+Z1jp8i/0AIDaAJY
xluFNo6Zi73zPEFK/Kt+hlO4zb6gUkQBMNC69WYTcLWEb8JmNPDSdehCj4LqYjEKKy2YD1UQEKiq
5/p3HY0JGLmdLg/sqGs30ac8tQVRw6Br67hsK5G6YMz3lVfT1YSjSAAA5cvwIIWItMLQXFpHZWZ0
tyKDfPd6klYc8gad7d3q84MwID/j6mXp2S/o2Z3maR9EQ+1zP3iZwStNWSS7WKrZ1uFquuk9+id1
3z560ogIUZN1pzT+7V66+A4wHrWqsOY20po+EiUGz96XKYWgi2xKA2wh0TRP0KNE7JKZ+Huft5PM
bCSDlBBe9ozB3uP4L8/BVAvCusYAjxrF5FmNYCzDHaPuGFRp4a0OQh0m3zqxAFS8tvehw6SAPRdK
RKtxLNo6t5nO+qvWeLlZKD1Qy48ZEFAHzRzaTStABhn/UGD4u6WVOk/z+7IRDcZo2aWdDIOrVUNw
V6XL1IaaDHgM4eu4P/ByK85kDZS1XGQeAbqWu81nZ0gKZY0xrr8RkxDb6LRAd3a6cRxBYLTeQdnj
3Qra6GUehIq1jo4TkNfX8Rm4ZJnzmFB73+w6o7o5NPpdAHiAW3xlIgmPOGke20Du5nr6Jhg+og6I
sfA4zgtyxs30Rn/E3Zl+Nu2YyZTFABA9eDi12GdSIVvmlM8HgPcHQJ6cWZL5lSZgAYTpqG7OuBrE
T8Cpa68My514TrXYozZ0zQtGI9QEhC8eys7J4tv9B6tcYvDse9B/+gjTURHqmIBg4rhuEyJfTyrG
KWG0d6lUdUpm/2yswmWpXlyN/DyKr2sPaHREciSMGFfuGfJ4cI2tzyfSoMGlFUsmMWdJnmq3Yo8a
1wJouCCnQJg2kIqYlZ63kwmWNdZnqTgzmsVtllkiWlc/uM4p5zHhC9UN8Z8JIG7xMr6mjoZvuBmc
WG4ujAx5lU2UbzfcM9sGDQ+LssirW8FvK+kTqfFyivPD79+ElTDxFIUoZLw9njMSreQViZue3vZm
BmpTircb9w3Tr9Hhn5GqvxbQ6g3jjGi34fac/KNrtlz8D/dCXkyCMSsVlP1XUphDWubhdVozkffe
hIzeS7MrNRer0gH8qRga3u3YnRg8igQIz3zKqZJzb1apWSfULY3ps93BmcvpE0HUvpgE+i4CAOQJ
BouAVGy1e0JitzWX0sZyCl7+F3M4SuLbBffPFhFl6sJFiseCCXq1hV6cAqqjJ1D1NP+78FiHDIrO
owXfJ04piOhzsxKdkvH7M99K5lksssxXL1mv5MbBm2Kh98Ey0DLwjxt/b0mTyWJaiQoCzlZs/gcN
jy4cvHOk+6k8TVzuzM2eJhrPLVovt7eoGAWDF1JUciBJqIqquIELtsCSFYZdcx8h49e5AkSICeRr
9gR5fj3Bp3ie9PjaKDw8mfsbEhfnClfDFsnYpCwjUF0Fr5zpkz/Xlb0Xw6PLpSUeTgy/V/6eqyVO
n2MmT2p9oKSmemjYl5F3cPMabWy6CssIzzBvJHf7/fsxa0uT6cQngWWQnHqSifKjhRoBz47GaYS2
bjgV0/PlHw4YaQcKon5CQXPykkZ5tO54XeWMavZDW8wA2hL6+M/WbuNPf5WewPFixlAfnUVgJ1KL
ueoGFjAfZSGYF+YLgZl8rl+qnWNmokK7nC8iYRBM9KrFt2Ih4iwALVe9ZhbUSU2VsNt698c8ZcXq
DI6AN+3g35FtFtko5/yJoO5lDchrzTouweSfp6yrMv1nE+28OrPAvmscvnIujQZsSluUF5p09Ttb
mshKSz/rQEyiic7BSIcRfEgLWdeolNcT3HriuhKxIrp0b7YerRrF5/f7QhQUEASc2ot9uaSsI1vL
+bdG5C9tzkLp3eKps7ULylqP9vSxq7RlLbltw0e2PfDbmza1b9XhyZ1wzQPiUMJYL/96y93ZL2Zw
dwDERRk5ZpT5L7lznKHDwf0LUXqjyChqcGVT4qZwPTGDDmfUYMqdsoUWvWIVA2X0VEsJCf2lmqwn
7XxcvK8lY+gLUtTAn+9MDLlFfOcL2ZQ8wWe2GAEOBVf5ZHZbFsyLeCxaGXqbKjyjLLFSxi84o90c
5u7wUOmyVfqKyIxBBDQjoMHzVBt7A1jxl6LwDwHn0bnQCKfTbsPEgTM+RNlP8mUC0XljMZYz0IYy
QJalrFbdxbW/lWa43yUixqRFpXfcwb7VaeZuaFxCqNZwr1GYAC4NqoleQkGqgoN5v9rh1h4ZMOCU
E0Ghxu41RrXnVXj4Z9ZLES6H3YpkGUvFvlMY9Q0P3oflpiQ5F+Y34ZEo1zO9HBmM23jQ6cQa9lyj
S4kzZ34/Irkf+aEKgXEeOKpXWcA2U4b03wdzhoVY+N6cFaEQqK1m4n8U+l4MlBS0fT2axRhj01ft
TL9uMEeXCXSdsBy/B7FZUnc6C6MULxNE3314/oYqla30K8hZRUX5YIi2cgWgTpcKn66MOwuGd65+
RkXCv6/5ciKl9+aVXqrVXGtAEu79wQvsSiy3EWkQdbp7Y+dTKJkLg4xllLka80oGcsJnZLq//9fG
1K6B1AEOEhPBtQ0lj4CokQCb0JuG4o09WHcdrmZmiAYycZ0khzfwwOSoyioga5tWc7xkTLXycSPw
jEDgCzQLHXmomelzdNSLEt+zX6veU5Lr4CjRxSwA2fvVDXCI6lu6WubtE3ary1dXLiTBPUIfTX0d
wFS6IR6PyAKJr9CvbhPxEEabqWKm6bAbLYpaEqFC693UqOJEySDYw9u1J1Tmr5OtD9WVbXcLu3PA
NkHW2Lt/qpmmogpiz4JWml79218xO9EG5E8cOysfbngVtbQBisBqV0mcuWn4cCZHhb7lK4or6e9Q
6BrvDjP/KC898ajk8r4tH0UkEN21E/h5h3DHGWg/eQO8SMw9h45eZBShyrfsPA9dZF1Rk5eFmqFr
hEbd1igajbTmfxRpIRpkay5xtfSoevN4WSz+XVUnZBfrPbBmkL7DdsFgfoT/04J+9BulT0lgnNdU
nFq2eu89xiOg/k/wjaGP/HT538dKn4ds+W+G+BJtVb6x+kn/pMqTExRUV55K0hsgnV0BJ4jNOvVI
j2PYhQ18/nobBwmp21KD6/RXxki7QHZ2Xbh/oW3+SRzAjrln8V4pZk6odic5qZBSkrpIPwK6ogUJ
jDmf82WGGiki24A+4Ek0A8I/h5rK6QqdKshcDna+Ny+vi0QYcR2zzKN2EIEuzaO3kmzU
`protect end_protected
