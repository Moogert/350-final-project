��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�FMP�I>rG�@��P�~�:��-îy�J��C�~L� �}V]�T���i��)9����xX�����7��?���B3��2��nj"z�p�� s�,y"h�z%�P��;,����UB%�=Y�A1�,UU�͖`��l��d`� �n�t[�����r�gH�co^a�4�v�G��@�J�7��s�7 ����pW�C��;���	�CTH+��0�6�p��sd-�#�ZpN�N�28*2
�5[�<sT�y�p��Oykh�i�8*��Kz(��d�e����#t_ҺX �h���b=iU	��*�}���=�>���X����>ur!��~��=�+�Td�un�,R���<.$�3�6�8o��Z����?�!�VU���=Q�t�����eR��a�A���5�$�?�˨���4㮚w�)gQ0���S����S�-ga%�^[��r�qȕ�l�`ȆRm�m�z�D��'7%h�g�|
�D���\#�qR��8�����a.G��:�S@��d�a���/���/�i��n3�y�i��o�Lڃġ�w���qq��xßÆC`�A"c|t�\�I�g�gy�ns���e���ڒ��Vs��z~4j	D�<�tx�C$��Tԝ�'���h�hpΒ��V~�#.�Ǣ�s 80I�6��s�&�.����h瑮�����Su1��=N�-u��7&f���(�JU����N>�i�k�N�t�ϧ	����uo�]�f&%s��D��7�l
S~n�O�N���a��8A,���W���ꠗT�_a�J�6,�$B��|{~��1��vv��*���?���GҜ@4c�������R����¢ ����ځ5<~�T���'k� ��J4Y�cy<4R{Q�E��VT�S���8�#e�¦�ҭp1��R�u4P��X�o�\�ʆ*>ÓC�Da��dl/�]�cD܇$N�����)ֵ�vZ3�Qt��x�����F����K�!}܏|��x� /wKC.<m���9_���db��T���vJ��AS3G���ݕ����A�/!�3�bT��Y�&��pط�^�*T��]�� �em���F�p�=�p�X�ؘ�F�u�n�%x�bl5��:���.��X��Ѐ�F]��V+�ɾ�ɝ>}�&_]�{I��,|팀z(H�;8��nq�=�A��|�Q^�q�ڏ9�z]�Ԥ����,��R���0�/c2aQR4,�����Y��[85{�S�����85�^� ~G+�a��M���g#���L������0Dȗ:����wG�V�¿�ʭ?�@�(����|������S)�c��P�k������u�ňd�'Rr�� �5u�N��SK�./w���+�}��]��Vw��<$�ח�O���[��1X�o��V�2Cv�_�����_%�)H/S�_=����P��?�'�h��>��h�5�����; 1A�9yCp�op _z�E|�f�S�.�ڰQ��ɋ�p\�!�|('����o<:�oV>�6�/C��BL���Ů��L$���t����M�?�Qp��h3.�2���>d��OD�<pg�b����f�O�.���b�Y�j��T���$�U���0*q4�i%}^co������R��7,�LP$��G��QD�� ^���~�@�)#���UN�������Z��f��e$D�uA�*l��Q?�
��)\�;<&�]�J�W��*��N��[->�酭Fp݆Jtq$%ny�&F߫��G�w	���7/.U��҈����P�w�(���W����g��1$��)�D��q@��ȟA(9�-X&�+��P���C"9�4C�4/��!5���뇓:������l���~�_?a�D:X�tE��"`�&�H�b w:��1�Z����si�<0/'8c�����h}���c� ��Ԝg�_�O���́��o)��_�r 5��F~y�ٜ@��5���Z�62�i�n\ ���̠���1�4A�����Y�N���{����+���fs]qJg9i�E��Dt��Q�ݘmw2ԇ�>Bc���m���s��_c�w�ޢ��Wz� ����~�}��X�E��T+�.*l�ln������&ч�{]�^h���>7�ht�Q�[#��݀{�8(;t}Z7��K�z'�p�ݖ�/��6�5O��pAY���1�w=� �x�mr��eZ�I�z��%�8�M�ԋ�b,�������PD�`o�-d�jR$ǉ�b�Y���:�2�� �Fm�ƚY�������~͜tl��{�Iwx�W?*�1��U��o��E�Kv��Ԯ��ߖθ�q�f�2P���
.NWm�>���m��很�s�z�2�"�8�p����*gj�`���Is��k ����<�l+�f����0��|�J#�=�UK�����qZu[߱oP��_RAċL��W���l�t����3�����p{}����]�j�^�ś�z0M��i)`�>�]�to�hs;�\���-#F 7������)K���n�')"e0wΌ��)I�"�ؐ �����W:����F�͐���D�k6*nJ����u?���2���G��^`�~��W5�E$��g��lɤ	��̘ĉ��\��NW�ߜ��]k��&V�u'm��xE��{�q�z�P؈dm@�o�	[s�m�jp�m3��PY�Ƥ�A�<ץ�*g��jqH��XE�߭Zq���\�1Rz� L�}A�<A�h��^$���	�&(XA�M���������;n��*'�M�c\�4c��xL���>����I�gd�	#f�ͻ��D_��:q���D��
SAfJ~����X�GZ2���#\�p��g5���KA7��WH��ِ�}�*j�	��!�f���oX��m�ȥ:Y��ϺHa��U\3�0��K��E����<��]ܜ!e3��n6���-����Q[���Lhs['
��;�)|��6��[z�xdx��m���H-�'�=ى�um �nA��"+��k⍗�������G{k���U�եaDvݠ��5d�#��i(6l~00E0�Z�dd�
?�o��s�0�.�V�0�g.�5ʎ�n����!�;VӢ�������^��/us��1���&���q1�3��b>�K�s���p�j���ʄg�*"�Mkm�V�S{���>�ݽ�ٗ����.�m �A�7�vK�ȫ<(�)w i�w�(t���/}��f ���-h�2]j�7N�*�[�ȫȋv���][3�P�F_��9�����t�蘙%����C`Y.o�'��_/���� >fWqb�_P�'�n��.s�è���`��*��'�z����B?���=�R~:���<�"Z�#�W��PO�[���f_y��U����5&ĝv�ƭ0���m�2ѻ��]Li(��e�կ�����Ʋ�VP�W��-e#�T�3xb(��������[��Х`l0��ك(�1AN�L�b5�Ƭ��6���� -�
��; Ř����܂�2�־%]/�����C!��D,����/��NFl����s �Ѱ�tǙt|좤+�yk�ԩ�1��ɪ�m�h��?$��k6L��*�C�m<q���,�ר�l���
�T��&EE_u.6���:�
��q8�}��� �b�`
@���.������9O��SNy�96_F��LO�C�뫮��1c�+mM%�ލtb�/���n����nb����Ky��
��B�L��b��d��= Թd��Z��Or��>r�b�kr�Uy��]�*
u�k��0���U�������Y���`N<F�c��q���Z˵z5��^iD���OK��,V\�Â�+�N�By�w4�)�2�?6�m9I9W��G�oK��PG���j���2ޒ��bi&p�g���"��RҀd.
��������#,��m Gzl7Sf�m��I�O)�o�c�sJ�g�b��ݤ�����l���c
>S�v ����l�懆cH�v긩�������J����b<5[�O�鲎��\���u�Kfͩ�:�Z�C�9��U�I�+����]!���z��tq̧)y����I�չ�<ـ�KoA���h`S'��6#__y\�V�0��6��A�L(���q�~G'kjy ߢ�[���z]�--,]?��>:|��}Y}2>�o�YG�!���֨�f�nGTH)�v��x����aR�݁�k�q��C|��e��{�s��!EK`�}͖eg��ܤ"��*Ѵ1���[e���p}���=��Ƀ��}��N���B���HB���R��d1��=?�|>��n�F>},����%��n��-0؎֜G�m
�i}�1�c��H'~�p�5�ߔ��蠔�p^�p�+rR����T�a�4LKv�'�4��
9.��]�k�Án��ׄf�ԅ\	<׍G�qI2��t�������ZG���s�)��'��~Z���@�MQl7X`��VR�0��q�9�yz|��8��������	��9L�_΄^Φ����Y����� ��UQ,����  !0�-���9�'�܃��B�P,L3A��|G阊`��W�o�+ٶ�Y>iOIb�� ��=~�'��M�1�i֤z��֘c�;�:�-S�����q��S�D`[v|���_�:�H�Е�ؠ���
H���p{�Jz�o/<Ѭ(�|M�����ÃX�1�a%���9$��� pہ�7��*+J��lo��JZ?�̼A�$��ֱ/����(��y���+���_�3L�05�i_	[�~�+�������g1����7+"h����;��W��4����Ϻ>�5#�]�IL�AW`x�b�T�n�A�����;Ɛ���	� �[������M��v�wp Րa�=��v��L��0k�O&�X���0J)�9.�CBG�fn>�{D����1��,��Ѯ&�qR1�2��Y��.>
�.� 1�u�-(7�_�B���@�JIB�t;�
�VB��pC>� ��aght�w�"����3㨏�m�甸!��+��D���V�:�v�U��[R1�qu̽��{�B\��X���g�9d+�^���[!��|��UA��G�O���뚐W������2�G#r�z���� ���q�5r@��Cr�N��Siv�v��? ZA5 e�2�怯h�wY�,�hy�_d�HL��%���5�#��*Sj#��oL�}k��g�E�a@BI��7�;AW��&�aR�'UɆl�D��>kC1�W�8�vԆ�d���J|�ZY}���q=A\,ϳ�n��ϟ����ߧ_�b��=T�`��h`፸��S�R������f�R���_&�Sq_#+ሩ�����!�8$�֏A���X��]�TA~�n6Ԛ����N��'�"��؞�<I�^�ur�{5۬5Iz��!�.%�U!ͿR�������S4�V��:���6��3	�w��/�jLZԾ1g ��q�]i�k�Z,
E��	VpԀ2Ө��n)�ް�рhʵ�@�{��1H�� �;�oö2���WW�m�)d�a�P46I�U�� �//��F��^��_�eȫ�ҫT��з���W:Ԇ)@��b��h��:�)Py���^A�9��cX��1��W�ilW��i,Dj�>A)g4@;�{��+�B�m&@5��W�ߥ�٤���>�a�-�,�G\LG�
 ��˃S�Y-���)k۩������m��K�90���D�C��C:���'&���fJ4$A:�ȞNZ@�:B
��{�۬ӡ�RS���DU��!����x4YOmw���H�͘�g���Ϸ��,��-�%dB��K�_pΝ��s����]An/���-Q	嫎��r�(`��{�x��_@����EF�"�Z(��2�Ԍ�2�"$��)�H��~��e��)ݫ�^~�M�e,er����S���@+4F�A�m�����D�5�FԤT��;}�SWD��En����=�KBy=�е�@�[LDۑt@2T]�w��2K$Iv� DD)9�XS� ,�\���m��D��О�L��ƜnA
l6߲]y�D�+9hrU�G�PS�s>\���(��2�ϡ��vm y���2d3��� ��ʱ��U]�30��g
�s�f}��+T�9�`�h�g]/���2'��:�*�X}�z��Y�:�0[�n��h�,�n� A�����5�#�ww�����by����G�^E/"�0%
*nrz�xa��R� ~,ׯ���`���$+8��a��F����\g8�H&�e�	V'Xg�2�\`��gFMF6�U�9��x��­���	�-�9a{��լB�4���������B<��?["���8�5Ƙ�7$�)�;F�	��Fj����F�ܽq�K1�Z�׊��O��j�빜���"*�mO�\��j �q�$y��*c	z��������X"�w�ݛ�ݝP;���~�B��� �~^p�D�C�3sblQx�.��}7�����>�d�yZ]2|�"��4~"q}������畸A�Z�!d�����\8���{�n��c�h%X=�,E(?]5=��;?�Fc�S��/�J0"�.��Ac��-��ލgl۰��\d���xr��6�=��< M��t������|N�������Rɒ��N糬�j�'u�`�So�{�XY;p`�SW���3�x�F�A޸��b�)08S���Jj�Su`�u�Շ V��Jp�$�:d�Tԭ�T�6o%�c���|���A1�����l�+�s[5\q�����0%�(s�06���R�|�܏'�?��\o�6�G��"��g\��V�D��Z.n�?��Cg���uMHȑ��a1�!�D��!<mb�����+�%�I���Xɐ��Q�oF,���K�ȣ.�B�m��FY��Q��$��ӽŶ������R���$ݪ��:��jUQĔ/%Z�[0���N�rS�1*�zI�VFibR���D��R?`�[_��z�-ްV��og��a�aA|��%E{�s�|�.y��c<��1	�^����J���v�+r?��O���%��vz����<���*�#E*�qx��[�)�Z�66*c��.��C!���\�K��D(��|NI@9���ߩb�
d �35�f�{M~:P^��A�X*�3U����k��F��Z����@E*k�6<|��fp�w�E�W�([pj	=���e�*vi�}5��&T����|���e��2�� #�]�i]��z���S��
 �\N�W��(�6KJ���h�w��%���G"��4�*Ùf}|�n�/�!��񻨪�K�GC�ڃrw�k�iPy��~�ǆ:"��;�(Ԫ���S��HK�G��A���H������PN������r^�#G[Ȅf�ܘ>\H9z�'F����L�� �=�{X�R�홃pZJc�.�
���s��H.1�)�N�^�^����n/D�ymAx�#qMqR�euƌ˔��Ĳ�)���3,G�)���r��:�6VacW �em�<�V�k^�%��X���v�1ߓ�w��eBa��)��>5Kv�M
>9p+����Z#f��|����;}\��i�o)�4���z�t}0�Y˸�߇�r���hW,/��o�'�'tK�HB'g���Խ@�H:��R�h�����B�ᡠ$�B��������ݿ](`���CI�E�U>�g$�y0�'
��9��?VG$� Y���`d��E�/b��$.o��̍H��������	nd[�`������\8�9���x�G\�6/+��<�&8F����G�
4��!�"}�e3�aA3�y��V	�2��xGhYM��]W�&�Ϸ"vC��|9@�B�� �bȴ=g!��.6Mq
�}�u��y��h-�U\}������	���