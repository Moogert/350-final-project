-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0pArDM0cvf1IWxyHigr7F+wJAhncb8YxxXHYCgEruEx0qTDMc9uBPLEkYbFyHYMX/sOQ9hHzKMhA
oZIXuVsKzQzu1rGBXguEfEJVUsMQMbb47csYjZSizWdQGiNKb4+oLCcVo3+AKjfNgIFcJXgfD8Pw
OPc+1wuz6SasxcKyZbwVl7LKa9NebRNZPwf0U2WfnkCJ8sXxOjeCrDXhibVCO3Vx/wtitsbBGkoa
sQCbO1Azsy01YYRvMBqss/XAmcouNJQzbPPBzC/BA6fN3NQASGyBrmHTDdo+7W/zCzP45XvrJRJ8
9/btXSEbIOeJFTz0yOqub6ZNO1Dxq+6c/q06BQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
6Nxjo2kPjIUi9g0b95WlaKmxIHTUX3S/MO219fgXnSUpW/mCH31Gwa79fss80oOsGOyWtSKUmMyS
kemFHdkaIi4WVmf+av7USM2HR05S6EBdgJa4kashViZVZ0icxes/vSJfD3CqUwNeMLn2Jc7sUEb2
/4yuzhA9OrluTTL9DVAXJZe+AOE/lS+JHp+bDz6GBZUi6nTG5c5fqCB7Xr5DJ29HzH6/1IwWnyJX
xwx49Vf+0VDTObAKLKBN+a/M4dFj0i55V4jeWqlaO+z9EEOw3pOp6colNA8VuoasOFJqf4ZBksLH
oJARG1dVSUmZSG7TQZWuIWz0t5D/BkLVQWjTWxwHDL8majRy1vbPT4qn9UxQ5URfaBrX3zptq4JS
eJ+z6H6oc4tZ5FsYvXSKPxE8yON+SmCQS9TrpNXneM50rTPST+1TnGiLSlagXh2peQPKVEdsNzGD
bf+RDEWQ0qoUg96ZgBQxgOOx2yPMj9rQYRqaO9Jrc8o9YhlJuypSkDjQ/dzVFC3dx5PUSBJP1DvR
nEh4J/gol98E0xFeFdQIhyW4VMOGd8nFyQ/VXUvm/Vy8u3gslElFMoD2zECtgnPeW75GbVoPOB/t
1xnR5A+QsIKlSJZ1Wl/b0f36oiFbJwPw64EbLwCULDQaoV9qtuENlVUA21CWCVUqtBj8OzzF7vMV
JVC8/17CDzq3psvySdhAmKDa3A9266jQzxe0y2a8Aju/JWDn28A6EdyQsd84gi93+ZgBPojzAuOc
78/1sXXZRjnwt/n9+vic3Uy1N4BjME4u6bnsekiyA2hniXnOzQkQYFwX/gbjBECZL7YHbcgWlx5r
NzSniylXyGRpvCBZon+jCJugx2oZvLiPbCBKOIRZAd7OmuDQOBoq3e25J2AVsAV2YWRkgvZU4kyC
yDX/UusAJCsptj0hMdtUvXFHOFZnCxOc4uUmZDWUVFS6RKqk82pChnn39v09c+mkQIystmTBEHTB
PdgHwfYoYLLbU66qLv5wkAdo3JV7u1KVCsvpDP5QHi8wUM+AtvJQ7pY2MtLfz3Oi9eKmwY7Rb3lL
R5wQvRi7qCRF50PjJ693/F7HqN+P9/m8W5UMwT12TPQR25MlLStX7zlgFnXUQmwIFmhtVDC+Ubem
j023pYuiY4hCB/lFWxjho/fv7gc0CbIxnvNgRr/+TovAAKwGYuxvg08CoORjefwQTJKOF2g4aQvc
pH26OkEpk8AXgawDlJtlWKTsCbOMuTi33bfvlexFglWNHb1aCXleSBpgPPGk4gyffjhQECJdvSMC
IXqRYrpDAHFNDscknOXDNMn0EVa5itBWxO1WtpILQGhh8XAJvLMe7BWB8MRA5pSZ5DHlk77zm9XY
rMMfoIPMkwDNG2mvQPnemLMqEGDm6WxmkkqhQ3ySnm4kSfwCBXAkUsc/+Qk6iur0sasOevXd5xE3
y2ihOMs30GrXLovTbB3F/6Hy8ia/QtxoDFe6L27lM/NO4erXBoeyLpEn2ysAzOpoiRxCC6K1u5Ya
qxUbMtXLyM1IMS0sIXUujE7B0URDtS65Wuw73xxIWIWAkAW5Zyi/isa0+MR8pBGh8HhlzUIsUsBY
+dIs5GsZZKj3SfEWcm+Kk9vOPlhu1UAIl+Z80hN3AMO/oHsBEgg5JwSCqv210EZPjR6FGrSNqk7i
vce8ejjUyoVUHvZ4wkU/nidQq8kAXVharX9yCtcxZ801fKesKSmxTVW4VnRtkNJUX4Hzwojtt3Fy
7P/O2th8qFa6dZJ8L/oWT9OcnkkXhoWMtVoacyVEhNUgAQYW77IKKd7ZYATcYwAkapHw9l0d42eS
8bAyPiBomVHAcPBo/ZiHNJrqAKOUxR5wjt9w2XMfmhezGEnyWv1bgbaUqtOS5sf9c58egLLEhmFv
Ce8TxYQvWALsLWXLVflymx9l8zuMtXTI3Mc/9tCcAYIuLiKROa8Ib4nPhGVLpNnnbDnz8VHR/19/
VT3O/9bWfyVzn8HKA5fcoXevAYBOO+aaL+7PdK0N1PnvkY6WakL6LbG26aAZPgL8J8hYhdwBhFkd
YIh8F+0M1pNx2yKRfiLgYxLSlYAY6+czkt5rKcpLYPPf1l9bNl9pGvqxA7mYNaoA0jzHjhcvGGYG
TZYZdvSAJOVgGbo292ROZMPuXSXPrYABTDOo5WLosEU7RcoBkSUx2EtUbLXDvFGAwzED8Ym80CKT
bcmq1KJpPkAie1znO0kuByYdof766XvtO98MDOgPdG29MTEAsIDV3Dk57Y/uMTdLPOhm4d0NlqOb
XtHdF0TSd20s7cI23kBzrqUU7YiJdM+NlW0Ht7iUE1NcoXzWAKrtYywfTug7bNjdZmiT0WS5HAwM
HFnuC3Q0u8AcvVjBFsZXem7yJADL1kSEHyUbhALeF7bWmVjaPAoa84yuly6ECKdUuzFg28zxCoJI
PtByLjATHMvs48DOoiJsRq7buhU1c89kXHY60HVhwBwZzDbQW3U2ZQ4qeGXZgwk53J3uvlLyzSsB
Nz1M8rL0ctMeXGscxISEaPncybC0f7tOC0QM2sUINLuFL0dv295/KIo58ujqVpEPExKWDVsMlUwX
SLLkeCEhk7WfrlkItNJQdIPb9q/YET+fBRqtMarOzlBtpilw49CfqW2IZ11Yng9E3aBgGUEendxM
LayqGixbQPx74k+7MToodKyvTM3KteFC6alj65RU4fOvyktjgEY74awWXfQ0Pg626ZGUwfWHQkXd
6Fl2jQnLdxKC+vFt1vHUWBGL9L6Lzc3HyOIglACSSmggzHtIJtsUUuAcg+LxmuXov+qlY085Vq9S
0gvd/FAZt58RxhCPQfAIvMClPf0ESs0cT99rwCw7xBfG4lqsvhDmKTNQ/dTB+HGMHNmzAPddgKVq
l3XpzXOT/+3AWEu11neyJ/CTjQvY/QzWoqX6dy98t6qfiW3kt71hieAAUkoA9bzTjEF7P+6s20QX
qknp9/XnRTlyXZR2bUAyr41ARDtINPlMn8NSLLY2a1fYS03X3se0tAH/+S5dDdEX3hcp7+BEMa3x
yo+jN4lEvKwHoYbjO0WjZQoWhXG+m8idYHZYJ10EiNNpopFO59AtgEarT6WcrQioxmwAClsRQSeN
lO4okkXdGakPNOaRsDvu8FYgUxfPKzp+obrHftSxZ8/xkncsjxvp3hqRTF9YGU9F05W1EN0w0GVJ
/lrxWb/g/1E4FUSDFTnpfN9u4PgPyTJ+gUWLUsl4ej48AdVdJNpesZ8q09vdCqFlKbg5x6mnPBbo
QYtxP2uMc4qPBc1CU2jWUg0jeV1+3VZjWy5Vc5pAFRMR+c/TOdmPgXKpGIrkhpQ5wnBMNlCxz8dH
uRQ7WV3m8EGY0PFwmCJbStiI5NaM35ANxazFyGm8NpaUJBT1mKNgpRuvw1Z3FrZWyVdADPYRILeg
4eZ8WEbVU/i27qCTCabKYKz/l4Jnx1ozR9sw/QHAobbtln0OWq126jaK4OJXsswxkLaJsgaY9IB3
5BKn23TDeVWDTUvPbeAjiClQvYwHgzpx1nWhkSHjMnsxXs3QPi4kGpbgqXzHPmv7nkDBLFIkXdHa
+7Wp91wgRvcEyLmK1+Ro6OlDGa444cLgjDe1zvefsd9UB6lQWnRaf7Az0SHZaFr6Lw5z+VCkaQtn
YiFnwuCqY6ujo4P+WbtmnvHXkx0qg/aMI+pWhVxZUjzF1YQ8JNb3P8iOa1x4q5bpiXyr12qAfFMq
5BOzHj5Y9lBa64TfQOJLAbzNzop2KTM6qk638yd2SdH2CqZ5KoAPlRe8waomJMYDVrg//jzs7Mlg
fUMD3Q9dI5sxgAMwfiILMJylFC14YOFNZT6kCwFRg0FgSzBRvCJGiGuksT9S4XX1ORSY9D8hZKPo
hLP0kDHRQFx1PYiEdNHWd0HgjuT60+CO2E6rcwkPeiVpHawqeTiDAl1ag5NTwlU5NH+I8grNYNBh
Aa4lS1Fv/q6YJzX0GXO8llQuEfjysYMTab52nF+7JLVKn5QX2BHrQnGBHCxq2TD9n3eGOQboE9Gy
62fwtWPe+kBue+0blpaLBh0THTvwvfDKy3xaOR29dAQc2Zj8jiNhTx5/rIK2Vn/uTU/sIqBmGVVN
z4wM/YtLYa3iEqNpYwaSi11BT11miOuYNq4h89XJ36plfQ0FHfaDqiWsVQZxLfHoNqyLYq4EBZHy
cFOuy9Dgv6LINrl81Sk0Tt4j/NX1y0K3wMlf3M6VRSl1rrO50ppVvqCsuucv+M4cHPJqcpWRXolw
DMhzsMgzLaGlSEFDOL5ZPUqGogEDDKF0WoiqUByfwQ6+AhLmW85GR2xiPScw079Dd3t+9DHrID9J
YggQRh7NdXcxy8OiqZBzuPPPkqlM4UsYgQl0uv9bjFIqliSJLpAD9kFCNF52SlcnLkD9BHD8/Cxk
TWmfS3Z2CaIJ5lHLd6u3qPEBmvA5kS3b+EDh8PmXUo7etaXZ1WKw4Dh+Z8CpB3sVq7ma3fVJfSmr
xIX6F9vplkydHAfCDf0nqzK2tLCCTDl0mV0rd9LNSwuZ2b8SLvjvtn0lap5wyM15E3K18ph9E835
6Bw+scbCxkXHK42cJ2nJMMxbM9Lrp1VMLK2e948eB+n4T14+nsraPW81AWwsIkpxXh2Bj3JTMRVb
kZDbQ/Xv+YzMPuvBxFlfi34Pt3IWbSGiqV1JL/v0SqJ9HlXpaQxzfMOy6Y6f3nrfELhTbZBCTLJM
sx69d1wyG5ua3BCxLxxp2ConmQAY+cf0o+vkE43ifOq3hPZ0bVBDs9Xs/oJXXWseszWF4zDbN1z3
txGDtbvk6OobSoRxfoY5BHcla7ijTPb6vmKozk/e7hvLYtspXoy1XydpYJbz79pbxqpibcO8Q0Gm
XospGrbnVGJzMJvtwgTWLtfgXvZxQYFB9OOiMFDuduzze8Qeixdn2FcvdgaSPUIEBG/a4uYH6e9q
1OAIRdQakvYYLebXLLuG/GY1zHydfAypeSZK9XRomfht0wMMaHi0XIHDCpIwVAr5pJrsc9+XPrrO
53ZMEVnstOYIodMfDSy/Y9ylCCv42aWwaS/mKAripIxtG4kiFhTezbQq1E8weBnxhv4PFuZ+jdXo
IGtrf0neyJNspe371ODjtWGHUoJbfbFVIc+6OHGkkqCFPFzfEE6baxVcJbUgq24oG8+VNMUmOwVM
fF6UhzmZ4aYEO1Cci8r2S8TFDC7jH+/V313asFtqyaE333V1HfNc+TkY6fiIqAM37V5eL7uObssk
X4Rlmj9Cpt3qoh/20Hg0iAOEfu3gCrUngNIypKbGOI6kPg4SwiBbfVwd1hfkmapn4DE36/okA1MJ
CLB5ueQpA5ieWZN06VeJznShTYb2MiidAN03pKi5YiZRr7il5XLCtdNWQpHHGLS10os4FpCyuJdi
Na3ooA0N+Y+zWHtxURxKcT0hJV+aIHWhBuLORC+yDqZQ+kGzqOtgf5rZyw0rSX+D9fhgeGSU/4Ii
LS0+xiuOhlrfHWUWyAsenSEizXlLbSoXyzLcIH24/zFkph2macH2tNRP/H1/Q9oLlq2M7D9VayV/
ZFm++NCtumJQF32EYpLTlqPgjUb3IuqERlCyb8j7qSG3QSpe9OA8NlkMmTKid4Iu3Jk0/+ezN1uM
KvgeZAnDN4NuHXAqUbjVIIneSxob1d51LiGHhMXBoJYprCdgbCsnpvoZVFTdhEjm5M4D0THK5zHG
EYfIHu+pP1ZaU8hv3PKlvo0lcz1C6g/Coe+GkoFirm1xNaaku/9fKCxo2YKOLFM5h7GGU9RbsvlU
4n29rGn70A510JH/K393hv2Ce5BO6qxZl6KrmkhFdoKxpOK67W95TSLxRGaF5jH700OilVJTVCWI
BUBva4WSQzBvKsJhaTUKmk/o3i8KJOFj3/kENs2lfWAalRNCWea9tVgfPaPlVT2IypFklo8RZ8iw
sitqGyPeoEGBOTUnKOb+wlztdXcdvxeAGTxk7IjZx0Yi6NP57oaABxmg/7ehwKYwcBipRY2ClfH6
bSDQN3h0xjLIKK/m5s5YG6zx8LKfRWnpBqaPLdIFrzhWKzy+yTfY8Z8FtgY0PDsAUwHlMB823/Mg
JuK5L90kMhLqW/h2eaPZM5tBWAdRzVg9k67wO24BYEYIwsOLgNaqAFPiKA8NPGIC1PyUJruFzvum
/4SV2IQOumKiTOmdc6RpDk3nsAiSh68d9/DQjYppIpue5zrDTXDq1fpn9o3v5UxfUi67pEDQLqxQ
FIURlnP0naGWaWsxhpAZEOkjoRQkWq6v5tWVQRhAm0i0RyUJm3FK0OZmkd8qmLFeuwoLdUebAcTB
JjhLIg8UAh8CDcGsDQFB6l9RA16Biq+i6lHj/gmCMEcjyxJx623TVMWs5LVBSfkY9bSvg4ECFB0N
xacg3fz+3W70fMJuvmfpns1+9LC2O6d0YXp3V5NIaxoFf+395x/eD/n8NBlFeUFhDf2O0LCjTGZF
LIXb75Ok8qU0+vwocNDv5QzEdyqjf0vpzh1bkG7kiYZzufqBHwspff44y0yTZoQV0JJFuu9URbDB
DqznPIFVsGLt8Btpdb0aaptjFLWDlUcIugbUX5NhKU/VxcDP5mMTdy+0UYHVyT/pdkkdhdVVeTEl
i1f7PbI7eBn+/eW7dh/hEjWUquBG89W6jiGzzvoEmBMxvnwaJX7DM98dFFvOy6eDD48JANpWG+Yn
UGW6bVk1SMfa3ih6mhO6qujCT14Hab7AmwUsxkyy+Rew1RCn61bzXdt1AWb3EjogMK08AhLLJ9r4
d2Q5UZJIaZQT5A5MQZ0rXP4haezLLDBqy1ji8xOf6bim2/G0inK2gJxi1qFt67HvgyIMr3mmh6+C
lkVwJI6ZozbepXJqYgdQrQ1B7r5gwAoXQb+kmYYU7yGdRzRBPyKVBTMx6EP8HCCOscexi0PVW0Nm
Dwu9AC8fWweHx9S6j4LYL+RpSxjIZSiu4sRrLprOvGEzRWUt5R841hT80ifa+oCMMOrE0jBq3A9W
etUKJz5p4Ythxl2aTe9Si8Y2WXEM/zxPwJM9ZI2GZCXt6C0jClXJiWmkATLAg7MsmmNoD+eZsPqi
4qQlredeP7BPy+gNI/E5K1fkt2lfFA2FMS7B04zI+Hyc41dkmygt9Pza8EvHKs6dmR/pS2RONXH0
Ac8sJOkydkU+d+xusoWv0vLy51GYHn5GmgBq/VaSGXvuwCaptswQw5gCyGF0bW3vLd112P8SVGBF
JS8JycWfw3loDEQxH67BQHlXTVomkmVB48wRnXF/nAP1aqXHAzWBAfKgzK0cueF3qiLP0AjKTnRS
tG5Tkcs1SXqVK+hAXi6qxD1rdN48eae8w8jtxQ7K3UGLH0o7n1yo69yY4RHARmAUfvfIo5p36SME
64EoGcOU26hp9oz43etkkumUUbJxQb6hrzv/Gvq1PVzXkoYFGhVibGjgQ/5KZZNGu8RMpOGB5vb7
jtOKqgiRxk9bH1D1SVFwS5GjsCKaOdy1eTVcQPtc9MKTAmsh003OzXewLJhQpgFrHh/eF3rMXxxo
hhwCMlWWttRfwJxbAE959u4hWu3UY1g9pq+NgHyRrLdnr+4srgcG1uzCk4VtGHs6Zto6lxYIP9o6
eeXN/5Ml7boK4c5JiSfMn9F/m/JpeWQ9kDRWimnJKsAzjdLP6vVlz7f3oir3arvp+2Ixc7kgKcwc
Z71DM8ITZQ1PnCJVTDvz0WfcGHyM1sVt7OJahsBgcECcO8+sdoZn/uLO8jLXCjmHmvrYDpZqGWNm
/yuZXBmWBJ2zZxJFeQaIzLseYejxPfHOlh5GsX49pdGX52re/N/NgrGUf4cUeYrfshY/ss3uS12R
15xRr/JFGYAihpm6I7cafVVlAW4ABJtxkRmb17Bgcv0Wdly+EZx3Wqvj2cLZwqbbIielJG2kRKV/
+NNbRghk//ip144gaQGmaOmG7Hbe0UFpfMENPa1hTYVSLZZPEHAYGljY+CznVaVqcfXtGLLwHyJL
N+WPnU+XLtTxRWuVRaOueG5vQNuI92b43KmZIwxXom3InJsAwSMuP8iNYYfelNq2Ja4JCpNRm2KA
sgtGAb4FPUrxSgUAApKclhbYQtDSdqge3+iW82Iyb/iQeoy2yqrmjKlRxvkF4iqU0sSGkYDBqwGY
7xbtICB4huirOjtONzLMtgkiJYkPRVsmfbb8hccBOBj1LXieoW3md5fa87LASxxVKsToHNFaT1Vf
CIH0opW1Y6X/ghDG1WCGOVOjs2XtV9XfZK49ckfaaZDBFWQ6FCJ/n7xp+kkJ+kOqLZf1dfsqA8Dk
xotDO+TPtIEuKF/MlNpF/kNwCCEaSkIIhpzcc82hENKQVpofU4t6IKLRjKsda3B4wKDZ0mOHydTD
sgTn7Fj0zNE4duS1kV27t94Ew0BZrFc+JWHaAeQc+kMboDuiGu4L5nDXMBxGBpAADjtMaWkTCaE8
eD7cffzDwacKqVhQznxMy/LwHCrUeYsn/tY1o9wDnEwygRuxJLNGfsqaTNN/xXTAKx2HBQQBJI+J
ceE9zLIrpoFI76jmcPwtiiq2UWHkrzEHiHXenDZoceByXvAX3guSlyTLFufjnFw5WG7GxHvtkD6g
Iek30ntse4wUDlRTIqZNjTuZLwDieKQK862oZxShA+1sqcxkb9NVqLHSPdn+9c/VgIrBQAFmYHLj
z6B7KXSpOYLX3L5x3Vexde2vt40ErODgwRz+eKBufpNUiD7YWPuJ2K2gAOb4TlvIQHLpqGQRZ6Wv
MSEkghY1YY24eDTc88eueACbYwihRKIR3QwOD8Fq3YnnbZuIDFDjTYmQmFg5eug7WTaaD/gcSt1g
u1l7ZeaBnYekxlrin0yEZ8ZJRNYV7/BCNGysRIBAZdguZllkHInUYXdTx/bsT4l+8WsnLNGbp0Nw
7wzGCqoAa6VFBe3JlyPTm72IE2cQPEMBMzmCbBdiHufsd2VUE3gjbwsrtAcWxCX9PGaC4CbIIXjI
yKxWlrttS2eHYYqq5m5mrqWwqT/P6RL/8Ms0BNGKzSsaVyDK7S/mnO54iYQK3qxlb4LqDeMtPkJN
kxyf6Yt8rQAZEB38pEGdY6hOzw3vG9HhvrO0M2Kfjc1lPviPZdDpWboQy9uNLNXmpvAV9S+YYoav
35oqQnwQX0+oW3WGykAwDGA62xlMux9sR+EDMvV3aK/IA83hLBHNV5f0dxFEzcyVekBm2djgBYCT
8PxD0P1ZC0tElURsVDQN2Ohd8ltFjYXphj+PesWhgSk1TlADO0tuHSm4lXsZpEnU2+tUTOd49Q8C
H8j2FoTXxn935AT68J+gY9sCx4ttZCEgFZ3J5n9SS4CJHtJN9bcq7TMVqFWAbKq/SllVamgVs9+b
zxl9UWVEfe/foCrv/VWivbqWGZG9FxxpMNk6/YkoinYMDx//NEtujPMvz/NVvBwAqpIwlH+uopO1
Dv4L8QycAH51eaT9fTzRHTakqEz68qclfKqyylV5PMSGZ0kJrai6GsYjJ+2qhy+JavVFsdsi/faK
jtb/fIH2/mL7qtQvE4yR2RXFRO1BepmIEQAR8onsMmTSJNXSL3MbQMpJzUd/mrMqZn7K/qyOhBfS
RL79H+UZnBvPoaOCANQBAvAKD94iTnM0O0a1vKW3jNOcTxvJthMz0odJnwvJkRKBp/qIP3O8ctpT
lux6LQerOppG/x0y3TBb0vR1W0U/UpqNCQ3MxgcNmK4SUAt1XYN7u5igQAmwsFLRopIw/8HhYuNl
JsDhEgrYaVfxuXBXYfVGVh5LYjoXqzyHw6MIH+fb/XhotCRLUUC4LkKyOb1sKMAKT6fG/t7lmWem
jJySyIocJRYbuEsu+oD96gvk9TFfX/fCW2n+lv0/Ha3jc0fEbW8yI8oQ49DbSuFvftNxU9vQfT/K
0NFpAucdFFfAhg4oGlYAse2cWo/V/idZ3P1uSgd3gb9UGMDaGRFvK0dPWFFEK3eMm+Byn5aByh0t
O7q+8VR5S9W8pNTHAKK+avdMRubjQh4kQYqXeITf5NaKOhIgcqS6gl36FyPmDVIWxT+/5CdFR4Rn
ReiocwHCPdmFO0Op2yfjwBhhvLolscVQH7r3UgbXcOqDCUfL6k3wl0Xv2AXqPl5c6OZR4xfxuzHP
RR3Q9liZEExDwYdL1LVg0Q2vTBcgU4TCw9GbYvSyyCLokS/+OuvvTxEbaVZuexXXE1Ek7kWn/1PV
cUcTU+Sritx6PqpVhJUoA+ghXU2YHHonh/8OlQlOah7BUMI1Dy72TTsxjOfFNRPNz5sojDgVNFaA
gOm/ZHTjDXOPP2zWAUFY8SylQs7HVc1eTJ42fG350TB1LFUX173PjZ/yqYr4TwkyyzVqdRL1Kt6t
kzxL1QokczKUp7Q4oyBKPVFEslmgvM3pS0+xjgO0OfjnjNbMDyEStjyBSSseg2EYfK4d25L46RX6
UV82H43DxNDVnH02PC6/II4q/3xIT6OXYgSjTn8W0AmJdec9xzBQOEwj1FiBd+ZM1XUjhBLhp3OU
rkV505o+RYMNMcpkGLISAJAaiHisCBiR8Df0zPqW0/STfaakFdOFIk3EO7pNM+IBS0Qb/8HRPfv6
H9dJpDl6H33uYNX9vr7XNVkxbFdCkdmIlrzXCaa2hidAqEW3Kt7rKEQoJtEyCsLQuumRABTM29/9
y+LFRyKvAQmpEhWum+8q8+Ny55rwxBS/0FUX4DNzO+TvcZ3CYmL2vq2YPaLRzlrT5R6nzf9fyEIp
Oacmn7VlA+dYvsKQ+9ZLeUZEK+TYDfKMBeEeRyptUIp+RmGCUbvIey9c1YNN/CQppY9/rD42OgFr
CbjeZCOYD5/j4V3sveqADmnBoJrrC1E8NUhZ87AtFyZsgSSf3Gkx0bEiHucq6f82OnW3cjzPMw37
P9zOp2Cc57alb2oFlSzYjURzNrmPFo8PXMj1LdGzG1t6Ymxza2kHZmnCl9c2/09YelafzlncBUO0
W7bNKmwRrI4n5QyKtXy+LsCyZwLBCN5Vg0w++p47cE9TjppJeh88Rcxa9S4fRMPgZA/lTCmaRgl2
6YC9IjXha+xuEXX2C/02zSvXnAwIKCGiitSbLE36PGJaxI4i6RWUNwTbu/au8m3sOHPSYsF8k0ID
2cdCuEb/P5JQFxrJAbGh+c3CoRNUaz8yyefmjWLowWMbXapNxuqi3C3va4+2xWVbH6c9hAwH6AMt
xQgrXHYuxN6gd33oXeq0BrDTBb8IUYPkqfC/CZ8RWSz+hNslBK1hFuJ9mf/Rf8ONC3/nt5KExGLV
raD+7CfJKeORMj6om3lU1e/cvJOT+ivIeF836IbIIUHNA4JnoJ/55ZanC9oMreNy4KFfOSTWtqOM
wUTvt9fYEhl+wYf8BY0FqjY9KrEvWpHyonVpiMVf+9x7P7NdZhNyF2u7F1OoP6ySedObBuwjV3mK
nk42L4cBEdzsgb9iZGeVR/geP3wm3RhMDDR+Pr41j4e8/OnetZ5A/IR0mKD0Enyitmcke2z1SwK0
Fhpg4tI30aLnPStw9yuMVWd6Wb8295ufPMgV2QRlzfEgOc7117hwmiwux6m+4QfI8j7fJVIchTbu
7YpZynQV+PcD/Fu5BIkpiHF23e09g/NX82E/Crd5yBK/wBiNfdzpSHs5OzhnS6BioEx3T7ecmntF
4lwGz85yJkOzHczMoSV1VzEVbY/gfCRCJiONq4CpLAO+T2s/WGdOauhnhhsy4rmNyKAOGfVUKBIK
Iloz1vSWFIa3lwDjIplTS5PpMZ93Oq0oTncWMSEjXMXfJohHpMcbS5G51J+0qlX4a/A7kE4EUr0A
nIPoDhpGK1zrkWnvIffLJZaQkoUB2vrN2FK5SNJ+sgnAtloGpqyXeb1EAU+V+//06omhAX5a4U9c
myZW97/QkFgXQzNFWE0CsSldv4HSqgdaNDr5Cm8zsOW5kxy8mvAAFHsQB4tTEDTM4syZhxIbRXm0
f2QxvQWterutWtmfy9C4bwnwX2dVlAu+nkpmU4zFuaYh88a7ErlmFcDpla58x9wcbBQZNeJ6wuzU
Mp4qSI2HUMNOMPfwuWpe1ysK1vjChNdg2kySJJGuWm1mHsfViEeHZTtHfkBYO1VnaYxL0NPXpEP/
3xPYR4Askqagug1jT9419tNvTMPOXXZ7Bv6OOYWohu5ufLPaefxYeJ8pAjjh6UKbznZ7fnRfh2j7
Ai1cHL1z2WJb8tjFTbdp/UwM/p0CpD5D0Kw2jP3cIWrm8y67+u8d1ru/l1gNFGbdOF3C3t5C6FFn
XLqXjiAdhDJselqgMRlZjBmnjtDRCNcUOjpD889watqSrR093pHvPt/CLV3MQISZfhqLjFEwaCmN
f3YmGie6nBIpGIbHXDUroOKy38tABLkesYYhqqhLv8qvmBdxqVoLwTjrAzNYv+NMEVdao15Q0loq
rMzdMqDly1rq2tSo1IA+w3SJGsQyx/MSeaMCPUUIyx+6aEc3lkbWA2EcztQGxF8uLjQLJ+CVIfB1
4XPUq4BE7b2+hMoCqwddVu0E1CeD9p0YHqBbQ/3j9CGdp71g7hYk7XGi5rGs4qGZtqgIBXzFfCTg
lZZjCSkiZWy1ztqAlqHB2d9BNl8iDgrc42Nm+fr3TaZ9Iz8w6lHwL0borqsdGB7O7+rlSDDtS6dR
utWYRNIwCB5ilaTczJW4dFdjw6lwtKhRubWIrqabF83NZO1ajnqra/njWs4ZUHvAXf2lAvEzAYjt
s+/+yqzNugtrWWjTkokI5Ejswmgx8WkIs/rir5J8pXm/osF2tFpQLARQPaA5+dnlle4ZUA/Z76ph
zfBiQQ4H3lkGgG9E0X2cKTvJgYVtSRpssU1RM5bGH/YRY+hLybNj2rO1WFk3jqZn2vymA2+K359N
ZpKrnC2qFOrHAACn9wiOzkBYJy3jqoGphS1yxV/Q7rfBwAX08Auf3xkMkJfLXn4JVn79htZ1ecT6
WIUzdZJtBv5NpQ/YttTnb3nPupInbqmg0mm+TCKFTP8iw6h6HBr6bQJGylmBopoLp6qRH1v9Yykw
Rutgby1qpLNoalL0hH0NVv39LK0tP3dIZ4wjjEV6tJH8Obh4Lzf4pE3cgy8SbcbnIQGzqDskai6l
yH6gRv5dQynYOjBJEAm7wh894ESPe1mZVj1iqyZBXa3Bk3CoX8Br6nD+Ps3e8ZnbFWPOEaqNqDHA
/jsIzqkmWhtd99Um5QhLJvJ4L0VB4yVvdnTa+0kNf9fUcYTNaor0aHVWoDOqzsEaNRnZgwRAU7yY
Bah+ePLM5QCb5yxEOi/ueJdhy3mUQ/9DmwucAeUxUgNJ0bxB52ey723QSoYZTkJyf0qWiD1pA1hI
NghBhlFFkQbWForVvOL0atwqdruXxKNgGEhddNRBKsS3z5PGXuR/p01+eGeDNm9/kYXOzzbG0xwU
TujrBVPvHEYo0Yj6J5DR5LlfAx+I0a8XRKp5NNVmBLSnnmqrzrPLZDvmJv373DJ/4nzo2jtuWIr1
ESTTeZbhaTIkhOKikLO5uvtKzbmxRIE1dYmSkaXcIQXZPJLzuG6LE53tfCUa3pBAArhLfiLBIFFt
LTWjPryySr7uV4WhiJ8UvvozWf1CkdTVwFShWqHML163WU5uJNmJQtKzgLRKf30+5JZorrF/eCQS
igcfj6adhHAMYTdTpEZTiA6IToBf8hq6gDe+W/47Sor7Y3I7gknh8vxiDWUOSM9p5vScln/+hj5s
xQWQiDMAjOER+xpoYXmT2Ush78s6c9BSULYNkORAR/P8qOaAWgR5h19Hydt1YZQjkpZKWWtrXh6P
9sS7qjJof/BmB50VlVKq5D0IfbHvNWuP1ue+/J+9v4eu27kYTIaVtJ6EAJKJCJpgkorxp0E3f+5Y
pGS2KDqNjP7LkR4MnqFeYEnOg5ZeX83gtYqSvNu/w+9J4R3NVz8X+bzhz3MWW6ELcwsWTHRkavVz
MZvtKcKCIzepljGO1uGL012+cOpyOjKHJEYDIG9VINrKjEM+s++J+lFBkpJ6KeoVvpE7G+SuqFZE
ekcC5PuvLirBZIhvu/Sd4uy3/0C6SLVy5L4y/szDmROfrMGK7UUgMVuB8cUsvKMc/pXFf7xL+w9T
hOp+TP9X+Q+eNACO22fuMiBMZS7pzuEwlCv2RjdN2Hbkd9tmwqepcVU6m146G/1twW+5KZRBI7On
5l1THc201EKew0RAWCA5DoN14wv/4ZkgUUpxYB6NrC9+RNExUAlW3asFHqkmBo5C9Qkm0WtR4fFA
NQ235Kro+0L8V9SzskA8KHUQMlKF8fmwvUuxGenN0CG/k77aWzU0r2LiDafaDnVEe/VFKoCbz/HI
WfZjjzuFkseHXR5F8N89em1VHSNRkmv1trJxgY7urJEClyKUIzeyyRxlCB+k53K9OB7exbMnPE6h
bfqMInyZRGsrW9PlPmH9KhxDRH0v+x025dTxSDp14iVx0ZKJn9+y5K2rcNC0ngQsn+xpcaI6VTjP
Ouz95RqUJotTvlqiUJ+USbAD2dfkvER+Djv03VCgqD80P6LU67NZRtCwFFlBTg4zcGy4fF2EzTJL
Q8gHOGLhiGueig6dYolRbUYhdIssXOgroxv0sgEX0JstVcuR3FacZHuL9tLIS7u/RgAeA56FAMqh
2DKtFfBXJSOzXI+ReT9lwdAUumZcGbjbUmVdwrhLSBJ/nfaGhSEQqoDy6bJ/zlQBEGRK5QLILvuO
sdkcfkOdnhDxMh8H/oJRZprT+MYSB5IORPRjKqvXM0+gDCfcEUzEoUTZ71TKpDvieBZzEucPzjfz
1h5TRUJrEXDXfL/91c133kctToO5Q2jZwvDFSEm7ApYJcf6uFXazkioqtDsHkjemq8myrpqF64pU
70Td6Mr+PeuMqO5iRaVbH7jd6Ev+Rre8p9ALB1cuC1WpLZuzC6AZ83zmT0/WtEyf+Mwz2MvZvU3U
H3ru4Qc2OD77n5Oje42+Xlp5vwVrqii2u9Bd9VMdQNm2k5zaYWVdfhskRsGADgCRQ0ur+eM9pB6Z
0EKeJ9x061xzEWc7wY6+tPPR4SJWf0wJz7pB/6dtR7eIcRCBVtXSZd8W/FyLv4Z9FwI4WlrFLyvu
EiV3uX/Zp9i4kHNnH16P5rz+pQFFNiiu4iwSXGxwIelXk29Iacc43EGOcy2US5ZgZ39HPZ/pgKot
t0r/QIUz3Nl67GBE9/e634Sk++GzAMaNRGVXNaA9Q2f7ewqEPC3lHTxCzGNsFGoh1ynb0/V0Ny+1
IEFjZG/aK97uUvKfYnvsrdrTMxKEn9PI8ytPjL4wHHo0r4qYTP++mL/4bSu6LbNQk8qn5aIPsPy0
tFVAxKaMaJd894bQhzE66b6B0Q3MUC/LmE2dma9IBEKqZnGn1wcxw9mz62+3RwYNEbu1ofdMHdvg
86vtUtWii48S9gKWJnmU7e4BGMRgRkNE72RXX+ac2YgicF4opnNIGL/wbxQGVDKT6LNf6LKRZtoy
3S5Bonbo3IGaF2Yn1U6I/mbZOP88LoZEugFHcNLly4WnKRpdmEtWetIREYd+7sYjdVppTj7zTA2V
+D9zhAeWg8pPnvOeFj1upOzHq00enZ6qWY/MlYzSaUQIS9IEo8RfCnIkmK1iMNRA2fM1rJ1VoHKl
qGelgpekiT6NF2LaesV0n6Ut1O6Fgr7UI/qZXbLvpTHv7/MAM1a4BBhQMe4LtW2RBD03k67NAATX
Etkt3R8Cn7OyNsFQInCkMK1qdr5Rg4XRCF3TWGwAhtVtZx050mxbnYOkbVD6kQysxuARG2iYpseD
FAxkYDIMYeR15w8Bo2KCyzwk89FuDfpZK6XxbAIYzPd8OS/dFkomNKeddFftX97NZuYkdqhLZWvx
A7qez+ftvCbBqiLosGcT7HHgOJ2gvBxURfQHcY3wILXXzrZVUGRBfa9izw63T8SHlJ8QaduW3j+0
r/yi+vvitSaDxC5mkuvHtBd69HR7yrbj6LeCeg20+ibpzqr16wUcUiHZrcSrWluk1jLFgQPyEmlw
kBSUEvxM3WMlYMS4WWtO844jJLxj9+bcXkwSgHc8BDZl6aUohd8xlRSqyyu8isdSUxylYE3Rl6cm
RTPnIEoBy8wSDzXnOppXvIsOTW0s9J4/40VoA9AFszZ5y7Hu/kAPKG+pO4z4HXusBQC6EbmhlXpP
42pU335itbu/oW8XjuZvbhu9jECsdX+kLdEnN+MYHZc0VXEdCXPkhLI4ObzUH8366ivHRDmhMBqt
TYZkBuA9k2+LHAI13qQFmNpxKJRG77tvAiCR1RC3k/1XdTDXvoORq5VixwWMd/HXdt+a1Jd9Vzs4
DvVLeUjmWFv20VJMP3Upi8ZgB0GF+NGwI+QfUPywmChEeqRuIC3+8/zoLLiK1+zpsfzaLQUCg/jz
qLGbVyqpXxEEBvC36YlGelPox5Maf/0CJD0568aC/i0vpI+CTGZvOnERqXYu+/r3VsEauQIzdHJk
wCooJ3e43bePV+SqiP/w8qTC8IJU+o30adpHYFT4XneOvz+7gkKyn9i/8B2pKaQqwVvQA1YORzSf
d2rjt72/I7cr+kP0Qi+jtD/+XkS7LR4DPrmek81YaQPhx7hgn/PoWLaXHobM4nxP2XTplHLLNDRX
PBRj8POLRAbx02gSkXwvhISmLDC4DNo9ffttIIiwiUDY0+v3a7h19nkwvDAWlgDiL7RjmF+UIClL
gpux58R4pdnmVIcy8utIGJ0MaBCHn1pZTdwiXKniQDfHzgpTygnoBfSMezdmxi4rLtoejresuNu8
OQ8Ps3Oj/0KDNp6bFvHNe5Uufn8mKS52zpmLAO+IQli12qX1ywXDw8mloYTkXtnM0G9P9khfQwik
4WHTXYvSYSMdKs3uml7fyc+T+lRjUDQjzfIzEApiK4dCMIq2LSlFAVKkInzYVfRNYBUtCqy8wepU
TxbrzHr7qPUViMogC33Pk4WcE+OUzo2oUF05C5xMqwy7HeN3C1XtdzLSAYuWQdA+Q+/RPmML3asg
vJY9U6SnSnr7Tnv2T1VR5KWFHzI4nJPJ512nMlMTZUWxdKAip6/aM5xmpt7UdMf9yD2bJvCDN++T
XsAiQPfKdYz2d52ukk54bmN7e3dwu7ZCkERooCHe7UhRGrnakWt5XJzFAMpTcAmBbyJWE/Hv7Ao5
Z6I04ml5VdBdQYzdfl+Km4TN0O34l47nKpxbnvvd1hzkF8Zi1It6gRjQB0avc1HgOkp/S+5/Tp8d
ilLaUF3uMUNH4iOaH9T+kagjPe4BuJfpTmwU2gHnwVlMtKdq6AfmX6V/0w029J1LD9RQf/yhxLe6
h8LmOi7bXEFhzJpYAH73FT/GBOXWerZtAJ6Xyq9Ki3Nhw3NIU/a1pDwBl1qccr/iKeAdcww3zj+Q
LGnNL3svAimHUuOxrWFHBXaXJ8Umtq09EUfRyiYTcEl59UIGvg4j6o9G5lyXL+pFYKSjft0862Wa
GMwI2NSOyTGcKfXS9MqsK0oXp6haycLv4wAOKUcj8yvPM3ya1uFoLpNEU1FEiPtR35wSev/XaV6E
svV0QoAcIJFxxSW28CvS2c+e8MsaobnNefJk0KGaaicdi76sFNGxLxwXzDI6//4+MbxNAKRESFJj
F+3xNZizJiDBUVoDdlm9bKDHzpR3pybATYRNfaPGkNG67qT6kWjfwuDJd9FocJfomKeZM05a2cUl
/ZJVodKdfjJZEWYJ8b0o/zlTlsORghAOaXG3R0gHcnQgz9A70PVgLOI7hfRpT6QIiPVcq57rQHQr
SDJseGBwcRpP5fPoBIiGilpw+yU/+6KwjwX+Y9yzzFxH+CMeuBebCs9NNM6U5Vy0JnJaX6MUynBf
D4PY2iKs1ujRBe4dI9MpFOdoC9/5tmMf7TQKobVj2kXKsWrwxjczXG8am/XT0spNI3RoJb84v+kH
awC4vdsAN9uWGBD9rVONI5wDZc3LRsM/UME42hKDaE4VupWn1KdOCIMIck1hheuR/qNS8S+SKAVD
SXK/PATreGMYANb760ID/HLhdq+su7cQeB9rIorkW5LqZ8I4wXtUm9IUlp09y2a5bsX7D6QJ/tx4
2xFWdL3/wXBI4Lc7PmMeYJikW1ct47Dk1LkpNGbldHmVzFu/Tl6BM/Eq2rTmXmNaK+Qw7bH2iyLl
OK4mMec6VWaMvFwIWYNjlY38KjjKD7rgvOdA4tYffW1LbUr1jJrYfvHGb+vqvNg3xfZKYHUBpjlp
eDsUjyAuysJcNf4BPLDLnRGs0gZB4fdShhn5GYuSFa6LyrDgdMHbLc77DpboXX+rfaBtDzjtIpJd
fSeW6fNtLlr6IaGI0jYigmNruvJe0kE1ItKw9jcy142rLzEel7zGqTkf7yOZuzGtHH1eK7ejwQ5U
0bx7p04/hyFq8F/ln4jzbw67pDTnsNx5/bKBsltIYDkZXIl92vi8loVyz3J8/mQ0QbBaobdubZSc
z10KBw87J7CvTqBYjBs2PQH3aYAzkcwJf6hES1DKLMnmMob2iZquiV4x5yCUayAoYzjlefq3ua9T
gynfjQzk65nCqo0FAusDa7cN8Po7Bn6xQeNymQY3exc4Pl/lrr0chIqk1i7YalAI6QgK2HNZAx6+
5O8D6ARQ+vvU25pumWBbMUmAqlsMr0UOxiYbZIGqOIVbXb8p+Lz1JMfdaJGzsRgqPRzsHePro7ho
yUMAqcklJ4YPE/bYY85kVTCrpaSlzslmO22FnKQOKzCXGHIJcI5YCUGi4aOsXY3mVr1iz17hOlTd
xLRbsw/S3dTd0WurK/jNFTSmVZBDMRM45DotLKepeG962awoeVGQcG2RXU7qWAiu4oz1NNaErEq2
EbQqk3Un7NZfFMo8kMD4RJGpw0l0wO8KLQNK27GPI3mSsdJT+UopNxeXbMiMSSjBafJ4b0t6wzjS
PtnFtJBTazAYhFlJoC28ph5mhp/t712LN3ru+RdAxDphkOrRm5ZRcJ01hSW87QrhuvBmrB4DcSHH
+keyQJ7Nnvx8bumURr/2dUhgpzRXUveyyPpHFgq+WzNwSKmLM6kmaMaYMsYcDjz3ln9zxVOhzF6+
PKNlmaBDPDUmixfwiOlyb4zUcFijt22d9cBGI41NqafjyBFy2qbPpYg8ro6YqphVDBQMIk2B1REn
KAZ4bWGDJU9XdMweM/JdFUWVoOYBjIkimCMqIdPrPZZdw6ip6TuAJQY30WKxVl4um/f6/pCsOnMg
SrW2coDZwkHmbm7lsVAgN9rczMXNS/rNnoXEyfr8jaRgT0Kh83CycSATFL1kHnlg5t9owWzXvFg5
/KowE3vixQ65GeAuNeI9bUwiPA6bWeCzCDGmg++0y2gx22nrSIS36nhWe6E+c12ouuCNBdP50EDd
CIz3JN3sViB2jrOwytRYhVGzsEU8bq8n2Vmy0ZpJDItSkDtO7VF/NJORLjNT4msMxsH+hwtq+O/g
fpf210iwoK3aWvV1uKsjBY+pvs0kXH6NC/qzbulYU4a7cBwBa+YIWm4aqFxJZf0HBaXtAZEpPhp8
Y1kIlOJRl+sQlJHW+KUx1mgfcvbHVesdBCxPWNtrXqJQVSLxqJxvSoM96y235hZPnO1KAY+gTPsf
f0RijZDjTbwNZj2rn5SrG1TcvBuLGNRRVCGkc+MpKUfZ+mX5N3BJHXAclBmGCtpC8K5dzHwBzkMz
dEMOdcsQeCl72TmNKuGnSeL8i7xo46KwAtDeqU2wpzTs9AN63SF2p5/WCjFvASWsoV8slXGumUVT
+4FFu8AuB2KW8BzykKwEwpWrMonNrfWP0usuIFPWioJmuyqLids3bTBAtrDYs0Ol2Qm7GINoFHUl
G1H6/58KSH/xVs8tFKBnu2bNSXLaU71J9eCGSnOkfe4nHcR9rrPwAwzg/MdEVeRieVt/mjvlRhEA
xoPu1XVYTGIyq65xjQWmjPL9hf+FKnPGgbXUnq8DBX43jZlH4lMunN+wWJtM1+NOjliKYJRACucF
VeqaBgme6fb8TT2V/KPcUJ44zVSVGz0gGpSrYx+mhsGb7WyMmXhZjAXnYKcgb4nIrYHO+HHyxzFt
M+AEw6b/nLQZ2dM5hNsRtWJxGG7Ypecx4wKfUpuK2JKhI4Lzh8BOTwB/1O6hI03P7d2vzLP9iEYE
amjLkffz/Hmu/I7R1d1IMquq4yvBMMe17HCfCN3+Oo2BttS3cxi83/vt/A0d/DPfdbSeFyAQZIFc
qNIJGx50WPmu5C+orbGGGtciEeqHitV39dh6/OebbGxH14iBun+JNy93NJdntqjODCrI5vm1TR5t
77vRA57wALCDvFvLBsolklGXkndUxe+VrUwGiklf4fNLmdypc+HJ48t56NF+9lkmAH2x+xiEvYyf
Ceny+JPRmVFYXDhjwLMqnE/3btIukTq67SZlH+76Pi6TWPw5Tngdr8LLM+jMQ9OKOSsAdM6MEiii
3p0XNGH+Nza/fFJiwzikT2Jj0bUc/hgn6/kSF2fqLGiLj1dtbqOqCNll6W9JdNEKWKeITA6nGiW0
00c+GSzH5BG/1e502ZjbZi4Fyp2YoMQFvNI6e67W0MkxQoGO8f4Q6DrGEMZ3gy8mvzkiPZdV+sb2
t/u+fr4aDwIRr6gcHIjpG8c3YwFahItcDhV43mZ4XboadG6JY8DZT1akeOhn7hzsYffsyl4vMZE0
f3Ptz9fR5sVj7pA6faU8zrs86Qii/Qg5IxU7oQgxQmgtHdxYQLtfdwFA/5b2aFksb4ZpGfHRRbM+
4imfa0fJ6HTvDzBt+rt8ptk4MXmaMydsyZPV4B+lhSvwz/mkGR6tPKLjXMwyZSSHIiluXggGQPxw
l0o032OpKZHpQs3Si/cEgkRbwtx12/ExyENwdhZKK7UE23UhncuocQht57Trka+t6rQbs2vVVHIQ
2Xai/MQjWyMK7nnuiIvNcfMWXtyICilXc5lDpFw6/nR703/ECdiA7wWuuKQOF3A3PxjfJaTRCa2Z
1Yue+UnzD1QHwD5xyh0gBBzhgYGEqNk1wIYhDzcmrXs+rkjmtF3i4D8VSnJR5r3tTwstmaieKhbB
KTnwsh7EUowXAIA7C/iTW2S/SLGYF3txyZ/q+Q3lZzQws1oGuOxf5p8ZVIB8jBtmJwUfJ/gwOxdO
9+A2hST9VoH/WzleNcXX0yy2NpBqGocWtmNDEdxPsrEjjFVW5C7Hg8BiUgdoa9y21If2nnoHnEuL
jYPz/75UacCuWmUesWe+7IqDN3kvWwiFBtL6td1Gj/LWP4J8Ozmh+UQeHizSyC30evbwNIWihGmb
0qetlAFwmsZiJRyJ8pBkyQ1x+O7mGyQEujFEk0qRxetVQcajRqU36F4rl1UFMRI6hTrW5iVokenM
H+EYAEh5nq+lkwwlvNyopU5pB/sToQvFo0a1lpVuUgAu5K7cIoVkBdpqPrLHjTYJ4F+8s3KNADHD
fBSo5vd/X5G3GoRplYERbIYcjvzxOFSfVewzYN385H7aeKQeiCn9FzgJgVhhJJ3ymkOV0BGWJD3G
vzx42Y1buuLR1cby6a0VQtSMJGg4Qzi158fUdE3lAoF+ewwtH9+/2P1znxnhEG6VXxvzqz+UFivy
dZP1dP3fz9OMkBmpdr2geBtKkHgb4+QQp9ummIbzD97fZqyxP55WyiOC+qj2Mgs+X1A5SzOMB/Uu
jLsZnN2DDqYEapfeLR7u4UiygYf9zkyE1Lr1Gopl4FpIy0j2I3ikss3Ajk0RoGFaCH6P80zOZQkg
PF2kHmvcUuLpDfMSQ29uUzXd70oM2AFxgGhtvNbILwMZ2evHpc8r+trG+ikvRfcRv6mH5YAQiBIq
Yblc26Lh3xrRnfXfPdSLqtQVpl8PzWPociig8Ecf6Txm57YEisGCwCiqaH5Xe1P4P6xDr4Hktsh4
MKJrGvZVkISsUnNDotUHTs7Y92RebuGUm3ZkIkn2rQSqGc6YoyiZA0w8AFP6PBXPNPD3ldR8uhBI
86AHSG9VVTbKh1Rql5qjpWP2E6fh2UM5oQG7Gr4hJwrgpQ6TDz91Ld379IPdw4zlk2D+eyHnhtqM
K9zRWYQV3rMu5+NlvCkMR8KfpyYj9X0QY20/Lp6EGXap7NjlVg4dlQpR3GgDIy26Hd4awFr2Ps+j
9iVPQ9+7J/GNctxjoxUVjQ/Cj3HPgM5Jzn5gVUJkHHf3Ek7SY/dJUG7TkyBg2BcY8RRcZgr/d1V5
jTJmC6N0uyDaDofq+m5IZ0+r45ueSZY2OM6ViCkh7CdpDjnZfJ42nsh+mKV2MLVPbWPCt/BaNnFZ
ZwWSMy2qGq0qPcZDijmuSrCPviGxT7ppjBp6RQ3S/IM+el54f8ruPHHK1uUDWtwez7GRWTLkjyLl
1m7TscqyzgxIvN0P6h1Eq9E+pSZrK0FOQ7td/pQZF1763neD7mrU3BwH3ZMamzK3KvnBGU1K6Vjo
b/sKKy/yzxazfpafQ5S6TlFOxB9Fg0RI+9/qQVV9Y4QKGKNMZWOcum9CCnQ8iQsRBOZVZwTShJly
+D+W0AyQ2B+CKThkzbgLJwSFhmfdDf5WrU08wS5dc1S4fBQP/EYq0hoR6KgKjzwmXG2AJpo5x9n9
EGkbmP6OHZwVTAWfMNZROOD5yoFG2OsMWKHtS8j7UsoIeR3HE14YL/ldjZPlRmjx3DyyxiP3ZZ4g
gR3MQ2jLW85zmQD4I1s1GYWMEQlKlcr4Hw+R8JoPW0Mb/cxi9zHrImw+qKhcyVW3MbP1RnYVKqgW
wkt+v3Bcq4lAIU3otLaJd5MGi94L7rHVKuUOtOU8S7Bz7tq+S1TYTOhp7ygpplTiXqDi5ykOntMq
/c/nXo60PefX8/svYIwVP98MIm16AZXcnLBPI6DUodhBSQ8OjFCZ6tQkmxM5nrixYYBrxVho+0Rb
0n6egCOrxgozPZXahuxqp9WBig2tu8g2vluFVfApv1Gh0yR0bjhOXRk35kgOlMwP1cku1X5M5Gkd
g5yYKpuf2c+y2zlZFF3eBhy248ooyg3rWBA0lPIKphHU/+3albYfWqOtDcHwVtjqw5NATsLw6f0C
BgsN5IiACf9vvXm1KWoc+3tU6aLXf6+GzPG/iLmJAkZg/9ZSEIJpX+SAB7yByDrUg9fLIRV1n0NO
PR7zAOxwk3rrmgRhDDaDxr6U9f7Cte/j/0qBOoHNypjZPE5vKt4xBnQfBny2pRFIvkpgAiY/b25J
iU/5ijWZf70KsTCU9r3L6wQ43FCWATce6RXHKyXQQXz7uU81zJMT61Kz5P98/PZ0xLsI2EC5lB6J
vE1AxWV4BoLpi6jjWVFaa2YuJue9Tpqc3HluTsedE83cbAGLGniyuz5VTGOAToWJ1b95WJhTkL63
P5Ypo8ZvClhV8cvINTADJhGQixIr+Eo9UTsK6zrz2d8xnpO/QDQSzPhZWRr4ziRMNpTTs99vYI0Z
K3lUBHjPc+UrcIzUx/dhteeutzXCt31M0yjTVT6tsG8a4JwQbG7Zk5X7FIAUGpxQRl9UN5fiP87R
9feMqDda3/FI03M1LRS9Et6eMaQliA7norvCvmb0KuoICxM8Yc0FgQLf1YZhOrMrOPKmRFsXTD9z
AvL2PORwLCvHlmLRWrUNoEuOO8SlqoKFeC4mT2DgYDh1l4zMZnyPqdSyB0ZcyPIfgAPtAfKO0oGn
8QI+egz/ZU1g0mluJb8PbQIGn/MCgewoiCI8yIAfgd5MNLGwIaTVveF7dq7KpKnBSUczyT1xa6QJ
1xinKnOkeQIb4xQs2AqqdJIjxxxAbKG+CkZbB6iGqwG81W8z0otEhBNYL7eP6BR64cJ16e8E5KDZ
VJ+G0ebmbGziDX/eJpWtBg+uCnPV5sNSQK1NLRwYUZRK5aYRTEWpYcfbAh7wfAaD0cx5F34cyzEo
Lst2e+Jz5OrGQmTPG+Dav8dC3DiZn4culEHWs2G2Lj2WurVg8aE6D3TFK4HN7cK6nVLpNh4pilFZ
Ri9pSXGSDZiD29JuGhjJBhRO7+DIzqK7VEucEm/b9aQRycsdoOoLLN4dImbUL51wba2R8bvBt4dx
gMKWVu/PYRtauGWB21Zh23s7F9Nm4ArI2H/Mg3UZxMSQmHiFEx9PJObW61W8S52snlhJO3Aj43n7
YNiJL7lloL+5yq/1N32tf/TpzZRY459CZxS6ck5OjshgiBJCAZMgVrxBHqRDx/H+03sI9wm4o1QD
oP4BSzhd0mPuIV+jyN7XqdnBvhscNRt4cPVSpxMD5FjXxcXVk9gUdUMk9khC4SlFGvn4YJfqIfKb
6V0C3i1tlz+85AEqFOawKjlu167WTiTkVUkF9OpQWBAuKe+Cq3D13czD8Q8Wkd+R03ffZGixmFDB
nOzB+jVG/sgtN7xF92Ow9C3vwkeqF+3380DRqLSwDY6S+nHiNXnY+Wx7C/kS6TtYsz0G31ASVXvo
IyEKWgExtftP9qWPeJZgesGs4wLWoX8gGCNYKfeyifCXFxhs/hJl6Ct6OnV3GXbGDJTjh+8Y82DQ
iVp0X/a/M37ZnZsOQTxs1bQ3zRCAWBpo7e/qZnfAlSkFe1LuTQTTMf2k7/iwvFGm8GbZ6CNfFxcT
sKTOHh0dt8cdLAfEod9JCIbTdZmdyAbyh/b1b+WMIMJnbpljRAmTDDIVd3QPKBM+BR7RQwXRAR18
fak0mDYIspz2bXHpRf6umAAn2nWBC5Y7AmzFVTw2XB7NgzJOUGLncLxpqX4nnRInTU3YhUHd6qJS
7rxOttPyB6uESy5e3euW4TitFwLZXknlUQ4uAz2D748DLq/67n0dk6MuoxhVGbh3tE4ThL2riYud
OUjnazvv40BOrcUJIUvxkXWwValg5f+7yNKW4nADv1MsU8XkfMYLnKQDJ7Z2qjn8q/u/AmAQEmJL
5OhAeljPfqxRlp27bGhhLoz1X9cVFdOLoVlmemg8FDoJRXd7U3jFVjgWzIj3v+jIei+9ejCkaRNg
A/PQNkqZaQJ0+FrynbEWr8cs/GKQygSpvJ6OpRah3fStyfnJXVRI2g77WEd5z1C/k/uE82n1QBQc
IoU7R0CLu3pbEvw1s3nZMM7+rlc7lZKbaizu24rucIJtauTGwdW4oJrAWTPpFnxF0GGkD4dP/VF0
zxQNPv8VKCVy39Q/ZCwAdVKdifi4iOWczckP5gY+bJFG0BVjViZQyH/EFjUslTlSXTRq2R3jmPhQ
0w9d0BgtpkByMWSDwrCmL4UJ7WyN5wnOt+UUhGQ9EYNUW7qRgFRjbCP7BbUgPlLAxRylHXUc96AE
a91/r48z4mA+RpUREWqwvYRUDWWIIY2+txbdyCzQyriDaGpfkSug7vNGq4VcqFj18XbuSODF3e5p
o1Wq9aUqGEKw0AGGp08+S4kpSVon/Nwc5zgVnuU8yWRzumBsgWN14yR9oMjtem0KzVAn43jC3PQF
yFr1a4GzKwUdtOMtg2DExWyMHMC+GpbBdF0iOgMCrYmgexDt6UfB/0at4FwH9owIeG1pE2Zed/9a
KvpdjcZ8HfvqGJV5OxoPTSNSAu9o0KkdRM4Ne4ZLI7yjg3j2Mv+7Hz1QSEUVz0GjUd6OZYcMo6qM
3Ci8rY666GTjm1EwYDWvB1HmNiRlbWndr/381p5LT8xJy2gmrG+Yo44hYVyqVmR2SJcKWOH1xGd+
bsvE1Cqv+ffaEMrC/2qAvuHrQBOBg8/NuU3PlEsoZv5oWYBByAmP2oT7wJ3nQJ9rTPqrT9rcff94
lm/jtWxCO71X6AG7HlEJmAu+6gaKQKy1QRhxtLM/75Jto392B5sge0k9USMYzOg6vId/tLGCS606
iL9vwfjr6Iw8J3Y8xPNKkLAxbAbK67ojBgyI1ZRCTMJJzsxRE4IGXYRS/+iKXryhGV6VOFxfDPsL
HV8tCHvR0ubXH54ukT7dhNXQg7jr0DRwu+WWMVVnr0n29lmiDtRCY1V1BWNfTEOkhSxSDdrzQkfv
CBhOi8qeBXvKdA5hx5jWwIpMkuDnOmNQorZv0/JErEtW33whQurH3TU9RMcZoXhjrc40rqTlIy2H
2vbteCAFZXu64gGn5Yrlar8SMJ8W82JPbhdBv2qyLmh/F6I6blUxntFUEUNzAkbXZ29wSY4IqIXa
HM/8/JAWAs2PSlEB+QwRvsZbz0YurmAAsnB1RukfMSSx8Bgkg6a4/NeR69wYHJZXXqKITmUS1YQR
GSG3bejd2l9T+96Zo3H8g5NeUctPQtLZdVSSOfv5r5r3QB8K2f+K0qSR5xyELNwUraRXjjuhgefO
d8/iGLHcOlvlSC+mpluklP1fWd/HDIOQemIR4FQM+8A5AspAY2FL/yf5idhTVXzdlCnMZyN8/naV
Q/JouNxeJd9Y8OkNdlVd65azei0d+fjDOXOCJ6MrTTtEc/iBWvX8LC3BlmC8gsOXJrSBobid3cDX
j8P1zAKjkRuwumvYexuE/hVPMSOwXdf2SHrC4KhbhugGhzkZcqBPeYu415kThOy3fm2bbXPWXUlQ
W89M7DkkS4xOsmWIOWYcT34Cj/zYIaIDNjCwq2Z54/rbFx6Dk+1ddiG+pL+UDHbyEX1J9u4Gh5dp
6yyTt7kLfFzA+XlZRh+KbtJ256QdLipHw1LXoh3HYaAnUBow0hXvazR7da7WhDYA2WzhebqL7Clt
kXiO86OvsYEL35B+kvBmc+a/yfHhK98pLwB3dgH6T/bMj2E22Il7cTlckvPZAXx6VZkoRpk7c2fT
PIwBKo5eHVBASbUOAuR8bkFe/zmjDqNWJdBHOgfsnnNO1v1eqmc08HOFqzmvZJbg2VE34gCexglr
IpWxx4k7bn1bdQhnrgRFqfe+UdNtDEK6qEsKdnv1YVHWlXlA5w/cW4xcYGq30eMNW9yXSsMfamoc
RwYFqeQDRMwkshYa3ZuA5mOS9ujSVgDSqXrcmMzplEtbGvFFDoVHgrlNVSOmmjVDLwXMgPw8Seo4
CP3x3EnvwCGIR5aJp9sX91CtBZ0ToRP6EqE0+kDnHV4DXLc5yy/J5jozZQoL/dOJIe28a0SoezcV
7vx+p3leKuGWqPZMkZPb3rPKArMrw1F2PtDhSaI51OS/ZvSQEXLWoqlL5wbZnQO8j8GspVaQYzIC
v0Sx3oYk/qzYtHdwXSP9jRC+B169JelSZGvSd6IhU4GH1hFNaAzptgHc9fTbPiS03LeF/IPmlUAw
UwVbGTguptR2OjXb7QWh/pvNHhjjJTtgVWtDMwRZKJqDVyV7OjUgwzoXn8kXbR9S2CnpY/WLl3HS
zpjdDx9CyrHESlFVhLdChE6iPlY5/g74r3eYRjotlUuc5WYJWFhoOxE4XzqklbgWzXklJlEB+IgG
Sd7U2HCNFQuKbmrMBSLXGauchNP9s4AB/8gtcbghMsQIoVZ5VL0PgxJIADskRMd/6RdpVdy6y28g
vni2p+oFa8uE5jPBesYup5MhELfPNEIFiv5CyzzfQZ1cev8xbPj6ZKyEbkz/FPhCio6vC4i5Liut
n7iDWad2BsBzbE/bjufnxmDeRLqthj+wFRwDBEKI5gSUdDGPaV9P0LqVIABKVNJVM3kurPZ7no23
a7H7uWoy5FRcAQes75nGIoLV1fEvLEojiumJWkl6OM/sc5bbuzvwF8FOnfY998GSQhBV3oSDGH6A
GZxEQenny6zB6qGGeOSPv+VOFoUAD3jr1QK92pzi2MYCQwMWkq4ZhITXGnehT/k7cGJ8al2zx+vS
BusccTXu5hFhdKD7+mJbimR3RtUv/6OHrjUyYpyRpSGkFiSlKvYQ5QKfNdkIA2AEILY95ne7kRUX
/V3/jgZvIiJgL53SRBa7WRJKUtJEysP+XsumFjTbmDdrLQxGU0R4E7dD1eh90g9HLpClEVDGV+nd
LHqsIK9rd1rKmjCUWfje7xCwD05lPU8DtS1Gn+qWEDHqaW74krfunB59iAROkg+GvxRTqU3qaem8
VxQMroC4icgY1Q4BIFO+fOoexKbY+CVDJhvSX6CEw0b2dcxzsmPFM4edlSwm7goqwfviJbAeGkmU
aNe1LhFzllGkKHI2oa+6Fc1hkslwgQGB18PxWFW6W0Aau+tEBIZmCeCv6iG+Kby1exStt+bvBwMS
vCit5e6621dY79YMnj2Bwmqnx28b57brZ7HdXPuUOkbxOMD2SGreSi87Pgtc51/xjMLEGR/PUp4S
gcenM1RrRAtSpHGIKC7s8y95mKhRJ6Pes6M3GCxxCq2FMEfVSSByubHDd9xHptWLGMzvPSfru8ih
jMI1wN32Wvy+RlGzKpJ4Kpnav67pSU/wJVIsGt/buXA/DN4qkFgEtkkGEWFx1QsZG+gHliS0fqpv
63/xqZip9nXgL6rkhM55rylS77sKyZHGU6URtd2eHEpbWYYMJGUaMJtPcylddpQm8qXmMatUN9kK
4ZFAx3rIQXdT9TVJsRqnB0X0lohfXCjd/dMmjbSlIOTKcIiJIQRQfP9eZprbyZ9nqvwqOMlGEsHt
Ll1vLcvZc8dU46SqGb0Q2007F5JbQTp6ZDUlAWkfdBuWYzGWIObYZjR3lwNbWNb1OGwPew15WHeH
B+jhG2CK4wYKo8y2qKrMGX/AAJjRt1HtTTNhTySfyBK2aCe0jxOHWFhSITwTmE4aYL3hotpaprmX
qXX+sapJlueRdVb302TXWJVYOUQHms38K9HXfdr8B2goGPSpX3EM+eHGsypcQVFl+yBrsLg0CMTU
hYA9o9slWN44+7FWVPHE1RT0BaOYHmmaF767npzqsVInb/BgManbysoTA9HjwCudcGq8afAe3n18
yEDtU5nm2D6wYt6wVN7aaSNbohPXgkR4G+N6CICiczhSnHkpH5ZII55aGqamzLH/3NpwdZGkqsPL
7GQNuqIGZr/VoPVGiwKPZZI8IMQcsjUSIo622S0sKlq5LhiRbRK9NatwlIqxDKR/ZaL+JeWO4Yzo
HAeFNJE5iyIc3BOLL0TSO/YWqK3y3Yi5bCl5ijrrDp4Wd7VA4zhGR1JZHJGvpJ7AY3c5ooa6//3B
99YUFnyOHA+WQvciEX7Qj4P7GTGETC5F1YTBu4/QKdZf0LOEWPrETygmpCScbl82Lc2jbzcZEVsq
9L1mapUw9wimnv1pVsj2gwfou6wBFrt3kQ75pewcWuQzl5+ZxJ+BItIZx7jRlkzEGD2+T6ous/NF
1QCzfZ8vIkk1p6/LtvhgzfCLxXXwnBwjEUs7BUb1i4H6YCZz5EttB01ZWeuUYlHUJmmGsQyP9U5L
41SRSIaHJ4y40r8CSnD5yCvcB+6Xk8bXZ+HjEuWJpaYg8A2Z392sL1ZrvRGwtFKlf9wP1K3bpxNP
GTbqbsq1+oH9hSgqnc2xcmat1vyEDS+nk84C5mnJug8E+UvHFuFGOylZY7JJuIVGZ/EuGY0SSKiO
EH92seAvN/5WA5sxc79SF76Jk+oiYn76JOnh/hpTLI/neL1qKYKSSF6T6yDUENfSnKJTRD7js5iz
uB7i9IGfpzUzB1jwS6Z/4ELvd/dSC7IhdNMB5U8WXZd/+lgwiJpoTUhOJ0IgEqymIjcggNlZOKsQ
qlyUOvAk0Qd842Avkbf5lXDVMwE0C0s5XZOFwDgLPwXTsK4FQzOcR9I3VaLAuL4zPEgemMa42Odf
TbkukxFO8ST7RaIdMMsd1CTk6wwTNR015AISFN829z+vJVSR2eU4fRpk6sEohXOeMlkyJOtV3PD7
QCDyxo7Qr36zp/2RfvTx5lLU7dURiuIZKBK3Pw2vY5mMDYqFpUY+JCebXn6GNKTHUcmziCJboF9z
XGRhOsoY0noodGpQqxWsWUZfjXwbHzJM700BN4kmGc197OOJtWuG7Q1YE+n5gAdsiR6nF1UstICw
0HLw5imLcN9G6HC1xFtAX3GmHp1Zec0YhCeIO1jTfm3GG40xV80gZxYOjpwCRlxJbF/2Eg84K6jT
AKcFLrKKmUq06LdOUTVaXlh+lAFj0FckQU/2ZXOZNYf6uPfeRNjBiOcOwOuKtSYPj3ySiGpZgfAX
odsmnEXRlv2wwKR3uODrVzWRiQc0F5nr0GI24gb50BVXVxJgOfl575rE9l3kmFUJ/gtK6rYtlk9n
f32VvZkSqb6Hf20FUMSziO2dzSq6uAFBkGxqDrk0R8/CloJIelH8n1Yvyap8BOqN9fGnLvAZ3boa
IRc/AbO7eKC99fvrMM7mDtaIiF9HTR5gPWMUcaaMHba1P8jy9nFS3XmhhSvUVCauODzbDY8DlEdU
SZj9ZZiWt5ExbE/cTbPC/bxd97sqsOVM8/9b2Y3IJZgX+XCZ7a4r4HV2kvRg9zoAGRcLLs8jFVoh
l9nVr5W/Wafc2ku77vxCf/v0Lg2AKS10MliKDiwAzCBQoIq3kgOpotJuFGIrLlc2OOJRZ5S8+uo7
xaAsBLnZTwjIbqSILSKNLvYUxeEYhrbm9vyo4q5ZPq8w7hS9pkquqIYwwWjvEVMd4HS5EnvHQx/w
QK3FP1onuejH0GMZrp0ygoKTXrQNTNgaxuiXcjkS2i/o92JdgPGJcE3L/wHLjG0XzLqtK0bkaDwL
DRwR+GFjpbesTOHYLBUOQbFsALqqo0tc24d9OHk1isAfMxYHWvlZluNpMYfV5knWN+vXhoUURDtu
AWUK+wOW0Dl2IOkzZRB1kP0j1K29T0EjEQVghE6ag22ElTzl1ZVgNUh79kRrKCymNSEJjQvnTSdA
HPxrBIq4TDD1BVG+kjHPEOh+xweE7jvM+37FLG2a+Nep65S9ZU4nTYGwGzEN+aKQ4OJQOZXPcle5
Nr3P2lyT2sJ7S1LUlSunPEa0qyYNwRZlG7WI80rS91xiBZgsClEedK9jclPw7FrvdCv/LNBW+42j
1CPplrAmXXQOnCvUoJGWwhPiNeyrZGqht+kxLMKezdLZ8GAd736WLt/XtDjwIFXbhHvtBxGOEFrA
qr5ZWbfD2ewsDJ2TUTOm2PS1HW3ToaMZ5yk874YxvviJgFufrMr1y7zn2Q2jlbOtd9rgOFLdfYub
3sJV1uDxLHhGuc4frVKKFV2nC+ihTAb+6QN2DO7VDPXiqbcXTkXzOa5T77PvJd89rxKRO5kU0Y1P
9F6G/sEVO//fzxrhU4LnjLuL8HspxkxcAECTNYQ30iqF4HRIOD9W1nqh1u2Fg1yD1+4O8QoGCRrR
LZo4+pqJdzRLzs3MobdWJxtAkbLpWTFr3LrSMYLW7GATumLTKp2EqTtkGl7ukrvAA8VzQPd+m7Ga
Oq0zaOjCnlBovthY4CclMoiaU4YYHMje5266ZM7LPPQLeGamvW9OHn4amXHIpTe5vyZEjY+AD0xi
zmY1MOHK3HEsI1pT3P4xPtYvlCY3U2Ve/ZSNBszZNe8A9zQQ6hBhkpZBzW2eihCZmLSwMC1oQPX/
AFf0YfeUtENJTCTDOx5fCPxA5Kiqq5De4knr3qTto/fMrgWRTmfz+Qz3zQyTQqA1y4bnGy1rZAM1
30BO8/HwdssTRPjFXeOREym258dEZC+eXd7SfHmm5mxj08tBWX/ky20hIf2uj6QSeIevJZJ2xE9M
9xh+PPEH+sZIeBusmEiTeJjkVWpC9C8sDN0WlFqNWFHwwSNdAdbWPlb/PlzYnxg4Q0f4bJy5y0Hc
9Ir9wnjta4ASRKkO6H1WfqrqDB7YYj2e+rSKT4XU0V04rgtJzR1Zqm4tsi/9YN7xasSLOnjLqOEn
jtBXA5NdxcoQDfkSKIF7uFpkJ/M7tAc5oOI9anuRbj/MSsgdyW/WLuwTaPISzmQkE3Ms4WGs9h6e
IigpNVT7WQTb8LnL35nBLkoUYHDoGSNcT1yhDcO0tdFqalbLdhNo6VLIp/LyHtQ+xpiNhcrEvrRZ
hrkZGsY6FHtHuQnXJc/hVNqhc2bxwp1VwlMBFr/4y+XQ5YzTa+Nl5ObsuDiLezIMUlXabDmjPtnj
R4SwAT+62n/0jLAJJEFxARACxSB7C78/CebyASlUgk7EJUzj8VNVscbdhiPN7mueve89IQgGwqQ+
te4XU7Cx+EPX/023j8f/07wuFlnGMylegKbDhwHgC/kAvYWNasE2Yu2fFO8VU1dF7crqATrME7tg
HfaqO/V7JySHCL4I+fyRFqgJy+1PTD/ZyonM2RtbmfkA7dQIc01WAxaRKr1eOKJ2iXyOoa2yK1TP
PobEAS3TrZEwjcB14zN222fuV1j3qk7S5SeVNiSjKv37x55cw4BIFlkti7dAC+WWUsJTOcZ//vvL
QbHOTVXsZuo/55QHnOHEH141ja6LFykT/UZDjMR/ABsyFiO9HLuTt9pbDmGDCA7S8aGdUY6GwLts
UE05oED/7N/KG3nZvl2VD5IlQjhjQxsvPKQsyzNCnAmWlWLqb2ZQusNRDd6D8TMvjKcXQUx8ePri
GHEvcheLy3TA7UL1LaMKTh8i6r7hczr/R0ZwIfiBJvsWLCy76PBxNKN1sXTvsl5JZXVAg4XymjUf
IPaQDNphVXQMw6o3Paqqocy98nhprGK5qo3X36otHYVL3i19yTM3wm8ehw484xo3zDEWND237jla
aO5Wy/huKWPWy3x+JoLHFUQo4kd3TY+xOdqV151iCUrJADWRmEfGqReMB9YLLzO1xnEd4xI6e7YE
UFkhZ0LRFAsx1424R0vTyybfqhinEAtlLpRT1CPjZ2KPgnJtyex82JlynylqA+VrtOW8hOHKwfkH
14AmmHHMTh7n9pibmiPXI71Pw2Vll1XlTbYDu3czA2y9eQw2zFtNpfi6jErFzkJ6sYNIDenkxl6W
niyWOLL5N6TUu2/y86KWXasUnoy5zo4EZtHK6+D2dQBc0pREPFwOr2owyE3mNg7f/lFfvC8ertKk
h5yJiQmzXh5SWNbcR3wXOguTAm9lVxjZxBTQuicKSzzDJp2YReU74hqyLY19lr9vxR3GUe/hf4Pb
qN3atVFVH7aB/yIMqW+mr6Nl9MYqT2KGGbCxvouceH69nyvalPqwVDTYmQBCEF0ShEXmCbN/Wh5g
5ibEzjE7IXiD2yIqhDucYXrDXPCZf7v0Qb9jUDZLjMVeTOfFteolKDcuilTdIw/wVGYIs95whDOG
2oHX+Xspqu1yA/nhbBmE9Sg8y8avg+Ps1Pw8oMZukvSXTKsSG47srtrzx6tXmWJDY7O2VP3TNNvW
y2pzqx6vEfuFQKdnEj/1KW/e6QUcn8tVUSE24qyDuHqD7i1pqBT216inz9RWa9N+6JsuskHrOoFR
FfrXBFlbfG9tOTGimNNRHC910A5LCWsT1ijyFcrKfcw3i/N5m3rqBacI0DdG07QAOtlZGjdUr7KW
3pszJ+IUrVBBIzJ8MexXA1Kk/e1D/s4zaJ0Frv9sAhLB9pOCqcT7bpw5QlU7IiKX+h6zgk+rjwjI
NVRY40747Xo6pVNcdguM+Da+7D1oiaTrhIg9Dx5b6yv6lI5/bS+r+k6SuWBEF1WJSbfD1V9N5YGV
097P96dluiC0PbqDANHt8O3uzuuSYO78RciOvJPJqA6JMl73n2fz+GHKivL2aLPRsVUI/1HdK/du
imxiJOy8XSQMtk/MVL7ZyR3/nBDfAUrM+dTSHRE9hnMZjk8aKonFV6JMeQTKDCeDoCUYzW905gRH
jKS3B0qpgDS7pLH8bSXf9eRwhsllGSA9XoFB8Ul8tCio563E/qedfSJNF3cach6mWg4LCgVwLwuC
gR+I6vgiEKN3PZ/NdO1nHpqyMommti7fsNB7C7/f1q9MN406GKAgykiVOb99UhO6jlse0IryKyXK
O4wLANKfsJPE9H1kkPCAuz8dh3ECjX/TpvXuRJxxEX+gpgN6pD95fi+R1WYm//HrJG+5vysXly6b
hCXELicArgbX3rVfTIHUTwvUFCq36jVmrdyRZXN9ErtdNbxPqG+XCum4u6V+phvMnV03KFjoPFn0
LRLc5uD9ZtJnp6rFvej2LvQs4KRMzIJDKV+L7jDzTMxYRNceoKALoZk5JUFIyoe4MACanRci2nnh
LvhfXNpZPlhlWlhcsssqprVmgdMnXnh4dWgle9FTbCjl8lo5544kNzsQ/8aUuULRCkELExCldWhq
Ir34JJ2HDnrlsBn6uTMohU4Xu8Xzfb7OvCM28htB+2bq2E8pZTdhf+p3sXSdMMNH0TkA8Dohcf75
OHbFP8Jb2bv3VjOSYQDCjVvKt+1/xljAtrGy0TKDJBBdR4wg0j4WiuH9sUB+6fqJNanGTwoNzcla
Z8xtwwjcxsiJo43T6bRrNopwT8LZIr8K4Ti6cZatKOsi3HIZnuQ8OZT2PyN3poyjoeQdog+dE06s
ynwVro7Cff0aCqD8wNqIRRJ2kFcdgkQLvoMchAr+CqQX0D69ZE38zU/4m5zQAPH7M7K7FfijaMQS
4nVtvBHwd5EI2m3HirpbOOyd7tFnwihSfDjOaf7/R6M0K/bXIFyjqaWBm8VeQBdAUy1JM4pgzjkJ
oTzv1coc1ky8r8MCv+iQ13qnzvlFWhImyXjpaIUEcCWjRmyDUcgnkg3CyLtS2afPE5VqA4JQbJhz
uP3cIlD646/aWA5fWHr20r7XIO/G+67IIkxBHzzqZA8GkVVd9417g0GqdIoBBzrzQZN5a/WPoDlH
KYc0IGtO0g0tQRe3Wt+PvRgqvp0vhtUenRiGZtKs7AWWzOIRuMgfxWpsP8yr/pB1dzN9nLFILW1r
u7bWINf98eQ2u23x/IXkjUb/5mFKJsyudrvI4DjnIL+YLkKIzPLxjPmbOnWwhED1J/B66LrNtFxs
TW/6zJwJGra+OpZ736nn5i5fw4sQy+KV/CXP9nL75CEc/JbZvGkPlV65nkVvPzxQlskNc3keDZ+p
WjL56a173GoMyTs8izqi3vDZzMuR97bVQ6D+ChbnomKc7bYP3IfTbExRpFhYGLAClHYfSEA3lK8T
tIS7WNXM5gBXvPJSeDcGwgSe2UZ+s26bj4l5Jjd/9Kw5rbvKqGEuOoJyDqOHS3YlQ65tzXh5ewqD
xzdqHdAu9HnA53gJICO203Tnom1irPXkAec/esafQBvde2nnWyQGoawym6WzphPG5lNfhaHhr23T
CK71Gu3EaMg1TRSVPTNv8Dj/02jOMfqO129HhCjWvPk1CXayFnEPFxcHaCD6AnVdcDKkdY3lrWxT
ux6k3Lpl7QQ/qiB8aIkSG0a+3NtFc/O0grJQIz7zIK7AEeACXZJASNp34wvGMhS7dM9lVIL8aGAa
ioHdAsU8nMreGsYOHvOPAP153QV4Rsd66mdzuuqu27TvugGe56rwQF5niFakz9wm0jTy4YzVYZ87
PSthzGX/y0fDBTBEuNe5Yro22YdtXg38lMCrq9qKetKykhrBRVVxxfU7pqT5rfTDWjnzVA/l2+vI
PocGZGddMRrXsaqJEpCFUQ7I3UHRVkHdT2nVB5oxu0tNHfLt9fydWPk8QRDhr1JbFOz9UUbZY4/H
+61snOaxLjndDiAkFlP+WRqBzKD1EqlqYPexIGHX8rmNFdfrlEqByvqFsSaUWwNeQy/o1ruG6ndS
4NoBFepvllu2NrOcOLmevbH4XMbRvAcPZ2CAZVHyBH1pnY2wpNZykSXUPwPrdoC2Yw7X59xRyNtV
Z1LTum69/CSOnoOZ1BSt31yLfhSIBDFYmOMHZLtanq92QTY3+Z/YfciE0kcvgzkcJ18IHx+whHOV
Q0S//XCLtkR2RXXKzifhftqmlBCAVqvLCA5il5BdM+kKnbFbpwX3R5FR0D0Iz70nrGF/BkA3N7WZ
xKztwblRrRcwgGiNXTpystGeRb46LD5Et62bIVUsuTGcEhC/Cs2bikQzDq6hyqYnjeNsvVTxglWF
BkCvz37IPYUONn/SxZ2ZS08r7hQZtjtVluKQ/rs/ff6Ycgc0luT1yHHqSThFXGZP/ge+o47LAudd
sORfxIpdZVwvDyGOW/ezhC0kcaQ7ccHXPLz7lR2hYyD/xfJaWbP5nzDn2jTO7GSvFQ0G9LMH65or
27VgJi7uTTZTvhQN1CopiocYQlMzrn7/7SbjtzFIROUoPh2Y8HTGAuLQhzQH090OTWfrjP/GccQg
zKy43UUbwqoEJ53dz7FMlW4ZHsNgO3KIuLs9b4Gk/Mbsbrczb+0+APbsBvVg8FBQNPcNiwE9ftSy
gMY93/RDw1mJXdJa9OrZZFltiH/r8Bd3gLeDXV5LgAGO93ZiNSXRVpjFaF+vA3dni0Lwn2Xl0svu
uVJ6NCB2i4Nij0D4/MkNupH8W+FDcinANyJHxlFIqJq9atsKTIul9r3CCFjJaQfIqe4qXkBLWduW
ymzEhhol9IeM9bi60U8UKTH4wFWwHdfrKtfaLmAkjfnC7IUxWtLAxQKUWHeqAab7Ti9eTWPv0PCz
nb+S9xSeg5mugEehbgSRzEO8LJvD0FNcstVuAMSoIj1zeD+yXuADQL5EF+DMbfKKubG095ngEqyh
z99xRXn8BwmKC9Ek50Hzb5pMi7It9RRRdxTlcchStBLRPEcj2p+LaN7R8x7etZ0bPhCx61mfA09B
E9JYwF06+KnRAACh/cVPl3vr2PN1WeHfNe+uwjBkyAFKskQ6NJFCh5n/tXfTMlq/OtXf7usCME24
jWd9tTfUgnJfIgzUpJU21jl8Hr+zLUB7qVQwVYoDh/iNDse6Xnx2yw8iBryhJwBrzQrWrZ/y5b9A
bgakTzfdUdSMrH62VzVJPQOl0E4zN1w8pqBu2ayCOOKvV/wmrp4SXt4zxK66RA6N/FXnzuUteUFU
pIITjs4THOmh89fUlKeqC63iHUmVSwTgGM1twNncxHuQszi/RccaqZFXHIG+Nds6xH+CfFMFSYXA
apHJvcw3uO9pn54q5aN4I0MQRq93iVStki6cGEDDGdAG4cBP3DP+ZQzsspDlyPWFF1ug/yONnBa6
avZVDv5P4uLA4U1f2Iytly79R63gADUV3iDD15tkgcMSzVw3aqurSNr5p/YnOQWnFhEfef66+dKI
2gEGFYypiZuPDQvH1DzH6snp/yNzV+wk73CmP//2PKwBjEASKA+TjwyFBI7mOR1djK3gh7/BjN0J
KCOXRWcWEQ1P62PFiNw/7jvYDcq5hE/Ki40PJL/C88oXks6H2KpcSWdL9maZnmo/r16EM4PRRw58
bB4HeBsKGjWVou8UyFgQwc+Wb5sLyHtP0FnJn2nM+t/+bslevG1Mio8WwOJisadkQ2AdJTqos4Ph
58PQ/B6kS+jGAf9LLqz8HRRDsSB+jP08V+jQJMszRcuJ9mP0U4QL7KVQIwqXph0NcDJBrli+Yq/F
vGhyO4avQhtpQSa5gFRQ/LC1phX4KrY0itmiP8LTCfwntH3F/W7GRLkvZxVDqrTOb/VJJBn2llEM
oJHSZkwcRLm6VVKP5+CvmZeNTB36v8q53FvioYRPbMEeHiKZNK8cdyu2uCMnxK/Uq3i2Zq2KJraC
OEDVwU03r+ibmC3yqvvfljqzBbVuKzc8I4XXJqVjdlmw6v/lcLScq7I3Sjb/zbyd8yixSFL6bivq
zq0QksJnDn3OMkNW7Rf7Uvd5Y22av4uJBw8JLTOgW9Z90zUfTP9Mi8Wy+mqGbOEUUuHUdkFclTQa
yWqs6EEXmQMVRomnKp34HgLv883avTqbr7WGyG9GXQlwc9R0e0+cB6EDB1XZR3UEYFwzTKTvMURx
Nat1MZnRldpDLsjF7gr/vl6UDoeF9671OSyrBnljqzwMZZkzmrM1g1zgliQ9UZNPZWqIoR6HUdT+
MQkxItLcjeP7G6BebHqq4IRS6oRXh/NZ87pu7YkvxlktQp1T+xRLuy4ND6VP3fP4V69SWNCMAXHR
wOEYtcvE6QuDe+339gEWrPih72Vw0hMCBZDk0rYrQRwy0jIAogaZhoPAtIQp23LAyEWeihcB528a
iCpxj/hMpdi/Qkc3QO18Ow3wvIUijniYt2WOB6y54hXuAj8sT3kL8NPS7AeVxPLIVW+PHmADZrZH
BU6z2Rm3awTR5HVF/DY9/yBYWe/OZppWqkTL6AuOb0Z243qlrwF8XYpfKtZMDj7IqAR7X39IwVHC
JXk6LVuKtWDLZzTwy36bp68udScifuuOutlxjXS+2WVY3mux3qcWQpTkywmucC3CVewMLWgWoNUA
/SksIrNH3H5jHvc40Ol/59/NoCQcLY8yazn7q5lq3yF2/JZLAZKcAJdk4LlMcPGpH4Zo/8GbzjHP
6MA1KjJ5UNkMrDwTeA2R+IKHMneinl3YrS9msQgDejZ45bwWe9diW7t3Yex/WYzv49AveRXBLNua
hAEGA825KPJPoGUlnycT7Z7wbWF+moGxZLBkSliuQ4ybAlW4uvrOvdm21yIkBBL0gh8ortw08q3/
DI1vFoq/oxrEUXFXwStZMdg26TQKwPaXb1KNlLxNb/EzmcSJFx5ReW18z+lgMiu1+VFK9tiLnACy
C/nRoRi9DNZJ9uVbT9CJKPGt0wdFCWadFPpAKQXr5Rs6j7SF5wIGBc/+aTsmrrXFCcrrl4PYv4oy
gNDsH5HFu8q97HSqe1lk9ZBeTlJbv1dW19mji7f0m0uonLnV/+/drlNUA/0sVwOVehZ9ZHKqPg2D
/c2Qr1aTKSOVDH482VhgP68ntimZxNpyaOuK3sZrKG6g1ARJFJ+mWA6/XP1WXcJEug4sGKPd+a4q
qZlhBlEmISIzd6rFk3Po7be95ZbWhMIkRKuNE9Rx0PW6fpzbnsKM62YlOZYORBSNWCoX2HxnY8Ow
CspBzfq867k3sjlA2qbKwrghTe4PHgwk4dMxgWchGmZxuLxLBTdXjt9CqzikdLnVovOuxv7yxf/j
zH1XauFRBrq/8W3pMegK7FCpYqZDZtGEeNn6p4ScwopwP71i5+v1N1IU8KCtidEgb45t5G40VyPs
7ORpLfizEFkOSqtEIJYWdsIpxRbg++sNmUKY5LxQnE5BgAw+MOmXluX12+hDjfZXlrTticCasIeW
25ikptZaIKOCW3JMSeiEucmLXIhVoN6tIfflz/KRrd2bqLMLrsRHSCs2HEASF2ELTQj9jQzroQxM
rJf8U77FNnQF4zShPke39PsoTPuaxzGE3iyAtEPmRtE5eOvx0madMlPNhjcFuoLdiPZNjPpUeeyn
Ri6YnZDcD9BRUDM3RDXiwoyarLbwU3iwkW/zkgKedW70XquGJyot+W/SnTIi21SNt+VYyd1u4gni
Yrw8CJQGG+GQZiJBH1dt/ycUJkdWcB7fLBS6UJsXKMDUiXBNgyc+kxTnsAVAA4GmwHHMFBWtATh1
Cv9aVJwgXd2f7DGFwEaDLUmFIgx6O8kBMoGDNaSZkA0/KZ+GIp4FQSxXGpvM2tVep/TnE4lT4pWR
XV2sOAWykUzoKrVHVKOlGiZyJpn8oQEBW1G2W1fPLP53817tz+nUZs6Jl/wRFO6M9YvlAHD8nnPb
eV9k1ViUZ/vWpCUf+XHijtbD7X/wkRZaOww5PWUUneHuhzx/kIRj16hnB/aBFi6y/yNqgQzhFqDF
QRI7UwOmiG16O2PvmrduQhKxY056lLakCeGxT20sfU748RdrkaLU3DSoAvKgY1IXxjaMM6YWz4PK
yA8Ms/9WfQ/Q6WGDZaHMyv/vMZM1HkDEMEpw6mQA49WOfPw4R01AUdhOET/CmuhcAoDP1Ve3JIT0
Y76Lr51M1Tic3bN4VOcNrHfpQi4kl4BqRz2rP0EOX+lqbjaMedv3oTUN3hUyrNXtG+JMeeM4qlcO
+Bb8rLs6NyzXQhjTs8qvaQC+OSDDqKm5YLAIxS37nRWWTSyhYiW6AzlUgLIhVJp7Jcn1oiqBPTH1
FQgk0IX/NZ9pzYO6e/dLN6KKeAfXhhRjRLAx1/h7/yqeEIPsQ2im04Y1+qa4Ig10mP7nLhkOWiLp
gnJv/CAW587MDe7sy7i8sxBWZM9IEYUCYo0r5NdAzJcAfAmvoANypq0AWhTcARAY30zohv+/sVIF
4jsZsxVrbWJ1uPm8DK68vpa9nqI5z7104j0c8Adtk6nRGlIV+is898MW2leBPbmvk9EdvTd9K3ho
RGc65LGH8DBevC+sHyn2+nUca5NMZPOil0VENmOirjCQdcpXDF0wKAypyeGJeIYwfC/vBQncp4cf
soo4gHneQKIV9iJdabALMsEEZeODxspaBjY86bQ4qhIprgp50oVBYhBWElRqozDC1hCv4lGV1F6T
O7J/aUklymxyRPVHVK00WizYMmnMxSz+xkYx8PwftI23ckflzPleQ6rk8bqx4uf0+3cW2pEkg4ZB
8vmxJZrA2U8Oumy0XAENzWzdPIOlCsIpF39kuS7GTyXg7litbtMGSUoJFeIrRkJk+H4qHksEba8P
yFCvbElGf4GD2NSN0MnbZuKYdMR/ubwYkwSmmkEj3pRuQrz5wrSo/t7DJO3NG4hoRhKXQdH7kZFD
T7LM3syEks0GclLySc0eO3+h6aWGwW+m++vU6C8FB4cwmX6osSOnKUY9OudCyo4wnfP6ZsSQEWuW
j1GjLwK9juQlUStQI1Yi/bif9PFpWfDxdhcfoqTxF580pV43Z3SKuYqoSmSjEnnXf5DYdMZT8eO6
2t+Cu5RsDyUVHoNwJtYSnyNVePKXjFHVj3fp+82kkeVhfoaBeslg1gQJOGIrgV/aMjUqGmEu1VCj
iDVTA+5RRF1dLjYAUAIkrVajuQ+qgE88ev/IXoHVaRbrBNYR8ESLWEXnhJ09/lYQfwjfo0g1EdCG
5+FvQrzzZSb39hM0t3tN6z+7QTn1SF/2fp7b6IZAR+kufob7Y45fC1qUZ+H87BcfClrtgcp2U23T
cuASjHJ/ft0ch5jCd2yxdrWV1JyLWMQ4ETOx+vuyeMV+FinpL1BdO7r6VNfzMPHfN3TA4uInG7AM
nYePNrxmW9VXF7KMr5RPPSkIAuEnFZFfqMOdmT0CkpM31upV3rOiphqMgHxfRY9RldDqdZLZUYUw
Muj5Xulq2OsVUrnhTpMhOUr6n8AC1/+ifi914TSc5/oyc2BpNe4GA4auiiHo8MhL2ztT2Qng9MHL
ug2Qvf8zvIVi8o/EsZvBk7DVYp8nab9y0j9oawVemv8L3NiNuHTL7RjYHonnqzSgJfu3MaNklmFU
bOseJ4gySs+RB2qJiieKCLQkKYE1Q1I8RUCQmALRFRA6GkkdBthQSs5Oest0j6mlJulpOurbtvit
tDv0H+bqYXSFFFxm9fBVOB4o4biciE2q7HUkUiUXW5/qsG6AqooTeujurOXUBMWQuXmI6Nna6vs7
4ECgHRMOB5z8EFa9q3ANQelovbAmWkEQzjSRAV3ksSotgdsFriTWq+792IxdbRXGPMa48i7cQjM6
dQ2eunL3mdASLmBhYFoTmaT9KKpAr/WT6A8d8YDkkGhmf8ZitjjDzuA1mj8t+ejexPXNY1wXVJWA
mxod+8zM3LZ4UWVjqrg4wmkBxt645xMHPn/H5aTVoDvcGlJMmKCqe5O4fofCLOIIogPIvI/bF5ul
P8twH7re+u0Y8haJl0kNaRAkJTn5VyatLOb1c6Q2DmGB+pz8N4grKBwPWgSul5VfmwuuhGXjDAhY
ekCd6cHwqlOcknnGR9WgflsjFRpm12XNvRt+Xs+inVIzLSSlB9uwRrAVoKvxL5w14rUGFjh4TRVU
pNASROQ4DKiL4HK11Q6+NDD45Ynw+duyHB/5T6LCD8D7uadIxqUnYexjV/qKCe5xtKxe8rDberxz
t5F5oAG48UQppMIZFEh5EY2TlfwZDW2NAYAyT44/+112yoXc/ZOQfNpqdyeTAy30riWwSxsVNAFv
eE3iuptbEw+wOM0KhB+s97F9pOr1SE45tzd0sYTuNy+Z8o3STY9LWx5jZUMDFoYO78Xv6CuiC2pg
OTJqlZxg5w0kPPqHGlb8A3ImSHtFUtV5DpZFxjuNQ81ghWJSO8zW0znV8VU6myxk7aTW2QR5qJCA
LSS/Vm7BVCTHMszKA/Cx3Ukn2kxvR8rhEYGwCh0lFF6IQyPTT3E52k9LkBE1xsDhU1kP0saAskOX
/bJi/Xr5rVs1C/S8PLNMktEXA2pHNFKNaaM9T1KeWJmAgD3y5wsP5W/BlAr0lwo3dCOCwll55JoU
yyYfzFuDvWRNKvtZxdXNTkIpK4glIAydASobc4bhmZhskF6U76iei7jB3zpFZvWSTrsd755dj9x1
lid93XuNkglyKhTwbr5ahZv2/U8eD+TUiQ+5fi3uolS5ZcvMvEmwMh1ofKPJgiVJbWCw4591F23m
KEe6qgc5Sv6UZSIwE+Z7Z3O20iQqgggyHDedXzOH/iUFFO/hJMcZrb5yhkfqgQIB7SOsxiWK1dc/
wSJZkffk64Zrh1ha0NojZNNJV5XSgaeKEV+WRehWQNfe4ZOvvdlyl1Mqy0drvg5ieIdTEtpgrEZ9
zN0vVEZjD6ntbCtiJXk4aHr7MJMK5pOi+Y3osnTvbW7eo6U8vclAr3Iy2AFZy5dqmLo/V/QU/mpC
SP0H822co/ly4Hxruc+DewD3GikDNlsazwFwk1TyV0dnrl39mPdt1WAFOgaebxUoiV7SIgVFnK0A
d6AEiMntoLqHV1yT36kGZtOrKSDwv31OylPldBE4BybCqzRwmj9Na6mE08gGQxOiKWRiLHB3xEFY
cI3S94c1md+wkwlrFi7nxJCiN7aRTIrl2LLR+FXosy0niQPZRrvnnxxi0dJa2FwpLa5LHhj3ODwv
Z0x4Mnx7w1jxVKi1rimj9HuAlH8F255hGlDrvejAyFFCV+1WUSdaWvqwxdhQfbHd2b4rETFQlKn8
KW9m0vHr2hcWIkS7O1Cq/0y1XyrjeAc7tc8FEdivfYYFgQORIziC+DfGsd0PLH4FcFk/4qsz++65
vGPqZ8yxFlhZJYZJm5dbPGlvg3iEz+QZosG1qM576C1MUbnrHq1UX5HF6l5nQg30NQ5xib0FUV8w
A9gaw30LEEAKgO3Vz5mPaBJPNWgVq4gBAsnYJYFnBuxW8bqHvRVn/j6OYM1/dOE2AoI+jKqoiggA
d+WN2W6YAFOFE9iyOA49wybt8XbhrimFFYxzhDNcklIPHLqGdY7LdzWKBz6+fq09btX9eQH+BLuF
4zots9INdiF3CNMdWV92eyhP2YAAsSFqDpmCZW23tOOqKWM+GgdzWv3wSeKzecHAcXozKEUZHStj
5Gqhn6xgXWMFJ/DbXse89gmMfwchFCyQYe/yXfRS37y9CxoQ9Oq+NN83FFw8244JkrroFECZk1TS
DmKD6cMkfsuLUC9Yxc1w+Tj2WKlyx/xu+SuSZnzkCj7+fq+5+DkumXdop/1/pJmdhd4dK3TKE7bg
tSY62ZFhsbyTYD170ICpnyb+HeTswmQCgOzZsrh5FY1inhkMn4Vhky822bb8X4hALYxEfzcEQhIF
2fxXqk+HEQ3a4VHRzK0OP4uJ6eiYTPzkX/ZTC+jdVlCZIxAHuT2AXbkQgAG5N3lsLi0el4JnrpX6
ouFfadDqf2XWVNfIIl5I1alI2CqJcwcihRh8anFgEBcqpz+0BiPzOP9LVyB7cM28ihXqNUb75svO
lKwANZH5xloCWeBKSecEzialRlf2Is0FwwNbzc05Uxfv2Uf+Rx9pdiSbfWgnRf7cWHlxzb6Mzx50
6FAu6Xp7hqqbaGJSJ1kf/gzu83felzwpSFhQAIHCkTs8DbThrmlavhrZGOcVWCKYykX6fbhGdIU+
9r2AeAcjjd0AaAgNO80VP6GGaEYX8bYXbR3wZbnG+b+5/UiSPQ0wnQHKbeIfAeD1+kaDLCsuNx8O
mMWrU/Vb9EENXtZ620gABKEmgl5LFDTEgk6J1ZVFVmwyAxzXu5P+xx9+EAjVSoL6rjLa+3M5Pv3d
NdB6xdtZUvSED59zLG+XBx6qfvcU0uADRBFSM6YA5a0E92iWqNtnmF7PsRH52q27ld+JGQV3YE+L
U7cpbPjsbokRnaXgJyTaLtmZr3OqXI6i9kbhAxXd6dauvmIjHLpF8TTRXCWTlUufvYnSdtzp3dT+
x3bjwYnYV0/FKbi/UdmSJ2T50Yeu7NlPDPU/34ozZQUEDNwCsab31lky+8ujw6m7mea59gYnnZZZ
o/XQfhRzR9GE5zr0H66Kldm8Yc3/0Cou5x11HMHAzH6LRsHwCwW0AyGgdd7yc/0neNlLdmSoLvAt
N7YY0l9N+omOPNHukimqrQm6w1wdmdxSpUnEHp5cb5fiKuwyEjPnDJzmyOgk+NRJKit2Rjai8/73
u/9KWh/8dfeNt8OwxvzYRHHbBWooTogg+UjzMZWLEBXhunNncSih5urZ71clz4XO8zMz7SXqvnja
eDFqetvsH129ZA/UYUMWUdJ9i9VQjVFk+7AwvF2AJus+tzf3MhzDGZb25WCm2i7jI9MwpevvTIoK
vqbXvokLR+HTDIdwkwPlN5uM/JYh20lV0xNrptDAaYgHeCUlOj4daGsvBalZGiTaDzFoSdzKPlsF
zd3mWNJemQdKEV741PMgWvh1BoMSH4cobCv2KEy8jOK6FgbDkJoxOYPjFUQO3b+EnAxp8bZGTAdo
jwS/v0OBhMYTocSXB7XUqKlAWf+jIaQAyYAvMz8ktoAqTYzY67Wh3a8dksvXPvI4wbgQsDdnHKzL
n0NllC9NkHNPDYql3eCOEr8gztoy+OzV5RZj7vA7UnP3+teXU2r5pYr+PMTub1tyutETQTDJEK8J
SYZ9KRts34My2WtPEcmNmcS/SJuxgyD1i1HuqXeOodxyoCiUFESXJpuJgy6+yDoo5/k8Qxz08af0
Utejscugh0JOiFLLsU1RR/P4jaEd0gjlcfPS6+ONGzF+cF+QC3g0mVI3gcNWNtU2lFzB5qV66iks
QCHSm7BNsiMzktJ+VqJpghK3xPnTSJjuILCf0dScmAu5rFHu8LiP3w+Zg981W6+zVpgNvnq4TnAx
NTiRwjU0D2lEvYEYkq14uCi0XS2D47vnu1ZAQswxGoaGo0ng8KPUubgP3l2fsXrsy0xTvC+3hwN6
6QAqmp8xv+NoJy6aFeNL3Q/ZpHglR31hB8vrYClf67mZwvBbPVaqps3wtfS+tZI1jogjYGly30Hk
Rmna4ts+u1djqbyWwNeuhZiS937+PdzkDmU/kH3fFq/HzOayw9xoINSmBWHK0ZA0ULqevzHY8xeI
Bbxngn5U/K0J4G43RKLkoWpxJ8j4inMHlRPK4H5cV8Vf0aH0XPz96/j4h5w7j54TcFsW8TtBX4Ky
Z89atdz8mF6fMhY4O3D5knqbwx3k7XX3dByU3+SURMRVeA7Jo8xeEwSvNX2H+uExlEXu/ctXNbZV
kANqZID2CvKXCeLPcq9z/YagZ3UUPIHTtfNn61glSzyHKQ63y8GfXYMuQpG+RW3Hc563RiCb5XA7
VeiB3wlDCeyxog1KMo90bKDCbdqdjF00fU+VAk7qvHzZYHdTUnQSkA6pgJ1hMUS+xDJsbVE7oNH7
2Y3CKjmXTo18YPuLboAuTDu5gXqrJKQVmOz+hdMDBc8AcCPyhsKLnC4+IWkHZ14FYCWFLNVgigJ1
TPpxFSTB3uEL//Y3ClztrcRTUM88HuRD3Ej24MB6lJ3EuUYWnxFMfFyxLPFR15N8Pl/SILQwke8K
iPIJK8vbLoPGGLrvpEEWwZsLrGQrWizpKU2g8mnGCF7kcyhxCbV2QZW3gN626mpBXMLunUsDKX3U
wQHi5Krnp4hOIQ8zC13a2F9OQiXhMVAe/qm/w5Mk1VDMuYbKGjyycJgbPu4y17IIhALjz75qIRfB
YYM2VBHdJTm96e6FlCneqWBvS8Z3fVSjfVtelg7xuArK0ajCyNhtFE/74ydJrqUO1FpNAU08kuph
ASaGqonVDofrCwc9LIi1PSjfJLfwr5ofJSZw6dlaLo6Brx662lpmwuoCD7Ye0nWYvvlzax6zUn6u
V87iqcqT7pAPDqaRa9uBQufRzlaA4wlQEQ6gVvE0VRElV6+TkimPEqVsWyropNskd3oEQRzhwLtY
KTK3XRMfhgktx/9yQRohj3WkBJ/QuVcr6z2FWwmCBkIzfcJiGhiyD6SmZsp+d235vOZk4U6zckw7
ADFNLHaPVnHQ5hPmVbHUfz0Gg/U4e0mSMftSdzisroN94y+vGsH/zg8Y40DYXabSdixNH3PGca20
I5VT2PCUERU8I/EiBtaWwPJYONUUULB53vcTIkj+fhRdmCS8CJzqC1HkttRkvJueA4XY6/CuXpgt
+b1wZLzecv39AIr6IwdARMoh2HZ/uzha1GciUJefMyhwmsrLybv31UPWWue8uAFWvzch6em4X438
BdPVWaIW+3JHiz37L3ACF9qowePSGRkzzt3q0XCiElc67N20hWjgPHjQuY5NqnGMPLOM0aZv+LqC
6Yx8rX5Xn2b5h500u4NKnUnCoIDbXUU1UO+rETiEjBCH+sg1P3TEhppL9kuyOff4AY1O/yBF70Jp
n5X9T4gEl0T5DxQOPdK4MReV7wf7j2OGG9GO/3Ed1O4nsRns8nkCIndbTj6qhLsdldcZNwcoVo2y
Y8bL0r/D0aLTaoke135QnA/GTJQXVIznympj3ZJpNqQpo5ibFNl8U6B4LSDGBP0w7HjgcnzLSLQq
WT0S7Wk2bn7FVIetd2lV3RZxPAnbeFS+imuSR3Raer4QY1J4rqWXcScI/FgoAgjsvCg2Dgr6/AQJ
7rCPNHbJEIWeMZCl8Lrv54TREiJl99h4tLPSRr/hgZcl/J68yizvi+s7X3Cx1YYv+pB7k5g83uBr
vDRywl7P0/DhZgw81ySEFT1bQ2Aufj8tPjYzSjm7LWhiX5An5U+iz/cWNQfowwssW21RB6EVSFl1
/lLOXnk/PLIM1p2xttZXDUZ+ONvJt6LAmvIsKVG/TTRpMFR0whFJYHIkvmDXYrdd/E1Qp4FdTnix
0V6WHq9sy7O47oXxhjrc4T3fPVbiqAu/MXlPpeJvIJE06ztLPwDT/WYYs7ANvGhuixNSJAqaRKXl
L8LgdFHGLmbOUP0l9Pl95hIOQETESqyPtbNHmyjJ2GEEAdYlmEiSC7Oql6pekieuV/c7XlV8WfFI
CBOLA1jCqFSmpxOxLHWkyHxDsrGBd4ZLzAA+GJbWpizJE0H9ccpcs4m9NEK+NNNlIplT/QdT8n07
ZE/tvVRtNyDY5bjEHWAPAeHpWTUHp3joQGgZfdkXvvd2QoInGUxbQT5KyWiegQqOQ0W3+PoIf48F
7VStsKYgk/B/Z6WJSjkczLDPRh5/EitWOTB6kQ30oSQVU0viZOHnnlO62hcZYvhDqbq/C8o3Y5hP
M4HeHjb0N/3Ahzq00giA68GCq0Z1jH6B9bOlYutFPLgiTy+RkSfN3wOAJgfo0d+X2hGon/nXL7em
/r6LjNaRvLIlXgMJ9BNyuKey6lQBIELZ0budJk1YtPEaEOudMltspudHKwuT8Oos3vfuyzBvH2FI
wWI6grSjow5ZGBNlEMxTCgofGMnvGij7IOw47LoZzf1zwd/hLeyN8jhC8xcinrFkeI3U+t/6iBdS
RbxvGzvJMe31dcEhyOvY5LKGXmQbjsEnD3KmRRzr9w5HuwrGhVW5qxgqo7z7JKCQUB57xRvakuW/
M5NLOvPrvfkWcdKD6Jfv/702qD37RnI6lUqRmqATkz52ipAZBNTqWRnmH8cjLcw5sI8DtRFvFKkN
bRQ8EUFG5eqIGZm/lbtsKNcgCD1lLeFMV9P5x6y0U20kdG/YkjfOrjWey4qT8/3z3fuSgd/QYC4h
Eg6nHHCOet3UzNuPWgzmQYP0k3cKEAYxsWgDrfXUB5rgY75ipNxeTIN+z3fdf2KgnDNiNgBz5Jht
LURGQ2riFc3mRPRsSbmKBABwtHevF+W5nkedr525MeH9SpQnNNPw/+8wf2skUOiO5QHT1eQamEGm
kyX4ktUzCsUFgGtFLGpVDladQetxXpJH/C4uWayjslaMZSJRLU6PG9gXTU3lNNYBWXd28HUNU5qJ
yfZzTas91rQAe7/AmzyZRglzGciHoCudwq8LuG70bTE7wnCgsSlCqOOzxEyjn/fNVvB6RDMl13JV
XBd+60f0JKtJjDrcld858wutcMl2NCYrB03sPxt7SCIsEFXSDS+DfyZOw0hIFJcffh3DjYM+uUYE
pgMMoHRSRrs7zjqrEUCOPS928n+ChWD514Az2qFSQDCrv+c2ILCL1qTElK68yO0pmWE3vkACnWy2
hf0TInZY/S8Se5R7DgfmOmcV1vjhCMPgAQSvV51dGnBcCm0rbvGY9anNm7fQa/0Stq51JXypTxNa
NWzZ9XSOUowDwJbcM6nB92ahkkHEaxBUtfk6EXE4IygETA3VrnmTrCUN0FMorzSvaJnTkUsRDpfA
Ej0uD+jLBqoKH3IkaYIJgY3p5D0AJB1zQehiN+9/rFay7YxVQHPybF/LMZb415mli2IXote5Oqu9
Pa4ICIo968OPdUaN6GvLXIIBP3pXwO07IV+uF5wPK7y1gb83Yo96yz9J8rLXgObqj48jvBu3/hUl
ASzqf/+hdmOUC1P32g+RMOKJ9RFD9kSGPj08rfJyfqKt7UigN9ynVCBDiAsesbi3h+fS3RxCebld
mh1F/IKidXUKuTsGZv3fmQ9XEJdZvyO4KkssgzsDCKKZBp2iP6l5lWw8OKcWbU9Xki0qzfO4xfBI
16X8MhUYEMa+Z2RdOr4W2f67bSO8Y2ynkz23bHVGwhRUFpiEIo54hp9LE0iVY7ZvjAnyARXBaOtT
vk7pOmh1gNYuAGVamyiYNp6L2deJmxMiTO+KgsxUO+I+MioE8kUbeZV+byFu3WMKt+Xw6n7bGsn+
wZEw1XfJ0glTMpaPtMOO344RnPxe6dN3Gjob8DVdd+rqjCZ/DuU5+1wfU/CjHBve+jFup4E7GYaS
cUm8PJubliTNsSyE+xeDnVqn2AFZsjmvBdsx/ybFo/wYT9S1vYYL7T42Vu0QFPsQ68L8gN9tIUEG
Vn/hzWRCVukQ8WwhvFf5C/XUvPXM3pzCnXEi1efdCGOjv5SHjaol2ejzpvlxQLxuC8JfcG07f1k4
5P/m/vL7utnb9CreqhGVEqm2EEfI7/v6ScUMk36LICyZwfn5WvTWJFKd38ZXo3qx8nnPg/nZ9k3V
FQwSKyTHarqJ91wXkZkrWDZ+FcnYAYbW3ExCQUKcxHmHZuWNWazvghFkAuu+m399BJePjtMTzHjO
g0J8ItkxvIelJjiBoaRa+DN3HTSLMvvKSciGLfsqdMtQbN4YWDZ0mwxw/oJyouNhz1CIDOdWQNhn
R0bZlCMSmMOJolw6vE7A+heWCSsfPq9q7/fGqDidENplvCPCdfHZVmVVJscp/PD4eBPCAClfgmnl
4pZW8lorp3V6AHZ3Itx2M3Sme4TWDV8g9Le01hkD1D2Aw4A8B4iOgHl/0rKVwLZdPEqCbA10yJgp
vJptX+rcAbMuMEvVfASMd6lIwTKRVMTmKdL+LHr6VcZ7PPTSnrvDFh/cEgWuN4WOt/NRaRdeXJGf
14x0pXVn9dO8G+muo41XMqaBCom2jUNaSXlJogcfOqWHuuQJmO2jtnpHE5Mu8HF39vdvVZlQ3Lq/
I2coYNms+J2YMfHgh5roPyow8mV8CxTBon+zftpC47rZy4ml7NscHM5B2s+vaAoNUwHjkIMWyFx7
wpK4gpanQTAzi0/WCuzaAMFmL9BlXdmNyh4LEganktR4bjGMm++SgsgGt2LP18JKZkrACMw4rUyG
47oHFk+V3BpnFOJsVIjyHYOcLlaS/6D0Ovzn9NXTQWwgxjK3iF+cEE/t9T28CVyXnj7xPYj8ucy2
oKGuzPc+YIzUUsxMr3CrhqJCPC6FYir6yeR7JmM+zSElChUx+R+DHVCuo6CHrKf0fnN1FWm/PaNp
nj62RPO4xTOTI47Iwo5iV8OSMktJYP9I1XjwNDz9d8CrZ26Pkgj8iO9OaqfHz9PreFpQs/bGzCl4
EQnilnqMDyRWdfwu8f6MO/YU+K5tRQNg40McwmhqsqqoDlC0P/14pi4P7hj1bzBawI1niNlk6xrX
bgmkwkf6RCZ/z7VDsvkDq8aNiANdvtsW8Qnm/hs6jjHXAykkrrDLEg9ALFjEl9+gQJYNR2PvUcl5
oYWEtlD2G0cwoJLkF7/2QSWE+nECaYG0QRCrzfFa2DB8IBu30EqJ0XrZOeq9hVnXxCI2V9CQA2Do
P1FNcbfaS/FXfcYZVkrkSZx9oBnJcWhpYyBeSGslm2Wjt6yKAJK5MnZ2QzxUIW/rvEqLUqC24QAM
O1PWNksy7ecmGO3nkrj8J+S1i6kkZCSJ8dBy2pXTZJuxBcMCS+Rm84aCGawhSeKsxtYfpU41btuN
TEJgpmBMbvqyMPOxCn+GylyRheC8H7E7Xnv8dr/ORU+dXRVREIjBo7tKOwjIoW4dZQspYnrusG0u
F5YQopay7F0FG4zEv0g8Lem0jWmcyCMnTRx+LsRVOdja2zXcHSC9ZIQmrk1AYMpBtVDWXaLIAnTV
UUb7NJl4OrIVvbu87R6XwqDF0oCQIUJY5NXcNcXleqNT9lSxyts/9QR+Szfypa2+uGk1Wv4Xd1Dg
Q/EjhjCR2ArahymY24Xk7orPBtpwHYyPrI73ji/CPrOsgG2gIIrkhrs+Ib1v9zP+Asb8DV3+3vSg
925hrRDyf7IvpZOuMUkf8w5yKCJKsrDwZamX0qE4JlJWOKQ1rJdSd+3G6urBm4wR5zCXpZoTsiNX
Hp/DBhzo+3HGRXRhk2ofara35aDnBMGZvuea0T8GcP1mo7o67ia/W2xBKgpvI1DpmDmI7RX8gSK7
pxe/Ssvr7hhgHOlIvD6ibCcy+6JS0/3+aUjo67H7ay/1ANYnYZL/+QCYk+jpLO7HhE4QSBixE7aF
ibStVPW0BDeQpSDJcMTDwxo9gJApEVeRAuTJzzT2gaIojOCkinS4Wu1tuP7qpDmEc/9Bdk1mfV9x
w33n+VdfNeTBmtxJMiThs26PypwEIk8mk4NRSDL/2G4IZAppdEsdVMRanr5mTSNVVrn6sq5Bpu0V
p1u1jBuTi2wJnt9ozVWXc6ZaXr5P2XmYClQ0JPJevHJEc/sg60iqd2zgEkUASI7Tbv9hfbg41LuB
RISj87jTCvlQ/wJhUStk8NE0zkY2ysmD4kKz9e0tQHHJNvOd+RRPwZBPRfx48roSquSlJw63/JJ7
pz9W/IXwJJxWoAOwmxiCadX0BysPX8WOPcLpqL34ROtCrK4ePq50u0UX/rObGZEfh5IEWqyasxOs
bZhXw1crE3/Xbh8vVcIJ6YoUjKzhdL2kN8X0JTm/5gt/UOioPC9pe+rxh7zfcEuX8cnPu449A4/Q
cd85/HrTnvgrpbo5acUdobjP7hdlT33ion+Sghm5xSI/94K4/RfFzyp2lw6hQXDn+LxqGE5gT/Xq
J/94jAXwPV7SiEjXNN6VEBDal8dxA0a7clIxOa9WaFeqwNqOwjjslnV3hM0CGHNxNdtdpvvbqI8N
qdUp0Sr7cVsQ6ndJzyIR0f+6wj9wo29rx8QodV67rzgNunVMjk60av9IpM0ZTqt9vFSVq5gtk+jx
1QloABJaATqsvnIOnYSa6QTegOhS0NQWbH6RtVPQ8mC6DG/AiNqPv69CrZxql78TMlrKe9ovNjUB
/nen/8fyKkuLRunkHnTbJxsP2QLEikUINafhDTNXsi81zGPk/6+7Die68OtZRliqx8UDi/dF1QLS
6CFvkVmpE13hGqaAsHn65eMTH6xLeHF9u1UHt0t8P4hgPenFm5cQc7UQFiCq+B9rs7TGmDiNCZeA
P4kGJVXnJIPtdyRCj79h7RiP8T/IJYDlsEGYR51PyVbFDwNOSDKpP1SqgnK1t6mpllrUZPTqgx3q
EQifqJmPOh6CT4EVxum4etaZ2mOYQ7eadAaBhb3mMaMo9mObFtccxwOv6/nTCzOMlk44RSgQtU+i
Er6CeqeWk1P/0sPPA8criTwuJd9jOcImtAy0tl9hQQ1I9e9mk2GBI5b1LpdxUhWByS1m2nMTFBRw
dHP+8KeLRE1cEngLpWx7aaJT5nau0t+2YHX2YxzJyvMtyyoipOw4/noZG9JIJHOWFYh2KdNYR2n8
6kV3g88sONCawId4kJdzSBKt1lOziDsDcjuKhrhUSIOstq0t/d52mf6BN5oJc6HrLQO3ws+/Fe5v
iP+FyJgweV+WtOUJsf3oBsWUwhCH30I3g0Q3cBJJQAgaDhMkm01gZ9xZBJTkpwzKmBaPAHj3kiQH
MBbfFdK8WJerBQ5xs0TlyHA2yA5pagVU4sZVUSqX86T7nMtvGA/0/Qh0zU59o9cNdcf2n4vJRFKV
mT8PGH1wYZtXgIrXvcYwVf40nxt1kjfOnTRFB6IVkZodfuELRZd8ZxADMkeB3vBPZ/P1U3MPJzYp
niUW4w8LzeS7pnKnR5ErTuyvqE/yio5jHYKGu3yQiXZI/Qq0hwECIaE3UheAbfhxgRQTyC3Zfly2
a9K9Edn8YuUqyzzz9O8Jv4/LsTeFFNW6KqAj0ArGNfzossgORTYYqykeCLjTtKBC53Zw6ff7vP36
N+lWxkiCpCuu+fZZzGY9gDPTY5eFsUN6ma+I4s+yn51611bzGKtti95URrupXEw++xKO7FpFWoh0
tJWJWbLsHKoZ/QIjHzYkVlT25zWJ9/lrJUI2H7bvgGJN6RWMw7Jm9HH2sHqrkMYS6SsEPVMnzSzr
RDabbR6wF6jN1Uqcpcgb2GIFib/soZ92ZI9ySyfgOV7U8pSLz1gd7P/sf5qL4hZrjWsh8SekXGzk
q2DCz5bsL+9Da7ZRxLVQAHu/lOZio3mx2dDGcDk/LKu5+sidFoVS7r9PGjXNIC5+pFapAdbEjK54
sacSY8Fpz0IzAVJwXSWITJb0L4ppxy4DsjDvf3j1aM9/AmTO6hJUqfcKr3ZdzkcUc8MrWDX3WJg3
nIesUaXEynluoOfSlQlUNt1lzXmeO7lOc5L/ByRMALRG0v2Ki3EIH4YaFgPCglzYuDgpPJJjqncR
6Tc4A6EA9dtDH5DgmJ/CZi2wnGbTpRQVO53DTTE6YTqWZPIjhP9uV107t53v6ZzDDzGiFSggySAi
q9gFZIbaG+/B5Xyt9jB11+X2kSjto4DRiOKevhNzfUC4Jb7N8VS29e720dD2VMD/1PK00f9PTqCz
xu/TOPVCSusEYpFtxxlzvyPPKQuqD7SZq35J5fEKxWWmnIpKuqGUHU2DppLDdrFVd6Rbf2OrgxbF
MGPfFg7E2sXU31rOkPLaFmd6W76sW+wF7iV5lM1OdUwIFb7/HCDVx2jtJUFDUFQ8Oc7/duu9E2XZ
1wfCC6gRZlgxZJX2bTBqQefuvzvy4vn0eLporPGrnMqiSRMC4Aue5E2saFcP0pDg1pLr50TVfwQO
YeHjlzJ+l1i4Gs8epAR/fb+dgmlM71Gpqip4MHzwSbNyFVHW0uhKLlrb+Wxv7aZLyeu/YHO+I6WS
iGNRSZVEWmR0zyjkNqiy+rujFW28k+163d54RWvDMIJfrzUv79PD6yJnH/KdYzj9vkVjouY1Sd+q
lMuuy4CiMJJCFrKYoy6kPRJ5r0sAnOSXAHxTA435a7sdMXVwWUOjZV+wX19pQmy66PjgruMmYZ70
rELjfppcR3ZMN695ieqj7QvRPAK75lrLhgUNcLgedSFIx8M0ptnJKFlfr5oFU31AcajDVQvHGd82
A2X72DWOnEG0CtH6OK3iSf6rT8zKLyEQcHoayPa0OnoUEu2AAm4sKSfwMMhAJoSeXtCiOGvcI+Q+
p8wd+SBrk5DSo3WsUvljF6CwiwbzZpk+EGbUnQLLI6FgsOKt8w1CRork6S+nqoPPEG7nQRmtx65y
2SxzbQcAlwYObCbdmGTQSCU5DgGoUI516lvHVED02+aYMlkHsjC6GAdx7UVOdeGpNogMnbZREVG9
SUMLf3Q07e1EsCDs7EIc07aNr5lgz/6VvaFZSGT/npkuxXfpzRqGT61jzgnp2duybQKfbnuRbMcK
QyxxewT6PF1b6WFK8LLr4rflkBo0i+U0SZCbjvroI7/EZQz7ougsQNCRv6PK6G2Gcd5qnZakoTA8
t804NwqgkZWiOz8UY+7A9R4AkCbJIhvdspa5Z+7USZ/xXTwm6/sXfw8l4gkBLDy2juUZVPIvbEXv
FGmEf54qwyLeWRvfh7uN3GT7gQMiwcmBI38I04L26v/nne2JsJq9YnWEoVqODbrI6/DCRwLB8MhI
uEEX6MXP7MlQ99KOUPwR+uOVRIDWydzaozg3+R3N0hWQ53pyy9Cpd02ftx3iwxsGPLRd5DjSsvc6
l7UIXIfKXEMRRoC96VbiXYrFiRg2kOHNvEJNlp2KwCGayQ8Z80WmiKaVu3tKBRMQI4Dzl2smOMQX
Z8MBZlz4QhWtSpgpnRxG/9+b0FM1CmnWyEp7ko0zAZbQOgja0mP1LxK7OT4/7SCHvBpZqwr3988H
gU8kMtpaeCSw6sqSlqeTdcwbE5iXuQmm/AX8HBPZxhqaVRl4iHHyq5brUr2Zj8+Xe+piQ/M13uCh
8+W8ZI24cBVTx4jaUCz09gbEMjAIiUR4lA46dcEqQ0c44H6tA3Is6j5BDuL4RD7J6RM+nYGB2ad/
jApR6VrOcZvR4+4kDEzxI2YbQcwAHRVEneAIpZqwVKlKf7FMNsZbNBVcm+v0eJcPukLlcGl+3nje
P9aOcyrk1JZVaHWcz/zcnwO7eKGt7wqeK7RJLx7IyW5YRSdOjv9VqDvGgqsdlHdQnN4l6E1fGudy
wUK09ds3Nasz7DxW8R0tGSOcDCg+44zTDMLeLUmLfv6sqJO7R1M1/aDpHz4XDL+HOYPV+apAQpdI
snPTz0VmPPD5PHn0axByhosrEmBGTxM7r7/Le3ObfRGP3L4+F1myPXEyLValrVJ19mElSd0QRxYQ
mSRa0DKFRQ5e4YEznDeRRoRGMIjSujTlq2sSS/dKKCBFQCqLzXNDhuO+Se/UlLl3LLAOMRqGYXHm
bZy8xJik+gPauagne3b3lQ5Mqg59hJT+lJehFiboFG/A9m2qb5gYt4wDsLMp0DAmPbgPnjG4+ntn
sTQrVLdi+8NInpf+ZXJ9aN/c8kTP31gCgHXamrmR3KwT1A38vIzq3dzTYoo2PC9wRmhJAioYrAc/
mu2ARJROHUO41rVcGPhyweJ3vBe1imxAlSHM2URmz/97M7ZTIxJj7Dm4rVKBfpYTv4zp2wfKLVt/
TRfnEQreD2eP0UpazFGo+AqsXt6oIpb6HWbBtYmEO4hmjLOjG1X6DtAhgr19quJQI15X6tHuxCju
m1QnPNUvZd0pilcbgX8ABB7Bf6oPtMtZd5pT5Gz2jit0ng/vqyAPu84z4dkj/cWv0oJNAKDQ5dYB
x5h+v/uVsCqtuOZZEr7E+EYR7gxlRVR7Qrod7zJJZkyaeNXqK2hfB/BLQER6WgCFu3TKR779dDif
sHAS6iOe5Kl2FuIk2xd/UbiVbbZoDBjFab/Sy7M4eI5qs72v6GvAm7im0n4V8Oe4ObD3h6kgk7lW
gNnqz55Ksgkugcev1I7qR4SGh5ygw90fYjoynMWHQsLwoj/Zn232K6DyZ1eR4RCqhZ2jVH7tnere
KFOqPlx7x4lC9piquH6IUMARC3dsR9UMKWYzEZwYAK6fsZAYpDp3nd3S8Elo3K3mAMS/wuM7aXqI
iHcYktxnE5TXDfgg0qUAHY6NUDmssNPKwBw4Pk3aLvOjN3Gcrpjtpspx0A4X8YRgO6Gi0B4Zn6nc
SOQZ0NlcKGloC1+M519Wm5uchGOqbE6ON7pKsmcTshHx1wwyfvd33UK90WGMAgvv4c4AuXlQghqW
IDik7XQsnM3tl85T1hDJxldx8ItCwzhPCQEaKHZn1QDcWCyIVRaWpccn2HGxjlgBcaCQdBNRvwOH
aKn9nUFGw4ICg5RXGxmQV9D1h2PkC5tTS0cRC/zA/dXqSvBJTbgWZXT/kJiT1+gSPfeMtFvQbmq8
4hICFyNZHzhZ9S3TjcAds1CcaCg6i6wiD4rReOE02hF7kTYS1LkfhKJm/CbgPfRf79f6djRhW27x
A9JUL54Mr9xJt2nzRQ0m5OXewuqb+33ISl3xGnnHNdvWQN83Dz+Ufs+R3r7ryJm268Pcs6G9JM8W
zBSWty2sEK6DBeAepcQ2zHyC2KrN/tJbj9j5rGQjjTbncXqmHc2iHgUT43jUWpsIoJZj2hqK6wob
FwMS7N31lTL7QKyyzqYLDmp121Xdt6YMh2XGPjMqJC98fQJTJeXlUvJ31B8X7FAI2qvqWOCBaiR6
JGNj470ivoCNkPpDBOB7Lmjm/NiznHgOYTGQyO7pGPD7BJyxfvjRBjS92forL0lxdOGX6OPwmOvW
f3LQ+fabOhFHXGIT8q+HwlX8G0V1Rf+eepLpOb3iDXnumHNWNeZgVwIGjHQh++y7V+Mpvu1sl6Fe
dNtu36cY7Fs8IORFB4q4/oLfy95kgRLSf/QV4NQoMpBBYapv/W9O/rnmnQR//t0U60ImoJYzizwC
MtBbsIItaPVyraVJIg1in3iMf7zPBuioZgQaasoy/jPHsp+vQP0TfRoZLl/v1hedwPQnRLul0HCD
uUX6nSW415WQ7kJxytYWvyYoZdrwMXuz2AcNyBsQLyjBndLKYXV7vQ6yTZIp74bjBNm/XHbb0dGO
aHlY5MhldPb0bDoj1W41Smag0Mwpml4w1q+gNpNPwGX051e3cGDuwK81AyfTaj8/vP+MhakXaNlk
LCOHureL9z0oT/1oRcL8I52HqRGJ5mUXOo3z8APnolXskycGVn/JOidEuRhrSFJmu4dqxb0amw5Q
uoD4NNpZjKmH8KDTS1uFVHpG6xdytilbGYPVuugFIoaj8yZuw5LKfYKUwqxLy/E6NhqrriHZla03
Oqw8Y3zoFYgiTjDpyFcseFXaMBALJZz3PDHk6yPIP46kkeYqKqkumCtmEP1j17awZbZG7Ux6vsov
kbdBZ5RXvZNN7g3Pcj6r62PLDhveoK3AtUNja0/ObSv1rnri8dti3144I0UkVM8bncgIHZsGJrsC
Wa5zyV75q96PKr5LKUYmNxqEzOQRjynCVd6ogy/Uj6L6JwyabDYaV26ppRlct6z/mMshs+3Gxyal
HiVLK00kxnAkNNKd34IsZfYnXgrkMHg/AMj9SGNTgo9L+tJHO0hdHXoueE+U7m/v+MExhY0Uq3GU
fRym36MPc4UlMBEZv2y9Fl7iS3gvi7IR7efwgpc2eN0PLNBbDQdKhNihUYyAnnRL97DEWd5sz7/w
lXQ1onGAFOQUvxx0tKuLvQiBxuHJPwYRCeuJ+aH9AGA9WgVHYsDgsAE2z3VrN+CQ0eZvDBT3OYpB
j/9uEKtiPfatwUo2hTCQBEUaITzIlFtq4rYBAz6whCwvFhhCOJcm7Y7+FiJgQfJUL9NaMwEYfo5s
kfwhPMw3eF20xjy6/TPx+YLWFyT1iNqwqMS+FSdYt/2w6g+xkJNOl6buU54ZXmnXJJlmlxSKzkFZ
g6uM2faFPnaqIEyqxo0HKCZ03lg+tiz/5D51yf76C+oKLeWJfYNh6oUY58R1+8Vn4S0HEvfrXK6Z
P5g9GFlJ5aijPddBZg6J6hNKOviiq1eBh1ufzicmrBxe33Ttx3yigumn/z/6cd9Y9Q0ipeFOhcaa
vUZ+TD/nJI6eGVgwHAtF5EMLL7Nd+oqv1wszVX8+7Ba7ClwTdMIy3zKt+y64ew5rD3GcpSi/TF9+
rfgFw58H54MytaYY3lwMb/WCQAHANmB5fvb1XgLefBcplxO3SiGEFcH780qtzS8iF0e5LU6lx9PM
G8ICTMMAvv17ZBJy8qH0+9vPcfmBTHqtxIrROwRO56LqO83lFbm5tU5+ZZXFzh65wv1VxTEZL931
ACtj/S2nGYb0rfBqdVTyW6xS729itGmhwWHyLOXf91VJ1oAeJQyZQ2XM06KzdMPD5/s4HdSJF1uR
urXD5KTH1K1gJaCOJswOoz4fqAFQ/iXhN7Ej/2SR6jrYPh+ziAX+Yc2C1f4lvatoS9KNognDFTl9
2XbpUWgylpy0lh/7Y9PlVZ2Xxduca18kaYaNL8CsK21tsY7hM1AqyTzRx8PUhYoIUmrap49KZKML
X52ChhBunonVwaCGDpbTi+6mrtfKzLzOyGce1lR8/JJpNkY/cYHuGpTb36oQlbwJgYxxDxOpICh9
YyolOzdMkMhiBEE5BqC7xzrX5VmXpL+y8XJb4Qx0qLYPPaUElYI4AlLMlVLn2fAWuXtzDvY3KjOq
8xWbOE8q2MSc91euL1fShW+6Y6HlF5kmv2+pgwC5HL+HOuDofb4vVPr4YWDlk4DidWvnjefKIUKM
PW0B/MTLqhnHJ6w5joCHbGVXTUDdlSrOAYti1WTc04ejBNtG65SwAzj8tj1WLR2uFSI/7d1YcvGM
r3s24Dy1icPRRmsNobb2Yo5JmRmZlIEgodqejaVnsFaHAYXvcx9KnTDqf5CQgzVWlaz0XT7VmVtz
ebR+TriW9pIkxXovEONDbRtMFuKhWJheW2jI2AErWpuqPEVwMZEeKyO09Z6e4fhzVt9fnyBb2kdy
FDuaNvx1JuwmwL8Dm8Gh45Zu1WWOowSo/Pc6J2Gunmc/+gJrbsauWolk9dni476N8+lRG9xUzL7W
yF+0osBk94g/ILnRseAwk3FOiDaS8GgTUUkDvtEdvqkvgyFDZZVNbQQDHJq+P3sBFFAz0TnOrbDK
RL31AlXhnCTieKFxmurWH71zmgFDMqtCIuVK/bn1Df6ulTuIq2xUptVW9w21sZ/7jRf+0b759utw
WIPKc/3TXTSm10Two1++9uOLSP+zY74G9/nvg+iAQtcckmk/SyntRkUVzKTvzJzz3Q2M5Z9g+STC
uv/zuN9YL9Ll5Lw3v/tviV01kw/hGD1+QOxG8htzQewjJop47WLJRF0Js6GXMHZgFppsqZ0wXp/d
5xQyGIx0vsY8/9UE7shk2Q0b6XZha81MZDsinAPeTgk9NexTuZaaVEq1zlWqqHRo59iGVgDcoe4x
ML2rqjhjNBme7pf6mlOtwQTnxI8qY3VDZLrhmjLbSoDS8J3fegWUpkWzCR86oaZocZjQpEt0UXMh
qSErIA2ZVctQUdLUZ5yB3K1gb0RWCa+QGhMasR00eW409mQK9eULf6y2nFx174YEmD+b42rK5X9O
ONjmHHMhwKPsVOPTAVwIUDe/k4EGUmPHxKhFB2F0aMfC5j1pPM3+JOq9P6wmlziLMjKUHxpUp/lY
CrBfcWHV/mj9L/c9WHOR6y4lEosrg5fbFbYBMq1n7VFIuMGqNG9Ehc9stNGLgjEqE3QrDtVmg/TX
FGsIeQ8b5LXfva44BcWO8c0l9Bw/pqf1R9hj51GFiPrrkUm5M54cIXqBR+cuGklFAEpYTYaGsp6t
Ge4VDRDV1KJCZBaU7tlEF+/fQyL0OcRZT0jLmjNKVP3cTQ4ppPMLhbZdIz+IPqdxFeDFHmyZTdz2
uffMQ4vGn9PZbQG5ocJGV+Hbry3tgx2XtR8UMXski421a7sA8Y4sIf8bH1VLUBOcZwK9H6/NWjoJ
69M/NXkHsT7QF4uT8NIFkAjGSjYXiDHTyLuZ0BroXlmwsAtgq7frF6hjXWhLLkn5PCLy3Jb1bTxT
uXE9IMdsXHtJcI1o2Zo8/yRe9bBp4OHCysq2N9qCnGc74hsc9qh0iNo6YXZKOQnI9+aE9YMcEDfj
X61O4eli4kwhb2zTQikZNQ6xx1bqoclNDH/jWdYYl0HHdE+GdaX6MBhCVJxOm/ki2EY0BPlTqhS9
ClK0b8gJbreBdnbkSXaFvM5zZCoothZaym0BO7bZoV6BrdUnnyFZEUx44/55qvUL+GBoJpE40Ir2
TfmMLlqE+becAMqtOTTqoiB8ec/GAgFWVitfRMmnv6OrpLoqep+chZZvFVM6d0Uv7sKmKGh+BfrK
QRIojt8mnfdGRpBy004b56RipWbX/CrE+1SfTYJSJHYSzROmHSc8azqZ220DpRLYXjg3WAM2Nf3y
+jbomtVelvSCggzgl0L/vcge4fBb7AY1+ME2q91w2Qwfx9z1REkEezEiD6YYnmK2Fx12uCkR0uEl
5MlifyMYYFE2N4vx2pmRIon9JzRpsPaYGlhrouetOcn9AA8DJ11UrmfiBbUIxfnQkrtUaTsmMJ81
+sgFgmQ8ILB8q2mUCxsjAVlB/BGj7ZGtDIZHGfOvF4WT2nfTSK2Dd3qaR+VpQbHihA2m92xRurtP
bMe+z5dK+Caq+dPnsUtUypCuKrYVH2VsmF1+/rRfXFxLalWEYqCg1lzb+tWpZRrO8Aigi0FyA0uK
UIoqKT7RiHo2XuBwNN6DayOByO6obozkM69Azt1zzE7u9ZHJAmNbGGuZeYVJ0PqUqdcgjAWPqRgy
NSh3R2ecewkufYi0GbRZZ1Jr7x3mdzn1lWbEkXILvzm6pXEhZt0Cn9dtMoHBXJLzNPQQsXmoFkQB
KTY4je8u2IpCK1q/0tr2r6qVtMAFtZ+wDx6jH9MalvL0YrYy8cBY9FJtdMwlxPmqv8SfOvF/yJtR
mY9V9Jvfr3ib2ucyo5T2Gj3KSN9xXJFFRGyQaeCqwFSLB9u9puKHU5orGbfvKME54EUsfMy0Iyn5
ARGK867Mq7ReKOOGVJ5WI57HKCI3osnyWhOG/O5CkvM6KDUmn+q93+aIdtHmNvlcKw4/SUWatO5y
7jTOwM3+V9kNYXSWhfslZ1gmW7oC6BWmaep453Sqwyit5jdD7Fz1/HeQuFcmkx4uhKAszRxWZBD2
CXbvA9yOjrQAgroQ2vTlCXyJJ/63fXsMT6lVNPzAGBPw3c2oZWwM1nq4LvFn/RDYWEl3gicPolgg
uewKHqtesogzbpxEYfTMPVfzL2Y7W0568/fe8Jj8IixkUbDk1cENozh08cpQ7zoLoGi7U7+6ak0+
FiPfFd/4KT2oVlok0C4jqJ7wFqcUkl3Y5Abet/3qTQ/ViqLmYZxgwWz2CFUqK/dOsx/MLrmeIK5E
qlcAg1YBbAv+mrCGyozrlPJgSDmD6UZnFwPx0sKCzHMCHTQm12b5/L6hHcw2NaVnjdZ745a9xzOo
VnYavJthFmXs/QzrBJdC3BhPDc/kmHdahLIAOgRZ7lMkjPorjsyW6BI15N4teAXHhChzFaeWuSK/
v2JlN4+mKQCkUiKdJpxfXkBqDuDxPFswQ2Y4rcFPOcHkrs/25M1h9szOA5ut4Pg7ldnF+htXuF5v
Xy2JIFlj/YxCH/aAbnofgPcnu6wwosDUpTMM90oRSbhjm+zn33d69CCvGIhXTptOnN/61ld3MeD/
4dl1BPWGXE9TgVD6hYl+8YFj1kKoIVxMcCHUNuuMLIMlJOvzOby0Bd/HE4PqFfvIjEsVCKVX7Jgk
oYdbeZYr5fBxZTr1sbBrTh383ytV4buwgjHf3daP6CRcPD462hPJ12m8BlhqvNO0FmyLFzyz3Lsh
e/Vh3GdoHUwGjyn0DWzSLXRj0C38GXcoC7p5TIJa/DfPH742IS8SBYZYdCxDOEJVlMSlczD1MtQv
uijJdgSzhefdleaTXAm9hv3oatJkBZqCBCkPhtJtMf7BuN4S6QLFb/5Tk1Wi5cyFjvSzcdcQU2Or
9jH3w3ryPiyeyf5m/4n1yqBjkvb+0MRAcoczBPTNdkrB1ERZjgO0eoQ1BOCcGt/htO+7OPo9Ptna
tbdkwMQwxrOfjbKvtUFoPhBoSnh6llZYv8dn/7ymUlYyf5rjsLWEjk+yRAj9vzDuxohhZUaP1r58
F3kJBBeRWbyrI698wFaUDgtCNSLar4T+XIyGGUEMoFWz2o7lRPKy96FCOIXRcw/Z4YbbcE3BTgS9
XzKYsfo37pn0Xx3nWxDTIP9/YhkeQAAqTrZ2a8RdFd2Nl2C6mXYum8HlXVFUGjnwwHzViJZ3xKcF
EuBGCwYYXd5nidwrN2AcFhNf8JP4857bfX3RGA6AypEvwnc1GqtGKF2Hvg6tsJgNqtmGLugbU7qf
QLC2d6iwP6gaR9kcS0JuIWJ8UF9LxeJS9Pn0X42SbxQrsJEspvNG3EF3AqC4I4VIQvxar6UUJvz4
Y4Q1gZvQ4xXhexghui1BHjoh+ZOZWL/ifsSF/OH/3+2EtXApF5k1t4XhQ6fFuv3RdUczBpfVNXa5
hsDDnjF+ACrfFnicUKIgP6AmcYnBAFh2H80bfaZUS6kjilwouQ7raVVQc9SSTqWrGpkwbrBbO8FA
zPqPcL3RADdGY2HldUJLtxaSeW0vSh4p1bEE5d4UmnpM3TdPdqyuWbwjQzxHX/+Me4cA6RNm98lB
WZlJXert65AbQDWjpNSwwPFewmRcQa037U/CMERvEltw+uD/XX9Ocjk6H5kvIpH0nVa1+4DADfwo
sjOPi5FZ4OH58CRe+MxsxB9J4yG8hbcvnuW6+JhQ1PDaNG7SOeggLXOyIeOGOevrefyXu7B1FgtA
/awRoGc/Q8VoK7NUEK5Yne4WiZxUfUmI5iF4v5F0qjXe8o00SIeAQ6/heYccYZxQyW/NvzO8zniH
Mq8BqDHKeJ7O40y8YkXAxxN8v/WjVpl6rifB4vbf7O3233w8qYQafWc6TSr/9qqsIRjas145rooT
Ty3jNjhupQA3B9xZaMlguXyDTvYSmLJch0I1N5PPL9aPSyfN2zu4V0sEUmMEECyexqzr8QkjY/Vb
f5K2qr14s5T7jnyvTSkfaRl0W6CTVs6hhtsqppTKWZcY5vSTkUthNb9LFoF0DoWHxOljTtS8c6iW
zxfVSp0RgDH53LPD9cqidxOHII8H3yPIY9NRq56ph/2Ce2HYLbKGP6T7hMRtmxLLUP2BHegqbe2s
Fa/Mz9TnjW6jRjD6WxQjRttyrT/G8V2tl/5bdTybq3Rs6hBhjVQRhCU2wK/b+4e4wGBvOu7UziYZ
SRH0J+VYf+LLn73IoXTL6+wAdjo4qUg4y/gAhKSasmv2/vjUpIQZxyW3leANs6xIqrbo5+1bwW4D
R4fUp+mQXf0nq5pThICT2aWfc71O8D26hZK5/I1E7iWv9QlIbRAq3uE6avah5k4EpHUEe0JbXpex
NVSWlN5NL7c2D8Eoy3WSe2jp3wj3OK09vYXSmZa6a3WsIi4TUCTi6bEflvCpWl2np2q65pk8VM8b
jpx+s2n+h5SSCPLMd44w9A/0VUM13WjXTTDTGq6hnQQ05GHYn/LWCG0OmdNO01l6sedzHOyJxNrx
c0nHnK2HFCbT4hWUaxZ+/Mp0J+vMkM8lkPlkCD2F1uh+FS5a6jl20Kq0+up5WGSIWzCmuSN70GGF
OcmWvau/TEX69npd7MtD/HSSozYKthWiSh6pHMbrW72/jax6Zs5YAARQv8K2t7F2MDeq7IWSEySX
V03f3RN4dLT4VjRaOm2xLNVQKsJUnS6NTbGoukmZ1gV15MgH8xDxGjw+dIIWzOS1fMp8MkW4H7h+
ibuR9Bk156MYFkI8V5vdXZNybCx5B10uw+JKH9e2uBBT/DBqrNUX6DcUizKGeYtxhqYGYFJ20hVV
8oWyKmUIBFFWnSxqTLGw+xn/gL6sOePlpWrzUCQtmJVlR4l5cKa3vbv+aPU10acOhdHjGeTnwUsr
DU6rr1Od0iJRZQImHpSKgfFLndx3L+dN4W8xFBePF7RMXzOtp5/D8gmqpg2XiQthhm5tEsOe7byv
li1bXekEG4Yv+nZe/rm30GKSveiH1obWWIm5VV2rH2ezfUCOCwFr0lMWCQzrh5ekeV5f/++DTiJG
sKPGmLkyZh/EIDSVVrD/E8bZMJBzVqY2qMcHGIzga6o88l472KBbNfWVZeMTbRS0V14waKKwce5P
6l+UDgOWthFp5uAt8JBCI0bEwkInCl5yFhzOfJfONHAkMHaOlS2/kcLHMyIl/HgkgH5rRiCjlQlj
gPOHtxA73o8wbGIChTZx9w0mH/9hFJjwlCXNdcBhad+NDJfVxBOHshNqZPqoezGMBmHz4uKYFuVo
APqBvNiwutWwAyCPewfAoZ1O05yyWlPrTWpjbOOuScWoLatgMHc3xIIbQFLpxq5rqfJyP82f5vqc
16GNIy/lIVHAyGlnEp2zPVJTHt1Qzv9mWryoMocZv1J8rd+YoRXlX/Ejxcupog4HemmnI8DZDrGD
jbzi5MjBs0Zfrqsi2O+I0joHm9R+rM88YSfy3SV7SQtsSpvfAWm8kt3/JOeH3XHlyfDL35Y56L4g
q5w/UJIdS66pjBPR8A130SY0uFYO2rFrmnqIRjIFfUCif68yTBohlZWBaH6T8gt2q0TSsmEnPNmP
dBCXfkln19bv2VkQE/MfB82ah0dDN6tBmNdGQxYmdiicSYQjl+vhlOzPGViml0JOzRukojHqLR9R
TRtAqenwcpjgUwtwWEu9xADwk8S1pj8iOaL6pgRQqP67C3oscmc8b6ZpDlq1aNS9YZdEsOAF61ec
NerKME83MX5snxPxA7ilIA5UCuUkWrNcnLpmQEtNNDcPEWXf5RF9Qt6bOtEU7j27OADh7HTw9P2w
JyzOA9o/PzuiLaTucr07ZJCK6pWcVWWYFqzhgu3Gvb/61ENua8wFm04cggkgjbZpbA0G934cE8LA
KST2jhPIuFQY0pRqjYOYEPwrwPDjD1ryoVd4iaJheuiEZRYxMLhjb9G0AoN94+QPOReI8CfhYGb3
VLX+H0UfFiSgR9BYFeZiw33xi8EUaYp11K/NwX/YrwZYHuPIspS+T3Qo3w7q3Metc+4ZHi7F+LH4
Wb2rd3shRAjlS+IjG8GcdMWk9Y20IZ9ua6NiB058AzXKYENrzQcHv83Wu9qdcgEPh7WyZxROfbpc
bgi8RukfDZoi5KVFwcNR6A30X1qyWgidy+pPev44mYu0MMkFwOHBLCdu9NPAx8lV2SNfnG+2VGUj
4Xd5ENsTJtUGnAuPbX5S9GFvGIVENB2rAPGvpDTplKOjqCBjo2eUR49SROAef6ndaXqganCq2kuL
vAe34yFIVYJTFiaMJqUE06fwFtIMhBa4WrYev+TV/7yyqw44OvHK1lqytnu08hTS/lGpatoeJ67x
m8uNx+WY7vksMBtSFI7Er/rKAvQaCs7uJWnwCw+lXdfkTfJtAV5X04kMEGrgftzmFQd+gbToYLNC
3Z+nzMTforC9GftjQs/BM/pzGNaLdSI7PriZVm7JAOwIwQ2MC0l1kmhXYsLdgPojU+CLHur0ZtIF
J5UGPBSEnYbnVHPYpfgf/12vGfbtN5e1yjRuUWslNQk4tP08JAd4HJe/OGuWebOavoXVm2hNvjGP
zf6cM7t6sOHe+H1dq8rSypulsPhGgQogCrrG2UxYKBTzMPsQp83jbMKrLChLJHUZDIOIq3Y2bmdK
O4NCj1oGz1nC2EEbT4kNdvO93qLIJgKTk5UvaLtHAY3VR5tCUdjrKY8x13yfN5uj4h3Dp2nnvemb
iaXNBJgD0Ye/HpCcByYvxzPt2EAWNVhz/d+jI7aroYvWEVvYqF85WinYxL7TbrlqvYnZ803H/rKs
m7jDHVT3EMvgiveckVgy1vg4U9eyjxCn9EP9FMc7t0NmNOcpDVekLthD2zsbS6JNtaSoQttqfkRG
pOAb+kAhlAUxoD0lruxJRlXjF2zwxeCrw2aCQu11Bnq91DotOdUfOzglpb+rrBzIbaENmMS4og+0
jSNlhirl6Y8T6ABhkKLAPYnUl9pPLNokrRSsa4Bm5q1mU60MxqSWx+4rv8uT7ApjZeDLxXegPUc9
iZrsO4FcJ6YQ5Ei2mCxEHXaRHnWtHcX8b7yzzvG3lja0sgVZqura3MBKeY0WgjrILWRQFKIbPcnf
wSIBlcrDWGBuFF9j8P83Ia/MxIfrC3bZ+eTiMCc0166PWANzOhr0Gp05cnwTut1BzjFq7AjuKfwI
mxTc3pzxM85PC2c3KFlCjW4laH4e59dCpGit7glAdA+e+1kL/cErFPlleujY4lGt2p46YXWrbPk3
lppEYN3y9OzaCYOkVmNJJfaoyITE06TfZcSJoYZPU4VvWgEh2el/UZjLZ4/DDdkwDiaDqsHR73o/
ygcrdJB/MqzLMlOxmvIMhaw2Abadmio/owXz1LNqqkUsuWxKBV9elh39VahPoZ4GBYpMneF6MU3Z
Q15DloD29Ekj5zZfhs6Ys1XB4ypmbeDmkQXsngQoxLk71lzhcEQV5mwAT1YZH3GtPnY4o+m4eyGr
5mnzRWpzfNGX9WL5PNEkT32A59k4xFGLmfxl8jhZpGIqDMAEFHN5jwM5XWHu52wbRzjHViyyHCOY
7VERGuARYS0KOPdI36i4pCqjCZikRDrG979V8FXcCxSLbOv0fNpYdoYMs8x5te1RpKS885nqDOgH
7snVU48FCyXjYE2Np/b5FYeqi5zehjzh/AcyqvhtxJp0s2vQ8WUCzngIxdjKIu0bh1ldVWzRT/jq
i1IRFsqpi0dsV82NeYY9oPxHPnPEHHHYqK246E0TRln6X/QLN48ZMZh3PE/cjnW1RYA9rOyQZYNy
9ORKIx5wfgKC6OFInbGJ7qzyGih8hmXOTYcwf62JlJOy3ODD9YkkJzFT/mLn9ZHUnXt4p/CTp4Hd
6OS1TBpvcLC2orlCK+dwBYsfCaJrGFuheWtrKrMCD2AxVkzOd/e1HYpjF3acfWlTbn/DvEcE2ev/
p7A9BwrkwyHrdVurlkS6LFIFOvem/0d9cve664vAqL3Kc77//LmS0dkcswnR6GO/OVBTWfhzToCl
6gUTjEo76k4yU4X8NVSS7Odf9FFB4+WYgTD/2aCZCuHLdRDd2JmzMpW8So5FPARM1qruJzqxAjOK
Dg7nkO0TVoUc8+Wl6LUGebuMgdlMBIR9X9RS7nJxq7OcPNazdKNk5H4cwQE/OzUTKqWB/7DKp327
B/N2WyrLf5A8iONX4RmR6WNUM1vvOPW45+wGWRHVV8zgDo88PKFHZS8tkIxa9JIM81CcYAK5M+p1
OSrtKoB9e3EuTpZJRYyxZmL3Lg7ki1UdouRMvGqi7ZCglgVASGJc4rOGxy7xkl40sffMYfG+lKNw
oAoEWvsA05ylF/mFNjNHTLwmwjlM9x9CTejNac25NVmIWccEJ0/j2TU9TYgIGPn4KU2rw4/KvTh8
Hfhd2LUWFapBMSvJosCbndtqjBgQuPIknMMgl+rOlMhBN4Y+hgK9nHhpw61yVifSwrODW0frOflH
Slg9jHX2271QScAqPnzYnUbrT+DNCGnTflB+hFxbf7fberX8w4dGyaoBhl1YZJ7r4ZlGQnLUj2gr
xO1FKMf/uM+1G5vt0XtLcATAefAQtU/TApinUmI4y+4poCNAruF0aPE2IdhYj+NN0fnpQv2XlBs4
7Z1FmpvKE7YiON5WE8dRN1YVABlRTQ5VRHztzXg6NJ8A+cc1Y5VncS6EqoA+0vFSuQiMyuXB/x/T
7i/vSorOmvYRQLR+0nAuq/jeLeASuEJ/+L3wQcSE1BfplGFkUqmv8lyLX6VRH1U6UBt0dTvyOmm8
1jr8OJvaiKnUcZJzN0U8Z6z0PhI5H+an9GSgLPFsdOheaPvjcpbvOTFV53CWpLkSgtHAy7O2Waes
YZYP4VQsIipi5LUsJ6jqxqpsJS2Md8sPiVAGiBK8Rdr791b6y4RQUdNu2fSme5QzkQgF8GmrGdt1
WVv8752z1GIkRvzVdWMTbQK7l/pDl7SY9bJ50opaYiQFyUVLOlt5yjjsVL31V8s9LCuiXVAw3EgY
0FItAuqXSxsDTV6g+C9kxp3vUIeTfCO8diS8PF7WjNBOIPQqDbTWWiIThRDj/AsSp32vnWjSitB0
kY7axowYdIWuuUuo6lsIGCZqzVOXwlhjfz21SbqewLKcKvmz2fZ/ER+AzCjG9j3AWfnccprd0Md3
uV6pfD1TKH6lcAlAN9MfY/A4E50DJV6fEBtm0VThXh6trzdaGUF6bDEkVVpbbO+OUEE3iQruu8bv
DAy03E46Ve6f5/DqCR8ljImYEo3Mrr8lezdBE3Ys9HwCBX+CHt2EoIz/HcZ7RhdkwJXBNFodeAIC
b8xK57fEyfYdQyw9blLC5yOCwgNnxsuSQy7nDlwjyA153ZEdSp52qt9TdVRTDaKaI2V5EBGOkM50
BmhCPefZaF17V3MAWK3/40PkuE7noHPEQ6/Mofh24Fsh6xWe1UllX1b/FSOOwX3oFLCTIZMr3h+k
odwnZcQnbkIYgu5YufXGnHJPSoPlt5iimcmbLsCBBY9itfwivYJnEuDRx6IKxm8bVLlCg+s9YDvZ
rmaP0fqwWCsFanL7Ya8qYhWaX5R24e7TYSxXTix/h7lqUO+e5FrgHi6XfsmyDwF4pQqvef7v01UM
tzAOQOfg6oAUNygGaMnQbuQFpeRlyrQiwF37+kj2YiPjbo8vnJKZaXcuoRxOXEM+XUcwpFu1rxYb
TLoo5DyTy2F43yj5A9lDV+4v7clJNfbbFtySy46ajnjZaIqSOEa3naLYGLwIElZBgFCruY+WKF63
liqFFRqxj3JQZug8cAdlwA0zbQvCEBBXowFn3YwlRYTGp9ggY9BNhuLMYILo3Ec9cs3fzkbHnBqL
mjCzqQtQmHiCBfZkJa6Iq5pN9z85qEwEfuGrShgfJmNY1mka32xff2JpJrVbza8BoW6NIx40ERKb
nE8K8WMHuT4ArSOWtXg/zQc4dxS8cQp0HWVi+mW9axK9weASq0Xzga6hz8NUGSinOdaem+nNexhh
LrBXMNdeQApYm1HzGBLT15UTWuiEMm/6wu5XVQt4EDi9k7lJgrfXOIn+EBlG7XwfOP8UMGUu8rD9
9xAjc5GMNBA/DHkyXv2orBC1lP7Gk0Ph8uxt4+NkRBng0nnv1ScSnsZSXAuxb/rOTXrWFdA8egnA
0RhtcYkjW43NiiNcDs0yTPQxM9fqcxrqnyh+acIN58Q/trNsto1LlCciNoEPCbtkJG5qj8okAfTR
MpO71JssjokylxoC1IgJ6tvME6MolOSEdJjBLoG8W9mhT9Y0SC/w1aqfUIc/nvk/eq7ltICBocPR
j33DBPeb26aXcEZ4IbxbMPXW4VDRoorPWqTFMOSoP9q7ha+E591EjfU/GYEg0t1D20pUptDdJ2Yt
lfFNJtlZTahuz+sK9/+vSp6NJFula9ErSfgvwxjcbq2qqtQ5caqulE090Dao+ua8GCoy6QpYiAW/
NmCgBdB/MN32Ph3zTKFEEjD72W1r5HVYdf/rNpcHEo/ltkDRxOb+kxSQYQmCJ3aciahD02yGcaeR
2ggRZHe9zS1LJlJhForZwXywgLF+Us16W1GUBAc8nxl5s72M4KIuNR82EqsZduA4bLEwbr62ycSX
47fV5+CMIdthssNqdSLPEK+4xOmpmiAoaSzXCSbY7YiKQX3c2XkmhiP7hsshhd2ylsQPm0cETgUN
7vGiu/C19ULoFq8ostA4zAluDADv2Q4P4RDEWVTW67hAOeKgUvBKBiDqUUrKnlXR1HO2rJ3hEksS
yg5BuFpe6kkDe3m7uTiOBe7OYUkmin/YmGFA51SqS+MHfSccQAjkhB5kbYqjig8aCUNBiNwffdY7
sjICJhOkxxu0CvwSSDzPn9Ox8Yhas4FDm2xfi9qRRNwd0IRVTxYl0nbT1ulnMzjkXY7ZrjBik5Ln
4mh3EUa3v6u2q8gXiAxR0cnM4S49oQxzl0wsGqmRWmeQ0Kx+NdDXOx09XySR8WAvOXrYS3QvB1nU
1vVogQWT7DqVqWoewpKabSGRC3iH8x/pSAOPlU4qTDQ/wuKjSnq6QHcm2ZhSn02KmIrQoevfrPdk
2gUiapRzuFoqmaLpc352miI4SyUyxJ9jES2llRw9cYzeqMe5DnAsFYbTc/S34sEjboO3k+Sy31aj
6+5bc+deZ2/4uqHXrr6/N0dzwyzDaVxA9NEsmvIFXtqEH8RtIygxkT4ScYyRYm/6odU9gz1Gw+h9
cuHYmC4qCDv+IQ4aIwdqhfKzzpHDxvHbLl0eDlyIFrHBuNnI/cLVQIYmuNmdgHS8ZAyZq3Dq6iWw
eEtl9mSDAF/hE/AY6FXxubEqcUch26RABFvi3pN3vIvE0cEgwyNypco3HB9pIKSIXFCJbDqBfQ0U
pJfbJYEiX6hbCPmtJZ/b5F75UAB7ErrjsS0yri+1bJFl9V8zG/tOk0yPC0Jy/pzm9IMX3rzQ8U+N
guKLQUBUJXhRrWdv8r2fJ3oBeNHcqycpsGlkRegwaiXAsCF+JCJ+2ILCPRh+/82QX2k0ll/QIYFf
CuLz/6zxzzy4jrB8nuzBIEmqEvvkYAoJ8xvS1QAdpAXCylQ0obvk1jVEM8DhzbXpqNbwCHeSwS0v
c+zj5H1NaORdxxzvc8RN3uTuV6mWeJqQTiMZc55UTEz0UitCKpjJkdFWv9TlbG2f/lIu//loicgV
SOz194QgUXNfCsdpZMLSioqnQyvGGZvHtV93TZ9G/O66SSb2MKZF3cTUqA9Ri3WQb5VAioiM8NBe
mfx0ZlBsaWWpYgRuTi/8JVa2gbE6YY+0m1as0pDIcILlronOPR/RcpeLwdkA295+NAXSPDKgQKS9
hXecKbrLCZP2PS0/S0U7UPsc4IMRkDYXE8YtTjkVi5b/bZvgWF/xb1TxMFM6mipfqNC/ZKar99XN
8pIVtw8F+W2fboIHgfIecwo2/Au5RlpHuBIzv+UIpY7tzk8IBWjl2Rmk4oYyhMLriQ9B6FkoJb/y
4ge7SZf/3VfBTBICAV7Pg7uCQdTanj4G+HID45MGotrm/bUUVvoKk0SCaXruz/WKIOSyhWYMg+gx
9fUEDCukOMiXZeEBoZ5r+Ck+szKUXFsId86xvHXkXpIe9oOfQh1BDh0wtskVscc4vGunMLNNCWsj
QTvW/5+b+CKg2Rv8Ui/dKYXeucfvt3FSvhefEjqDSKaZ08djOUmI88DwLOS6ycVeNi8KLEgUGKHe
Qa6gZml3X1Nx9hT7c/7xIAEaiRBQfESy2Z8HM2bc2nx2HmGtX+79S1wnfo66jIkQb5mrDDc9fFNh
bxNGusmZuIFamPvzWGM/Lm8/F35mt7UXWmlaO66GYLxnG7suOJ3/OtXkXQVknCoMXQJX/F7122bP
qspMd91i2zFLPfJtZGGQczIVu7DaIHZOTyJ9OgpaI/B+gz2l2CMC2Dk0WiRPMmWpca9sfoRr4L5w
N+9D1UknWBSx1h26JL8S+MMo8GqbUBvsRcESE5S3ZCb6mqBYbYV1BuFFZ8BPvbam4ho7aUNkRj86
FrQNFJvzZLrRXDuaVJ2YJM7V9nexF94W2HIQlhWw9CxL1dwKA+DIW2iq/HeBbITqsrN8QNNt2bvo
mlIdIrXHokPvjWFD6Ox0jkCk09JJADgjXR+z8UnfL4lz90a5noOuDJjWc5hxHBVZibHAVTJUJGlC
iSWDOzLCuhOjkREHy8NfzsnY/woWRr7N9IdzfeiV+0gitQwGk9pJKpC4Wcr6Y/gjIBXhCopQ79Rc
+BMPkP9M3QIISB9YNDg28ud5llo9lGIWCCXMW8O/q8QJg59quBYO7KhEMrduM5SSn0uM5IdOPcm0
1Tj4vCFOZ90B6B4EWT5ghyEWCMk6KPHoqlRIwFdz2griniMgOwmts5Awga/oiH/4E3/cHOmYGphX
0Q+EGdbJyPd9pTUOe/6Aqc/D9JHDA8GO8/ydtRRsLYXL+9R+dnoLEe0r37fshW1eyFUIXcGjgaDP
nO5MD1hO8E4jQ89PuzZS4sVnHuK3Ur4VTbBTwGhgCP9JFlDgzs68LAhH8CHccSsSaVzXpllHxDVU
LLgeO+eXx3SaN3+6WSDcPocZ8oycrsGTI/D8Qn2LjR8EWlWhlkiz9N6IG2RgdjfO7y/s+GZsV7SO
18JmjCnkNHXsMU627GPu5Z6rAvt0eqjOIfReZ2llJUU4zJzHt5LO6O66tVx5F/y/OpCSW51qA4DT
yMzZvfj+69D14kk9tWzVSPuQtVLgr59V95398QiLdPsdJxYFwRq34/ePFlkFRyBCRRd14R4vDg2J
fV/9hPV2r/6dPhIdZ2jEjnJIk/+wIjbcr4BmQpR9eRVgzRQ6sXv3SUYsJbI/mzXBIprD1fjvW36R
rDcwFkVXuO+/VvPRD2ZTJGGTFuNaYEOUf5pYICVHf8JKt8JsmN90RQ8dICs6oW1PZyHzvl85nzE6
MvU+8cOwBNexLyM2aDQji70M8AeR6AVRRULoW4Ilwc5s5MrcPRAFg79vxCv2tKC/iQieGSGkyuwB
Kng0887kvCEZcLz818gsOpZYUz9ySmCJwlSncXY++FMv4YFsVeJia4qEOVL4WO67dfrn1oyJoLJj
G/jaMSOK6Isd/9u/20PTNl9xvAqdb6YC+DMRd2QYbERxyQDFCulEAQgbwRzVplpTvgrgVZKtmtSt
uVyk9Bmp/XnANzFGs7v8TaQvBzLh/tS6CkjRm5rp11B761BZb4BuvyZcXVXhcyxSg00HkXtkc/kn
PNA8vNGgLRDZ5ZxLDFvZvlaE1SHQ75nPyk37yNTKo9uh5dft8VHJDTpfeUArqZ5xFt3WnM571Kdi
Ms5+lVXZEXETxyt7Q1f8ZIr3XyglCaVNA/NZhQ/7qEP9iDmEpTkgcdaZFTC/tvLbM3qGNq7osT8F
q/rZHAqnJCUJiKoNHk5KItl48JoL1ANr7BMbB3PpiA/PdVVwu/TE5i6o/raTyjPofk8Y0PVmLmwE
mXo2iTMpi0i4Nm31Zexs1AEa3zx2ns2U7z6r/9iAIdmCJmgtfjRy/BcXxqGHXskXS8NCOJ6j3rGp
hylTjOFkc8fy1kKvEHVlsYXJrJcidJQTlCbale2Cp09F4DwALbS3BxZeXupVkX9ZXAOXBqn6yCC/
kfxZ7uyCNSX0gSK3w4iTeQOhPgpufzOa+E6/yn+phfsu37vCASysKJr18wLJj16tLjLKPXBpHokW
yD3tWUz5RMdqA2oMCQsg7ZiAN9MpYmqiqc7TGhyoSgEu+h7c7sxuPTrcmPB0zMwNqgvwSYwEwrmd
MqcnPbbtKjkPLPNj60WF6ZCeJ4HWnnNCO4JZYjSowE+/Ly/ZNDEUxnH96g2a5K8CRL4fEAbe/lmn
x11D5nZLMVpoZXeSOsa+BFibescYfm+kNEjhr3MKguP6W5HegcYlN8Vs7fjojQTdJlHZ95Rw9y1j
HZCuX4wVoFPopZ1SlfUiDAQMVDGjVqlViF3wn8a2RVWuXC+e91Y3iBV1u98H2mq8VXA3JMytILFp
rrmN8K9VjM0LyZ0/uwZ2RymemL8h0gZ4SznAFk4SatMNMPvDLdyBSz/wFMmyTkQcT6PxaxTZfUum
7IlzTUGki1g9oh5jYOJqlg38ZhwJox3vAtTS3MHL1DcIXSA0WBfWaEog5BvePGAfhE2TK14rhhCy
RSFP9/bYh+DNXaCJdnPuk3bgLP7BvdxnxdiWIJNCFPFt2QlgS2vdVsKnNNlQY5M2U4ATHPOo84iT
4591e/yiV1/s6hcM30K7qZ3QOesItTtOdqfycdf/b29Zsj6hHgaUaS7x10HwH8D8SCOC8kMspSrm
VE5Z86rtCLkYozLw19WQ9uL8EmSEaEPbImUpWXUo4tT15irk0ncRWVdzZJtQO6dIUAAKDV2twYlD
7d0smTyIZPpQSFkNo01y1IS6tu2wJ5KHH/pxfgWEau6+R5VnoOpcVkfX5cFfTB0LBH18yDBvQ6up
0nFJRHfnSC/WAaDIA5i0NtPkqjwhDnBAeYqIrdulldTa5NES8afCKL0n9vDBj5I+0Y0O4avbeP34
CeeHJeQVrDhB9VRO9GcbGT56chELNt7mySpGeuE7hgv/MBmPr/MOYvMPEIu2WCCe56d8Tyn69w0y
TeDvMiFXti9JGS3QJ0HaTBbdVb8x1AUeH7FYC72DKeEsIF7thhLkzI8olNUe8N2/j3NZBiO2Wr5a
mnISNpYILhEoAEfljiQvMfZfq4lJgobcr4cVfL66eaU0w2a66IRYfV8X5TdDuDIzttlDmC+w3G89
MHRReiJ9V+qomKMpglwkfYk6Sy92pw17SWKiecXB7S3lPNLpMYAxT4yXjl5rBv0WaZbXlvjD1NQi
3cj+9YykU3xObNBWtj77c3Nv15ya0ccVwbfxdgQ48KQd8ZRlaG8tYj5p5FUc3/brM9qCBJCAIy1v
9u9P7i5MGB3G0ZHY+0bZtoCT/ilW64itcCNkuEwKN3YQuGtBpg4tUCmZjT2ChaqZpzXZm/hPc8fB
CD1UsCcJdMBep+6ar6hKjgp4QQd3BrGMqQpiSWy703jv3UnWrIITVRWmO57/ESrbnV35SLb1isVG
fOQL3ptCnTa1kz2+OuCh/4Ld3bnUp/xxUnEL9v+4ExfT/+HENia3iRuy+bdmauLSfEgTzWV2zArD
DLRdlZoXeBx1O0LWn2HddO3zM0OKwa+mySIZkkE4zvq6XHVSsRJh1bj71e9BDeYTzz2mXVrGmUsM
Dk2uDIsCtLGJ0SrgUzGbS7w2LKsPusw604iL5kcf23YMk1hMZBVDhAgu6FD6Gklb3MCyUCbNMSRp
kgwS3Dor8246oeVgWiIovBU7Ni7wFDoM4+m4DlaXpdMC1mcvcLrlnCaURBn82Un7QGP5ah28stvm
WdeZrU4a4jzrRSPX1FfKV0gGq3peD5ZBwi4P0JydxY6DSH7bvSkVQskE+ozqJbm1SMrGsn4g+nw/
JgAdH/dJf0MKwTEgS72kuZ9W3g7ZirmHDdaiqNZXb4PrUZIqlghT2JlNGkHFH4Mn4pHQIrZB7ynb
c5QehlsNII4Tk7InKzcxNs3Syc7LofT3C5NYH1JV5ml/4fCGftW55EsCYFlzXhHIh9pwhwRo8nX4
TlAhMpCHxuMGpUIx6IRLrNjI5I65GBe1lNvlxigCWv01IDYHn2vRJe7VD83A41xiNAKMm1ZXFa8D
mr6SATbdhgC44fLDaJW6cspNKoM4nICEf96qawS0M1fZGdeXAb/qNIQbjGWtdpxU0xZplms5HRHB
sP1Wz3WCHpKmKHtWYaHsom7tNniRiQtUZuJgcAVA3lTcX+iTiqYS1m7RblLWlNneCE3CSnOlpvax
N1C08MrxEowrOMvQ4svwJuGRuOy/lDk95w6GSlR7BYlZzfdwyl0FoABTXoMcu7h8OvnxFk7+nwWS
LtJOyGgghDoKStOuhztFo2c87Domi/IwiKUjHubR8H/FHUdhlYWfiuIsxXH4ByF2tAOmNNoNeJr3
qlFT0VrSdyKVzpfBGtmZm2nE2KXZDli6oQvRAVs+KKR8hQeJVN8WSAMj/8hoPD8qvyXy3IN07UhC
FO6IdXd6Sc1Ui8hQOaKLMvjFoOQ/LbwfzGrv6ZvppQlx0M8LM25cVUYgjIUmunn0CYbxM9S0pmSI
xgOrO/CU2eLzk/BcmOCcVSC9jUavNnBUCinY54uay81RrvohZfikW18odh+OUmmmimoCcrfBeORf
tFod6SxuvrWkwN3uVCgVmv8ZgBHZnO2MdJgSao59K82pTwyKx5dzmJmeO/uwtaifXELuNHapW6nd
+Lb2GSznJ9X0v/db1RSurIeXq85FUoBC3qBoI40GDRh9oM/oCr2GG9Vwqr/vzZmFxKgCZiOe3TlF
QWfXYdsO8m0Fd/X9uNL+7FySgBU4+4CgL22AL6JeO1acZN20RNOgYqyYH2HdqigsGQ0ohNKgObl1
05YZHscRKNSb664P+ofU2Vym7t/c6xSsnX6q4waMxumv2F8KbUjzZ3Fb02r/gozLYwRTaTrj5Ybo
SnlyR+OgeGmN18j6MAHt1EYOk6ATUcFjFSdqbZqrmjBAkUt7otXzwhE75qlye+5krMQ9fbW0Kd9H
VkKjevjb2zHMKnyPi5XJN0LFakk3uX2eIzX+J0JDeMlt2oLrLjex6A3n9SBqpITQ3FMbytiv09A5
nKIVKJ6IffOOrrkBojgApxVlBkkF5vhPooGnmy6Bn7d1CpCTuk9+apBi7PaJtp2jwQPKkzqrt6pG
ja708yt34RE6f6JHDSFySY5ECYBNYzBulGne/yXDiDzpJDDM0YavdUoH7duz0jYw7K8ej7ap85Vu
7i34Gf2HE4jv8z3YG0BEBnl7AfQELYjoCOlVHdlVy9wBWmGMJFt85rvZs6cUckagjpOt+3bGGNbD
+QZ9qNr/8B6dyK2Xu4/aE4DttBW4DyCsO8cNF+VMgU/eTrCghNbHTQncus/x2S4rrfWUlqj3hmxw
JMDwUUTun+NJseSkgnKQ08fBTJkTw3mrwxrdgpfhmS/KMPWi5yI3defFMgSbvn+8/x3aI8IFkpM3
SV4/hwV8akmozjLDAaXKRXxfm363fYQr0rEnccJqsff57l2/YLOkVfuOWGScVxG7DJ1eJXodkG6t
3Y3mt6KpOLRnVDXvKLH9F4+15rd4+4hY0UCBgJduOCeZQuaL1DWZ+IU1SkKXnBGOMSYQXbpqi4ma
0F4kXQcPez7Q3BhjJmKmbDun3oYsNq3ctdggJS58iPEDG4BbECXBaZzxheUmZn0OotExn+VcwljL
7NsBw2E3pcWpKoMSdcm/qDVSxWsJyuu3VBlPs2Ht0il/OSQaWWyAtYV9A8lNmUKxvZ/Hl9wAjTF2
Jcvi1agE68AgCXS3Ro0EildTFx22Nv6M4glFw9dkmZSJWVUDea4Qh2Jli/JEdIh0qTXTS8lbiJph
zzbikq6lwl53XIWiMAD6X1rhwIKIHT4Guw5gppMrwsJi6+j7FKCf4GBjWP8hfGv2jNX698RVlRv0
Vy86LZDxHDYSk+6JEO26Wjaj4FOkIoMUbAld/e43ec3TFOb04uL+ow4BaVcLizplVvlENVlgDts3
RjiK2J35MvH9mTUijAVbe1K1xJNIwiXYiwpc7C8rwRRNPeZPjE3b4mCUGLmFyPF8oAS3fzW7Lrdn
xDG0NRzRSUg32Tbc0Zs8R3AmaBEr7CImccaOkO9d7g/IU4UcWxCg63X+vK1lxciJeC8PRAF8M/CI
3L/Qm69VJeHnTSn7d6VTp+3V3HjmlyV2tTC67+xMMkJgzW5zXqzdcXJRDtEmEn9CPur2d+yWcDNm
DIcDIzA+xiOjXAtdvcaMoydypH0vepvK1k7hfLNsLlayvaIyWOyeoXVj4VGoqnncK2L4CJ/Y4A68
yRSuijXZ8rITwXyF79Ca+fDoW5SNrl8lPB/WPTyNw1x4H0seQNAMeNzqR/A4MKOhcWPD7ziN/dMD
N7rfWd76CqkP/KJhztIus1m7klat0RpHsd7deux7YCKdv3KgYaqsUtxFqOeOsv0K8syQ1UNpQYPZ
P5WWganiQPAp2cmwVp/90/OW4HbJtyqAgwVMbmYbjp7KulNmzql2a/sEgPWMHKQn6Mt1JV46f9tt
SL4i9rIbwTgAeJeOA3AOHlhgghpfaxVZ33hX3souhfdj6LKEX8PekBSytrseLUZNhkZREbZwbyrC
FghyV96JdCedFbjVbnk7PqzWxEPpm+VWmBzoVCCTX8BPk/AfqwFLzwgJULUh1DcAjInAoFXZhtTN
gePl6blVE6juh5Cfr+Mzqvdl2CYPKZw73K+yrpmHfqqu/8J28rKEXX11cIWNqtHRYT6EWd3iAQTT
VuUnpDjE4NrkCn2snyX2Y+ezeS5yOG0KoW29GoL5MTEwNa2HxuSmhsZxHLpG9FtunJx7LhvBNrAf
HhruzjCQ9OGHkqcJagEldtu5OOjChnl/WJo4RrjFm3faO18utbbDeJXKc0v0myQaIZ2Eb1O/cR5B
zInsjqUP4Bna2922FoJgAHN08rB8aml1xmqVHvppbQy0b3Y80RZLxDgIgd10uP4J2761E/zNzgDK
aS05PkXxKVtOC0ZKssDegxW0YBWU7nDFdZW5cmHDYqeGKfHy/lq9HQlmpC44ROogrV5WvQ6/nDqD
zF9mKQVDvKiqejvP/sLXFv8bNl1BqY8a0RWs8V5NnyYfe685d0Dz1N77gJPmcBvyazryodCUoJZ0
FhYax8+74lTXvLSraJVKQDTuZY++ugN97ojqqjBTTRp4YfQWOwHLrAuMD55eZKSpr/G1NK4uWj1V
3LNadoner7cw07TwT3kpkch6uSfBYt4InLhP48b8Htxk0Yjjqa9/11va/UBQSrNeeV+wUMJrp7BC
Zi868cZq4d06jcAoebY7M3RFh3+T575fRVLJkOdxZwjBq8njPgRS5kTrDYDuMqGRzuOEybxsFVuD
BhLTnpBbV5yVBeusjIz9HcAyjhN2TjwViO8uvBC2SaX2pmYYl2oGct1fCNSP0nb94gXz/I7buZBe
IBTUO7nZJDY5571B7tIp0O0MqHmreH6fk0BTP6DrLv/MW64Ok+QhkYaE6MISwcL2jBHdfVmNtTqk
y0wE/lO/ZYdAteJsGkIdHNUmh29I+eKBUEyHWAt7exfMdVaX8j7zId7+VX6E8z2bwAxdAu1s7GP3
9zbKJevHtekRdTxSfPulU4D7LSM81CHCDCDNvEnahOuYqvdMYf6SzF1d9XN1/FbMGL0YW0EwkG6q
SgAcojJLhw1+M3Leqtb/DIAU4sr8RRXoc3XPVfNMw99ycwIAs1qoW93TaMGcZ4jwkBY3RAHGBXWX
eFww3daljIrKjSnto2xlisrnd1g0NJQyNaGhdOuF2B5B/i55wNZq6uYepFZcpOnV1Nvog14qd6Bi
DQCFJYZyR2ut1+49GkLJH4N1d8/ON7O1pgwEEApLKhVApHuvStn0Qq9yxIj651rKMiOgOIbhuOqJ
owylioEIJNi5uG7tNHcOw/LKIwX92tEMlFqOHz1ZwswQwnHXcJk+vAHY0MrW5kck7obOxkwNn9ME
UyLuTRrxe/LRCkVQxHe7pycLS9W+wYrbTG0XegocckuFeOSROy7DOs/WkeDuobCUGAWwzROB1qbg
9j7jy9EOMxof+apyWjQc0/9DKP3lGSbpxym6lGVcaSoohcKMS+bGGOtY7RL8EINLTOUn+BqgMUDU
DxbHbH+f0AJQDQOlXy9/1qnVgH9RT17GDgJk2WY6sV37skxxJ2taKBc9s0leXhpe5XhjC43Wdhw0
x8ENUjLQ3/K9AD3jfXRMsqNOj/XvlnKagENDRkEDUq8OgNtGBszwrYdibGRMD4XppTNs8BDEt6rW
/ONcfQsFrSe4s1m9n1wWjqo5pXCRenFPY7x5fw4/QhXfgX/dBXebON1SMq7LS4KbzbnKQP3wTzUA
rVHMA9x57E7OyXQXIW2fVAYM+4hTIv3bk42MrD6C1lMv4VFX+W2a4xatkmEbHCt6xbe7gsTJQzKU
sKOh8Tj8u0rDWztRpe9jjAQpHEHCGvVDpJV6fZLMZljcxKuWFccMQRisPo9xXrW6Oi2hNZHouLvV
Q2WtyuJn7q045ao4/WIspHxHGHW2B3OiLSrXYrLnbPcqwFAOBdTEy96vgM4BUmQ8Jxfe9Q0X4qFF
w4FfVPBvxpmiho8LBVhxhpiia31+ZaTl+KqCSLApYIPstvoGdfAXu5JY38J2QhRq6CFA7gDe/kvI
MTa8piqzpoEcmwt7VoFat8bTdcpG6SI45ylGmOCx3II3d2Tls50GwXE9iH0ZWY8yB2Vsv/22fVEC
mAvKIM6yxkm3MtlYpBg/Hangpq7Jq596eaElcINYjfRxrCU2E/wKYwaBgFxlZIx84svJsyB+RQLp
9oUKERq7mKiaxvFCkxH7ZW8cpuVcDB1t+Zos+cW359/XpUN8Ay8v5zgqNKaBgJIzq8XqtUBP/TF6
izHbAEUf2g7AR9O6wdFonhdaJwLKbazejs3aeoD2W+yrReAd07o7rpHK9EfDtfWoTWpw4lpF9x7F
foESNcgPIUJDX7iGTX5cHveKHGgk3hHQe4R7v+JENhIOiAkrXUTvac4IsZKv3tP14S4XtRPRe3Z+
rk67gG/vdU3omSqv2h9RK/DVqtGTnbPhdBOVMl8AtSyi1jKmPLKG3aDSRYnPgw7g7848CNBIm8Ep
hHstSuv9OcDLudfLCDh8tXQdvfEgKAaLVfpyrcns05NzQ5yBJBbRLfDWU8USxo1dY+2816UWWwaa
ZlDiB4tAgPIaN1+OKarqF8vYRo4xBkoWzE7ukQ3dzus4ZoZF90rFObl9LjB2QdFtHzH3i3dtBy1N
qY5/NN/AAjr2bWv0vZMO0uenxECclDue/HYHQPAVtSCnOLO1LN+0BC171QQ3KZ4ds1x3zph7cQl9
fDiyM+zB/Faxd7jEQOby0M4eB0benY7Ir8uraGhWQTrXTITSpNN9ugJzD645rFdIVwi5nCPVAskZ
uJeaEYBbCY4ukFW9qDFzaZ1gGPA/EcSrOla+kIysWk8QHW75x4Knf1YJRSiQZCvJfSax5SlAQTh0
FHzvM2y2960ifW/Oi0lO/RfUwBsmSC/lM4zz+24zHbHmBFyOE3F273kTtRdxJeuMC0l851Zg1OCx
NzC3nDg2RXjHhVxGGwU6nkTYZS92D0HQQcuG6UPuWoQ3KvpGBjZOy6VCxETAhZnqKH9OTc2sIJJe
RHAVlEhV05ddxULsWz5qW1CA4VmthjDvTCKAOVZtdGdkbo/kv6EUn0k3D5H76xAXfEWurUm7+Kbj
2Zwyu5ZdERCz6y/0dSMALJLb0obmDnSpn0WnKRHrLN2/CSnfbb2HFc6XO0CPwJpgtq+RP2QG1wK/
piDPzEYC+vmGdeUR4bGanjUXoID+skh5a15r8yWCj7+DVi3MduXugImuHipFYdyFZsdoB2xzFiMM
xQOl5xtSQrsBPPzAxPS5ZEFyYi+SlqqxuYqA0hbdVun5zN/YhFN0h0KVmTU4HLmqMaTWFn2jQtb4
8+CQWpoxNx0L/beqS9n7VYU6U7W48BrhffkfYGi3sVTM7EWMAZs+VkJ9zmLfRw38nwDZJBE8ZXj0
7mrZTPeF+1a7zctAq6WY3pgggrAOec4s37gVcZu3V9gd6QYfT3tN3VUGSJq+gWtJgJgoP5EZHBGA
rFLmoZK5/iR/1wgcOolYksVjY+jIBiQb+uTkwbyjyCg/X+tqAYHYsAUmH3gv37zZW9/AzW3KidVB
255nYWCE4I/g1ITBLIbrNyoOWfFvXWqqJ4AR/03tc7abtAglq4SF6Yjoo2+v/Hn7hmf1XZ9qIr63
fQUbdf8FXYRXQGj13YP/EkyoZVfCGt0t3bTZKikomsFcHOgrz4N0IM09aIpjfS70i7QJWKkZkrvI
LluroeqvX/gCSeaebN6/OND8HwTTiEaYrTMr3yUIU/hHppGt62qBYg65TsCPCW35wYQGqZPQzJmQ
8jLaS2M7nF4YY/LqVPEkolV0ND1dA6dqEpu5OMX4nUYXuf3L4L55rSDLhvWL2RrlDWbVeRxBn3Si
dSUmTV19LjLS/0YnDSlc1xljwIyzNbci0sW0ATL0MdjS7k84JU+8zFrV8OWvxM8Vt5y02j7qTriF
NS+LWBtnpODmhfv7XsgjmgzIhtoSBHHr7LFkK5eIT2gmqaji8Z6b+zRNm54AAxQOPBi+XNp9oL1e
LaABqy98tXCzL5C5uMnKMoEvmn3az8frXg9boz5vXGxcC0Yh6hJf7Wr+minKmrSg7a1TuvzTXzZa
1OHxXpqzib2xrfx2vl02FayFuoFRJyugtuExMRKExEdyteU0MI2w01aW7LjdadV8SImo5o5AKFII
Rj3FHyObWBOIybQXtS02iHuhEY1AWL9TeD2wMQ5TDPOcQhgCV0SSI613IKN21am0M12agi5eJ+f8
CpPCxuBEHnMnPwf6PsRQZJ9YgpjIVF2AEq7sIySSo4pXcwwXEVa2zxS+EnMij3mUQjLhSPPocoFd
78UtP5tennq1canKJOgUBQ0mcMXLGt9/nOxtxECWgUyE0h7JhyJaaSQCh/IzIGIY7yo2QaXE5yml
h74hkn0ou+kn6Z7goUIoF//kC+yx5wRVBbG7g9/2ESw3XiCk6J4iCpP282nBR+DsDi+6EmXk0vcc
+SoQtM+k2mCTZqlm2hW6hgJsBMGUM3cn0mWmfh3EiPTYyYns1ynAO20t2Zl83SDsrk3AAXfepUBP
rpkaOskr4kkqmwZ2nP5C5+Dur8LhEw0wKcAGJp739/+pNYoFa5QHob16i6dC55B/5rtf9nJN02BC
bzd6dzq85DOwsX5AH+TeNRVGYFzDeO6PbsPIHOR0+dBT7WeqS2V9tu3p5ven70JuKDJsVe2cQf04
thWT4fTxjireV2gJFPbAO+7HwvkKAp+RFN7veHhMTDm3Ed1kqYqHRZA6FdTbmy7BlQA8QDzlafI1
vTjPDNQDAatjjQdyZL28OfImuqe3qOMm7ExT7Ms4pjvaDsnq+7RNlreuyQP71Pxw/EiRs0/XOBh5
SGK+yBYOODfPDTxFRNqTCo5cHSz6YQwxY0ox0TYQ4inwwvpIBRHHRKOKfSvJ5/UO7u9Wq3xpLLsR
cN4/XnsZkspH6vRemU17dUvlMS5Mq3ZK4WUP3RU/vcJCXVK6e8Mhf2lH9dkIelT14d8OaTDvszIB
pOuY/2dF/EICqQjc3Tm4GnBmSRcQysKNusbvMnC6niur0bDsQxf4xt7OZA/QldHzgJyvdA0VOODm
shbwaaDr57LCDDGo/p7KSBsdk5AT+6xmP9snrpv0GiS4js3X3nDzFCgjwE9oELiMOGF/H6WFK5zD
GuBxHk0wRgcIrt75VKtk3Fiz2ssmjEjAgxEv+Dc4YibDGwiPFKxDctTMBcNAD1G1Hc1CFY6f8XcU
TkzjV/0G52pWyX2f5QIsILUh025WFa12oyHJxxvwPamv2VSJ6DV4T45NA8Enm/rkUl+siN/4sp+L
Z3mLoVRYMNvHCJGsbHyEbVgRL3mtswFkeFG6Bk1nem2uSxpcsn9TJfvy6kKzL+33zTtbe+nymGqb
+sMXDY+AulMA3yBZruLv73xYqNCVr51+RwBdc/f4mYhiVYBZj7n9sVdI6XX4n6nbhxpOTADhrbnh
8yhZQNyusPULUsS8OqvdcmBy59wxSS+5pNaPWiRmoMz+NBWY3ySEC172HKJDCvdATKBITUkM44P2
ZnCdQPiA5uEoZTCxpeIFbX+aEq9tM8MKVJGvuIj2L7fC1dAGMXAzeaQHZyz0yt2HnQhYe9rO+gih
tfKlXDwgzWIVWmDTSD+kzjpeM0tklCyrk6oUUARxx6WXxJKSF9xzMhL3M3XfVLwo6mLIWzOsodXi
WCuS/5SYPqHvx0g5PppEuBVLgPiqNaQWCqjtM0F+xnL7clTPDkowqQvuBbbgVUaN4UKQDNLZfeN+
4ND+JAdpc1bAEvKrMdRQKwssA0aBBiDKJI7SzEJ9AqtFKj3fh6xIa45gw9hx9H2uDIlZ3CuBeZbn
dpkCtH7Nj7nSKdFH0XfSmKKvT3s2V4tI0tvhyCbHsAhXfvlp6c2WvCp/n2x9IzYrRCii3TJ776RG
O9ouUZ9+naH+7fbuD36lqqKMCu0TUPH3ElMiqDxfESzNCkENCPfJIx6z3/aTz7OsWjR6EAkjzL+e
CbVqoaA6DBKQ3tyEWdH4a6Il56+JnsWATzabP/WN6z3mtpGTZ6yn8p5ySLk0ks279BKDkZO4pYXV
iT8Y9pTkavgTjUQW3czkpws8gSIkjUHfk6Hhrhign/N+qaQvTwttUdsuYPchSJUHbATNPQpgXUdW
Qkv3e2p9NDWHrsW7WWXbesd6a8yi6MhCvAmMxcPCjAUZ3deRlAZHjHlGOlky6mQzhPX0m9z0UyCk
6UHc66ar1PMttQXmPuz8NeqTFDD+5bpk31JNEf0Z26wcukd26lWq07WGCXN4gIVZ4NVbTSyI0SMV
eCYh56i5+8NIrU6bWWmuV+E7sT9HojLq8CEpCv01DdGUs+XxZ20x+StC0PVLzqMucPskDqaQs5OO
LNYxehFW50h7KWXbjQwQA/8lOSBdr7qRa9BZDa9aucKSZ2QZV05qwq3W0PHneADtaaQibQ0Vm4tK
REDU9m+rrxftAaiqqkygt2+fu/5Hv3dBFLYDbESWOPYhphv2yOTdqyhfbxx6KbwSTIdxOqESdUQN
Tu3KGuMFwjAXxMzAF6q0zT8suFxQ7uVIs/6fD6C7T6Unl07hTMl2A/RRho5plQxuA1eVum5iXZlL
oh/G9X5MgrLf82zwv8SlJvnV2njd8NpOfiQDTZxYXguuMvwzWRlEribD8KxmO+WRTUHrR9aNT7FJ
go0mkBurH4C0Qm1f12bzRli9g0vT2l90HX8VEzJIRV0zQRYzZXcJ3Q4JJGgU9vtIEoriedvGKh8N
1X73rilCkvnbSUfZL5qvdzx1MXmZpidQT3Q0ci1ypXK9QcfYQ1kowAImHzEQYbuW60ugH7SJNTSv
R8XkCd74LgvTgeGj4p7YbKCdxMHit5HLCgjBRa3sfc7UXV/7jkQPFPqTBW9+zsJ8ul+IC9pKomO4
n1JOg0J8w+FC1WM1uDczhXGo4n2viZQYpqnAC5SRjr7hacKoIV9U6SDzV0HaX3fr7plT8o0/uBAO
jqjUqUpBKAGWQHLF6DypGL+RS932bbNnmm+U83cb+jXiXCYRhy7EAf47W9dXouMB1TktY6ImWJzP
ywhuFkhjBbQiDEIsohVa492Ng9ampgGY3YJ5n3SL97LbWW3l50st7mKI8zUnyVh6g5mSEJuSl5pU
E/X8VEtOGx6owDGblIULr8uK0ijWGHKbkHIJXtozU2D/7rya+CILk2pkV056j7VGH33u6KObOE4D
Qqozc4sv0HgM2KuznqJCOqfdoeF0mSc3LCA73/cgdxB5PFBiqc2FVDXlPeKnrfc88YBkGIZUZ9G5
qQQbeFqa+Ai8eH6Qh0/xLRpcIA4iKHfqxsAIBE6khaaM2DWFDzmenvQn1uqsXNUUwbWPYoI8D5ZE
g1lsYuqcNQMkwaSOvv4bRZU59DrnHX4jSTZgp6uNV1RA9Dx0oG2OFqFflQ0Jcy02L7+JNvzM6LC7
m1bukB60Wcl5YCSNCTRsVu1XA33pJYxEu65+181k7goJD8LqNRR+lfNtKt8/Gm9a5m37Ppt48y6a
x09dsejuk710Uk98aZfI3bxgZRqNhTBn7b/uzT2Z77jr7cgc/NWQK9SDw8HV2d2bR1u6Jkpxceyc
5oSLwgk70ViWU3rmPqlvs7bp7fOHFWgp35cUS80P4KwVOaGtuuH9avvTfJHVrIky357xnWpAq9eM
pclmAlZtHel6kOtNKu3/1F9RM/qzZinyAjJzrr6XYsV5OeB95gSmIANJLr6B7JUKXExhbvwEZGfJ
6KtJKrkGLuuJa66l/XhdpU3/8usMVO0/690DBAg72ZkLCUvura/pMrbiyGidQzYQmdVJkPW7bmH4
qFIsRQLoXdND0RrhCwIDcNnw/BWu8tiLNVaM7p1xRXtiMWF6md9XbpMQLdH+CWPWwRjm/YnkCcNJ
qQhOCCCwrlLnUfAMj7QVQEfrekgPd9EoXWhD9MSRhkcndJvA2g6UwfVeLq2JUjGAPFZK6AD4NGZt
OtMpbDeVzzwrdAOS3+ZXZyroNGOsLZhojpGMHXUM4D/W9CWX6R7wYq8lwJ3TQo55hJCAjyjVVPdk
/2CxHBHVEUFnDu8DVA62Ee6Ryf4+igz7QosWtzac0gRskbVqZU1my3dC/rzWl4u7vzYWrm3qbJaI
m4eHQ5b85SZsmydsZZroA6QEDMsCHV/EiDAYGhFiSmMjmUWaIuxHcx2e5qbvhlW46cP1P3045PZ9
eXoNartKBDmZpJWLi9pWank62P+XkYlaOa6/G5iQgsEIkj+mlElfChjs+mLMBoegytZkBS7rTx/T
zXZD72L4OYTgMAGQn7gryHyZzfNJHQ9+RMda6dnRFAwty9dI7IIBFIxpci4YC6PoGHvoALMBDfkb
QfXOLGA4BYFc36jGqbgA7WRBgxVGs7PfjIA0cR/8LdSFZ9fEc/gNiJoHTK8VN0/rW4XaVDQa3k6Q
zM/l2SrrrY/28QDU6qx7E5O01a+iChjAz98+gmA7VeiyB8yL/1Mak3OQlL+jEnRIyDZm+hFaKnuS
C/eVPk+SEgt+ImDIGn/XwgYmhKJvJ+nUcmNOdbBK03x0jvgi0cErKormL8oXBfAq4I4g0gkgNQcB
UAFzFwrYGOYMlwZEceqTt2iVOAh+sUr6R5LOHo2Uk83d66yaCwwk8unRN+3LdqSXuBbZVrqZiUbv
RiryGalacfeQZ7iTUa0NTyy7p5d3z06cZIRgBHkXGy+9PTvVzrCo2FMFFt4Fd1XlR3UW/pvjKni/
w1Jrj4aV1gNApdJh4/aEU6GyRin62nUdO561oKODkcKiXXuAl25CGHTSGrP4hu0XRc2W5EXVhxDM
jIywsA6R7s/T97B8uRXpUYpe11zKXj8AK9GZs9jp6zdPkjZgZydgXTnGb71BaticuhubwQwJgxQG
hyKGmy7UU2mMcapxVHmEv3PIUH+WrvUR8PLCsrpqeermtnHaMcdutpNenlqmVohYU1C2QMupYkCk
hWH6nMVVkIpWNMn650KEPX4HfQ19kZdt5A+W3BRrIPLVXu4wL12RXjbR6Le5fQrJuBRO7w+dCI+n
wsl0s+2FhOXjKePieJxNiggiBSg0X+DP3kLPcnBPmv9pHOryTRJkVrk9Dr+3nk9ii3xLjz9p2NfH
yUtj0VzVOt0N+gAIZm3KYUuPaSVjVXlVlFuLk2PChwr2qS+xXcnYrVxeEF2qZShdoQ/MwjTZD9Bn
vXuSuuS1xeq/FuRZ9c1L7AgCFxa29TuOrcHiGnwQbjhd84reM4R3Xg4EfOp4WCcff0o5pUiS7IPJ
SeUZWCcBL43Z8hgVGsKVdveGngVP4a92UN57qZQ28m6lJ+EsNiaues74U4EG9QJkp0gADd2rf8Ui
65EJI1xGoLuBj8scs96ur0+LHvB59vi7NLEMnsgZiHWzLSXpQgV0ksibTsKMCe9wiRHAiaHRdc9r
mzdgpOxjHhi83nXaMohPwaxGTTBfYhF295fLpbV3ypJQ7Yg/myifkO8G3brtWd9TIgh3ZrnVekYq
MIQW8rBs1zvR1CYwUWZby1F/NKD3Na60wYC6OkoHqKp2MKmsyiGzzPBQtGw+/3mE5at3fY7y7e64
K1m0QrUbXrSoYyxDW3/fe1TBLtiqDJ6zLXrge5Y5wQUFj5GVdhoJrvG6/OUBAFhyAvuycAJgeRYX
3ACS4wt7IS/c/RfPCnekqOcU7g2nJob9vs0yTbDQz7YyBKOL2e8cTMcZsBua/BHWedAbCSbxHdJP
j2OSce2ZE6sr7+9kLgIhQUCJe69XBKKtOC3ASeddX9iGPbpJXw+jTXgQXzvoaiOHsAwvS0X4wMB5
9nuxaDO3I5FiN0yPmmWKmY9iF5y7oVnyEoDNs25TN29aiBn2ks3nN5o0wzARHdjIbun9zcv7Bcp3
WVOsbfq+cOexX+roFsFoA+/DvTjEHzOgyn8iatKC2D7n9lTXcnAKa0ETocY4X19i4getkMBp+wvR
+6vhtoUxa4MU087USX3PubzQvDQQfzEzAoB7zsG5GbvGIPo2/o2DdgyzJZjMKo0/65qjzvLKg0RN
JpZeDaNBx0NUrLGzspW4jlEmh7srWuZwZibhhyYuXcyt827IS59JCQW7+ixox0uYWOPx0KyuL5sS
QhNZ6QdmCPoVzsLpN/sUIUKg99R2jpzTYUPANLQGB6ZJK7XScHzVCZc9K7qTtmn4/PFuZtvweJKR
vKbcsv5Dl8LqSk0+fcYLEo0SRit56Flu0Z3DtvgfGWINRiS5IzXQ059wT36jo2ai3a9VR63a3hHm
iYV6mXSl5xnhT95Mry8pd5iFt9vTa8rHd7Rcg3F0YwOABgSGiHs+cain9vmLVv+Tr0zFROeAlboB
qSoOxx5i6GV2GmeC5Lkyxdlu19Q83Q81wTEj9GTCL9KZXgOoxDtQ9APPvgJZM8c0XeUMRWhxFgR6
IC0P387qgKXi9b4p49I/ENjcYiIyBsejq+EZMvOoHySUB2ZSwB2YF8BYfafoAQW7vRVe/l/PFNC+
hXSi69y1O9NgezzC5wBj5m7MNYdED2tHkFnK3IVfmxXZVaddRcon2EOr+WuQwCto2GalRWo+9JRD
OvxMTe1Na6O2qoka3ymPKb22W3i2rq1pkmn7UPtUMEqZCBehjSiKzRhjU6lYnWv0hfjgopyQ5Nlv
JYdNBUnObXAjAZjN1X/YQEfJ+ZOIOf1apmpSz/NPXsvScWcTJhzpHc3fVzqagjlJduB63nUJSCvX
DiajNfizCTfxEINUsSpMoMSsijIlQDuml6c2llzBqB9OIAzasZtFPqBrVkdzOPlk7XZbP/1Tr2P8
1b5O/DoDQPYUxSnDJeOAFKB0QVEa9U3HbaVMt0xaV6jLh48ISybAH/yqxCrojgYP7mjUGZIkv/H0
XsOfouSUjr5sQPp8x0lcXOfjVCBtuklUry7Fb8bkHuioeJUYcNGGwOB5I1TZFArLLb/ZNkDCmU+1
SfQnnGQbv9Ii1dAmM6r7E5AiO8o7+Uaf2w3RPyZkih+PVxGcfmU3QM13ramOj4ZzcSzKbpKOik2k
Mh8ILmY+ZVbjALgIE4sUyUG52vrVF0IXHGLyvSMW70nue52iMIAUlOVDtjt0VyQDTyNPLi0xqNMU
FPnvGWDS0kPMxTUOa5gJ9OE+u4TZXTt7GO3mL5KOKKOnKFUyjlYsx2YtBSNXBNjGd5+IHzbO1Baq
iOfCNLafVvl/NwgKE6u2HHgM7o9N4v3UZXOYimjlbeT+5zxy/6TdvDjOnVZxznerXIGMusqTRbM5
XHWLRDXeP84vmpjG7MHPRohI+a8PjMXGaJhOO7FLi4O763Hu5nwYtr1pW6HtzD5sUlMF9Vn7A4kD
cBixsEUPPPn/7mKz/VmWXPpfsIGlT/RbgQf+5NWQ35J38lqXm0it9xpJ0exr7XkvMjuefB1iye7R
AGr0Vhjw8hqd0XqAiNTUTGSvR/0X3pZniV7se8hpQp7BNfDDo5knV6hlQSIS7XtKvKpi81EyWLf0
/xyoCk+o/8mzNLXdR4r0V/suJoyx1ua075NxrwIUEribHVaqr3+Z/bYae+ZnIjqUf+VhsclaCRTK
1EenTQz+MeD6jDI0r6FDRCrCPDaOeNNuYD85Gol6W9QCEIqIk5idHuWvoug+A7gvXV7xVW92KwWx
bnpZkxqZPX0G2VIgb2pOWOMhV0Beu0ZsMtc8/U5XvhBp6uHkbs+zLlF59DOdnFfxXIeKTzeDrmzW
J2o4RCnxJo7KlhTxWP8rz+uMj9cnp3SM2PBwhc/wCSXcl8KrBx2xxiQaFnA+QaOW8ciQM5B2YrVV
lwaDqLeMW0ibTm7uZp9z/QbdHWzIgoyBOOas8gu4wfHdowaTHMDwWLSwV9p0L3ajmwEj5LE5FvqI
NjuOZEy0zDazvt17NcQNKTYbQG8FNSvT0BGJMHbm2MN2q9dWCbQjZS03CjnQP7Uufo9wU9Pb32mh
1lC9He9v5ncTxfQYg6IdydfdJ6//ljXDm7InQZ/gEZfLrjt91xY8/RksQqckMKhygzfMLSmCtMdX
Zfac++aKyf+U5NFmqdlUSfoTOTUQDqLBo3VhDs4aa6JQgVL9KUhrrU0ZXaNLUNEJ54/zNV0EscFm
PUXLep9EV/EVLhDvOqqEuRV3sW3BHAXe2y7WrhnyWI+OAzY3zgwA/2I3accyJQyfl+9NdWZoh/vF
10beCx7iuHtGTSXvjv5fZEYTj6og/9+ZcMfyYc3Yz+biTz+YB7dr9e1La7oiUK/qsn23bNG+fxse
DLMSwGhcaebD4Zl7vSrKju9MxzWUW+oisRxbYolTsZKn0z8VMv+uVS40Hl/G9Y9AhM6XPFcRFKpS
/BDHmGpToZFBSsVYen4VJScXDXFu/IrNAaZolzu34Vbx2S3fKOmTJjthyCT6dndh73AYjjjdAi1V
m+C6prO2sT+n5xARzRNVdWKPOz1C0aCgjGIQNRwqDwjxhHiH3fHaGzaLCNO3XXUF39jUYAhtOUfq
whr4GR7CdJuRAZWNRnxBGcKjU2rpNJvpq+oXvhD/dWMoluy7lkEr967WNPgcjhi+XpXOVwqZHQTj
sdrR37kemQVgTyhTLsGBjTLlw+KfvLPNMWCTAR3xryd5TjWf1dDuXFCWmxoTw331vTxJ73bM0yEj
HXyxyiVys9c86oJ8a/d4TysfozeoydISSNzu5b1/vZqZlFrdDZfUKKb5yYO9RTQ/jc5OGaaWqNLc
gWRNbF2467FnEb8VVVlzAen7uOrMIkF/114yT3JgYj4mw3GUk3RiwR/f+p9XpwVyEUYSctZ/mrBx
uXrgGxU90pxU1geD0zYBZ8gYysUfsCESEZoWxNrKDF5Wfcnp6KAsA0pULlhE3uqKzH+mKvEAe7SV
wlPEb9J4mU0PSpIaoxIoq9/4PhNVmT23vj+8BqGz6UVsDk+hujnT1chF21eqV+IHG+u6E+eHyqsD
P8YzLF364SLa7lOfO95Z+DtQyMYAzGmh4xsPllKNIRRdH6isTt/6kenCzVI6b5PlV8XB+oeKihcu
ElzhH7bBZYBRvY7qoEPF/umd0Cz0OBiw1CD7MXIB7MyFcn/OA5j9QqpYW0T2NAuxuX4NgAl0MlJX
vdkhTGAWprvEG7LF3+fac0w1ywm3Nm6wbSnbdG4z2Z8BMRK6azHP3ehOth+LeUscnxFZ2NKniAKW
sBGmGgEHlIXoIP8ro0b3SHidkwOxTDoK14CP3CMrZnoWn5HXa2dUS+BIM3aRAPiUwjC0XHKCpcFb
bg4k0COx8jAIZseHvtJcnEiveBlRtT80vbxnJpNzk2IH5qAWPtdqh9Pd4iKqA4+eeBT3ZFpJENmZ
+sCnj60l0eIepo0EweGN4R+y21K2RGvFNV8tcuShSj24LBvu+VoU/wLtwh5aK0r95C8PhQhCFlHH
sHbzezW41pxpvrmhSZBtRraH+lmuqXop8nU15eXUXjN0X4/OrbBUpdUg1KKnbV8OwAj2C0VGVX0O
xLOdTpeA1mQ6qwMfmBseRn6SqGPSceh0Hvt+vsSnflHNBbml4DQ1lQyF9j/SaNPb/kPuc7kkoP6Q
SXgkI8JyCLoMahR0JIfsS52XEqb1Yvd5vh37/wDNaWpgof8nc2aEWaItgF/t0t9h5tVjJL0SULOd
S/x3GF3kXK4W3VBzT5AvLn31EHdzeMyaop5Aa5h+8pGIlvbC/v6+Was68MPImOY9Kbikr1ixkUCe
4QDAVqwIHeHuvoWmomeQF76QYAtNt7RXMNjU/lBX1EEEdozxdgOaJWg5fCKKSY2gwtJZXlZYbmpJ
ArwNOCswNtn+AeAOvk99NhQ7Q1iKvgUtpz+qB5Smog9SKBiROWG2+LI36a4GUC5S9jIm/lFC2DOK
a+rmLTEvk5lfNXu8e7VAYkqRQsiZuIZEWpH6p0undpHxjM3ylkvTnGi4O1Pw5pGeTURJdw+jv7/z
dDiI4PWQpFA1S3v/759Ugz0LpAXrAzewdG3IqEaBqGDi1jP1/8J3Y4J/3uvsg9PGetZYyPcYmf5M
4/9KbVYBIknmQOd6GpU3lMdwDsWzpYwFT6MkC+3d9DiCvxfoTxWE0ClXFfDDOc2cbDzxBUEX5D8t
2A1gRw6tFcjKzvudBpJTcyzrhkL5/GvH5fAolyU2frCtoC+Ui4FU5k5LFJN/npZTKasi1AE0tibk
5Ms0L6m5UL/6WN8a8KDipzGIbDgLcMdZ/kQTntXOCJJT0CqhUT/fbCqL3Q5JHd6UNLzujFYIIaUd
2i87yBTrQfqUiN4o++u8I4i2gu7977rAK6vaJXfb5+AvjNR+4yuZrqYFFcLrqGz09G3L53ArqET8
bW9skbcV+BoIM112sE4LMlBFtq+A+8RktG4bBt98zxAv9x6S9S4BDU0bWHFXDcQh+Ewq/xW+I6SD
2zMRMi5cibaxzOhbitNWqLzXagq33nWQJSCmjEfLh8VPFASle0BtdFeeaQ6gTyumxXP4af6uEBfS
nHHEK6E4YB6eocHs2jlnFioZkeebp3rEfIRljrRn0V6LV0AeiSRQO+xZZek/vO6rdClILobMqq0A
Szz0OIhx+GkDmFYwVKXGa3dKevXP0TLNmaZCYqCNnvUxeKwggRr2eLyRqRkdMYORTzwtxLhWj8CG
YOpGb9TEUIKkrRM5I1Fu/9XW4SVI721GUq4Ez8MkEfwpKSX2M38kOwsLzDzG/BIaqdYh069oAtBX
Cbf0Ev/t6mffMZMQlUAxc4nbUeS07ItR5n9t/ZnqAZoSVZ63/9HqrlFI39U3qYNjCuUTF4y+OaWa
RY/iciaf6sOLGeip1lK5LGRuBfFphiphrqMT1VR4Imtd6NLZeDieSyRh5AEdDTeXHhqH1PaLh3id
nbODYxky88zQeuTbXDgE3ONcV51zQNi5pjFgsnvblywasj/Sv8p5a6F9+24C6IjT9dX1Zh9k9YRM
eqM6nX+HKrwpb9aP/+3fZdtQeb9HvSjWczXFCddpfRoKWm+O300+bupsJzx3X2wQvkxuC283y/9F
/Jam/IvkG9u9iSTTHSJVN4KHVaIY1LRjqmNbEd3RG93/giZQQ9SApErZSy7WfrmzfTGM4WTV3nuG
rSSD0+WAidfbs41yr3YqeUWqT5If2MM+MtBqi/vMPthHU+YZz3sFZVx1FY+/0GHXofEHLY1A3UpO
LDW+JlC6vS16QB5CK0xl+ifrM1AbZ1N3T08SFTnNkT+ujyAOS6E4AfMDw8MmGyN9ar/c44JvG+c6
H+ULr/Ld3/Lt8iDEi64ZmZrEFUlOp8v+FqmNvyNgp+x/EYv4kJzKP0UY1GUNqfI5cdSSeGwbvxxs
kaGvd5LMTG/K1+wDobLQ8sWr5+Q3khkT+DEdSqWSfoRkmlWePHVEp5m9gheW4S7x7br+tabNPxuA
0dSLF7xtyRs+vdvw04IGbeGZKAjZywQeZo74AqQbdxGlZZrBFs6Ltqd8rg8d0B9k5k4c+42OXIvo
3VwpUTx1C940cf7eupV9HbbiL6zl1LC6s/3R5l9iHXeazw/qNl8/LDYSoSrzzYnSS7sv0gspsTDT
1M+LRtp6C1rzoC+FbqJDATMYkghetE6n3fKootjrb51jsZvJ+LaF6PdvCPLvWaHERnaP/oNEHIjO
3gr7ZN02Tc8x2TB7mYJZPr21eS1SzneXHnXXUuF1gu5HsHRV0JIhPbb1VfKu7T+zToHecoM+MiGg
zdq3r1uuxgiqao/Rl8br8vCOxE2Nv2xMFbkhRG9Wzm3Q6xRwawpqxSIlgMNipf4SHdFUPHK2JJOD
3eq7H5c9+jxmHd0K4u7YZK5F0X+3A1QJVfj2JXOli/i/tUPEzKcK7i9Fj3g5Yooi6Z4tDCi835X1
o4+17V4sGx1TbFr1fQ8qSLmkUPlFnT4ZeNLuKv+mVlhrxRXKzays+IeceiEed0ugxpCpI7LFz1qz
mlfsqROWWanFdK2ZMxLApG6chNvKW9H4kVL5lJiWrNnKYMFYTn1LkmLWq/E688m3ESO2M4105xv3
0sCbOyygugy+uSFojI7cRuEzq7oI0woYCZVXIHBsFX/Tpl1R8lQhX5NrdR9e5C/fl2yEfdHakCdq
937WfrGBlC1ZPY58yuEBKvTS4m4otdmitfOgZMuV+BPlO77n1lDCF+4u+oPFDOPhc2tLPhZHVwgs
z6ytCZhYCkvt5lA4iPjDd4mRTSCrfUeK07h7/hr3RUubAnlhevUm6fwI11oINXII7ZBnsr2avlsN
79qbMkYFnyhUQT8e3vagw6HvisME/NsRd9cmMFodLmxwVu3Xr99snQdSZF4EjkZjTOG0iCHwaz5r
EDiM+0EsChhea011s76LWfj/oqDOkqg7qT0ZNm8jgpk0Fz8KQMPmSne4vclL87hZB4xGeXWi3HpA
XglIq0Ch8givIf/iCAw8OjDVqYvPlK5w7P3YRk3sDSjrw19SyB/T2q+J4k0jnh/NyF1PFDwxg5mw
vSIlJBOB3m8AajNTo1Gso+sXLGDJH5kNCLubKJyjRd080pr6qOzYMF9msX4/DFgcacxzJltn7I10
256rja5EnqeJ+ogQhh0/Y6YhMKqsYyNNExaWOkKKYgTPtOnQwocsa+NHsjwePNmNxcX2bSUa8vKH
dyg3cv1U62wa89X73z5HKO2GnZtgI8e1ygCiOyQmWhDuhr3gE88onqzllyg74iNiiv8BhN2cxoDa
kaG/GUsCB7bjoSuB9EEN3FBAoaslvA7yznVinS4fo+AnQ6QhqJX3nkJh0Ppw6IV3YZUkEVMIFPWs
EiQ+WNQUi+9zk08sDXZS/bLGw6l9mfb+4wJIDDh598fg+IkVmGGYXEDF24ViTIdUUsv5Djg8M3jq
PrGCOZJ/YzomjbVU78o/I7Ceu1AoIGxxxYgseb0YRHWyW/cA2EmU/QS+MjNy6ZblKFz+BWUlWyZj
4yeFrjpqLjzmXpds/LraqkgJigXVdK20mY1YNSeupZOlDsIRg+/GyP0t+Ysgk39PPzjcdteFawGP
+KmulS8FxfPsUVlNZJuYRiyp1hg0iEAa2ejHG/AiVQar4jUC4v96PMdyPz7uErB/VhuB/EjvO5Pi
UNF2SjQCbjs10ndzWKkVnHld/diGMuRrowDWgRZVCttPlgNlI//1XwPKYJEl3Scb6xQaKcUbz7r2
AAkI2Q9iKcmTFTBvfHhCHf1sbHCPGxTZ6QFmoM5LG247LeND3gjsyoE4cNbAVWiK9pHtFPYX3OKV
IzKSWuuDsqfOPKPVdBxynBweDAzdzs607NmJTX8WDmIaMdreUyjobPn8ZN9vX4Zxs+En3FX4sGMa
1vuANMqtJPCilEnvby8NwFxksecv4ouYl6ob7Mc8PXTiYMvIDD9DI1QGMlBYtYW57VM0kKItiuJO
aS4Y/FgTesvTd9UzEeCbjtferfKTjwaSOAQehVmIvW8WifwLyC6seTFaDscZYoh1qiiKq1tXToqL
kS6B1i8UlcMPqpxmicJtjbeAMUQUIv9OheUrTwyyoupr9gxwmaMY5HQRFSPrR33QBBspu22qOfoS
xTuGbGdnkSV4gjHpQ0m+MUDmTgmSvRZeaPmyEsfvMeW+5da6Mzfs/qyECoX8mDsKSIsbjmv2iO3s
6wHBVmzuyiuufr7u5NQ3kPg6GsbBQgeIjOvJ9V1Af7TKBiTS+/SgwWTEkp8CyT6tJeJPKYL3uIYt
HvOVmMn8/J+vkxSC838wEBUCt8O0n7Qq3KJIjTqTKy5BQHzcxG2EHnu33ZZ4JleUjMpttTtn0qOz
2H69zluPRWdzq3P763t+7MwrVhehfdH4Sccon3P2jIqfrb/S2zoEf4ZdqZ5o2hNzzpzUdPepkh/Y
9lR+6e8vnp2/PvJZXFGqc6gYhdwwNkYQKdmzyF3hC7cPiCYmZW5b8RLSUAyi14Vp3YSQx25TFRBa
mbuptI6nG+U0MWfKIh9T8WMtGWktMMUC5Kn7X5HNDYVzUgPEbMsN4OcpXG9DAoQKhzS6oEdbBIcc
hk+4tZcioF0+Y1u9w0V8IV9abuhVhYkOP5lVhBeGbaFaoo03xj06knxiVsymU1MZ9spLJHHMXRW8
nA2UjyEE0mqtjbJMDzNzp/4gIsWtLn9BqUsqDQ4vslllU1etyQhOjAomCtvX3GEUd1jc3UEFjJKg
fxCCSYesa50FZKz7+4eIHZC5LbaEmzmd4fffgcPituKGKqrPpKq9VTGdGi+DuHITyo7kc7zgpPRm
iVuOQxRw39o25WdftDVd0xyx3TfkZAAXxNhwVlbQoO1T3EOx02dKxfGyCnDG1+6UxjryBUpkr+yg
EEB8A5uWni7zIUqzCQOleX5upSPG0zHDHnjygCjeH5n/VPnNv/xzSns0SaVsyCl3oBvfqN5hxtDQ
j/fPxUCw0u3r+N75ysamD1Kzk3M5MpTmQdLutEOFgRIi7zvFFGULnsL7RkDWzgyE7YcmBILxrYiB
UQWtAFI4ZjRCAJe17oTxOAhKVvFmoA/Eest5pGmV1crn4vwBNsPEvMtuu407IhB1KpBPhrDdBnx3
qJ+DkVTZuzcgyAZkyLAtfYVrSAHzdceDHbkER8Vmh5D78eNNo4KLPPGThatmvoYN69a+JyqUYh7n
chZUncA79KFTTP3MsHgXN8rH3S7bCgQKvVe2S5DUAetC9q84YHCEnXsLCxL5tnIfkqDObAOD3+sR
3YcFgaITXyuOBnPGhzdzccCFOjt2douAvCqU/MagQn+WgoLvwEButEWUHdgwOfsK+QrEAaQ/1F+q
ErDoCuBliqMBjGEwHNI0vJT7qBaMT2GlJd3jU+bSJUPihlOIxYY7yiLc1+U/iSJ+PPh+8BoFtf5g
ZNaP1MUt6v/tTzIQ5RYfUkW13kccmI8QCuUUA2HLB4dAW9gOC1U3E4gBFcAO2zGtrV2x2ft/lQAd
N0C9Sx3KByAOa2tGPvqaS6i0vKNAfI76AFjvPU9O90SQJMQvq61dXveWh7eHET6MjO130OuST5PH
U2POteJr5A7VwxPU0zuA+f8+9pPZmYpCK/VLOwamUa6nqkderYaydnQ8bsSBND2Q03xmZN5N+6hx
4JpyEJxWpLMEajQM07Xc4jhfHg4CUP35T9Z6nZWLktKAEmxA+NaUjCRJnjTT2URiVZ5aZryWAbjh
d4XbQzQVvZQcFA+gdVdP4AOsnHdjdbhAbVFWKQLG17hnzCWRlvvPBZZnjlVdGUWl+A0GfViO9nOJ
InCqtCMcC9jVitpgz1qvGcCf7dPI3Nnuy3ccevYUtoo25zblS9OKreh8It04JjVygmwPW7iGkJgy
Vk2OiBwU3kst5TBAU1GvhmPQPE3bvAD9QMqtlYryQ2g6pMVXWwxUvu7n7Ho2Jqoqv04jDFPi8iC+
hIiWi07NduEojIQBd4ffokUOcWEYruwNjTNCCvZZ//0qix6Lv3bfg4IUbWwfXbcvvh0RKndxbaxD
BAU4VOR+p1jLSLaZTuDg1KKxjwQQDMhzA8J0Roizr/KXj9n30kT7V6FmR3GnHqILl09VsEsy4upv
n0oZ7lwHd5ul4kmD1QJNwIJY0yl0SNLdzD3v7tlFRs9oB5PNHwRS6dNcrOLCFmlRSkkDEEJAypPv
yDzXGnCUpXQRPW54W1JxyGmqUKoH7umzQsMUmOyM6v8eD2ixCZHwrIy8QGQFXTbUi8gkoHNw3amt
OChhVCrb2Ba0EhYKOUtgfiRsRRkKlaPedk/0H42yMCq+4Mvpur1to2BisaCTIWZxNdkIb/diwvXw
05TxAMEyEQoPywvTgzhb+cuaxeGgoZTXHS97grpXdjfJk1sIEsmRcTpyAZm8rCmFouFH4hOrYuzC
3xOOOWbz0ERzkf9RsTGJmYM2e/avq0ivjGxAAsmzhQ9sGGcpmBhnojkTYksZosWfRICCncq7V/eM
Ch/2cYcMBshXG/WgAAXN3EwT9VHs2oh5i29LlzWwHjAxxH0N2UKlbiGNZwRRi3JkoHaLRsvzrmgW
Xh7BHi7R63+ntvjCssqc3TJWYlM/j8tNWmFr2148igJy/LpKAobZQCbzsHAOTe8fjAcsPIL12TaV
yKb9RCjrBoexo2BFqRbE8Y/KFqxwqetYEMq8VNHqJ8FLMduVRssqDQTMXXlXBuFOb1kKl7WE6jcJ
nxwSDhaAy5vSjzWa/Vo9TNHMENRyYizicNDzQ5Pji/AJIPc8LsV43+uUgXaak6r0Xl8yx3UQ3DnO
jSwIKgqBboBrdbwM7urE+R+tE4vYymW0HcO26aTG+DPBta3f1PQBnfbK19H5m4wX5r0Z7aeGsrKW
+i+MN5m5nmQn0UJTwrnnAoKAUMO0aXbnyRDjP8ZN3+m197uMyWMNCMPacgsk+VSTx3h9Xct4m5dj
KGgLvDFlvm6EdyOwgPgGkePvqljMOlyN42c7XVIusGFYLJpTk0X8IGAwn+g/hf/CHtBOSzy4LJ38
Rf3uzCbHZXgSoU/htbZp76Gp8yGI0BcugxPtRSoyqIYmdFKz10jb0FY+OvBTBFljhHvFHP7xECo6
zaa2o0U+b4+mywJDy+vuQVdQtV4ic6C+U1ekhHqzyjpRTM40OE4tY7hx1/r/81nAz5PuzJXZqsSk
z76f5gWzmN1Alz5dskTSX4G6r+Ai9iguzRWCI3vQO7jWN2tw76gcyBwZYU71Xc6XuF3rrINDKWoP
kmzBJ5xfwPgtAjSWCbXFOL6oU6UFe6JTgQJjezPLYesQuqLQAN+SZZSkU4d/xVKWc75x/EiY/y0R
QO8yiW3QYw4kgUhPpIKZyHv2WkAwb1kJ9Wr3WaxJfU1qSuG+euokuU12FWHzf4svZW2Rd5aWcncs
K9VYz2F9cMJXHarZerWCFNNXZrsnCfdxWmqWmtSXGD9C49flN/RGkf4rinCBtgCU1af9K8Ldv+7u
DbYv52umXNDtca9uW2PnVDkcT5RtT6e3pDP5AROF3G9Za2JhsLuATrD0xPBxJ25EaQvmCZhSMdz1
cH2S+0PT8FyDYMXwRWOvY/xEby5rhZDi7NEJBUGjVNOCsSkH6KIsipsYn8fOnYTOY6p9FBEoURQO
jNx0KTdDkrkVu51y8wKN6RQUt7r6OAYGnXzLDcql4crGBgvwkHFX+RUmfETZrjTvwCBPE+krWW7r
KhCBe51gFxJyYTp3qvEM1VEhlgrCZ81XlVLjXbwjLVEDX5KprBE2YfyM1Z/jBSoGBRIYi1jGb2+i
DQ8iwa4WJWEN1QOuHNZdM7HCeCd0wR/JPpVBvQ9vmvFb/caDH5P0LmAFjzRCbZQMEVMYAACMKXaR
mgI+LwD8S1t7DKaZExnKBpoCtySQCNeTiA/7kaiEHUJD2yRN0PklVtxWYsQKhl8PQxTbMEDqePhH
Q4nzI22O0y8zl7udx8R+mQA9vMVBuX+BYJrB7PUQ+oHpeyDczm4K1+BAHjbpd6NFGYgEKyPj6NA9
BVoLul+05zMXJsFa3LOc4lp194UF1LC506BkKr/4SRsmr8V1ZVtl+CpZ6XLiDoT3olVHhA+QpvZ2
ybYShED0NqXFi/0A4qWhsK6j4y/ozrLuKYVXw9egJFp5gCxb8pvk+x3E0gaysl8RJhHkXLRaaF+b
lThKl3uyHpQ3NJKxXpq0EEN2SUgV4k038zvCyKBgFvnvzRSzto9jQEgj2B4QyPARXICP4/ljWCgK
JhtKYEUnwDSm/gURFkDOJbahz13TQy26dyTMk4G+o+8Wf71C8iXCodMHebSSJk+e1/qI/wHqCigC
c1Jni42zwGxroKYDiQLHKQD1Bg0WjWfLVO95dnPvUMZUfcweH04nAnWK/wvqmt0tjUJ6hv6a2SLT
cY3UvBtH1aAwxwWY5YTDkcSVwHs3B8Cd9LImAuiltKI+DYELysA9tR9u4qYpDNpwIL3T2jVb/AQr
BlI4R6IJnkSxfqReCSCvQmHkMEmjl33aoBypPScSFJw7XdXqT2wuTKPeGHaNUTzLob3fGOz0gcQd
IjDyy9Di6HdyjuXo9VEMg51LzpXx+SjVhZqihxa7/mbjj/OcfZ1fav9TR7S+qj96dft8cxZ8XGf4
eQODbReLngd6YGCw08YRnw5OdL+gmuivP4RMRwA1HlbsKq7obUahtPzPBh1ITAmZ6jEyixg3y5U0
hGYsETo9Jm40Cf08h5wRoxVcRuvtn4snEtNTNxHkLu2FyK9Ypd4uMwz47cFQsEBOA2rfkuEQ0BiH
owVXKNfyjykSrxO0yvI8SsXne5j1dVS4PKlJOvxMMX7KksnN4A1UEBufCXHNhHhyFaFJTSrdoUnh
jXkTur4fzNoIalxdWOJgnhrxIxj0rSRfnF3zrog0WgGdvS/VsiTNTYmtUY2wUuqnQhcZePoNIFgU
5wo6g/RmbIZjoHwbOURTAcrWDrcApnUt6iiMgGvXZ1GrNTAhM7b/BotEAjQxYI0juqpIPF7o+Dky
bgZlAjLmEuY3twtTNQ19VVOf0SKZbQ7xcssod7TqJslrjeakxARo+XrCJPYDWcmq29DA+oU5fZgX
MiOWHyK8Bxfp2+VqzFhiU/c73FqF8HF/PEBB76PAEZrfKjlqnRcLxIBWb8tr5UYG7zaEh0TMDqI4
a+wbjfmKq/ckqWrKmStH3S4cSzmi/lB45sa+bet94XZV19mk40S9f+a0AKQtBBgfo8FZR1mjkzJb
wVpaFJ8MLuzGGtbgX8Qju967C0o1lCPV+EMkAcmhIfxilzHpDtRGbau9rRqHf/rTh03ynstV10Tm
LSHpKaIMuSZtwoDe1jp3qh2O5pgvOSoTnKNy7bkUkiw0thaZVJk82Hh9i8KPaV6ubYirU3O9OlEM
aMxD44xdNbCdxKq4+S1rax7mxowW49KKeCSkTZhmyGAZNHldbC80df93+McX90Q1DfuaCq8WtEwu
9DY0pgbnoaOveI22YZOQnMazpYHv+N2zXS71E9ViVwzB6AK3OmpcMx99ljO1sZEtQ4+BCvZSHNs+
oZ4CKjKx/A96KkTmzGUUe0Da4+5dhJfEeKif16oDM5WW1m5ARPKLUfKvKgtsDscqpf126xQ1ZajQ
eJImOvSl/LE0HlRJFhw8LZPNIslQAEUrgZwCqWjqZPpJuYgiJgS8tvUGdSjLGfzWzf6nA35OfDU1
BSIvXGVwLxDHZ0IlpbC8EzVqzkUPtub9GjlPyeemS9YJ9VRt0A2vHyt7nY0VHy3uOAogrZONFjXI
jQzWfrc9jxYnYGglqQVS5CMA8u5QQErLcd+boU6tDHyXzM3AfHOE9goUQw5anSuuZsafGwPSBad5
jIbVRZe9UBGRsy7JgLasVn/Cl0uhiTpJ9opbevJeq/bdcLvB0xBlXqpfKJrZqHhWIhNH8SxntyIL
6796cEwySXHA4Iq6g+1+Ztgzt32daeWMLI7QjMJfNvCSkiPx6JfgMLmPA/Tn3IIvl7wxRtGSD1OY
CB/7V3Nge9lxNlk8Avi0shWFQM4+hNRIemZVCXYuvxDEOreSaPYzEc0vsOH2FxQORRS+3zLgQcn2
PQuiaDWK5WIkxVas3hRSKphYq0Ytx9edOdPIEFU6q8vGpyw2UKJsnBW4xfGc49kT/R1vENKveOdD
KOCQBWRz/dRqDlHtIa6hMXRN7w++XGkQ/0SfYNx6SbJWHDnC3I0wu1s+p0Yw9YjIHoZ6na8H1ORK
KEqs2JOvkim/9enfxeSPS0uHlSEXDrjH9jjFrKEjPVSRFRSJWk3wnyWCiyv2Xpk5Xyqb/LblkVbD
XhLOYonrpz9NZ6RonSNFrON0l0qDzckfftD0mfaM7P50+zWHZK20yVP7XXtstLgTz2tWlSfW5t2h
8xcD8kNctkc+NqklFNO3CYy/9jZKk2oyslAkWNKiyiXEdmSGpaD7GaR4ydETFZpwgCIsPK9BW0qJ
K7V2uX8BZqsneSmcyRZz3AO9gRsCZaSlK9V0DzRg3eyKSbg7oJQ/DEMtentLTrpP/Ol1M9JotfP1
tapbKz72kQGGt5/2Mk7leMillXJpWqSihPcy6fZZiABULGWWHbSP0/I4RtKCvM0ymWAgVaUGMqtg
5XLtKIZkhBYAbth7w7UbQNkSaPtWFnYeHuPFhLRkvsePI6wBe2gPuJgeZ+/wlirovscjg9SwERXw
0x6eMqqCuAc+NYgrjLbup+huHoeogAvgoWZ1evWvLO2HuiO4HH4imIYenjuq6xWGqg9Bv1EX9h8L
AbGAkxIYORWt/uTtXEagRZVp6jbTFHM5HTsMWn6NI2O783LWei4GriBcxdWQTtM2Bq/CxK3jZL+M
5umxj6LYK3S86lc3J+FoWvgN5MTF/WBwciKDpjdbotjiVoWEieYabA80KFT2/izA/qe4Wa7BYdE5
F8reyavVA0Wj3N8r/xDuFjzNE68f2re1xmuWbP5WiHkxzzbZKlizT01RSgAbjNawNI9MaTIqcwXT
HD39Wf0p3SFMy6tsVuarls09saiYjIlGReuwGdHUv5HOnoUcL7Dyqfmsne2Ls69tlFqzA7s78PvA
h/M6LTDqmno4HAPTq9tDRzS0MKuqKCLKZQCDp8aAMzI2Bzge7xaI1PXq8N/6Q1OgCsYIWfBAi6TL
Y8LDUNfMiicABErtLhtIhaYnRBupuScEAFN1XOWUobZtAwktPpJUQaZ9d0oLZDX9+hgWo2bywDIQ
BaOlcdcSmMgSPEFEyd+hQdx3l+el6sF6Fm5+fzTT5RtuiRX4XrOoG0We89SKSTSvPlNu6ZP64vCE
lFZOG8h6yx9RYYkqzUiAmUFr2Wn3LzMYYvF3G00JuaZVe16ekQWgxTtxyYKjFMPw7IMKT7CLlpp8
njiVUdNX6z8VKetFKAP6B+cgN1tVpMsh2HrY2aT/vYe5WkkSbHUAtTtyx9HkYuO5G8jQpl0hlqQa
NEJ6SUjEIpVRbvR/SotvYbot9Xb8/BL4TvmraArsae0ph6RO0Huey9cv8hcvDSJroTgqNaJb4g0I
2n8XWf1ZraUxKGXfCmjKmBlFakIwtKr42862aKrS/mKpUTgI9LAqObglHHwgg8jbvwmVi9geRLgo
feCY7V/OWWSFGo6eGEGz6c8LYOkzQppp913Ch3tpvTOAe2BXep39VmhvrenmONLB1F6IePclOle+
M8edlthiw7lSxRW2cDaHArACAF8ybzCJrdEssaDkydqGCF3/harTVLU4elLBLxdPZnuhTynxn4ZG
zQw5CMokMapdLE9luRv/cPxJlASTp7gN+MCl/RQTKbADLC1om4gpP2ok+80qltTtolbRnOFLpRRM
8sTMkbg/iq3IUl5o2QD1fetTYUvx0pukRSyBBc0lFHukOjAVKBXZIFm4vh5Wue0G5kWJLGmryFsF
nD0xgtOM7nfBBVTQCQlYAnxMkV/lt8eLxWXDTLS2Ou5zVEKPORq023Kxr60ApsoubqNVwe6ywPry
BZ8fkyKAkIS1/jt030GAmrHVJ+qqzMvqeU/vFNk7VZTgQAZRsJ05j5WAXpQnkLKGZ/24/LmpEU/2
MFEzrC2dfCPDTHxNL3ar+wSN00mfhaahf4FkLQPumX+Oaee03wYNUspP7bWWZ0L/Tdc6EkzQQCB5
CXSDXTGitxuJsFxJMJJnnJvyXtazjlt/xhTfvrRz6rPQ9u5T33IbB3UhsB5eHM5DJbNdHaVKyxuA
ABiApVDHB5eHNxr4wQol9B7ofx4Kc43jPQ9QOehAOF/wog9RaHolG3YpOUJg8bZtCJgETazn2c10
ZR2sx/NvbdMcCcmmUSuAxvywlCbf9tHpr8qPnpFPllUMRohfjoUMXcJFsFmKUyGl5zTxwWeyAXOn
S8HFBv46rvcoE4FJSJHpjSp+iJTeorot8arHNUiNyb4YIOcFzbZ3yAT9z3iC3z8ZLu1iLAVfEXJL
SrGJKbUB/6iUR/t2ojJlhO6dEDoTRCG5hH9pWmqTdGtBQ9QPX9K6EPlZpECrWGlxwOBFphIMoCxf
6sFNsHlFqCkf7cDAZTRspz9B/ckcJw0nFdIvFxqvipdMpGgVIIhUfE/oSo1ScHhK1Jf3VghrrPBf
DNtFtDKr94OnTNvWJRU/5/X2tdiTSHa84yf8RsB9kx2XQyeKFVMmaWzjKr4hi+PeZnc5Y1QNwaOH
6RhEjO9w7F0LIE79G9ODLS8QCjjyxuYwvvD/G4z0N4vYshWwU2RS8Yix3v/CofqoisTUT5Di1bfg
T3Eu4XUx9Qs13Lul6FRIsH9kDxMpWrPkQBphsXLv9E60FBzT0LiTD26DPwy0Zmg1geYu44ZRRFWr
s1a7s1AmmQ6NpaL0ayg2oAiLIYVxLawoV9YjkgAx000Rlm3VzEX6Poe0mvxIxh71jAVMbVZsx/by
nV6d30EJ9kwjOnCT+hCn6WwbGm9UwdaYk9a92kbrZRVI3/yvAu2FnAGXutshJs6dynuRqmIh1Bmz
ebtYIhiU/liRSGlkLR7SQnTx40AuYVm3Y5Fo3kk3lknYauwXQ3+Qwm58zacvu+LHqq1em7vfujUP
CziWb7EWUuaqBNXeV7K7/qsl8fmNeQAi7cGwTclrKCyJUESN9294cPHdH37wo0VnfH1GKnKa/Qj9
d52RmhID4nrKYMGS9C6wVLHmDx6Yh42zDLSo890q+vanErmGaWKiujXunAILe7dtY+0HVUQzLfGN
fF7CprJeJz4qPdHJ92snPJyzgVNMV/e4g14qyMEaJDu8nA1QsQN/Lp+jIOrVREgOptr3tFC3esCZ
9eMzbb6dV49hrqIbfdFlUF39OMjLrHCiJuqELpixO56TZeO0sxw1VMG0wW0bHjKwiIYhHWdSmc5C
znYexU/AjQnKvBY4wSh2uphCSHC8A/mfdLoAREZMwg6c4+GLxo0cqLW8Vm8saH6S4sAESwT03ZMs
8wIBkD6TXlUXWHxtLQDxMrT9E/2bTJ6O/LMIxz0AOZv6G0E2CAnNs3yFu65uVDYVjXwHvc4e6wTy
x/PSZ3+xDbRVulYAQq4I5Ol+tJaTrr9IUvlH0001dEMvMEOUupdmOFCoMIJDBlPjWSIWyBYgnJrO
g2VCcxpdVXfws3WzL6y7mgjW6ME5vwVk52+uIJGELJbMJl/iQEv/9Yd6krdliU7sVM/gFko3H9SG
RAHAZV53CMrONcIXvEEHhtT3vSecWEpxtBACGxAnqt9VNiDfCGUahekaKiSZtx8wODIyr3aYgZBg
BqH3/BhM+ckG8s0AebtX2d55cnHullASO8lnQPNW9+Lzl/qnze4YJnzm7b9UlZ7JEX3ltFcLqxhE
PlzLe+RHkqTx2zNjUQQKqaWeAvr126yEENuoQtYUIEewohAfLnAZJ1nUXU0Aoql6ZOPFXL/opGP5
3V0gG/ucR1Tdgz/Y+SNxNLFHK5fPg62BnIfmhq0YhjJ7shRNSQbEfm7iNROR8aRz1CyEcOHXb8vx
4pKYLLUnuOC+Hja/ZIGz6kWZNIv7qiOpQvb087T0+eLF4evymCL5kzBS54GFbos6tokKhG0WJNK4
r2WzsZJYyjCtFDNEkeYgUbxnlPOUMP//13qie/3N+2HKe+04V/kxZCh1nw3pd2WSelvRunXOlqPh
XVUbFVn5LETX/Al08Y7naKic3YOoJLmr8UA5Uou+oExW2MzGMJc39LB8gFOAElDzpM+96lgFKmk0
GgvIOOjV2AqzerfYQV22T6FY5DAOX25tME4FWJaQ9uhJKKGbEvtQf5KT6efgif/nXlBUODIHR9K4
NM4ifTMe2CvMBB5FOwxwx3ysdyOcBum2mmDhsrFna8lkgoY7K3iblQNzMm3akaKvgDqovzxMkeOp
GPYY6jaNxM51mHr2SfRyR6qfiECee95CB2nIw9+0XXJqw2bq0v9fp8ZhlCzyDlIy16JMHv0ZZ4CD
XqDr6v92csfblvm3kkPtdh/7qxZlX3o1xYG3e+H7Y4zRwEEe3tvWww3UtZEBlYuxam6entab8DWl
ttP2lchMB/M2ysNaWP8nETKYJPaeVn7PlmqXoVkj0mRHzmRMLHL0HdNlVtSaZnQZnNI1Gc6fhSux
mDzo1cevcr3iXH0rZPyQj7AS7ThJCjQhja6IrD3v0Yh1AOK4yFo2Av0PwJekqsEUEawIvnquprT6
7Y0kfHO2qWL94TgLKqhewd5vS8oQ3ealDu/IxD7sTCCTRqkOOPRQN56gd6Zch2K9rl+eg7Ox+8z5
hc/cFMGn21Ep8QPIMG/5xP9IDDXtUsmnCHbatAni3pHdsoVkK57J/n2X95CeAS4hQN24kidRdhHH
pxm5+NnnGlhHtCtSGKRrG/5ysJr5IFdH3h1l6IFFvgojokdgzQ4ONKCtERcg47IEZ9RKKurbvKra
Yp9bQHs9gz2gDH4qUfeeatuKJTemEoucTjwZt7O0PfeGFGiGxAzF8wtJgEnMkHdsHmJxiUo14mde
dHnAfvuUDnyuZucrGrog111vwrarka+rPEZU8g5CfoAe42PbgoGoqrDNk83+fQOdjnhbxFl+iFQN
41FJLEwkcTrbyK+3nftfPx3whXCCSWpiZ6cqLC2fSH7qc6XaqM6ueo/e/6VFtANQ89PxjuExBSnq
A9ITozBMFjaUSnZt5uGynVmQ3RBpqRuitrr4vkbRJZiRQhuwarZNGwGHjAEDOK63wLIZl9v9hzOZ
x6u0pNL1yoFux/uYG8lz+dPQZ/8YxYRDBLk9gHBq8GaDSqdO1Qd1GeP2zDD2C3H1F13OVxQ3GwNP
nub3yZZpvNl/Sa6Bhg41MuyRC6l6HfjIwWXWVMl7VnPDlCGUj+HyLdnq9TT1bLnbqAG2n81VyYTd
yxPvYdHi6Oc5HkgkxdeWbawNObYCHRWc/jVB5DnyitCKk118kA76HPNNk1X0elKXRfplF8gdbVZZ
AgaZfbE7CTuPAsO14E+r15dDKrBcqeYS067pJJAGNxHDr7ESEgCIW9AEGQyDeG8myfI5KqEKjB3i
NM03cJzHO7MMcdUngyn2DzyKgIouMDBq/qVsQh19H96uL7zVKhiYCsErp975e4TZQADO2tgTodTM
THrCB0YZq558bdan6amrgnVBtYmrQXuwIsMdl5kqAThg5HkH4Ou3WakoF27K3P7+Vi8KbuTxsdOg
stQsVw6pHR3HDkmXBx4ThFKm+phTUTqRhkOw8qPj6zXnaM32zmD3nOxsyy7+OyBCNw8mdRQCaddD
yzXSOOa9YvaKugHDluUQLwJot6xOJqNSYzEpNjdN9M3bPfIajZOfZ8dQwsggC4fDPnVCa1wp3+ws
e4f9bZqe5gYyUBC+31Y+cMjPkRjz0r2awhborRU/q2P5PyUthNi3hpLobI6WElgzDdfhv52y3iM4
uzi58YlnFokGjSx91CYr59yixS3DcvL/830KaCrJ9BpVG8KtT5ro2jHrB0nWb06ArInLvO77H66E
4bMRe6x0GXx/DXt4FieszmAbOdUOB33EUUcDP3MjkWoW50AbC3sLOyp7EU0PtKgefnMVRFfA9MV1
njqweWYaOQUKRhv1H8HFB4G+W+ZdxGduUW6oShGC0fIyMdNzhSFAxWOJStQkqSBQ97GfBeW6U1zO
RXRyucuB51sc2FlgIXuzRzf1VDaf5LJfa363UnzmfY8aG+Q2EbS0wZpGEUTtgTqmMR6IC7qUK79p
QeH1UeQH4cKpuP/glij39baEIJws9OVrjkXaPrSUPVv0UIdTnH2zS355vHv4eNesN/yTmQ9Nhwr+
V4iTfP3vp2VTpVi0KedKrSeJTDyl2e4tRqwHo+qNwqIkm5sK+PqOazxJuZZlnTOXCgJZrz+AV5P2
JWU++OX/7YyEEeoOVNQTQqXd9ZeKearRo5EzWsNPXHtDTiZWAAZ3AoFCKR1zLzDQx1aZDhlWWyz/
IKKfqUOIv2zvIW23v//K7a7kiQRRd3iXRYSLJN8nC7GNJBSIUy/BE622Dik0bnUKv4wCZ1PWjzV4
UdogrHOo+aFtb/VgqZfLFPUDXV7OfmQOvp5OVAd6vzwxCZb5TgFErSft0cNu0YKHKxV7Ln0pngT8
LCYvdpl2vMbn3WTMFFxuJOwaS35Mt84Y/6oWLHXVwx1OnuexiWLmU8rKlQn73DMm/9y7K84VXoBq
CPLeo//Df9/sB8U6EPUQTtBs6llU7e7Vq+XQGN5TCbRTNnFrdBduaqPkRYSjCtkksur+j41VdLOM
fWAzEC/OhYxfDcrTgOFHde7NhE0nDUtNY8UDwGSPPGj1+vLLkDYYsxL1jkru/KGSPPsRUjsGktyG
ii/rB3PAo5ZRh8aFxCKGKpbb9WB1wa15JvMQvEAIVnifZWKjak0q5sbMxzAgFhDn/nyQu+xMlC1D
rc1kY6Dgncgkgj7lU0EmFwPrqtjHRfri4VIbcenECFmx5y/7QY5tFpsxhxOtEiP/9mnm2wCDsfTi
VU+a98O62s8GFI9OcgUHLmeCENcfuQU9J1nBit/h3ZFFbaDewwB0hRO9A5eEHhLIfkXboxsJ7Bmf
rxrI1ZFnD/0SomekykuEM4YDchOrs7qiChPQjSCoxyswIiGEEZvLKGwrGct+NS4uslvR8M8sshMx
Ax9p/OyQC+xks+zts6FSbP95PfagE29FMxA0EBeUt1ZVgY+BoJlHMX/VgNcbGubMbsn6dd5TQbFn
r1tLD96DIhG7XEZsK47wJ0MZz3CPyqxrO97xTa07hUMeE4zSMGAchZ3Nv9aEspyvYXv+Ujl/EFXl
3xdaCi0gPfo+qAVCx1KuMoNr4TjgIRaFJyOlPEqWz6wk5ycuiDOF0z+5J7m/sdkNAMCe2OXjeXOF
Vtl3FNlQHmir1iuj8cBBXWtVVak0fli6Rzq2XSTja3duXovz5sCcMVUcbGy6FeQRuZCO3VjkKjQO
2CKLfVq7GhVG++93jk74JZEcoIBFnH/++RLo1HO4xBYH3f9BChAc6X9NTsS+aJTtuEfXvR2L81VT
fHixQQ3lt9uL9NpqoaPvcHyHITBmttCxE889Xeh6XzAIG6KfcYIcTlhCirmLum04888/v5zEMUIx
oSZWoy0lUaj88nrs1CRUEoR6Bv5kVwi9+Dc3Qmq7VMrIbG9Dem983UqA4iotUYj8r57MwhVPv5S/
7e9d/UFf2J3iftNeWKtxmhnU5LQCLdpvgSc0kvIRutzHX1yWuZC6gskHtbTW7Y+/ddejY95ZSOwt
M87R3YScL8mvywEsHiXMcGQ9yP6qUQlMBPFWNnlWT47cAHWJ2192RAaXluc8MzKUPyGdr1KexJ+q
6wkXtd5quIMCl/6i9DwOhkOHetwXSmq8QQPwhfHl9nE3qVR+qQioLtL80IyZxKa4/Z1Wt+dP3I80
EO6nn1BDRixS5fx7SWwLGso0gHj7NH3/CWk1jgFau9GiO68rGC3xPZU+0BtpCwSNRyYkdIu8zuc7
Ll9D7agYM+DNnCm1M/9DoBm2E2GdK99Cn0OfMVfFZtdjzKTYiudfqmKuXLOKrfYWX8LRHp0JiTWB
5EXas6Q5CH+ndIxwQAu46eUxgtXL/XTmidmavZH95xtKHf8qolf/9afrx4uImPnE4clEroshCjNp
AqXtSWEUbHFGrPZsAxk/RMf7wG5v/aKflwGvcfQOuYAK8ird4ARxvjE+rkAN9gwLMvLzXJElIm1E
Z9KF68TIIDxAyjF3N6Prp3F3DXz9yM7mtZrtM9L++qW76gAHnVvNZVtUpBu6cjhD4wFoGRaEKQ6y
obU/UKpRwvFV5M6DPDTt8g2qCTSQsppWwWf1fzUSxUOk7BFcHVhDJXyCnfDDvdTbC48hVQ9DQMUI
Tb3XlZxwC+jXzUVRee6SferSvmjOgMV66A59Sj1w1C+zhoNRn5x3SQQ7mzmAHN/ZiqVwRMM6jdz7
0/avILTMvwy1A5gRyO+72zfGAQBGxUsxCUvcavLW+PU9uID+fwaNkTHRgQ7ghksQWgjnxdtkvxso
vRb0TuZyLu4DZJ/q0Y0YCxkRfsYX9N5hgTd1OmdsdoWuXdhyvyl0vN+grhOG16+jml8qARYu6cO7
UWBDbqCcvhL2GuUBeAVHgpYtSlZW8Weu054t+NkN5igVo5fCLsn3M8NX4YIZ/MMZ2+lw5QFkumX6
jwQ5Gw8msxAIL9h7Bchy+yd4R/8Htsk3RL4uENvp1By3SCS7qXctyS8ogtXaTHSdPi7e8vh+ET44
WQaifssuTaOldnm7uoB3dryq5TqzQQkJRXEp+tMm4JNocNcZfyCAojh0bt51jhPITC9omNHt4glH
+wvPnjAxbwN+JAcV+D5iVX6leHfW6oAkFvOeFsTzY3St2LQns9DgKfTLx0De8ot6xUn8ZXKN3Gg+
nCf8+ZBPQHOkoUaTlU5EQdZOPw7FSsBf0uayv7PApBO1kzOQ1JXaZ48XcudUOg7x6LN/VLJ7BHUR
0h5Jdl+uqRKFuWTdgTv9JwuSeFEq2+T16p5OZzl/3t8VjaGdGmOmLl1X3nU/EVnzPnrMMzU7vImC
9DxbNqTUsl5ZEKGBZ1Jcd588wScWhl5oXUpa+M7NJM7c5tmAhQI7EzpGk8e8B37rhJRqWt4krWmw
RPyP7J5bwH1LXW1NiMF2SDRUr3M1GF4yi+O8vxEhBAsyL2U/TUBS/cVjrvCClFKZKr6TFOKEWOgC
Y5YIB4rte11VafVRg/CuznEUJt+xwgH2LLqJT8n5YoSZecr9Dd8bJ7TtDPm0bdZ+zH+Vhqy2iAuS
wiKP5lsoW2+hjwzUGazDnDhbK6zG0MIll+WfxgkECXWnjlB1lTagOhvAJmdRuDaexFKyFKciflmM
iXLfuV8VFNMs03xmKY7w/4gszAjHS41pC/aFXYkpsAeSzFAzvILjabA2Mqf0Cfl1fpg1neN7+ZOf
rxrqlH0kG7PqF8mGfj8V3w8XJlNn+gV09SVa1H0uqhpsYjT+RHZu6FPvZWgWZ4cIgrYEBqLD9Jbg
UPk2ypWnRnb/HttLRo/BDiRimod6jGgLgOTYD03VBgYx8jD/1uc1eSL0pFBgd+xNlr4ZWHffEfYz
yQVY4CbvP8d1kAIqpL0yHVPAeUaJqdPmwPRW0wwR12RcAyf7HFi3ccFEJft0D2PD0r2S6dHB0+Xl
Kft9R3DnlKQeL4l59In1SFe+Bf+t6EH9FbfF0TvIc1qtI1nfw3xCaG2pfpcGBcy59aTNPV6iCO2X
kd2IqcmQz7WD2fTE/NcO9hlu5gp84PVUITUUmKCzzx69KQcTLZFv9Zqgu3yJty/+gmnpBce7c6ex
P6yjGXoEeY0TxMsjTkF/51x4xLz+BN8E3s5L5JO78DOHpCQ86MSfoym8UnXoruj5mHz92Cb/bnuj
rpUqVcZEjVvZvHOc7cVurLTTCYA0HhhP/dVGcNrZCJJunkcrBm7k+y44LYA7psD7fKtdrZ3SLhpt
CiIIABklQ/HQh6OkpfG3qhnTKpSMO5XephVe6FIE2R6tzmFSTg/1zuKesuGpzvU5/86qbOMdusmj
IHQoz8jq7JwyeEx5teYkj/FAC0O0xYvPUy2eLGjvhhxdFFoo6sL9/7XOhHoC9pkWcIAa4ItSYBVY
bD+KitFOSBUwuIbhxz1UFHfkobgoRRW3/vAq+MTRYW3fP+id7F+7f2hrGpZ6SBP4y6fLppUMUW2h
TBj5CNSD/8Lktd7AVmuYomM5MIe1+58aZXuFBz+9xWIdrKT9xa7AZH/73pohfu0EZig1kUVjUB74
5wX1D2Fs1szu5sE9Zdjuibv64Y5oJnPNUPkWMe0AdRMlYlzc2cYxjeOCWnwcTbNRBXq/LWYF/eYp
abW9FHvPsoQlct3GQ+e62vT7miUl+GyBUkmz7d2frNSbSCD8sHJasdsX3T+Hr+OF+iytSnQ3WLg7
xmGMhUTyS+kk4P4HO953oo88iG2A0bOJPAGr+AOKiqdCfImGcJukV9HuxE/uqcudZexSL1WBxB0r
9rsHr5kk6ET4NYQLzkMBMSnpU9Sm/Myqis1FfvYzOxA5sP0t9HtYGOI7AtGOt36PboXi6OcOeJiT
30Da5DX1FpITMp2kH4DscBuYDFmWIsvkvu8hUXNTyHDoN8hB/64//qmxdDOVQ1MopXlpgzsZp68d
wNmuSKZxXUF6DSwnLt2VQEQVGQXINZdwskcR9Sag4bGSxsQhyBa7mdCSzTSz39JK303B+qqD3H6B
LS1g3gIAFHQkhuYa7+87NdNGpWYizk2kshmMWHNO9vvIVaZ77qJJxIi2IwdwNkLDpauiCudiS8iN
pXFsXlsF7+2ieB7GUgsCt9/8eRp62OstXFODFSspsFuJF9/O+aw9kmB7c6D3sOwgimlT7Oi9kWRE
sQwK1z1XUgcOImBN1zQ5JQM5yXWPnDK8cucIrq5pQtfYFY179pAvyCWB6BEWFSGMTYl1C2t5NOv+
6sEqyg8zZ24dbwOK6QPcnGHJR75DxLYVqzVwSrl+Du5QdHDvUJVAqlhmpIy7hyBqInK5RqdBuGzX
PqGsDe8ZAVJn4kfTQ7/uRDEKCFPZvlsWgeJqLZbcvUD7NfTd+DoDDy6qw9PRQAcfi98IQGbjv6Lt
EP9XslS0qgW+lJZDD9afCljPy6+xnrcs99HlyDrMcaJ0VWPwfYG9gqLanBm1Wt8LIicG8dwrycQQ
DPLdefjoujARW0kklfxu7Bj5KE+6oHf7kMLcAvLTxu5UzO5VGaBmRSLtqOsvd1IHAQwDlDsZTFt/
q6zyr+67HWIrBA4hIHaHoOLzXBO1YHM0GmIPSLiKWkFYmH3qc0q8tTrx+f+zpB1wsGATqoqALTDE
mHSQV/qE6Ly2vIYvKTes+NxvbsAhZGqaYzB0zM938Ki6QAcGHBHeyL6Gi1uLq7RwBNarp60S1Xs6
QksM88K0Zq1iganlhFAVyn4qCKGo8wC6ddgevKHwWp+4xvnmQ2IeGMtVHvt9fF24DKYI5N5s5E1T
OJOsmFGZSV+BfrTHZlI9gif551oNGVMN7X9MEpZKifoXEjnMkqlz1Y44T5WhVeyGmrxl98kuDhcM
If7IeyzzyBzeZCQvq8bDP6SX7aAMP695ZO1AK82TST/ERP38/T9Fzm+zvbqHvVJjzgyHuBewh8gf
TJjx9Y/smR6IWyieE+L7D1sjd8/h52FnT/vjqnC52dHPQlDFfWxuw6t1qR7f9BU81CNd5UuBX4cS
cg1H96MVN4gW0RqQwlFesF9Ga+Yg8WeSmO6sE5jAOPQn8YewmPwsGVpB66V3yOwEK03epAVcvSaP
mcx5wcmLoIlz8D/8vW7qfyNxkO7yZdIASNGiza7qS+Zr4/gv7NoPRV1LZL0tLHDDE1NwlhjYvRmI
IXJnEHISBVrmDUKr2W8y9FSDi4qmpWrocpq0KCngTyifM16sOppLIru6ESyWrVSXntu/6FwMeeke
ScK2nzJvnqTfzp3lQ6MsgAgSNXHh6FidgTYpdDlvJwlrJJmxRxtrpMZ1RH4Cbslpvw1KQ4rVx6uk
bW7BDhQATK/uRK8v24HwzBT/b+gnaRnTsBlaB4ze2A6csjUQnKEynj/bmNwuLVi6J/l7JiXiaYXp
KTa7tNtlpIvDP8eimXh1UeeKT2pHhG3bUmJG7tbWSVtPer+www3UdUs36i9uSNwkQlwz0zxotLXj
uWTinl7auI5Ok8z0wup05+xuhBZd9MsZOsKsoqwGh9IYiDt7wmap2Oap07LQBLGlS8F04fgdkxA5
beXVO1SPLxImdKCgs0WnSwXRTtVI61dSMxKIbq1ZL32qD/bLo2WD3cciKfIizks5L/WfDcgMxifH
QD/uwK+EX73UPbxeFP2hPrwSIGvyRYRteD5K/8K25v+4MY0PJpPlIFqMSq5jvkLGZj0BjbLZfoMl
Tt8pTGfZYy21oMV6iUOZ+ez9Axl2Bwb51DpBhtIB1lPNvVTmwPhXjMUtoaPPwVzkm7LndeRgDm2e
nv5et6sSWZASqLTKKy2x84Raj0YBUpN3xd51Ioydr/dif3yeT8TTAiTiyvoz0KM7knM3zsORUMJu
q2+c8duhNCuONoSK06VN0wJjs9+A8GUdQ3bwKL6AUYh1IdGCg68fYOZjcC0qQQaj01tvIgL/aSvH
BmmIB3t1fuz4PNd+nZPXGWBAC0QB/RshVuR74oZyYy7M0yJD0HLVTxo+p6PcSpefBtUjY1KR5hAt
8RJsD7TR4LsvCgv7cg5Ku2GU54jsNzbOFqv8HhEY/9Tr4Xsgy+wmx1vvR62CXKM7H8DHdzKFWMQQ
Y+ZCAXzAVmiHypxaAQ/sCrRu7C0kYCM5+4QVCiWIbX4tRLUovqQakDDo1kbjphJ/yAuFrToF5LTi
2GcPD/zajgHGVdzsGxRnmBcBrPZilnKMAlLPADufpprIar93dspoudbWOAmWir/+C5VQmLzzQZKi
FVJ9yWXlOxrXUX9J7IZEECngwd/6WV5hiY/xGzu4/F7KVO+WsXECMMrDA59jWw1hq7jArknAk60/
f59BMU2vZryorq0llvU8X/SGpNkKPZCByjTQutM6aPUk8YfTQks/orCn9fxnlbnZNJ/hCQd/ukLA
NHnBqnNo6mtv1qccYt4hHyDYEcoz0ZUNRFmem4zHj5lm/g40e7ARiIETP0APSkDLTBsM/dDL0yiz
VO7CNJT1efBtqTrDjQtGK99cj8h55IfPsJ0R5CDM9i4HhAO2tZyVYbpct81xjAQeI2FDJR258MYf
mZNJWNbQMcbJvaleIkmbEUXQEQNCpnjOfaYei+OeL22NulTs1uP5JK4fg3hfeZAZfH8jZ2Aamc6L
Z9oBdxPKyawessyJL2s3QfHGk28iqOQVxD+Yy+cCIOK8J8cq1kFpTpbEmT5lndDGXIjB+ahwJUQD
UibOFrlOlqZS4amsCSA8xiLmIzbbUVxnh8vBZKUWcix4DgU4NgoIKfGIFLQuJfvQYZsI6m0ejiwv
DFKfR83XbvzKz2Og0FTaJUlK/3j1vOTNRaEGS7YkGroTswcYWvBHaFYqTp402cBpgqOnPwQL51Jm
4Agd3f+p9/PZ6nZOzmp+6owRXYE59Bqtr9PoTmkmeEBxv0EoNYxu0IAKLwsRweEdT8fSb62+sanB
Y7ngxttmgLPVNa++bhMft9pnc7I1cWO8B4mZb1FnNvMrQb5bqtmJx5axZb0k8IfB5daigtpqnLSu
iLPHkgB1MljHqaCYINdmefpFQ3FizBenDSVBDjY0lnP3z5XYmVQYcT9NM3r/sN4bCg7AfWxReahE
xbfrvD3xPfxFyJ/pu76PaxdG7vyGk3Y+5ypGl+Y4QzflSbzv2eAjSC8ujzBupj9QYRF1cCg1E1p8
EfJXO00olUPowhPkohiIERpc5sSXkUWFzl5U6l5LPgxxN0ax7jXomvbs4q9T5HhzHAaWM1BvSCPE
ptmIIltAkavIpd9XHIuREDD8wH58nzUlh90AjKuhBTU6gYYQQL5XT91WTAiOuS+08AeLMBWIVbr/
9EfX7lUd/pCEZ9RN1lpHVQL25Hx6tTgucBdQBz4eLLrLbfcdx6R/Pbv3jqMfhmU4qEgC3Ff6AuAq
bzF1l/LmaNiW/dWJK2+7rqC6kUCv1nZFh6TjUL8uZ4YNbhjPhAwNCwGr1usmi7EvKIGAgIrRDfWi
5jhpzekDqzY58+zngUzBLevRe9cEhK6lJcgQQRiY994G7EUf6moyzwXxmXtm3Ns32nmJxoMD4cr/
fu0AgUdQyWPcXMsQuUAjFxjx8cCVHNpq2xor7+CSGg9gCOOPHPXfxVhDpil80PCXWUU8B1RsQben
N0EDIkZwNXu7S+xY++/aPurQlqI8P1HvZ8vVasotT2vz5oLtcyjbIKn6gUzkdNQMqaYn0+D8tSYT
yaV3Pw7549+m4czU68UVQCjquSEgfTM2sN9AIgr0qMUBSD9GBAEb6Yl5i9rD82H0mDnVYzpeUplL
INRn/z4WlaGzLhb7Bf52TlDVwfhGv29UttU+H30PiTiuSWfJ5MUTJ3QK66uSAp3CbsC+MJbPoLc6
AuwSFc6cdCWCpn7pPwAoddHWz7ij9cFqEFefVNfaPGyOWr1jVKk9vE8lV104q7VukEJfl9vDKIw8
xbE9LUeIdAAsedVUWt95WcEW6sTQ48ffC68YhqZ7DyhBhn8qZAPfRqQCCFNldhvC2lDWUTnKT4oq
/dbx59hMM6BzZc5ZNcE4ttlZOfkA/01wyxlxiq3Ur4DxGT8sFJ86bSbE6OIdNny/nv41ODsvXcLw
qGll7BTWqntrjzmXqUPzzipFbTtGyBUZ6mJvwcKd1kWfrmblzxqt2RVmTZAd3VkLPp6XYI89QsFr
m0ardgt1S9KuI7UTvsYPv07DsKksS0H0+cMa2O3CZyQMw++cVs83XpL7p6Vr6HOsyj6izk0zFrG3
vei0OVsYenvDuenWyVo4rR38UM9khFhMVexmmtpsW5BR6hTQMciBdtVLkIBVQ4hOFIV978TaOw5f
dcrBaBAyCvhubfo8lxz6Tq/20w6juRZAz97QYnnDcg8FHoke4GNuSbp40HfevFPovwz+B8YR/B9b
cHVvF0kOnvrNpk211WkFksaGq11+HdiQY/Xbzu6dd33Q/RNlohsVdU2BusjPWZIhPlYiSubQHDzr
5eo19QQrxDT1RBg1i0WxKt2akpFnpoKrlC1K0d4u9Ov1ym7Y8NPLZqO+ucvOobgpRsvgnVOTr3Cz
Z+lIn2bUpCGFjwSpj3K/htDu9vhQ6x/Ef5Z4l/2ZbwxXrVrZ4Ynpf5/nWXfUnv1HDxpkEEwtl53f
5s0kOAhycg5Fu8Mkc9pgni7x8FAEQlUWZdrW34F4FZ3vI7MsqBtmmBksP/FkOfCh1WY4R7bLL06y
L7AlhJoi6GZigKvLkW51oP5C3ztqVVhGYVCjy6UVBZAJXffjwuUT9R82dI1noHmMPKZMOnPWl3jk
i3J8wpEvU1CDUfLCgiofWZk11cdkWMvbvf3J5B9wSK02oCuysmIxQ4F2AHEx12a8y9BUWsZrYDQL
zsW9Lw5zw751+YOtHAwiN5pcS47ECQvvU4rXEYf3PToLmCqvMSAnj5tonX9nmkFJIqi07pCYHBTL
vtQNLtWsxo8sJHYrJfIJwU4P9dDTD+WsR6zPgrGnvZ6+LwCRHUBCVL96O/Zd4GMimT7xltaicWWb
uNcP3VBje/0CJIrbNvIrcnphsNDzZTjNqwzNbdwGZ/LQ+8QhBSD/OnZk0ldYKyEEi5YN08nLq8RO
DY4EtLdu6MClAnvy7FGKOEPC/lYed9PU9omMBQmp7W5Xt77RTrwgVKFo92Sn7UKMD2AHjO+coOOl
O2GYONouM6SYwZdHAEKOSufgYXCG05+QVIB6IP2e9uQ9GMYGZ2rg+Z9TPO5gO+irpXFs0nAUgD9O
a94JubgWdhWWAldwtBgEXjhhYLjKvwAI4NrIxnK+CHUOqLpaqd6nMVEpoCb7BhXnUe595bhp+uLJ
1FqgO14UIBmwTb3v5a5IvtsvmLHCx3+BGb09n/FUKV4VCzdPFvA6cZ9MqM2jYx9Vbq9cqdRnSflj
HYmgAfrq83MlhzOcLQDRg6E/CgtNmlr18fY3QNTENDuWwuaMjTRxporHvPQL1FWM+54sKp41H2VO
mOcvUymWk0o+FkD58gujk4khTPUCn75U54V6DjwYXVoywEMz5LD7umzvcNt4hWjnIP3OWkyJyivp
zhYYpy6jIpqIRMfiJ/HVF/B6i6tLQ8ScSTmm4mGqFBN5uzghbtAhvZwGhFWPzmwnRG1K3G14ty6C
qm244Eoqj7Zx+GubO2TprTBL4IciEjTub1qlklZSYxSiVFMQ2GuC5/UR/lZ1dTMc13YFBSKc+UZU
Zb6bacH7H5udmv5RPOSq2yzXGxxVEdouNo48sJORPhajEtYGNmp1mGKTxdgRSozKGyS+z0jZGFGa
OeNaKdy6/7FJMaXlIGXpzR05ZUs3PSSF+w/Y1JDIt2jqZPBa61ZBmrdCKke7Yui8L7D0KmELSF1X
iGAQwnfuph21Ykh77gwWUsiPYUZoEEqvAyjsq64uNsh2d1O148RFD69FHOArzlPLU5lCi0ROZmZa
pFFpxKfE0QwIQByiIrcr9mojnNIWHNyYx5OVpKc/kuo3qKRoZYi0iWf5hnoPuUr3NGtyuVE5v8S3
KADQZ3CLtqb94H218Hpd8VmhkoNb9IVbLPorgdcsxBsc7aw8QCmig/nJRhwANi28DYWLa/l0trpj
tJwvA6HW5oOFRoPAerWqnVpal23twIS7RMfYd1YoPVHq8oDcgrXWvHmnSyy6Hlh0JSQLHV6Xz2mU
konfWu7wcNSfqOPqwMzPcg6SMqQWdBeDrZKQIolJOxCZk+POfrhPH7pQh2ygZjPplmypwXUbdxst
synafCDcD422OEIeWevbRtuB5Ubo6oGRuu1nl7EK3/BgkeVcdb8Lduc20y888AdkLgutzV8ubL+t
eaLOHQsVbwWAai8MvGBRc+tZpkhOsJcuM+wUNcSYl4CDtVtr2/NYjQWXAFzfJE6lwwJLd+oj+PtX
OKcP9cUwEOHlU3kvePzgWL8hT+R0qRIlQS2J6JESqIv6Mkhx5/RCyhVjN4mZgoDfeAZP8rEI4zuK
eATf2y/lu1g0EcHXrLO1QpWAnqTu0ildu4mx4TmNIFksSsW15i4ijIWCcohFhc0ac8AXv801u3P5
fy/oMHGxGGzEk4NbWPAkMpEevGV++8iE4AuA2pIOd13WvMe5yj6C1lIQD8u1jiT5+vRBFDctviI6
u/uJVaWi0U9tFl6YBpP3VJqyE1/eRfMtBozyKxyJWAcv+axPGeP3waHFy7eqCZV6Nab7EF//dw/z
6S3eajQB8h3IYD6uWoQknDwzTGLH+x3/o/IFFb7JNXe8vfXn7Y5AmuQLjkPyb7+fjF2u85sG6+rG
hn7TV5fgY2mBLATwEFs3m4v8t6uzpSo2vsy6qd7Gd2XgBgXPcH9jI0FnWFGmA108Gyzq61fKFeEQ
kgOe653ygI5G5sZC/xGR85WGcacgplrR0/pwZ42DwH2Me8vLuO8d7TY+RJt1yl5UJBH0oQ9MnxtP
QgpP9QW7HoBPUk0HVZVRXdsUQCxhes7DuH7IPwKcChJze7SjlTaszASqeALroITjVD6Ew9LqLlF7
/9q/u44wtvCABTNoGMLEcTBDy5yAgSwd+StIZgB9nA67XcJXkCB3Zflu55GMbe31AwBa8sthN638
zn+7X69u2xmo9bpwj2ML//8UfbklVpzbTSR+1Ds7dFEoYzoSXIh+5kV+9ML0FK7XyBfcn/6ODwiG
gPxzL5WBOrU9ocjmd59vjnH5nUA1uVspMtA+mG3oneHVTaCAEZj5QWxTYb49pe5ykMCgnPRTkKx2
4FL55UZPKLGPLnw94pvolP8rrnEfkHtzGagubq8FNaWMBOdzrkVoVfvZeFxFFmz1GGKRGp4rpEVm
y0eZlyD29VDJG9fpAXrZl51CKND+L0aab50CjuIwYBgVoa38OpPU/MDLSRyt9d7NKtgVxNjk+HeX
uKw7FQnK6DuDpByIaM9JvdAgj1gynsFt/tKwsrDLhBCy38VDwUZCLaRGGWpc80k3ayLqgB224GGA
BrHoumZDrglWWM8aYcD25DMcUySodYZKFlTv5YqUcywaz+tGZVD5ReT3OqoUH+Zyg9eBdA/XLd24
kUQw27rxuvxiL+8H22akyRJZz+aJSGBZVz/MLU19m6gQe7dZPPcNqSSv8eUzr245ZvSJXvQA1H2p
sHtmHXC3b9qXhYMVdjZ0VMUqzPop//1eal8I9/fOoKC9EpKsKJkHh5tfluIMkESkHOZURv7lvJmm
KihzoC583TinN768O4aZM3YHL3u7TUOAMUTpFm4OIm3t1ZjjVOvOgTnoB7z+L5Law61pWJyk6cJU
cgpq89UtGJPPHp+yZ0H4WP6NFGGrzqhF1g5Dr9MLZHcRlMkY3TRJ3eSpldZNxtpiB2VfBzDtEA7J
YQlhZtGOlfRT6oTPopOzKFQlq33VmL/JbArXp9hn1x7SCyyAkKwFxZONTwLYyk7mW46F1l6bjFz2
P20/Olb9ZyeZ0E4cB4eIJ1Dh2Go29TrcLyULBAAEJiWyu9N5n7RD56V7BTRoTItQMXbyrIih/g2p
qpMXJ4NOMbU9+Ep7Ip+TvQbpfcaL5fXD0Regl8buqGbWNtYRQN6v1sNzHF6NnbjJfk5XIFFtIH2w
SJNXIoOlg0/+f0hqC7uI9/zbIO/QxkS0GZUiBrfEPFYRfEUBTXjBh+xFPRnDsj/uD1AKye6r0l6G
MFoQejBBTCb6hI1TJc1DKanMOKn/6kxUhghvFmW3TfGIsAYlITPIx23ENg3O46dI9VgNyRcS2Lvq
pnko6NYgaeTZ54kkTEAvOkNZMQ1djXI4ylWFH0cX8oh9MUs0ZSMh3zTLKlL9iSLfePnHrTr0fgYI
GqjXUT8U9ZKksDEBoRmY0rhrgyKkUs8Yo/iKkHyNb1waJ5RdpqHyjqy4hLE3aWxWBCRRTUfnyuG7
EdHA5Ml3g38TDsp5Uc8DmC6mCoXKqt0r+ShMBKbxeqGXVA3LqlKM4nQHPzumTz1Hzf5/IQbLU2XI
kXF2tI8EpoETidTKg+5HbxTdm0ogwHNDViRX1588MKIqg/9AMZl3lNi0dzrBzOpYzzf3Un5wMHTy
ixbRJFzXLQ2dCC5v749qEHK7F1OMfzwC5kFB/S9neIFBydnkOcypHb7RDpmWhj7teKUuaSmf+9pH
IXkCuwgQ/As3chBNrAOk24vB14Lt3Rv3fIRvQ7ETKEEOx6ujTP/bSdV+nPGmMXaHOHeU65HZv4XK
eqssJ9iiSk7r9f4uoOM7OLv9dAgj1MtviASk/Wh18Fa3uZVy20zZTBqyYk1uHaOPhwHr8vyPhRMz
7KJmGLoD4Lo5xSHsgWWAJjt6UP60u+K5qMKH1kXDgxn5+XDgjgclybGd9JUznEayN5Z88rWTAmHI
Nq0z5wFmIekUPZTRvvpD1F62jyrKeCUC9T+VtzbR2BZMLU9GgKCkIt2HXL2r4Xo+n1CjP6IjCtKp
Q6sb0MAC5qulklBxfYC8FKZn1PakgsBowRnuoUKqQz67HdDpOnlnda4xYzgxYCf7PLiARbXzH/hI
Jxd5H14Bc6AiPe55FIeXz3fLmkz/bp5jEepF5VMQuleG69k0FoU2/l6lNlVN2NnyFwMsGmJwCuZG
7qpcGi3bCBX4srp4Fkblde8gAWaEPEVtRVDKLMEhCxE/WiSwsapGglaelPsFHvfel3PClEv/RSgJ
FRg2qkPRpIOFVQe+yzqFv+J14Z86MWoqzzRm6+XWLsXI97W5w4EyBpLSK6S6FvHX9SsXnyNjKr10
mArZaFWgelVPHrtej41p7/Haq3LqJWDxdMJuYFEG/sjUQwQhaCbSdTQNb9/8nSZgBR/g3wyAv/t2
pGPYLDYzwVkw3X9vEKxZc2l6aMdKs3RS4vd6VaY+7WLY0oVaWu3sB8WwJt4GIgELJ+4jbVOMu5EG
rJ2ICZjb3wZFVJQAnNVcAezzCOwzxfljYCxV3IurkHAHd3CnuZPrtv0AngYB9CbAbeoWoCT5UjEg
sxJJf+TboF/YqKzdcrFuK4ct7QEIh/XUamoNHlDLIRZjUlvHVFUxfImJatgbhdV8LXr1nLnRu3K9
tdTF9vbbwstm2eZuVs1tecNMvEpts5aj3pHpju733IDyU/r4qj2CAawFvWP00ZC76z6Hx7A8FMiy
ZRDY2ySd0DesPeyrOJOMR8e3yCRZLfsm63vo9cVyDPCNaU/cZUZ6xfq1GlL4sZpYEVa+tJP81v+G
XTjsobilpfxnhwusoHtDDBgYM0VWcoo6nXP4yeJxT/y+2N4WSlzd7a2I4RZa1Eld+xO8FdJXl+J1
YgizEhSKUtTCNr2X0CH6aqW/+drxK720kTxSHp83mcmI6XK+FSUadWJBdFuShSjQ1Nr7lBB3JMzZ
uErCM8u3C/lJcyvq52XJda6fGDyvAYQ9ZGjpd/ybv0ET09AH3swWH60+v9J4i76zi6CGY7GELV9w
IqHTARl7bYkVdMfvqC4k7aOAlyCDzWzqk4Umhb4GMeKRs92Tihos/jFyeUrR+Vn1qN+PNXRcZrvu
glbrENJKRUzbQeJcicU5F9r0Xq/8VLQ3gqqGxd7n1z4D3uI8E/hUabziXbyooONt45Ue6s3XsiMk
3MRxcFLNTHW9Jvl/017ctWp0JXCUaEW4GqZiZMRARj84Z7+k2lFEH0DSaWZUGg1htGOFYrki1InZ
MJ/TVwtnJ8jIwKwqHdHUbTBpFZDmPWK0vlAGz9blHuwGnkntGLQP4me14XcKcjhivI+oXRR40GIS
rdubh1A+ZMu5ifMO15EWLabg5ekUGPeG2Nc6eIDsFUXPlkwJM7g+30w1BLH5mlj6uVKqnndTV4kX
60qYTURhRLCkOhiWE6PI9nTsog8+HVE23gU5UxVaM+a5K1LEkbnEadeC0Uk18q2cYpkDKZxUwARi
tguzWxoWctnhruoU/bQs5uxUW1MvBE50Trxmx1TwvZfgi6weBLLRyM1zRn3VqIYHocMUfHNRvWaf
HJ4zh1ExnBK1OZc+yksYq9Wx8SbOhNxFrM+5zYNPOs4uDesJ9kbpqp/qjgGOZru58lOy0V4Vrmlb
LAOT8IzDhPh1A4YKrN1VWVdzPbczpGxbbRLYI1UCar8sFugj9/lBs9XhPR1PIwhLF/Dap5qTEynb
6ByCaMI2p2exyHnsHh9jkGGP6+JFu22A9mijrsQ2KTmBImRKAWSqpi9+B+x37xytOKYUMn4n/Mng
yWx8SdCjghbe8+HfPzqri7WgLh0O3Y3WXEDbtVysfoBiFbS31PJ6fTjFve/CtAWZXxtO5V6Qwsed
yMJgqBDYtYKIzOE4XZNWjI6smTd+Ld8oMfwR9bbUncpMj0cczJqq1dGarZEFfFaCooedeqkVXLtn
hYcv0H4EPoARqQrf5eJ5X+5GKJWDRFfxzGIlmUER53boGaYfjZTCzMxp9q2l4eVxOJFpT/l/JAwt
UPKioSnX/ioMhQAYrN5T6zFXgm6J/TM+Q1aCfR2J88c/YEXX0/ErdnEol+ayJuJalJRHVg19SPA7
O1vAbmGVQYkNmLqisICYuxHTpxiNNYT+UC8dpIRmjlkywkA5+cT91EBYua5Tdd7NBarV8ap268cy
tHBdg+NFprJld9F0ICiy6mXoLSvcJnapLZt6hJ4MVBNjhsmf07dkPaNRBAmJFE0hgrBcmgCcuelP
uwxf/ohhj2gvAQ==
`protect end_protected
