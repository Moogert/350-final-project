-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QYb0qy+i3fGESd1vEY8JDBHlWOzU9y7tKF6gsFRvMb592zKlD9APJyEk9dSchTylUV+DNkeBqNtw
X0lAaNEQtnxSYbOE++h0nzIypmmqDZANvmliI8LpCYZaRBkLLyxCsnvmfkFAx29mGkbcq+g/EjVd
F4SCiPME8FX0VFRRfgypc0Oyochq4guTJ6ztk8M46mDDhSlIB6+uZImC6HrJcpXAXUqGBSF5XYSM
IKBiYBccd/Cj2K1HATKP9RhggXVJLj84lrQUuxOkR5AEB6nLBT+YpMHpYS2grs+B9+2ImVFOSGya
s6qW89TZJer0FoV1nWvbz33A7K/fN7aTYYjZSQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14544)
`protect data_block
Qed5JrXz3MH5R01RSa5p2u/kHIFB1hXMGYIAD6HiZ8RV81rtk5ahKQvu/V7i6PM1x4TugePnCXJU
AAo/DpAUhmaFoVi2hPCBmPgWfHr0h/VFXSi/qtW8C/zFjQjE2SuXOkbv7ZLx5sfuQWwEjUED8Ydt
eypFTgyLB3vIKXzHyB1t+kfOC+rmtWtGQKvEWGxw/4WaZHFKjKWBMyORXujag1UiAbeFJEUK9JLo
LRho9TuqrEPFOUpZaD8n9617nECkab8oKHsP7Z3touy/bz0oDLl+eOUwA4czo5m5q4m0xGzM2Ch1
gwr2TgVj33XfDQEwZvHw8EnDH1F13RYGLFz5DJlL3kdhPnZjTSkTOjhbftkENmMOSr7GG+WOZ9nV
7/9P2dLGnu/d9tOWMtS7+HSh7BKiKbzYsscififdX6B+LsLbDEwFrCTbEs1H0SC4MDcON56Vb6Qf
NtxdWgFSA+/4CujmjC+J9WI9+xs11lvzg4hTTITgdOSAm4VqokhALQgCbfpijL5zyR95jh/bJ9Xa
MJ63Kv5uODG35VyUsU9mMqyJPSuWbKJDtmYO316TjY3IdaT2eWfo3uVrfkKFvsc9E2juVCuPXa/u
JlclaxRf0DATasJygTre/2t8b8a/MjWOIZjv1PVWOrK7bBsJi0fZdMAMf3HMNzFqTa2dIOTIsewT
mTftaWw/m4g7dCMvMgyVQBukY1KGAXRyUlq6KwC8Qrum4ev+OYeEGy1PuJGkKQWmSjyFodOThxez
Qbnui4NtelCPhpDg6Wq9uze0tMOw0w9wj7fG1mnme6u18RXLEazL55dLh7ExewkLjo43hBEzSqYh
dbkz6N1boTNSHTVimnegB6udKiKbDSEZlSis6+cNMVMvR9KZGclu0+ZbMKh0TgY1xj+LyKj8sh8q
x+bvNfRA/HBiTcdC4JVy1ohrX0tPgTf8g3CbX0kn9CC0hXgO16CpnFLBt7JhQsFUFuVdNJxQ++97
ViMA2sO7z9laShpqFjbbXWlNKL082j00BVPIkI6ayxs7d4pVN/HSKKbrMhW9EVVO315YpJNFhOdj
t8o4N3n5LiZwRi01XzOVP8pYT08+5u/SE3rxj4A/kQ2Vl+SPu4iIqImy8hlKuUUqevCzMiQdRV/W
/Bwsc/bEUU/ZIyufe+NZ5TJFhBij+SUmD1I+3Rp9lZlv43SWGdGKAhlvOxBX2Nhx41mAwVsLfZ2P
LhTmbIjVvl9kUG3KBOsc4IhPQt0q6I3VUKWs/SDdEp4LVFIYDFp7FhJZ68Hykg0M+dMCK7tSn0LB
+5f90HL8zot8rNaOVVMq8FBDvgFMnYfM9h7NRKkRnl3bQjqCq0u0sQKBVDhDGwtTLqQrXPtg8E7z
kOd2XQRRAhBAkExPxz55T5zEr6F5x5EEuzlzLl1hDOC5AiQNoidObYfPRNLDWZnh6VHR6/mTNo75
a2++E2WJ6qy/zWufA5+SSFGQoxIPqD5m2A9BtWYqcZFApeClPyJHbbg9haqlJ2JbIZUu6EmMHZVv
bUUyzSvHsp5uyWvqoU1yNpcad9yP0tCoqxlnkswmu3zpHW1O5SRiZkF3muVD7dYH72v6SZWyhwzq
ySlSgE3CybFD7KtprsnedcAFTppcRXw4t1fLxNDaPBN+ZBKWWpHsoHqi72lCbQEFoGSbf/s/oYtR
IpHuOXSfi9kxPrDLo7fO7P9L+aNmEdtWIbrFW9UkV8W/RY/pK0YrHCFPA0S6ISYtLvmpVa8DNGj+
XdIdPH/UjuJPhFy7XA0bmbE/GzKCuuvLz32ZZIYmb1b8jdFDMFrMoe5/0yQ3HSdnrxvwRDvFr2sD
HD5H6/WKDpiGcdj19hTc88qA5OwzOcuyRT+uGrPzcvi7eRQKPtPDXVcNDao+6ZZBuPPTrkHq+akI
Pt2IFV9H/ZVc0II8uMGNnqQzQ+HCDR2M6y9CWYg4jXplt0gERfMNXrUKZLbrTFafj//bN/uoesfj
AeVk11o96oMpP1jz4YlDlJ/Am+eY9AuK4uT12g4NW7t58Y368UPzpBkqV7ke5hmHws2L/rP4X4xr
Vq6DOzQmGee5wXi6xuXrz9lc+qZF1H8RiW04blwpZetmNafZKXQAaQ0/TXjCKhqzM/dHWMzlQA2K
oDlH5VCrckienBgnd5ZsmezyhYCj7VQjPUcUV6g/zRRrRDq296cCc64oEHA8C2zyLGh9mNtIidrK
oPKrfuF4DaA5nByQ5GxXsrtBt6pXLLYicPONnNGF7T92XHpCY7Pvua86HkSmxY9n+QX9CmAgUHq1
np02Y4aEWwfXtdFJCNxNXFbRiZ5XEy+isO5RAYNgdC1wz5ePCuWqDo6USH4PsxQk1sb7fhKGX4DU
M/D7+6NOmtECXyconpoJRd/ttByIQi3oqZtJiUjNLAu2Z0pdO55mgC/fDrw64cdQt76N9FMsCZy5
fRRwFl9P5/tyjy4yC82C7rcsq8+NqSnVf7W1JQKzE0ZZUr3whZqJkCBPDAvVwhiZx8ES62pSsH4+
jw/rn0MN7SBJ2n8AERPHB7vbTY5sw51DsLjE1jn+OMjtArQRziZx6zSf5Rvh/swVEwc6VWNW/cQI
0LI1uXp9p7XqGNKjuYdTZG2ykSxzo8zlNgjBpkjJohhvlMcn/zPNAsTeZW+CmRndS7UuujlAzNp4
+5iVOVgsN5PiKnKjOunZa+P/A3x0uih1tJSi4TrxirsxnCKPsjyK8P8kQyV8R+J6cUn08fFhd15F
3zH/woil/0BE34gbsJDfnlnNAdBApvwySa3WfitI48fF51jXV89IeDEflelGWbBqrK779jdP3xw7
bcqEPC+AWvixSybz4flX6WeTN8y+srolg86EFBiIxeX8ZYxpV6wDFinFaxm6xa/vR/Q/O7YH+ZLj
QDTWDhqjhKWGixwf7W5n1ETjUFjQEqMyk5nVskC+3uitAta4+9y3H5zs8CivWePQtoYgWj70GzTz
beOKse6T56xw0X3LSZuuaJRd8+yxIKs/F+YycQju3bmMVU7hZysjuoeSVnOV4NY8NQqaMONvIzgq
Ike5OHIpf6RN5afAEjJYiY7CHVLoXjmDXz7lqIdtW0FBrnd7zzuXPSrxOEpE8+L0O8nUeL0oA6wC
Ve3ggNBHlWtgSB+foNeUULkq7oO9jpSjxGaml4RLF0PZxTtFuDkERj38v0wgNW6PMXQ0Co2pPSqb
GSiquj9mRMEll18uD0GTCf5akuTbRLaLCsRKMqh8THgIBaNkSQxSM/FNzFmD/wYpTJR8Ve89xmkm
39cX6GdJtPeUcReysOQbE7W+xV47t6UJA+8siDxqjq8ohxdwPffgoeGKmPL5my/SsWjTynt18bZ5
7BQqfAxINrZBJiGhr+ETQ0E4LL9MEjw6m2t54whY19YcUhUz7C1L6dQf3LvZsLHMPx6dELqRu8E+
PAx07cUwuJGwh0YgNsnCkm3tIz9nHCA4yBUdDD06PUTQ+IIOjeZfieNZaLxTvLDFZTQFu0wnIWBk
Li6hNL/xppP2goPQlcBD/+cCrcwAmjtJlDxNooO5NAc2NcPGxl4R2n/z0zuq2jjfKIUZb0OIk+5D
ViWwWDFM07TDmVIgvpwqEp88Qnx5cEJSCpmB2FnXjFA71Eatwohc7viIuWTEM7q1FzEsPemUAI/F
ZCBwXaQFnoMTcjeytWsL4VbVumb5EsSk4bkHgXNsg8zX21k3XLYKOss1Pbj0OAxT7cnrpF3LSy0O
iNhUQnEDeXSPj6eu7DjSGtjlvfXmkzmXRdXC+eF1lfjS+uyf6SLC9eDO5ahWRQ6IUsFIwb/CEkfd
Rb6aqrwra6ExsLmI9n2zzbIgn3MjrSGwToi2mzmgKXxKY17FsurltJ9b1y7TS2hnIAqiCfTW0iGc
BZBU7MBRLw/6sRmwTWgG8bO3Ahuf4yNc2QWlWgJSIbd09v0qauFB2AaojxughJM82SsoW1FfI0XY
DAok/5pepBB9kMCsdtgzMCqdKzxcSRx2PWH9z1IWolQ6vkUZs7vz0kLUxYv/sroPiBn1oPQzDq8O
W/ScBNaIn03UI1/TO9T/UOH7POAik/INs5xSNR/MhsxCTGmU9R29sY1IblrPN2v7uMolG/ITREE6
bIfXe3cmkXHxSjkBrqHUk5fpRyTb8jsoHvjTNUZM9+FWWM5EbyNhet2LYgZOVuEfKrS7rLA9MolL
M4aJlJqft7EP5pCwspfKrCZoJYz6GQgiYB8+jLHd4c9eUxUZSL2ZEjULezn3bho6SvEZyhsNBRKo
jgo1cLhzRRR81hlKKBfqytY05hAzqT32elgt4FqNTIOSNKaU41fHnIXqTRxSL3eV0s49QwkYu9he
SMLsjiNRvmbxXNf1d52Y6rEunmk9YG3gdoA0tcsMGsGCWwqqgQbGQXX6A0Z5ZSVUkveugLpsYTk3
WJMonNZUHB1x7EODHSnU0k9bHfdMG2Zou27XBnC+LeI8qMbI+cwJpJlvLUqZsgag4hM6BfpqcqNr
xRuqbwj8Fh9zgN7rfQ7nl+AbQhE2cRboMOqIeYYPtWj+s6zKbCHAR2yg/74EQ6anduY9M7VXGKTx
Q1lk6/kc+QEKE9pnxUiWiTcjWMO3EnZGuVI6YXtbkVB+kdOfoN4XNbG3GSKSXeMGHXhhV67UtWxG
Fev0tn1Eu5Gg6+qmzLeUR9lFfPWzolAWXeD/pqkc1mCYse+OYpf4OGo6ztBO5J5Ymh2jIdwZvZyW
/MvAL3AQxnSYepp3HtIR0Oi6lQDUVmzh8ITW9ioCh81M6aVLwCW5GXrlIuN6ze+VdJfkh5AXmFpk
SOf+SY9JGcVuz/Ge8UWvIdxa9chYw0IXynmuVDFC49wWRKkxOH/VTvPLADPEh4zcFGaLY9e5hGYu
4xE2S9lL5dwtJuMnc1FiGk7lJeig92OD9uADBfMagYp8Tl5sFPSVLYn104KLYjS3OZ5T3XDRa3FS
O4q36F+P/OyPhPp9pJUF0oAlk3YaL1f6l4J0sEkMbNK2ycEUa5P1cTCAEyoky5kPz5F4bBMBHhOJ
ZYL42+FppzWZOxD0zt7l3n1miq7OBoBYSVGM//FRADcpu/Ks89+hB1/qvNfzhuesei5W2nqayBoL
lpF24q2uWuiNOEiYAWOLyCP7v55j+6P/yVuOoHqse/9Ho08XYj6qWcK2pUvvEl0B2IwYKXR+iJuB
8u4VJo85JicIvnf5GZMDvRSYW/lEGFMLGKY6/ZMQ34p0tbW55Dv2Ykpn+01kHDNSY+XcU/2r+uzs
vVMb/NbJz7IPPvtfj9uiaqKGfA4cFTxMGwor/ILTyA1nlvQzMaLo8kfNXmEUOfoVM4kQqljwszvN
ftLfQnxaFUIX2YtrEMbVtOAWaucpZPO8F1xD8SoEADiNbffh2JmI+VaNQUTzKEYrdFko4LISWpAP
qV3QvFJJWbITqECrAEGq2FqByUYYMtJere73PcXQ2WfbdY8Pzte0Gf/+UkFCD/gLIEQ4ahiB5yDy
zh5k157GwIsKyRH2o+BLVtXpMzefUk48IHNH4rnidj5tYiNLvyZEtWgdWDB3vFjQHylzGmuWhor7
N/U15qEbnER9ASGksbcSIVNZit0/0Y6LoCfRB3FmX3AknJW1bkYtKDzK4ASlsLnQXEJ0UQsVt0tB
99IN3mxZnXWu8dRX/uz1CWMIn0my4UbM/QPzYX0nYCsEyjNvFV26p/hncIqh4HVDRF+cUDrl3R6r
Vkt47OseijLJRSz5jcP96+ALN26BdkLeqUbQf/LuXqiop56Z4zGPE0HriEM2JQ4OHqf6Y5ok1v5s
Ih4bE37LhgX8Neh3X4aWiAgs5qdxgkCJM2jEWZAZmTWEyuhUWXw9pqnZxuKmFgOHLUe2mshSdbkk
va6g5yC61BbK/9wBLDIpZ58s9rVlmZOTHyVQDSLXHAe/qJuanYCt37khQSPW8SxtCkm9PoeRBg1E
hOX7gltY7ycfIyaF4W8ajKkSnHXDe6AVGGldLH8OeH0/FveA9kRYLFuRZpCInfzVZb/zO4t941cw
n8Iwh1hlYX8FVXYlvDGnxTKc2qeEoONJArd+6LAFx27fjb4clR54qEAmLYbnrUxR35I8X3iwxvVt
QuwERVAmICICFMXaWuLxWXWOPtPI4/0Z0W5Gf9SHYPp6OW8DT11l6/vNZbNVxguXX5BQ/TOEoyDA
Pt+VblfwftP9E3NQ7bA1HnxOGjbc5KJX1nWO5pFBqz678oVhOoBNVTBWSsejKd6X0g1TCcPMGONk
lDgS+Hovu1ibxtQz5vguPkCi0VYqpE5y7ZJD8Oz2FSCqcNURAscMAvgn7hBIWOg1dhk2IpVFmmTz
tedKhISICN0z/u1E4910WwaEHiF+ykht+IXclDLuFL8MEb2EwkMK+yUXFAuRiKIS+36vxwA+VbvA
SIqYril9nYXyhEZhUMoQLBG49faqJfiIbJCd20BaIeE7Z45xSSLUyReNpqfqK/U9bWYVY+GH5TcX
V2MXxKn7vDIWywJEi3CrmVgTV075y7sHGkaBUgE2VwSGJs3m8me2CVEEv6rF8edzh+k9LwDRMMVl
trXqtRai7a1vCsB2DMfEMvKfIecV2I6j4sMRwAOYn4ma0uvN67NTk0Vjn4MbAhTUFeC8LjA/xDEb
ALsr8DfJa6b8a4v7i/tGGJrkzbnQYUncuHRr+n17kvjVvej1wnEDl6q4QhTYfrGGh2ilUmfzXJJh
R8F4vp+2ptpTlF6BKDuO2kbGjZ6fNcYw9NfSmgtMZDOVTuTnCiJ4mfSw3iV6MN+vDbMGrjaozDb4
JjyAqYr8PVD5MfZE/MBfT0CkZbfk+0E6wsuPglg/YpUGrwe5X1hyozaRi4jQRs9ZNcFPyPKlAGzN
QJBQYDWDWNAw6MAxMx3x3gvf89E55aEUTWYoD6DwlC1QilVbjHo9lwPbzDWoZYD4wb6TPQxR9vZ2
3cD2F8HbJAW7bGCoKR2k1F6PhEvKhDEcFxpIThbRnMjVVsJjcfuXEkGqSIyyM4zJ7boIW+yFXhlG
V4tSiJrJS4zf42dGEksfAF2FaEKNGWzMgpgTvDWY9RvFAkvDwFFWYfxvr/zV/P8mwwOtSfSsXBl0
YbfqPGwXzIKUQq9k5oAAcFPcG1wLuGq4QYipkZpUT3nEBQALewbU8zqLarAM8/K++L5SMO012u78
jo3iigDEJ/GIW742g4lr7IWsxMi8NpuQ3g1U/kGKZYhULtmEOYJY756phSddG2+VlH0kAeBSBbeQ
0b2iebKIT5T1Ko0Qg6fThY2B4Y8NVbIQIlD1KeAQ/tZRLXJreiLfRXvrFKnryw7SCDE2k2KOa3YH
Q+nNxy122V10hEYYs0qiwC8usXVU54p4sjXxnjONZSbMjca+7NnTpqessuWmpyGGnvxJJdNsO5YD
Q2OBA8h//v4p7gZ86XEL6MJkUfmvZj1ZCIVmXRyzkHdiQElwM0kCxxO4nLR7bIbv/em+HC6L8VC4
Ai3fhH9CRZ9aYB0PgsDdZOY1J5CephxGV3uvr2mQnIfI+Q8LQWmHMEV2MAlc0XZ3zYLJauh8+DyG
Vs5EIKGwJgAQYUAhxmYUCooWg3RLRrXueIdnmPphr1n+Pl82Q/BhhqkJ8dKL3EYfk79mHCoq9RQQ
6OjDW/w6PU7nwcv15aeOKUYQnTcKs5Uyod8BjK3Ezr9QpNFfzGWEz/tOPQC3gUA+iZFnT0CWjeS4
F0kTT1uOXCJot2yBIbuzPJVwHI3VqWe65gvKPpsjLemcgsb5dLD2WkOP7IU0HcvvB6RcdNCnUHrN
L8wVg6n9omiCRW0ZCCuOCvYkZlLpPqmC3djm8ymJR1+OQNSARWz9vgH/7/iyfAyoN4Gxy/QfqE6A
FchviM7SpQ3OXT1M+V1KnN9GiysKiJO2YZcCIep9JBFyug8eOFrezGzm7XcTqwsNMae0Wxvim1K+
dDmMH165hhPVS1zjYP190ORUr6zPOoniJ2pTQASg5+BT45cJw+O7fa1gFlLxjzrtDjPVCg3uVIcm
wwVvM5FN08cAopexbKSomgTi0dQfGuJIOWWRYPYMn3Bxu+956qfYqWfVER+5iIcTbwb1cSupJx0j
RTC7b75s8nq94oIAe64rUcEFeHskZOoMmp+27mbxTewIMbCDJDxCEELLUohTjFyVa//VLTPrlKrO
h6Rh0elBxIKF0+6DY+wZXAsTzBohuRWHjT51XXvJZGQY6oVFEuMtvPNtWh303nwjWEg/zy8rikqQ
J87nMQFcYqboGdn/hxwmeHSrTMh4YXacm/rUdoTgUjpXQ+9CwEoVgFto5M+KXG8jSqQMJIC5fvGO
7aojIhFM0GgHzywdiIEqgudDWAjLiCoOmlnpxAcTzzK2U4BIRE0cSaSCvkb9t1frX8PF3WI2cUc0
N8yUlgsOSNHO6eG44DdEIgJM+OrF7c1LmJ27RVrUTVyWWy7fMkIKbfum09JLfedXNqbJj0ytv4Rl
YzKmuXbworNpu8U9u2i3f+iOBBJvEzQiJaAvA69NnjSMp3TnKsPz8NqnREh8Ej0rcjolIpLINFuJ
njWF0rgeaA3AggIHI5v/7vd9zJ26l6EU6hizKfgBSXmPS79hhvbw+FIVvvqoxAO0t/b2f5YBrmO5
l6RK1euutH2QEpTwa9ugLJXAlbqooevRyV/KNHrdOvdqHnQcAuYoz6SdoZSiVjzhzGWXkR//c+eg
yNNVuFzb/rx7zThuB65ciJ4ADyLBKEFtQ1NeHSVD95rFlwzeAkVM4mfycmfKo3+/caavsMdUHn+N
pDclglEH1Z63cKrr9Ww5yZO9ghNdCBUPapwZyvnffKWJmtUItH4IJW79WlRZB3hdtj9GIyQKBiH1
ApK6+jlECy9r93t/aflRQee9TIU3AX13WP8ccGKzpr5D1y5P2wg/VGavq0QMvCLIjqRHKJrYbO2h
IwY08RBLADizG9ehhp02cUIW+Ref1A7WtEl/ZGxKHxebBpIyLVPmYjvPBODYT5tq6dZ82oLltdDc
BTGukyCmrDNvcr9SoowMHVpqlJqa8u9DRT1egoYIa/Dun3NBFNXS15lMZ8UTQI+XXNAXBnXej8QU
t1+ZtClU3jJKKQxu2iKBi4fHOrAoqf9m7u+gKqdIVSlauRAk/g+6tcsPaxfIas6ckW3t5yMyZdVi
CH5iVJIGq30bNZltWFYzj3z/4izbmIDhVOcn9KS+MhGZNDCT0Bnflh68Co0erfTodcJOtCPCB8uR
iVcWiArIluy1z+pJWE+C//TYFFIFmPLkm/WSs6xTSXZEkB3/tJpLWDezbyogxsobUkFtk8UyKs5U
rcWoX6GApPVLwN/Qcgukx3mnBGLVMUGVx8bcbjsjhsngL6+zxNIBaNu14/b+VF9bpIWJhU+dZsV6
DydtE6AnmR22x5mUYPIES8goFHnK4HEfiqEAeAcduJn9kn7Wfbs5xy63jGyNB+UkgdCJJUmyUVLi
qOe1aaq3St38ph8366X6mNozvt2+MiEhMaABJHgxRyBgT+xFPHoSgAZWNTcmFG9TjSFCRIu6A8ZQ
wipAmvGPl8Zp7B0Ac43sC2hRTdHfzGuH5LvIkQauSTVrnIOOb+9Po2tRl9a3gYeAOPKaKGMOUDut
W/CSz1wgR3Y1BfnIQ1P+RgPWCersbljW5rMvSkqOqsdX6mTSyVRkU3T3gLgGAntYEnWo0tSMTPAT
mWOO/I98fQI7Ikygylw2sXm2DNza9ifG7yqh3hoPeumXu7Hv5jBqkwi0X9BuuMAHMqXmDMhSvQX2
EhAXL7+0TfnJbTG3exeaJpGyAdZdUssuJm55lvAdxp+TSWXFVXSuX/Bbl1Fh9G65DsAyiNJLpEHO
u0FXyBkkVZJt3lM4ZtohMweGYVKIcxHowOfDpenK55uc1xg4sA0NUDYeDlSTBVByoP7tCsM7mxKN
OkjsINksEyt6/cUJFfZwB7SE4+2bsgpzHc8gvandH2aMfsBqAKahFru9Ci3orjNcGrD74e89Db8i
dWWEkKbCWdMRVuO2rqNy8TM6jMmX5as+3vwdfmmkTwKOgHtr5vYf+xeyEoCzeQV40cdFgqolI1Xd
JXeSO06RWEcm1g+L7JgCzET9GtjwzBawZMgREFjC2emRAxw0tf7OEe3L68i/53ew6M+vjjTARZ4O
VnF2E0OqPuWBK3ts3P+LFut8XINHwuJ2CxAwtfMEh9IWowMPRF3K6pyVje+1WLO5TwX+VMEZ6VuE
tuuYssLOp0tlDweQWBQS/OsPhoC1Jnwy7abcGZuRJKZz85xu63MZzwZn55frEPJ2VcoIQ8QFyiC8
o6OVTI2GlIWWIz5aGPxj+We2YHlSw3xeHKYcCURDJYIX98xYqhmMYsPy+Bos9yZBg0P2DX7r1uC2
WfRUUAjdzj35Kbtasq2vGn+nzMpWZeDH5ZdbtxgnJNVHbDK35uG7Tx1mBQcoKDcqim1si7MZLr/c
HRmYJ/goGmT98xP2xVLDxAMJV9o7m49izytFQex6VDaW/3rzt/6aiHKFnSCE+jfrvkdhMdcMA9CZ
kkVC0O2gjFjYNJStUi/ttBnBDOxcToOe7TcQE8/DBbiIrqlGV6g89cBaG5zG71sCkxw84DENbC2p
ZCcb0tuFOkvC+PaTlMvC9i//lluFnRlJPXtefvvxy/T64W6PBvkWXPfks5LEyQwfMFzYV8rUfyWk
39iIqjhvCuktA5YSLWIecCyA7hoW+UGaiapuwZEtiWtEykMHrDJePEKrGdEs8xD98UKYYj2SLypK
aA+2YDG4ArTV99mFDk/EPfRC2v0LiBWEVvAj7fJsvprcMtCjeXJdNGp+6E88210M7KVf8yYc39q+
dgettRDVvK1+H5p71Px8Xx9YQD2/CvZZBT6IVuGb5mckGwBCy9jSM4bJmAyXZsNu3nSQ8UuHLls/
9HFCePN1TB4sUD+pwqMecNj7d1MWvH4PoRNSwPUpBpk3so1Td7NGk/S6bogOaezkD0q9fwNpoZG9
mVB356rS72bojpbhwqg/hm2lGj4yLMoXXumxrDoL750oMOCpLNuaqVnguXJctE7ZxwEoTxX4oxzG
aF72kFh7yYZFqcLA8vf7Z2uPtMTbkAx23L2kd3dbNm2t0laHl9Kd69ah+TwZgt05ajRV1mu7R3Ns
kh+iiypw6ZitTgYa+GrxDUSp5IeIPgYxHOyZ6LohWyk6HyEj0zZe4Lc6RUF/HQboTlGWF+pWt710
RReGKu4tc1znEGTSYD15kr5USKrEAkRR28vTS9vrrhKzfA+I0QyTuVK6vn56Df/qcdRQUhNen6Pk
/yL0SeJGmo1l5lt2CB0cJQn1I8lZW8PApNI5qf8HYkXmVePMmbJSKFG723HsvrS+ipA3sGK96azj
cclJ+ba0ZJCgoewgsO7DyBqYFJ26x6kBAkq2hjLCq3BaZfxVOpkS/LuBHx5uALCxVW8jJ1Ux3GGJ
aFmRJPdOhNqTjSHgm+LhBWH9jShqHhei9ZDhJLej3K3WihKOtz9bJ4EiTnd27yKmGk3TG0qBOCu/
zH7mhdEotKDOHtxbVCuJb1rZobAAIXFIiBkJ5Wj6MNbAPum2p5pGHdcSZmrZlZqd+qApIN4LpJVJ
CkpxQwnfae6q+Hk3GwMb9bH81S1OuDKSDo9x7aXJcXW4h4W4YSu+Zqt+K9B4ztVTdthNvDVSEswI
qZHO/w+ZufS1IREzMiWhhx6t8nXj+VbYx7sHlOqkE975Os119aEARqaCxUvLNNwDIU7UQ8tP9WbD
co4aHKhtDwO6uB3kfeGF6QE5sXSeq/YsI11Td+jN1ApxG6IIp4KM4A3YUnGhux/SC3DKKqUiHhqo
zB4v9lwXVJBmtnaCmwuYvLrhjNU0Sfgjj37Qi/GS5I1SbEmPgZn9rT1JvHTHZayEHzEF9ssY+lIy
FATDAUn9XxSr8d8b3K6GbQqR0XWDVSqKBmVIxoEkc4MgDPLMtVXZtkaq+82yIbL6EIJTHqsy4F/B
kBmZjSMONnb2addLr17m9iI2W+LFbY2S326FOjY3NTRlmYU23mJdcTggXSsqXcvl5wQ1jp3godQc
LxR+TxK4elYgoBJIYhrznncGsFcD+Duj7C1Q7kM08aSSEI1+geSVPlg/m7935Oc3rD23VdB6tgMJ
zUR4fbk8qK9BcEw6AlHUOfDgAwnPU/n+SfSMaO0ps0u1pwGKBaf4TJZAsdRsEhmnPJSq+dSG5egi
XlyqPkJs0W3bpAkiK5MNPU+YcsWFWEDsmdD0KdC5X8LddSmyVqJ1/uT+yIGb9R15QGpLLbE7QnRX
X6XIdB52K9zKHjRrzdHnISG3djJj5FqfhYO/ji6jGu9LMpqlEAXFkUikzFeif7dR/6Ce5kUm9LIo
zB2/isBeX0BxHPBjmQF3g+jOF5jpXRqWWWBFKwWu7ivW1TI6k/QGhBMw93NaSVoyWz3/L3ElQbaQ
8DANz07b439IaXqvyz69rI1M6u/x4qebdi5bZz52029tz+3Mn9OWbzqHvIFJ/hCfJvWmEezjCegx
eRpdrVuFCm0gz1FQWsHj7b259Q2qYFD8vSnnDnoy/URbqGgjPtExgF+YrWNXFQBtqezooR6Pz+VX
OtM5Mo2nTq1R/M3SS+veX8zCeAycVoJjbwhhyva7omZrIL5Nm3O5inVLCVJ6966Qc/CLxRiIe6h2
T9r3JqQVCWqpXom4R6075zXfsaoBEvUyfhNlk2V2jvOl9s/KeYXQyJyAmREpp/jb4I4QiD0ecnKV
CVTGEdMoELRRsy258pYeTefwo6V12ZbC8w23mSIJYH3aHjSG9efQdIBwnqINyr023NvboXrY4GXu
2/0w4k5VhYSdAmnheUP6WU67XJ9yhrxUg2186R7ATqikvk9kaOSX69QwoQeKpu5kEfPNKUNlP1eV
Palh4P5GQy6MbkrrSxNhpaqK8F/CIW5ZS8fUyLKk6gZXDz9ENEkE0Tn6XnAcCFoDRqMvO2RxvmVz
cha0ryAbf00DfSyMP2CPFcDRmDR9pRhZWAPwVymaDNiZBiYSyjwx5RxPIIYkeM/MaO/wLmYiCVIH
8IcZLa4pLaO7HKgvkFQMw5wKMVTPl9xfAKy1IO21KAfZ3QTqsKfTNPakgnOYUAoYmtBespT8/2oa
ca4QiULOoZw6ukWVDJKyoVu14fANlKY6SSLpHYd4vWPwI6ZkmlhwH6OORcTl7ptlObLf8G60YzK6
EqyptyMz8bz3RdrnMge7P4AhSWEPhwDkAo3s08Oi6dYiWKMn+FMksS1ACJRLe2OTjUffGpVQQrM6
mNCXV0ICY0zU0RA2ErEBy0iF3QL7R4fBfs1Mtv9vB0KYvECmFdr7GjWuCyhG+kXjTnX7NhJ7ZHZz
R9KijT/MUUG8+DrrTxFv/SX5H78h5kmfYWfrpJdasiqFdIizuW1DACuhDiQDbnS/6A88sWV7rqo8
iHajOCkLtpdzR4RdwykY0+6ppgDY2jdZC2TX44LE/M2SjVMAK7dL5adRb7zFPNPXhyCiQ/rTp4yh
7PxD1qgKfdPAs9hEr6RgO9ZvhLxX1cBzYjBRKv5PBfZ+ms0dMtwQBu5VwaDWMJmDi7aNZZz3OaJF
8adIgP1JkTIccmzzE+XfPaF2t5RKY2VTmir/w/0Yj09RS5o6gTIdDrk5wswxO4aL5SqH4lP51Sxu
XhzTsV+y9QX7Htw0RWJMW2S+v+xLL9IQQ/hGQUthoYHltP09cPa7wWWVA4mlrKoZQOiiiWa38g/8
QVQRSiC+L0QPQSARbWEa5OlTTKTVUGEgzFOV0WmfP2dfKSWG650G3aPPEyQvRdruYys9e/Mte/Qj
PKw9FQrhigqWVfDbtENb5gTr8QP/V/wRT3MbC3YtOpAAIfdRhQrCpvHW6io+8Iqjn5cmnv+pbZtY
95G6MCtx99apP+/LAuR7iVjoeO9WT4Cc0nampqEj19aG05EUZ2aDCvOIjq2HTe//qZeaJs1pggeP
lk52UIg0tPxrM4J8rHf/npkLugX7eYRllpQ2LP3+Q+x4M89022LXE6GYPYzMMda4U06zGex/L5RK
Qasdegzg3fMZlJmGhHOyPuKOznP04qmK7nTC1SOX25NSnDoJqMV5+t7XfP8rkn8qTpRjbSY8ajN0
v6f6khuUvfErFdkPkTHHdKMxsUZZI734JjJIiqj3Gl8O9f8a/uaq8gwFqWgnxA5sIffvkEnDF6NG
ZxTRW58fZ+/gaCkcSKV3Bro9g5ImUMNXa4Qmy//wpsS7oh+RKUFytSJDuo7TKEzqHlAGmhRs46U0
GDICEEnhvclKqptncBGeSvEXmBUcK0z9l1FL11raf/5HfpqbL1AohsC4q7DzfKkszQ7yrFAjT9Pt
G6soiuVBFs+b28+p/rEzpV9U52eojABi31Pk0f4UK8BtYB1sPNX7lHTJbWqhYXnI0lNyaJG29dy8
2FySJQhoi013EfFFkNClXoEVU+h7ZJvUbOGmnAqpNsuNMbqLuh2da3X9Ptk1HMtOVGfWTDlK2oCt
SDI5hhmXOjWLnqtOslLw9NJ/+6C3IMGnIIAL2KE1ndg3qv+iwEHIUFVrQ4CwqVySYcybqazv6uTv
AXSN+lTa3kmYN6XfJtgU1cDKeEFsE9qwHsNhzafVz2zN59C459Z8kS3TTMmZ56HOM6OJPOI3024B
vz0tfb5DtbmGRmF8pbSSss/E52JTPaGvQlbPnaEbMKMSEuSA063uWoTk9x2ajnDnRBZERkgz7hPJ
KbEnYFdZLjtpWdrzTy56CciEKqJYTQ/TOaB9ydKUJv8eGenE6gZNO29RqevQcDPu7rlaElIYbQ2Q
X4yS6QK4WmuhTJVlA65AvsecsyWcjZTnYH4t9CJTBOdtHY+aBuK0rZwXOeKwnuSdajtrNn7CN4Mi
GpLiyfXJd5m8942oiDe70s/8LuqxR8IUBljzNIz+DSjALAQirT9+DUmRg18UAa3UrFCKDzFxfg1k
YL3AltgBaCcfIQqZKeybUxnMrAhCb7w3yaNCSfO01LqHSRh5VBX6ryXVjJffaaXdcaTzUYMocVYV
gS9voOGtYiE/wYLga2pKTAvRqkiHpUpntoRzWFzcyFCqK9gQ9QJi7J8xYO8CKoJBQSl9gcLd7Bj1
2Vsl7Edd8fYbKgOXoWwJ3QlOxHVkj7tsx59aU5f4ZCZKNbj08JYAOtxlQgKRCpz/E+i/ocTEHSqe
5BzZeF6YDMUvrhAaxv8KQ6R0ERAwCZ8OrsH63tpGwQMUjuVAATrLl7IViTGpKxyUy+QbEFpypHAl
zpBR17CUIlXQlcpSjdjc+9CZGYXesTJyLFBWoPfb62EeVQuLJ7pf0I9Yg5McH+mOcNrTzuPzgiLG
MLfYtrpSBcScIXklqJn5I0re9it8a9pCWtcnbqXaS08oZt5x13G1yYROl7Yh4k8xt0d6wh13LDuO
258C0vOS3uQ//4neye+z+H4kJ5m8dNrsr7Ljyus6vZhQrueUwfGC5BAXrYSmrOuDpG5J9wFqdLqF
TrpBJ0FnMpBRb0xK5LqkK2pJFL0VhtVnHcEEEhscrPCTgI4O6WXXq9G0OVbms+jUP7R+d2qmB4JR
l7IXhStdt18mhwlf6zGYyYPiaOdxOOUIGK4IquOgZ86cwpJkzXWjIVcHw3/xxhndDx0Jq1UMrWSu
j9SHNePzItES9HWo867iVyWq1x8Q6Gw2qQet71ubLLIiVCk/uXtKJRwQ+FJu1SheY8VC7KuqCbPa
468GlD/ytl22UrDCxTY8FNa54Sih6Mg2WZqIBxYdEpL9mv3peZHymBnXHsZPvYu+MdZ8Zhi2NxlX
Io4dZEf8vIvSZqadZnxPA/AMfxGqib0AhhmdSpcQTbO9HEApV3qwGjz11VuaR8TIvVCYT4SlGSM/
zDggrJ2nt8zkTl9yZATunSw5LQQojaWt0B0dtwuOHHlh+PKbmg/AetsFjfqbrs1dY4DO/yW2hOhK
l54SPYioj9oqQ6SOhGiUWG5WG12AlyKszhYDZVkoY3/EPeRN7r1qEapGEsqFZ/h3uZrwj7KLKo25
ZYq+2BBQJzEm/cj5NOlYeGmHEiIh0rCGBvMhwamfajgJNSCdgx9SEoIdc41kKKt1quBHwxjnLTGS
RI6g2cUUrbjvF5Pw1xdDS+eIL8Ku+WVTonvOXfg31cK9S4iFZmQClQPmPIeH1RZ2zB03PiexaDKR
ht7izAm2frA2kYAiQuftLGbR4mMmF2Izjit4jq7OGd/+owvKac1kcJw2QVi7QDgd1qOzUwvrAcCX
Z5HOieYETYV4+fpu7Gqiw5jbAXrCneJ4A5V2SSYlN5Mf1VpINHnHzGndPg7J+vxQydyWgg07dhGR
8p4zD7ovyviLvJDwq/9I5x94gpafsLI4getobiCgyymv2d6Zvxiy18d9LAnN5zemoqUmwiBu4iOX
Su9x7B2YJbGqRK/UkzugVll+mf1Zgg8ncu9W/DoRhIgM3GFus/3w8v9EC6vFlAOY0r6J6IEB1+3X
HyI2Fr9gq1HroMKxARiY36/zcaDEM1pngz8hAl75INhRQQkY1gV9touBRZWTxpIbIAHvHh9lnwGh
BLGjoV/XM6lpVCECGpxdOxiqGQaa8GOOWPmbCTAiMS0Ljb1InX22Ek7CQ/MZ+ujA2b12BplmeOi/
ehEN2W2aQLPJVDjwZuOF1k/jpUDiBUToigsxPaHLvW40lHJc1tfLq9sA2ttR4hXmEF8UE8PE7TYy
LWgbXCmtSjuIDogPmw9JaGU+3PTeESNgIE07EVuAlJVArXEPqWzQKGF4vuDJ1GFaDavkhByjXGlv
VxfWRfUsiVl0BHfFVHNsgt6tTyxV/7pniX8i+rV1pjTdpbQA10r9796ssvCB2J4cMBUNe5kMoV6n
+1pGTf4M4IA2HItkdvHh6fKwiK2mwkdpIDz/6Nu6VznFnc0CDETyq3bEYqtNRfDg0CZbUjNNFnjj
VwddSfS4l0qMSdWiFCEuZv5xH7uIEQGLjyfS0YdjRWezNfbFQCljh6GxGSNr9mmjxzzgEP9QCwyQ
D/p3OfDWMl4oscy3C+//UzfV4nnYMOgVu4htjAUdq/ZKsl0E4fUITJMyrSk+qDxAovLb+DX24zwx
mfl3XYi7DgHAYH4mJqaT9rw5QP7Jot7VxWOPLtIiMVIAfBdogNIIjl8dQqei+M/znVOYQ0wXkOf8
9kNnhdjRJHYaFJleb07zC0Xv1yMnzFkupVluIfD+f2cnUS4+n9BUcR3Xl6e0ALiyf5QiW/xhy7k5
5aQhZl9fwXn7ZBL5GtcDR057K1xQ0W9RLHbYhGlilNJWE158S2DH2/S4l//S94a44SQkUkQc2R14
UGKgT220XfuxYNAfirtRBj1h8v3irP7xiwdKGuA00eO69cAC4A/aLXBawC7g6sbFp9aEPAjEOLEy
Tn5GkXKnRh1drb7lwVpdVs7hCBredgrjKI/ApoibwAIBRT3I1289yechuG4Dys0iAcPI1HRjjljD
O1srr1+KGUV6CurG0u+xiZJma55wMhlRzYzLajQjL9Tvq+sE9MnwiT2l6h/dzrorGgAUEFlMSbyc
mCO+3SAgV6YAZ2liV5tB1a3DYydQXTAHQBkcsjuVB2Lqq+fvEsRkXORkNzZahkrRWYtIRiN/VM6j
uc4fP4+br3Y15o2Wf0h7homQFgugPk22QSY2xCZNf+kdZRa6K6MehOGKORi/aEY+Go813ZYa7eke
QTLPBT9dmLH/CTjAgGjyf9KQ+HW2yUnIpCEEb+fshDTItjJD9UhO+tW4UY9CazEOt8dcJKNkS2ma
du0IhUsJ+HZ+MV+zXEHPPIWPsBV068Pevd16Tqrlb/p0I3w5CXVWkFn2fyb9PtWftKaU/zsnMlAc
8I3knP6HA+CzLGAnz5RuOAUytK4P3YAxxQdgqPGRDpjBJaXj7rCbNVWQrPaE5aBzyww6XvgodtiX
MAz0X3nJdXeai3zjuF0ue7fCVJaUB9ZL4gdIw2r9kv074EHBc805MijzC9jdjaxQ+YjkdnaAZYcX
2vaLBwvZtj4crkTAeesEcekI8tDL1qnx3aEuwgyZISlFebsdZr/IPf05Tdz5B789+keO/thI1M2e
EouDOTxJDweqLQ3N7ASul2CEJwNGWL8zy3Vtg+Tpnlxg1Ypuhe3KHtDruDNwUsqSjpNM+CnLYSOi
MpQV4GeAk01Hch07KZ0Acr5DwU6kjb6W3cOJG4L9NiD0236Amifa6JjGrtteeaSBVs8e13rcwQbJ
b81gMDWYCWnO+2kNA7qZJQrAUiIQvupG6fvl7ZtQUongjUR6t9s+Z38MF4RcQLKziN0RpqAZXg3E
yLxHYTxYILF2rOhSGZ4NT3Nzws72mBLbAxw8f09x2V5MK9BQJRHhRaBqX0eixDKOGyVMT0LFe4cv
0NLEpB3W45iw+cZ55nziSLI71gZpmKrQ/K8VVDNIF9ZEUmf7vCg/Ki52THZEcFAaj+3wRaDcRY3m
P6Lh1QlJ0duuVGBxkF22Fypio/otYLwqt6vda8lV+cgRMIE3/Ho/a9Qe4osOBCGIqO0QIG6M4gFY
mJNa6I4wA/LDn8bP16DXnCZ26GSiiTeYy2+CWYtHFO7enDBOlY1BHq0VR97lZNWqnAHKW6XB++DK
d779viIsw8N6XEWeQ1XSntygK7VCC2dOHs5XCSrE9yknZrd5si4iJRSxdOY8EM7V/VX+TliqF4pT
9PGfIpfjlpObYAUwylJYh43NIIeZYpaCRRQLmFoBDCs4f/JPBA7VbD3osU+UeUrtcg0tJsJdHBki
8UVjotHzSIBH+VvQcG2g2EOQFZgraB6bzW157bi4I+6NnPnaa8fBz3evgf0/BW3KFRCLrUKbfdDa
QNchJZayLD4eKn3JWiFL7+hQYE0bTkhMLFiYHDtmZnCngWaxz1KiWO4W5j621+wkDO/nXH6dUxm6
TgQQYtxPyw7GjInYe1/eqqhK3j4D/MdwXIWGXADbRU2jKOZeTfcbBYe7CQj22ajqgz4AF1AGFZGk
pGMeFshSqICZfhz8DRXR/YWbgnmuUJPSVE6gEp+NcDRBxTtLMTeWbFmONoTwLAxJPp5cfx8U/Hgj
co2gaCwkMg5sTYb0nBzYE4qeyBQIdquv1M857/nryRKuU0jtnEiu4BVETDhpH2BWqzgWf0PbYfsW
TazPMkpUhLb9Lb6hr03PPcrdvEoQA6WPw5iaNq6ilAmhPospMtELRkJVjNV0Vyna9SlwsSkTtSI9
ldXTTxiNBe1rb7BqLacmhvkbo01MSVShxLeU5b4ovkFcCle73LEgvD6B9mnku89KVOYxrrYyK2di
M04WadGwXYO5H5a9IDMZa1vtL5lzgzIz/oRWxvaSpmU2cRQyKQ/oIQWrzh8oKCMdIs9htlRHZtql
Tf/fdi4xHeuq8gtY/Jc9tkjGA1pAy0lVwEW61wqSlYsELiGAi56KFSOI4hMKmnBTaX1TBijnKuic
612qqnfnvx2a
`protect end_protected
