��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g�҃�f	��m�T���ƌ��"�C#~������VMb#�X�f�����|b���e���rQs��~����2����؋��&���K��٣�M�*�h��9�1��̻����d5!`�S�o����@Η�I�]���<N�����%F����0�8k<��~$��~!~��dV�Tm���s�@����Zl�U|{G�-?ҡ�(�K�ll9:߷dW��'!��ܗ��W��w�#W�q��ܬ���ݓ��Qy(%8jZ��{5�k.X*g���zۿ�@��S�k�!��������e;�����l9�&�V�����(�0mJo"PE������ט�w�.��e`������I��n��ӯ`���� q�l��e�A��y��˴�l�Ⱦ���g�Z����ބ��:�e��RrE^��'�9�:�qٶ��_e��cB"�l����s�TG��D \4�~������oRO�~�3V�]��*<�L{H��A�	��i3��B�Lh%!�!_�/fcA��yp�!�h����(�� %���'����*v"���D�R�������ΚW�o붑�2R�$�~IGZ�A�P��Y��#��Jo4oS���zZ�m0���Dyw����(��p1�Z��>;��~���5E@�囃��9Q	)?���Ů�ه!Qz;���)�X���[�|�� �a��s{C������k��B������-������k������W��d��G���]?�XP�����?�-���j�c
"~�O�KJr&O���}\W�7���0�q�j?��A@�C,�h�{���V�5��g�ۂ��$��S�Z0�m���a�+k1H@����0(��Z7��UMh[@5��}�Pt�s0(��v�e&����XgD{"����*�d�"stR���tx{	L�7�������'�����؎S|�r ��Rs��-FÓ�w�W-r��0�����&����]��H��?��R��Q����K�����A�{ټ��.��-�x:1>"�Տ�հ�<��D�9��^'ԛ����_oI�h1�O-��UR(H%[�N��Ĩnoq��e|�,S-���m�\�o�#�)�^�Jf�c����,�XK2��E��(�Qy�1E	�i��+]�! ����|�g�փ��eX�vVz�(��a��oc�.�j@�L��A�-	�~�A��a�����>�7Ltg�h�xꌒZ�[	�H����<P���#���щ	�$}�b�afV R�F0��"�1��j�#�,��*~n�U�x��G��/�[�X�B��ư\�f4p���d����}R!A�B�M�TWA_Yj�;?\`���h>dޖN͟r}wס�Mƥ�~��s��q���̑א��$��;E1=tAD�{H*]%I�P���x�{d�*��jd���������bcNЈ�3�=J������c�TR�%b`@���]:o���d�K!���E��6���J�<PW�A���nm�鲻���Zؔ[#2���9�V�Ʉ�p�xB����~m�d�)y�GX!�F:�t{���'�����_�6��L��᥼fͯ����e��f�n_5Ǘ�rfSbZԭs
��9��V���)/"�to�x�	':EF����q�H���fEV�=F�V]>Ｌ"Yf_�f6�� �è��ÜK0^f���1�0�f�ܦ[����y��8���i���93��?�Q��Kz�1n�8g"F�fB��^�uTD@�˥Ȉ�~��ӯ�i@	3v������P+$V!w�oɗ�����f�������1�>�>\��33�y�OU�uͤ�TT">��1}x�Z�*�ȱ3��-�@��+x6칆�>��3��,�/�nqw?���xx�nx�W��/D�I��v��
���T�딻1N~��/�NF�8 ��2@̏�����E��8� j3|]A�ߚE<��)9�����[��oD�øuM��R8?:�8aɛ��R^��a	E�Ʈ�	,nMu������`E�cxg�u�AKC:��"��{S�#yĞcѤ:�z��,f"l�t�g�$$��[໖ʬfC�N9�*|d1!�����MĪd��2���}����)��#�*�� [�%���Dk˞�M�u�:��@�ō��II\>6{�'���v��z���cAR�,�y�A�QW	[c��J�(�ź&I�͊u'D��xM��)��$�&xO�%��=��R���'����#�����NCo6Gn��?���zīqxz��0��i�[�T·��@��aOZ�F�N���&�nΓ�P� ։,�}�~��{�5�g�=�'�~(�	��XD��Ϙ�K�����y�,��2z�hO.!�uZ�Kj��w�45�^�%�B�+����Ӎ���r�1R�s�Rq�A���K�H%�>����j�C��`&��i�H�O�/��`���P��|RR�h���� >�w����!|0��urf~�wvŨ;�2s�
�6�Y���p��M����m�d�0xPI��^�����Tw��9I����`���Z�J�:���8�\�_X4[w�5���H���ތ`^��l����m�W�"V�^8�.@Ca�����
.eCtB���,�.��4X�2G(	ma&�xJv�����Ѧ?�/BqQ�6~�/�D��f)�ve-VH������~�Ev\=�Bꛓ�;������~��<!/�AT�k���ό�E�$=�ǅT�;)��[1�9;[u�_�U�J�l.��u�>����}�K�.��3:���ߺj��)"�6,c�r��Ġ�1]	V`�	�t_T�#�����$Q��A\��#jx�Vd�m��#v�.h�2�Wܗ�e@
�&�>R�t)y� 7Z�44 Q���g�HBi�4x�s��&G��/�l���W�R���`�>r/>�b��E+m@�ʐE�̫n����_y�bS��`�">\CE�J�����YJ%������ح�E�$\fV�ϋQFx\�u�0~��.g�J6>��7F����?Z�pT��������O��d�4���v�o�Z]W��Jtf�Rd���ؿ��,�8��,���$��|�=�b�4G,�pP�{W�
O��P���xn|>;�i�-���Wޟ��t%�E�Ƴ�O
����$~t�D�ټ����d�X�C��،Y�pW��DԤ�Eu����/_
�LyX�̓U<m�nw<o#���YR��$�QN�� �2��4�&S!'�_)@!S�&f�np���w�#�F��l�ul��A�'��k��Ck�M	lc��x��ѤG��)��eb�e
	��&���L��I����\��_͠��ouJv6��xy�VX�d`y���o�P�O��j%Z��/�@�T��Rg���抉���+�LΨ'���h�E���?hJa��u�0��x����=;L~]*MLa!x�p/���P��(1�a�}m��R}s����ʉ�ܝTʁ8?߫�@��@�N�.�I�K���Ud0�=AI�Ƃ���uf���K�lXߣFU��ô$��%�ʶ�>��K�|���fU3��6��&-^���g�i�ƕ�?�h��a����)u?�*IK��}��BL�*3�:��/h��{�u��3L/��7.i�ҕ'<G�"�h�<��Ζ��+#FHy~qpw���WE����������Bb��ڢ�g�mf�X͉���ɐ|*��_��NE�f���[g� b-	�_�CSx���F�$$�����|�q��� ,�l��o�B���c���N�B2|j�9�13�l��6��)	,*xDMw-� ��S��XB4\䚈�>��R��)��p��1^H������&{�`A�n��<��Q
a�$��Z=�Bd[�[��J4hC���s�}YDq`B/��Q`����1���Y�ϓw	����Yp�;�h����G�އP�e��[�*�G����zm}��ֲ.�=�C�b[j@���Ρ>���.�1F�^Q8"��)oB�,2��,�������`��>9���^�8D�ԈZ�&#vP�����f�\�7+.RˋZ	��<��Q�5�ݨ,@���PZ��s�C/{�c�9�� y���h���G+FG�R�j��D��s!��h�e0;��c5�Da��B�e'i��DU�<���v��ѧ�mHs zĨh�bi����׍���%�,�'w�I�r�lDc�
�	�th�7�O�'^
��w���I�b���L��(���-I��o�
������~�o���jEC�?Q'{_��7����>��.�e�XT�_|����� �/z?I?3��bX`�(�H@o|h�������r������@*ĥhڧ�®F���Ӿlѷ�10O��I���	z���/zmZ���8*>pJܠ��j�1����3c��j�վ�W���qM��g�&u���i��t1pCY� ��ڤ�m���'�n!�P���e��$^-���Q����w<��a1{�o��k�uH�ZrSΫ��`;TL  ?��E�q�/3gǯx�g(wN�J	1)����z�D92Q�#�	�ɅO���&�E똺@�l!���D�y�#)j%u�^���	f���x����f���4�#~$�w&F���-����"0I�&{��1��$�����
�}����'IA��_  }�����k�(���F_/�D}	�liDOS0w'�e�g=��A8�R�A���۫���p��d�O�3��􈭖a="�ұ��� J1�g8]nL��*����$�!�Fc�$o�·��v�+J(ʋ��9yx��4�Z.4���|�;�.�!�9o��SE4��`�s�Ag�@$t���u�N7�8Ն��{��a*B�9��e��m��~���ͪ��JNf�hC��?���Ѧ=YN\���ql%��o䉉�,��2�{VM�A��W�H� ��uԉG�Qw7+����5�a��w��GV:���j%Y��7�ħR�U<C�[���
A(�A`a"L��No=�}G:�9H��Ž�
ih��
����_�?a�m�@EDL�c��o_��Q�(�*�xp��P��b�Y�����5��h���e�wK����RF��6F�(®C���_����^��IN?<�ҕ1��R7z�硒,{8�xW�1��q��,#�c��𑞞M٭?��k�X����Wܛ>�xP�٤zT��{B��%��}��I~~³����D��0>OE�	�����K��w��4_?��͗d���2dky�QkM��]C�!��!��(J�G�C@?U�%!� %�!��SJ�e�(��K1;�٤����y���0i�$�/�R�����$��Ruz�f+ڎq��Y[���MF��kC00X�D<�0�c�� 7�u��y듇�&��j�2ث�l`�"�ryB����� �9���`�9q��+�T4�����ב4��0��㵽�b��ݪ7�XI�d!����a��F�-b̉\H �|�f(#����<����K8�_��|	���`�9P���+"cNY���*P�֐
r�?�)L&��X���a��b{�2tϡg�F�����9P�Rx� Iۑd/����h�O�!ω'(�f��(E������ 3^�k��=̫��۽G��*�j�z�>:��es�1!I �{��+������L�?̡�C�]�j�����sz�ڣ�K'�;n�VJ{�a�Ψ��)�m��a���5��'@�!�W-t��j�|�H�n My�����?
�=7��H����B�$�oj�;�����̅���[o��ۏ����Y�_���Bx��t�#��/�P�i��0V���>m�/J���Z�=A1�y���C/�T�n#s��/����=���5��g�5�����y�hqZb߹b�t��TJ甕B�m��+��V%�s��û �tl@n�*	r�C�
�b[��(�]&��|̑�{\�
��j�w_��gmH�T��l��� Z��PyYZ���`��ֆ��yƖ�^�cJ����^���B���N>ͭfz˦��
��X]��es^Հǡ����fea�����uQy������7���>�k�������K !��F��d��"��;<��ȷ�4�9�g�k=F�c#+"����e���6�jn���#��hH�q*�=�t��pК��RP�7��Sm�V�g�dr�"G��Χp{칀苣U�����F>z���qj�����x��1h���2�Z���k&e�7ޗ{�Ma�����0���TW���)�틈��qS���ϔlS<lnl�ko������x��_D�������W�M$1�/X��hx���or�\'Kj���� �� �H�q=#�@�a���%Ok� }�߆��c��K�"����٧}�I��	�oyT����E�3�Ӷ #ߡ�|�c�E~aena���.7��n��y����Q��$Y��brYz��D�)�;�	��*y� ��!��+H�U�}WpJTĪN����"���G�mCi1��h��� �^�d����[�"�����I�л2���;^�7t3- ļ�c+�`QP
)֖믺�ລ�_��)�orP._b�CѲ˿�v=,�"�ܘ&��
�iǊTK����j��@gh���5�(]_�"b[�*KۜR����U���x��ַxǹhH�.Vg�:_n�q鼶_:/��O�'i.v#0�E�n��H+J��/��[��R˗̆�
o����-�A��}7�7�J2�ѓeK�=w�e|��5�(���+�䂸� d��Hxߠ�������Ǆ�y�2�%��e��A��%�[�7�se"bO�.�u�x �MN�h%���=�Q:�J�ɵ%c���Q��)ڼ���}����2-Y�s�p��7�W�A�
�Ɗ��^a�N����� Dn�L�4�S �,�l���YB��-gCM���d!��E�m/Ix�'�R����MI�����8\k��YJ�Ӛ62E0�A�G�7���1���"�/� �~mNgmUE�Xj����	5�L�Zo	�#S+=��%�[ȱdI�o�9⿑�^SW��/Y(��g'�����,����Z��ק3R |VˠsR�I���&�̜/`5!���"��-�%��0X���u���f�뾕�rm�G�ƭ���"+u�OOA9n����Q��@�s��D���fN�CF"o�2�Q'�#���A��㯩/	@�0��c*S�>B�1fg7`'<�W��T��ϳ��{�l
ן̓~�ɼ'��e�U�54L�2�-�rbo�ټ���Z ��D�i�`yL�3�R�<~ �����(�W96fm��|.0��/c �z���me�%	�$!����U�9H`�r{Y�-<z30�j��b��"�+N�U�0��J�pT�?my���z�&�Ʒ=W�;��W�ŀ��Mh�`L�^����$-�=j�yT�(E����B�*v	�N�uXܶ�e��7P�6���Ij��?y�!�#�#N���zЫ*������L+���o�E�6-N��`3����������(��4���qKۚO�6�R��9�����m[�D�\i(�'y��0��GͲ��j�m�P��;0K�=O�+zK��`K��DY�\C��ě̛Q2�2�/����=�)�]�8R�����W�}r��������e!�����[`�o)r��|�T�P�����i
)����K�_�d�
	���@T.��X��MD���Dy��u�������\�U�(�5C�i�ܵ������w�o*޻m�K*����5�d�ō-�V@�@�y��JF���B��8jj�I��G�";�&@�tG~�EO�]|f������d������mtƼ&愷�ky �l�nR�+���q�o�\�f*�t{�i���"�5
��M���5A�/"<،�M���=��6M���gh�C޷�r����[Ȃ	�fb~�},���O&�l��s���
Pݯw�ʮ�J2���޹nG�+�)��f�vF�����,kܪ(l����+D�&	��h��7u�g��NLz?R����F��B�*'x#��&�����Y^�䄗�M-�E R|k@�����⾜j��lq}�Y����+�f�����7JX�w4�V�ڡ��u >�sM�M�"Dh�Ē��ǚ���l��s����/�cD���e�"�?9r抙�q|H���@���*K��[�1=�T�6_�/�X�I�{��YC�$^��&����g1p=���5q�M�GdL��Tm��ǚ��)Ǯ��A��C�h�i{1�X�9�﫶��D�����,�4����oU����2��nQ��uq���9�
Ћ�m1K��0g�X�	�Y�������Y�N���,Q�T�,\o��]Yn6�Y��%���^q��Au4w�M�u�(�`�l�m�J`D84�^������V��Y��3�@��4�:k���HH}V�	�TW�_K�7�R�p4k.�u Hm2��jtV@��\C��TȪ� �����(�w�����
��rm1��^���^H�o��-P�1�H
IVH��J(��YQ��\�^N���RQ��X���F�U�p�v�AD��hʢ�P��WO��1�M�Po-7����'2��*�	c=Sn����u(#�,�jΕ�����D���)i��;���(�[fy�l˅�^a.�T&���]�@&N�k�O)T���O6�C!�'�~��x�v��a��Ħ�����j�d��Ԇk�gJ����k���F��өڜElcA���+��°!�<��9��VA�H�@C-�ڒ��lC%rޑ��b�r�)Vo"�I&�DCF���I�c��2φ�?$a��1M�0�R��Qc������;� �dBι0Pڲ�UW@�q�e8c(G1t��q�E���M���������M���{|mLh�9����Uf5�^#p̓_���R�`P��cb�ͳV= j���hZ��m��/�t�ht:�lzß�� ��ogX�U�ǟ�>�:��K0X����������������Iw@�C(Ƞ���yڃ�:)�jT^v�z-�2�^����(̇���k��B�+�D���N��oY��L��c�
q���B���E>`�DV;#�h�A��G&�X���k�N$�X���N/_DUBWV_�P�-UQ��Nl���]�?��]�昖L�|Ӕ�Š�[.^�}3M+�ǻ�L1��������XH��8��Sƫ�mQŨ%�T~q2�938kG&8^�j[$=�` >ظLq/�aZ�1VltI��+���=�8�����\$!x����BSK��lp�Q�v�붥42�E9��Gj�k|�9 �|:~ι+����WBl��������@m�"B���k�ȳ�kOC�(����F�W_��T�jB����.�-E�Y��0���m����N7|��!t��(^w��J�_3&|>�J Ye�	r�rnFS��,�7����9D��ZoE�ӗ{hvY�d1��|���p@s���Bo��\*U;��C�	aLܓ�E��.M�LL���O����ѩ�G�A����L��"�����{���UU��3R#=�+�x�3��u��:�;�6	�����m��p�J~٥��vf������\ρ�BP����1��ݯ�tğ��<v�"q¦�X��U��I�Tt�̕�R���ڍ���މ����*ɓbe5���_f�x��\߮�P�Oq0A�FȮ��a���TP�����dx�6_:��������"�������9��#a�s��jX��5 0�� s��J�>
s5R��@W��,���~i �o5�n>��h~�M�g`������ih���t�C��� ��q��Y�#���W���]Q<#1�.Z?Х��I j��B|�����X=4T�D#H�2h�y�6\m -_��E�TA�t쩌�(ϝ-����D��n��6�q�$��ײ��XV1���ᢗ�+�n�lK�z>�����![q�;tՙ�߃;Y'E�4�c"[�"΋(�3p�8/�F�TAU��� ?��8B�ڃ����=oK�Y�)w���U�$m�{l[H�6P���_�ц����x0�m��̪���;�����pڬsTQ�`[�JC3F��l���9	Q��p�vx��U��PFF>�ı�_82Q)7`��_HJҪ���8���Eu"c)91�r�1{�*�����,���D2��*�ղ��϶�){��<|�;�����gnl�X0;P���l�3�<���fw6��Xl��xS�1J�ޞ�F#@�-6}��ޝ�)B?/��1n� ���յ�����fF7;*n�!���f�u�#�9���]D���"��ހ�bV����k�g̙OB��ت.���VX�sהD����{�E��A%��r�[ ӹ�4�p���,�[ʨ=I:p}jxV:t�gye
�ۇU�3�ZR@���V�Q)y-�����[�$c�
5�Hkp-�eքd�a�4�7�I�$��[��+զ�n_kڂ�,�����IT�x�Kۥ
�Qf�G�����_�i�-y�����f�[����G�ba�$��4��Z��F���ㄌ18Wi�VTP#ʅpA��)�i_2^Ǚ�
p��
��Qd�i	�	�h��`��n_1�6�wJMa_�P�>h���\�]e)��)3�rBL�3��	�%�?�6�F�o����1'U������e�9�U3d�ͬ�5}�l���]����s�l?�`k��Y��ث��p{sM֙-!>L��3�o6�dOd�K<8N�Ez�L��l�#=^��l9a	_�2�MsK�zkd��Y�?�ѺEC��^ؖ�f��V�+�rm�;/���^O�	GR���Bo��2�J�^6�V&�_�^�X��6�O��U��8�Џ��][��whl:Kt5,�ڴEԱ��;�U�����7��)q�	a��uH�ը��CQ�%��JSC��;9�l��?�9gɢ�3I�ӵ��L���k�^�{��!b�\�Z�Ģ@�f�7���<�?��uĄ!�Ja���Ļ�p�@���<�ȡ0tJth�4'��YWu����Ѫzm�lH0�/�}:�Z;�f.�����BT���˰�������-X�Ym��ƐաD�_�c`�,�/ot�	�xM}-��ݗ&%�ڷ��� ��9H�4|^����5Hz9X��@�t�l�����k�v>��pׇ}m�>�:.Ӟ.�A��&�i�U�f�" �>�<qp�v��!m����"��~��(D	�6�Ƒ�c%��r�a�MYw�,��h����1���y�[��||�`R�
�?�� S��3m�3i*���s����A�q6$3���M>�Ws�f���Fwg�x
`VW�1���9��)jK-�����8KӉx�jWL�	]��*�_��P���`EQ��݈H/-�Io�)(��l
K�T����~�Q[ȁ���]�f-�y�¸Yn��b��)��wib��Û���uן��.ש�Î-�xM1���U�c�ʰ\m�i�^x
�]��ڐ�.�LfiH��T"z ���h�����	s= �1*��?��~#7���=7��0��1�<��)��5�Т�ז��U�R@�o,��y,Hz�Q�_ l�����/�?�g�NK�\t��S���o�b��!걅���o��/�Rʬ9�q/"/�;��#	l��'n�c�a�*�843͜�LU�Ē9��:�O[r���W�Kv��E��܌(Gy� @s2@|Q�=��X�.��_����t�D� *��ܢ������v:�h���.��.U��S/s�@��Q�$�KI�kc5�����c	����q�O(�])b�۝��Y�b����/5�W��kB#\p��I�'���ul�$��nG�
X[��D-z��j��;�D~1^���#����T�o>�#e�~��JU ����	��vw
15ϣ"�/3:R�O�!vm(�[�0��`��L��2Z��A(��gt�POg�/ŝ)>a�aҬQ����ˀ�:0΋Ql�hd���
��Ȁ��H8Օ8�� �����b����:�W*���=%��*Ё?9N���Oԕ���6��Q��å�^� _�X��d��uYdl\?dDhȔ�n��X4��E�8G��0ܽ	?a��`1Q���O�떑1Hq�}Ùխ=� @�� �|�%�L`Pk��%����ZQ��x��M��O�풢�铘 �<���NM�DfZ������&�8�H�u����� EXu�	�9V�>�E�!&q"�k�$F/+�<�0���7��uB;8�����z����@��BИ��+>��I��8u����fڂ�W��&����n��7LU��S\�b;W��[Ga*X�G���:�t��p���aMe"-�ڑ�~D�'�aJ�����nz�� 3r���狑��o1�0^� nv�F"r���ǀ����}�<]�!*�7i�)�s��u-,^м�`̽J����2��Q�խ�����saa"����9h���_O& l=x��RMF��!��T�J��'�"[���L[\�k�M}m����*>e���<j=����"_�[	Dd����NVm����~�%:eo`�m��F4��8��$`+#uhGW4�U�$N2C]e2��	�J��xʌr�$����phG������x
��λ��8�gg"�H�[���Y$�]���:qZ}�+��˖�j���Qٿ�X����=�FCbP{���te�'�-��~�jZ[��>�P���Y�h�1�eR'��>[8FFH����,z�}Z~M��$�<qն6�`a���u��E�U��eS�Y/����E���ؔ���U*��?j*�ȕy��*�uym5c��%Ib'�(��h¢�QN;OB^��Y�L�J��㓯I��L@N����UJ]s6غ������O���];h��Bq���8v���7��-������	5�FC`S�x��y�ҚC�v�����tp��
���]Ƽ!>�"��Y˕���T%$>k��L:͗O%
M�&q^��H�}�l���M���Ȯ�!�����g(������̄5�>}?t<��Z|Ǖ�^��:�ݶ��(��B�I�	��	s�Um>�����u^��딹]��4_Δ圻PF��G�ы������f�s����B�L�d�9Tp�#�}�A&+{��gR��ƢO_雊<7��5sH�[9+��ĕ�G�I�&�=��� �֭ދ�K˦̥tGt��^�٤QiQ�
b�詩[��c�m��>"OΧ>�㚅?��e~B�<��`�'.��nR��4{��+huS��~�	���@!�U7�η�����12�̮tM)��y�.1�ݢ�ъVl�����L�+Z�����,�tY\����Q�C���ƴ���k�{�~���y)C~�d����Ko�B��B�R��}��1�I�Z=^b��_��Y;t�}�/�����,Kw�D���B�Y�>8=�Qx���S�V�*+���Lo��8�lq���?㔂�;w%�i9W}ʊQNɭCf,:�[�)���Q?O�V'W��-#ֶ�)�4����͟f��ҌP����T"�>8��ߢ/�$퓝9��;*���}'�ZF1��H�P�h�[�����r���ւ}�1��e�r/u�������L�mqzL0�%��{�;c�HdN̛�'eɲq&B�g��փ���h�OmHCq��_���`�*�L N#3Z���6-�1
I�v)(0�z�*�1AJDDՈ��@@�Ql)��m�;�R�f�9���O<?�]0�W�
7�:�������h��VW_�L�7�[4��z��#J���0u��mz	��y�p��G�$4�h���-�13A�5�uj/�H�*�Тp�9-�����AVYi�j�/s���A�����-6?L6 ����Zur��_Vu(ت�eF�|;nԐ�r�3�IZ
�4 v�qo����pf��FJ�z��Aʭ��;�.�Q����/9���p��c�{���'v~��)m lȫV�h�f ��β���L��[���- �щ&F'OOP��q�:Y+l��ݙˀ�ݒQ��^f�^�I��M�'���1y�����_��T�l2#zD���L�G�d�]��O�}d�k� ��{�N�oBVyxQՏ����p�����'1����/��α��R��g���4�%b6����,�&�T�J:�UK;��NT�~cIǖ���ꅏ��׻I��@3�9J�P���C�x�>Q�+!�?5�jw���� ���z����5�^��7��9[�o�+ƝU �p�.E�R��"#���rD�%��. ̈́���/������b*yKƯ��i�~XN���t�� � �����^ʮƢ:�;������6<U5;
8_V䳡'iR<��b���W9<e�vTy���.e�Ew����Li�E�܀!1��u�wĦIp����1�����;Cw'�4�8�G8�D*���X9�A�_�w���pϔ���f>9jQ�Vr��I1�mt3ʉ�m������聊?��	�~m���Q���vq�$�8O�ۏ�0�� ��e� �E����/:t3�z�|��ыg�뱰���7��ҹ���._OF�4���ު��A���;��/�!"��դDÅ8��{��N�]W���0�̌	�A�w��&$*"Xڋ�:,]��Φ�8�T�(�z��:Q�����~���8w��@�`�߫$91cIA�u_u��eYʡ;��1>�`f�"���T�٠���g:��*�&\��Nol�4tY,	s;��_<��%��נ	?���&�f�7˔FޟB�ݤ2>u�U�����e,^So,L��w~T������L��-s�r�!�u*HI�`}/ִ6� �|�Q��0�S ���%�G3��7L��?�e��5�����ՠ�!?�	�{B�9|FGޓ���6�sj�Oy^��� �x3� ���1$�܍*�V�����?ý����l����TP����@^֡�ֱf%F��v4�y��hA(�^�?ue�G.x7���|�D��VSRnT��z�-H��N���
�;X����l3+>��鶽Eh�=�[�@���WV6ݾ��!��O�M�"YB�m�䱽�h����b���8d��W�M\�ʮh�NO%����bz�I���Fw�2Y6��O�-��]��cg���ѫ�$�g��J�{����8?+��m%1�V�G93�~p' �1`ˮ�=��9c����*Ėm��Ct5�s�	M�)�;�й�6��P�*�eCq8r�.O�"�m�!��ɧ�P����5����#L$~��I���x���k�BT�;��ߘĢ��(�|M��4�A�.}l�x���li?�]��d���pX=��i��^�����N��`�<�<��Z?h�"�I�^N +�/�s�w�'��	�ĕc�����H'��P$�I�0�����	�ȋ�hO�n� 
�=���\q�����Io��M����p2x�5�Ѡ	�Y���ﺎ��F��b��1M"�y�1�+�Q��n�J�$�Ą��@//Q|����b���5�t��EL��`CYz1���/�����6��d���j$A�dڜ�T)��:�P���e���#��
ď׸�o�����
,2��YF�q���
iX�A��sY	�QѲ�:�v�Ѫ�08��:";��?6��蕤���A���9�m�uX��+���~R(G0�m�p6D���8���]�
A�aT��[������F�HiԿ������G��gNm��dn$DKX*�S<1:�^�L���9���\0���뎈QV�h�or��� �_��٫L~+#u�U�0.���,�\T��֖�L�X?�[���\)����V�ox�Q~m���9.���6�Qw�!�|^c<a-��n�J6m�|i1f�~��n(��:鵜"�w��X����v�-6�y�ՁM������;��ZE� ��!�yF��mu9H�'�~9{�l�f�����7���n���	��0�蓦rf��!��^���Ɏ8fʟ��r˜6���c""�*�Z[� �_]#�_��Ju�_rw��65�!�0Hf!k	����/<O5縵Mg��M��Аt�3�g���j6`��C�I��s���w���@�Ol<~4��i���e��,�g΋כ�Xn�!�2���B|=�|<�U���N]�)��ǋ8����~��ơq	���割YZZ§]|�Xn���\2qH���=~� �:����"�6�e["����=����NP>�HLd쀱����<ŇX���o��-D�3�R��<�@&�Z��t�I�7�nE�s |{��JF��n	K��g0���ԢX�~�Փ�ٲE��M�2�.&/]яd{_��l��2q&���Q0̗�.����U��*���������3oM��65�����T�y|<g��4,"�S���vK0ڂZ�P�bﴣ�	��]�*���v�6�N�4��yN���[�㠧G^1�H����p$3K������&��<�dA:�ރ���UυE�tW4�ģ�@_�t��R�e>���ڟG��ygtUH���8B�D+��Z����^$��DL{����Ա�_���1*o�Iq���**����>��^�@��m�)�����.C��Q�^�綮gS�3�U^c�ޒ��zo$���F-* n�D
����gjq�8�:԰�	nl�J
�=�t��'��]isI%ƛ�+n��;_숃�N����fuǳ?0~����0��?�Ȍ�̓\�V;�6p\ix��p��[�N����z��3~ra͡6q?ȝ�M�!���HCd)�D�Ғ�?���l1Oh
(sz?�M��I�/#,1��H�ɇ3�����ig��5�=����^i�!�e:D|b��ԭ �a#�1D�����81�}���Ѵ죫f�)[������SZ�w�!
\Ԣ��എ�l|M*��t� ��0�C,BV��

F6��q����e��i���� +w�����݀�����
L�.��0�N+�h8�p�!9J-@�J~��l5��
�Szh��������'�齘׌�ȴ;_ݎZ�lfL*���"u+�[���/��R�^���ųe��:�V��Mk(�
|uS��9d��Z'o�G�T��S�ؖ�d����}���q����y=���[E/��/��d��ҜN�K7��.���zS\5ڰ���=�K#�g8c�/7>d���i���f��!�߀$�r�A+z�t>���:τ���9�s	�.R�9�t�Jŕ5q�=&r�ךˈ����Ѭ�بs�_�0v4�)O&� ��~U�����j��3�ȼk6x7\%+%!&s�5.'��IK����%��ҧ��;t��);N�*�8�[u
&>#���ЬjB�7��i�T�V<�&P|�Q�'֚���� W'p<5v�&��s��p6�iRp9�8E�c#9B����f"e�=��=�TjV$TɄۓ�3�+0C��b	�)uH �0H������B��.*S۞�"~qӿ6g`]��]è��`!�,�M��Ԇ��P����Z�^�y���ϾB��[�W"��%\#^��n,9h�T6�u�w��o���2�|<B�����Ӂ�g"�l�YAY�C�)��y8��m�b��d�R��u���ٍ��3u	M��:�b�Q��3��-}�u� �[�n�>��I�LHjJrb��F�q���**����94�x���'���>��/z�Ӥ��̢\R��&"�;�q�y��%G!|=p���募�~Y�_Y�P3:M��Rt��{R��c�O�SUv,G���G��g�j[R���[�_�Ԋ� F�_�r5}�D�T+^�n���C�2R��{�!�S,��T���ևKҡb���yТL}<`+��;���%��?�Ā�K�< ��H቞����O�BiڌCJ�Ğ������R5J���w�8�g;J'Rh�������˗��F����l��9�J��xi�i&$��咈�n�q�X
������mF�K?�����]l~D<cܒe8��!�~��~��6���Y{�3��{q�nm�i�ĥ���Eə#�Ư  �m��OԵ�a���*:�R`�Z��y
�P������h*�������z��)�xI�JOu�;���Е\�X��eA�at���Qk�Q:��۪���H�eݤ�N���X�h�p��2C��;f	�qB�X�O@�ݐ��=�pm_\��I��W���+x�Һ� _ۡ���Ę#X�u�	��(����au!"����%d}�]��ǁM�*��t3��ad=�`�=*5�20��ĈC�U�8����Z�������V���8W�4��ѓ*�BL��?О�{�1��g$=�*g��>��#����n���\��M�^��˯e����C"RC����.���U���IT:	�l�{GdC���^̘�(]�C��\C�8�q�]bn��)�#�4�����o�S{��)�2ִ�:J���of$��2�:6m'n��0Xh�Dl�
_�
� !��;*���uo�0f�YP��lF�՘;�� ��F�J�!���<��t��?\��WOm��T�G'�c��c}�?N��i��I�����Q,3��ͪ˾�
S64��f̫�\���됂.mP1��a���Q������f(H�'���TX��V{�}��Ӏ����r���-8#8~��Q�y��"�8*C�we�9%�C͛n4KN:�(EYk��Y22�Yl�~���r��h^�d�)�JQ�N�č#M3B��"�fs�7x�Y^??�Hb��@�׊>u��Z�k�	�Ӯ���&B\��p�U=G��lA��n���OB ��>"-��l�r��]$|�n,�m[S�����gJOG����٧%�AA���=����8a����D��^������4���I`=�zC��=���GnX�fs�.����Vf�L�su髄%l�m�e��SM������ߍN8���6�R������) ���@�67�jEϸ=Z��PN��]x�8�O�֣S����tu���	��@ �&�������<���R.�뗍{�(;��w���_�@�Yt�h>�Y.4~�1˔%��J`���&����~0x0H1>v�m�Gξ��_,3��ٮ�o��Z�o���E��į�4na��0��+΅U]�BB�������E��w�퉮������b��t�@d�֋���/��S�r�ZY ��ޓ�+��R�3X��$#�31�d�s�"�ܢ�!iA�a��ɳ��'�j�54A!�"2��ߙf�O��vq 7ā��{�E���i�'��ܦ����?����P��C��7VK�/V#U���kND�0E�o �s��ؐ�a�F#[����v;�]���"@A/`�tBBJB��<�'hY�o�`��l���w^�T�'�Q݌�~�>a��Ĵ�d�i��+ռ���-�a@G�	���j~��Z{��uGԀ����(M�`՝,�7�~|Sӽ5����3#����s0h����T�x��? s$̢^���ھ���c}���5\@���P=N����b����!*�d��I�ۜǢ��OM#��;��Ͳu�SQ���в8v��K�I��f���|â٬��kt	�>6��)X�8:�KF/��#w���-D�) eYȋz��D�S9���ZO@׽����A�Xi�<�rSɬ�[Yz�� Kd#���P��0?Í�!��E�|"�ˈ@�.@7ڳ�����#J���_��7h��_�v�4Q�-h���ƒ����!I#�ܟ�G�q&���oO�C8p�K��y��[&z[+9J����� �v��h�Mh�����HZ����%��l [f�xn��p���������- hC�<cZLu��i(p#}u�i9琛�*h����jŀɗ^�jO��W>C���iR�����g-H%�g�5���2��`���N�<�!�^dC��s�����k�ILPB?��߮�H���	t����&8鼁.XX���"�Mi˚�i���&�0�"���;� �!�=�|+�X+?�.�]��9th�6D�.p�FOGoPd�y����|�Q�W�~��@��!!��i�M�~���G����M���@ot��)JЙ)�ٚ��ߕ/:�L��z|�l����G
�y�n	~q��U�}�4i�Y<VQ3�@ˋ�;�(c#B�I�og��tnH�.R ODZ�z	�_r�Jy��G.��  ����H.k���N1ڮ�@�i�nɦ�2ٌ�sn0��rk�n�$�5ȫ7�����_o�.PW��n~�G�u��&����zP���]}8�$�z鼂g�v]r{����{����%���=jf!	����N��U�R>KA����z#�=V��"W���T�dԑ'�A�/k�9��X�6��ADw��x�@fT�EͪRvq�0��Dʋ�� d��ɞ5��,�1�b�Xp =FPP��B���#`�W;­�5�~���]�Wj�#p�F�14��a_)z�ݳC��H��#��-�m���2���r�n��DGĩ&�y�>�M�̫ł�S�p��K�^��|/c�䳉���Z�Ӊ��:�SnS�ھU�-y��,! �_W}ݗ^�4�s�T��sZb�'�!�Bk�8�)i����.l8��f���_��V��x!_���"�-NS�k��b[u��%%I��o��KvB����z��:�䲭���g�;�y�A�Q���K��>(G��$����t�fk��#4b�������/�}_�f%h�yQRU��q?�i)*=1N2�N�/�r��$*0����8M��ӅȨK�ɊC�2���'q돭<�0�꼇�W�H�3̗Ѯ|�6�G�m�t�+(�DO1z�����X~�{X�*�4@G1[a�sC����t��1։{�\�n�%�i�u%тc��+�A�T�*��<F�?򢰿c,y��:�m-��,�"pϢ�GS�[q�	�w���AVe)Ae���U�;��:R+��Yӏw��l�X63���� h�qL�X�'D�!Jbp=�c�.�^�D�`�|�%Lux��(��8G|�� <�";?h�?	(����9c�'��Z@�I:�[WY���D����ŷeį��|����ã�*|���DlD�V��i��h�n��S�E Τ�"a�6��3Y<������"�5d���7�"e�ET��n�࿯27ߦ`I����Ű>��ۦٰ'���k�K�4n�)�&ػ����0��06gf܅�P�o&�H���ʕ��n��v��Ovǰ�ّ���6�f)U���6��n�Y�u�Jw5��4Z�ߢ4��A��1����_=!�e����i�z ~��z��_�m��M�7h��wA"UGF�2�V<=|Cq��aDޯLA�W�HJ�g�@����c����9Sf?x`lF�5#q'cL�l�}�°���'0���?��0~j���R7�FH���tӱ���R��M���0lƹjo<�8&/;Z὾�HQ�-������}ULٜT�F&�|����P�z%�Vbef�6K��m�d͕� ���W�ۍ�Ʉ��%\f�;�M�%GL#����';R�����������d��.X���z=_�	�$b��L�
���qCd���!,���B�7���s獡�($Q��Fa:**��v��j�
nz1_��8��u.]��6�������� ��9��x0�����kǺQ6��Xo��H�gBxͫ����ޮA�k���V��#)n�k�͏7��1-�(��n7䔉j��%mz���N�6.�z���ئhv���S �_E������4o��R&�!���y� M�5�8��vl��oպF�&�P＾d�i'@���F�y�U�y�y?zvyZ�����4��A��P��.4x��#���<�!�q�*rO4���6[(���A��a&[I����k��O��T�-�J� *�@]J.�	#b�6�ܲ;�ȰK{µ�������:yv�|U�YǢ�]?4�>`S�fQ2�H<���E�a�i�%�!��o�x�~��䪤��l�Ch�G̜.>���l�Nr����̘�B�+���=��C�XWti���Gr���4�yMϴ���kà���= 1�l5��"�o������m"~~���ח�k���'."X@m�2�)U��� D���MRsZ��5��k���D���o(�Vy���ρv�j��$��}�$��^���������]�R��]��ǧ�O�YN���:E��T����,\���}����=�v�na^=��.§���d
�s�i�N3��LWES��r��LҾ�l-2)Ӄ)��.����u��3&h�,eЄԾ}���sA��zo�K���� �V�~��`���p���=�����/V��!B֑���n<�hcs���d��e�iZ@�?e�o�((�𥂑�������8!<~���殗�u"n�_�=ֹŖ�$kᜨf���s��"��Id?�G8;����k��7`�U��!���\�L�)�}L��6��g�v�o����-��||����)���|6I4� .)��|>aA�h�	&��4ggq������fO;�٨S:&���	$� ǈ�~G�6�U���B�D�mi��ZI�O���<�`�s�K����,����tk�o/�|� Fq�U��Ù�	�O'�jq�@Yn��Jv"��v�㕝��_J6G(%?����*b���Z�l���q����2M8~��C7F{7	_\��F������m�QQ.��ݗѺI���T˽W�P@k��d�\�\HM�a>��g��!��j��7ȴ��3�Eڏni>r
����O+FU�w����3�V���h9J>p�`��*�[f�~UIki�[|��@/�3׀��@�x��Z~�ky��� �B�si�L4�%�����%�0��V��.9�$,���.b1��Q�l��Wa}4��_��TF	�	֝0��.֐���V������.�-Y�	�4���OO�������5�\���}���Ax�Z�^�;���?�ѴG[�V�r��q�<a3@��X2!q���,�@�6w��`��{�+Y�6!*�*�.Zb�ƪp�2/��oM�.��³����+s�m��E�aaC�<�C|�Jc��˒Gi�,H{ǃ�^�*snw��!���g`i}g�+U�wn����`W�˔[/p�����wMz[��%<:�z?�nt	�w/��3"�]�~;^��+��!���o �"`��D�U�l?�yT���u?��ǫ۳u#i�p�;!&ZFII�.�<�z�H�2.>�:u� 6��-x7�fu�洵 �c3�YLXu����s��KE�R'�忠
;��*.q���o]�@6w�j���rj܈G{-|ˬ�
&2�	�Ϯ^��H�6��+8E���F1�� ע�{�m�����_�����ix]@�^�p
�#���;s� �� �4N��6��4��y��K**6T)�oJ�M%"�a�s��`�7�Z<g��F��1�퀍�~���:��T�tFq�=z�$���m;�O�g�t�qo�@:�68�d ��:~��RP�5�T�{���X���m�fd��3;�u��7�ߌd�B6iەn���e<U,�,\��D`�������BJB�&"�jެ�-��0�r��|��;����č���K+�$��Fc�`�X�k��y�ܶ�܈���>�����R�ٽ���1������"^�ޫv��G���7=��11��v��I~%䢾^p�˂"
������=�̏`�b&u`NO~Ӿ��u;��5��1%E���%�f.C���YY��-��+�����MD����{��ir������=�-����6�3{F�<�}~��֜a�W!C�|�vkW�|��$P=W+�!�u���H�hU��n��l|*Q�$��;��k�����o�� �T��h�M��]e8��3,�,9b��9���a6oU�j�ʽϧH�rx$�,IF\Ct�H3å@�q��&����BdF?SA��Q�;[U���2����o��"��دm&�aR��͞Z���@6U#��$)���ol-}9r֌�C�5V����v��q�ڕ��rgDؒ�Ń��9_<�$&�DL������}�"�A�3��Ls���c<?�{ă�64�P2G�	�C�)DlLvW�e�dI�k0�&��!
{�o�D�� �<�!�i�_݄>�Ni��*i��ƽ�S�C�J'6I]@m��jo��\��̀A��؜�V.�"��4F�����kU��i�,�v�t�������7gm����ݣ������8�G'�%3��}�<�����vH�S�X1�E8q�璕ⱎ�a�&OvI��r���0j$�2���WZ=�@��B+�@�	��͑�*Y�u��zt~��E�p�֡CN쓔�Bm�(E���!���� 3�dݫ�1k%+NP5JwLE��d��|��;S�(���J�bQ?���y�o�FJi�X�'BWk��<*�f@��^4&��m�5)A�v�� �����Q�L�}��z�%����V����i��{!@��b2Rmʔ��p��5���{��O,���I���`�}�@�u*ފz�bz��j�L�(��5����Hf��'�~�͂Ï\����h'�s��2�a�-;��V7�8ۊ�k��*� ߲�u6��̇)�܇8a{d��&oTKF�1�Q��$��u1|-t�R#�����Q"q��OO�،�c��pEf]�1��u$�@ �!�1�y�4��z�/�.�k�3��1�Ꝋ��*�yiŗU��4��/*&a���mQM����8�+Ӣ���\��|��9���T<��S�T-[/�&��a�	�R����ҍk��J�fOo�
.�cGt�d�y1�S�ښ��&ФcP%��8޹��i�^#�4,�#B/�˗�s9ޕ��7�+�������0<��/]�؏yM'��}����ֺ��5glQ '��/��er���H�;u�'�1��eK"k��&Ĵtٕ�E��M]���\!䯈�}Դ1ft����F�ze ŜVmBu�+{�K> ��d�<*3��y@ �?���y�~R�D%�C�&�q�td%���DĤb���y�E�4�x��j2bQ��&*0�����V(�����u����`���id����&�[9w�%�8�I�!����_ �ҍh�F�G ����?�����A�d,l ,H�bH�D_:�{�Ĵ�3�+[��N&�.�˸a	6�:j�����0��]Lg�,���A����S�ӎܫ�ǽ�����@���X*U6@�:����n#�j�<. ����,�1T�UE�S��b��3Lw�UbrJuD]p�GD=�h���S��^��m��S���?9�C|�nAo�#����J�W^]�<��j"³��zJ0.�^���($v4�8v�}�%��.~��D�ț�"�-^*H������=�!,\N��2~I'H����T<	�A�΀���]�N%�wF�V��Xq�|�K�����P�.Es��Ŀ?k�����j�WJ�����>��G�W�h���r�]�T��1E*�<qW��@�xXI����m�l�a���:|����j���#�=B'Q*˓���I9T��r�(��m8��H�I_��L��[�u�m}���|���<�;�t��n��\�¶��@y���mD�BD��,��Jԏ~O���Gϕ8��0��|�re��̽*��������G��$�x1掼�A�O�xu7x����Key�<��'f�)DB���M�-����	_�J2�x�(
���m�on�����fOx�D���U�@�/��?�9�2-heM�O�E�N�lf��e8z7��0�@hP�B8�����N�e���+JN��?���'�cƨ����Ô\r:fC���8\4�``�8�X�C�M��
L�IAr�J����82�.����8ȑ1L��n��x��t�<�S�+�f���a^��R�+1�M\)�W��;�e��j�����)"�j���όGo5e�ǣX�э�Fe95Or�F\�b�;���������q>8dN?�jA�t�b!@��ȿZ�"�̃L�/���mͤ�;,�aš����j �#��hl�_��
J�ʵ�O��I(����DZ���wl��]tk;J:����F͕�qǗrz/�pDD[�>4郻�Y�V��m�����f�;m�@�Gl��@�ڝ����zЧ��*��P��U��{�N�W��O�z���]��W���b��<�Lw�	*����7;&����e�A֏y�!c���������ba8�CI�
�e�ݸ
����[�woJ�^��C�\Xy��q̼����j��SG���÷���O�a�-���+����ɰf7��
W��V=����1e�'�����	k}��`��/�!�4ܨ˒*�/X�r��`uf��3Ů�K��S�I��
��~��%z+������)K���(��S���8��:w���nQ�R�n׿4��ʵ4̏�t"��;��9��'�WB��ù�Q�(A5�;gi�2����� %� �"��56I�]W�FN �d�!���ZM�oY���r�8�T��*L�ً��E�v``���i�.��k�����SRB-,}�9	��O�?kQ��
��#�sM��p�a��}\t�{d��mJ�D͸d�I˹�8`��r���a��ouS�,�M��RT�/�Ƚ�@lp�c��a�;_�ǚi�l���d�Zh8��eLM�-��)����gV�P�L�*z?�a��]�eӹ�s����+~f�8�-$�)��������y]��i*X�m���4yJIb�[!��},�xD�c�qսv9g��|�V԰Ü����J|�F���� ��d�{�%"g�u3}m�����'ձ��<�S��R�e4%��jw	��t&�n�X�u uU}� ��9�mOEp�?G����/`X�c�h���t=�X?���'��٥�i_A��B����R9F_W�w�}K3��ή�~�v�j1�0�@-�^����@"N�6A�io���������x�Xǲ'�F�{��÷�VIL�m0蜏���*�@��cfe�y�<v��`��j������@�9y�����\I���D~uv@�BRi�!KhLʏ��Z����N8:��{`���]�]���B����g��q��������t-{���tL�$� ��$ey�Be�_���-83C
�ȣL�"70�Kʤ^wDc*IA��n�>����sv��<"\�i���.p���o�=�Π~�X�ݐr�d��0�@�ÄG-����uV2��r��"n�XL��^X��$�	[:��_D�7�QAEy��*>M��$}�c��[ȼ��^X9�.O���`v��y��?�~�*�W���90���M�VZ���p+��R��}�7���;���Smw4�ε�
ܑY�Mc8��Z��P	tR�:�K�U�H7�ln�׀�� H�hv�X���|�t�^��,F�=Ki�*�Y�!��&=���V���rz��8�
L�||D�W��mA#�p�#Ð[ʩ������â/���ˏ���)��&�j�����׌���W��틃�)��w-sr�%���:8�J	����4�gAڭ�7��F��wN��Z�]���^C�� �����"�Ǘc(�(g?���K�ow��q����Bֲ4��dT�����Bm/ٴP����r����dIܓ����W��v��ܛ��=<�Y[��w3̮�������NtP"������ǄD��'��U~݉"�ä����LE|h���,�\Y3��z�V`���q�Ej;H�6p`�l�/a�����o;�pH���E�:$�/��97�)���\t2�v��ovV��R*��B����֟�
7<��[�k���Zе��:sQ�LOl���3��<��?�=C�5 gʁ���-]�@��T,���r��N8,�Y�`wNԤG����K0:s�6g8J%�R����
��y�"�A*R&��]�)���6"��Z_d�U
ݰ$��\����X-�0p@�a�*$�f�q�.;�l�b�ft��Լ�LiU� �����*�ʨ�q�����x�u������@�W�rYb��/v_r@�T�{J�!�����а�Z���Z�(�o�*��ss��a#n�Ɔ}-oe�"O�Ե���钭��D���([wDp�b6����s�lܫ�G���p�ηK���0�#g%�~���v.�y�M"~�+�P�7�d("��R[���+}̲"y�AN朽�.~+T�;t�GN��'��܏]fF"�Z�i317�0����k&эL���lMg��$�#�m��ߌr�}M٥��~� -����j�$|�	Ud5����0��dc6�^I�D�3�콇E��y�$�3��}�
:��O�3��W9XS׈�԰͡j��G�f�t��-\�'Z��L�>&���*�}���ĳ,�o�����V*� mYNbiHL~t�	۔�����f�0m�-��Y|��Rr��n*�e�0e���>r��K��r�t���'�x���7ª��j�� ��n�tw�gڟ}a�Z�t�i����c$�T�Z1YW��]��U%S?M#������J@z�$2��mY��ӫϟ�i0k9m��ܧ��i���X[�i!'����=-�6��{�[���>��`m	)33�<@a��Iޗ0D|釮��ծ�7~�uNQ$�&P@j��yٺ>�d��������Ԅ��X�܃&�'^���9i���M$�O���5��b��h�(5��k#��Y),Y�H�TZ]��C���g�k��m��������e�B"�W)~�Y��(�p3����t-�����d `��xPTs����X�}cM3ǄDp�]1ҬvZ2�2$^��;�ūQ��Z1E�t�����Z�!+?����t5�'Hr�tDh��*�{%w8��fWÔ�Ϥ�#��͑:a�ic��_�2�]ڵi�j߂��2�>��~m-�-��ݣ��뒺��!���Ҙ�N�E����>����:�13��"�t�Ȥ�*���A�����z�H���סKp�R�<�e	��ș������O_�,!�x;�O��Q��;�
��{�s^sٸ����?m��~��l2��p�P���۠kp��0��+ǎY�U�U��J.5�RC�8�Wk�Ƭ�L'r�7�4�>�Z�D	���3�֯� $$qZ��V�8"�h���hu�a��ʍRuH�,x��G�`�4-���9���{.��j�:!� I�:��J������F�Ss����/��Nx���@�Id�OK�v�݋�� ��$)���,��u�f��]���&����t'�\a��s0XW�Q��r�25ʁ���m���~_�4">�:}4�(��k�?H�犔�h|O�b�즂�DEW��e���dT�=��`ntw�7�YCo���j�����~8P������w��&)b�a$��t��ou% O/΂}]��k�B�K��U�	}P[��?�����Q"�w0�����?�nuP�5��8Y��q#�=�X.�F�箁�!�.R|)�3Y,]�K�?�?����R��������^P Ο�/]����6b`�`��ת��[���xs��?X��3�3�SR9�H���\S����y�t�4��*��,�v�ϯ�^�k�\�%��1�ě�f�Q�sp{��Ҝ����s<�YB��#�ёS4� ޗ�H��qrg�-�8*@"w��ɲN�WA4�m6�S-�P C6�O�����c)�AuԳ\@�tU�������Ｄ�!fr�g�s�O��������1�ްTf#S�c�)�NX%�	L�YV�VY�\�n�2���yXXe�S��/����%wM��Cl���;�U|� #� �'�b)H>a���e�iJ1踣1�d}��i��]*�gszcaH��Ve��iD�4P�Y[��%C3K�2
Ь�j ��p	�ܚ��l��K�V�pc)�W*�\) �@��Z�׹����u�)K�|��z�m,\�a����=rQɚ�������'�痔�p{ |�U��*����"ٓ̍��1l������w�������p��+5�qA��)>��U�%�&s���7\����v}��^M��NcstX�d9�
�B�a��YGR�8��y'̩���p�y�àeC��Bw�?�y'�"��f����
�g$z���#�_i����(�ٴ_���D��� .�i_	g���9�#GTA�=@c>����_��np�M��n�>�W�	r���~ � �uS7��N�b^�K�5�����J�Ԧbr/?�#P�b-��趏�N�\���hp���X�)�s�7J���ޛ>�R��ZH�]a�x6�&M13��G���SDҗ�Ɔ$���c�y�L��U]Ep�.�/U0b����CP�W�Ӄ�����)�p#�U[�*	�i�ʛ���4D�WeA\K1DMb�z}!�P��&�am��΍�	��b��zrf;�d�ꇛ�kz�o���3w��-����ȯ5
�"��Dѵ�g![�=�S�����=:�ha���A��E@r�ȟƟ��tvNE���8xBn��˔\1��I����F�n37�ų�_$X���o=�?��_@ZTwkgN�Q�ݶf�_������:Z�өL������o��L�6O#�[�ױ�<2
�6k��(�����*�.���:�*����青��-%%�E��Wva3$N���������D��l�b������?X8��C������ �ko�m����s�O6��sA�Q�����1ډ�(lU(Ί��V�%�dk>:�l���5_a�p�X�QG`2��NI��?)�hgBWvA8���L��z�81l�ީ�9�Щ�j�/ajF˾�Q��������z�[4Q�/�z@����t�ޱ��ռ���μ����9��$�-J��]��/8��&A~����:{��^	`�1�sQ,�؆��Ί�>L:�AB��:��>��t������^D<p��� �}��B�'dA6u�m0��q�a�1�a��mN!
Kr��A�L��U<_��V��{ώ<�����5Тմ�b�粌*.�{�7�ŀɹk�}���>���]���A�ZQ�㪙���qj9��➋�"v\x�	����8xF��O��%*�?��&� �hB����+���nY,t,�T�-Bf���v�`�q�ר2=���u[��慷�]�*s�ңG0Lm^�'�$�Y:�#5Z�칈��/�DN�
�~a�^��̓O<�a3��C-���XYu�E��::�~�n�R���^1����;���H�ǑE��!��6���muI��8��jF�o������ŕ�����M�u
�95�}'�4�h��vi�Hx��f�#0�GI�y��3�����=�f@���m�8	 q������%�:VWk�!�1*�,��M�e�'Y�mҫ&�GI���/��3�%�����)�3��#@��f��%�S��!MS���X�5�qcl�1���$l�D�_%0f��E�&�TH���5���d�yaՑ(m��w
*����d�qV�M�D��C�cb9�~�PR�\_*!fV��u�O��Q��*�����G�f�pם��7v/l�gL�e�s��o�ⷐ(���w@��f҇τ,�z@��M?�#���[f���%?���~��d�XI|�{_J~���%|������x��L"R%��C6���C�������]Uw� ��Ti4���T�ǚ�L�t��ߎ�p�T��D-C6ts��[��1�]�O�iz)�~4ɆP��I)�s���3U'�K����$\�n#����>-���Ҷ�v���)��qy@B�SU������ۣi q�䃣�J� �R4x�}�4lg��<��'��=��ʎ1���j0>]�+�Ÿ��.����P�Ĥ7�Ts}���%r)��6�����P�IR���!~�6���g#��Y�VB���'��ʚGϩU�[�q弳;[�f$!��^[�7�b�	�y`�K��p�hՌh���'��R�0$z?���'B��T�\'��ۇc(������"�Ce<�e�E��Aq$�|2d��3䟫On�P���k��u.��j��Mkq90Ef��K��_|p �Wn��哠��T{o�����VxU�o��M�glВ�CK#��`�7�2G�L��l(p�eu��[58Ҵ0.�n�5�>lQp	�R��T*��G�&�᝘���/�W@�^'��	Zӈ���Z�lk����b5�:�H�r}O4վ&�
 L�V's�RŦ/�e6�!���b������\��U14�]&�9�/\w��2�*�a֋kh'��|!�9-��:�RL1X9�0C�
�?~�T�]��%;�YR-Vb��(�EbSHE��RѬz
�W;���ղxa�t�	�!��&:5�2w���/�����ǔcl ���WF|�fXx�5�~9�l�m�G8#.L�Y@�V�����x����n;6�kW*��0z�����V�a�;������τqX��|Ȥ=L-���L�1w���@p-&��!(�Jj��Ea��>'�RqŅ�(�F���;k2�-��❪�2К������rV�V:d�]xAb䬥��y�?�\i�g��`���f�Pr�9�ft�x����qW�L7O��Q�7= |��]���2#�o��i1��Zr�4<Xv*�x>�F�P��Q��f���[7���>��u����o8F3&��_@���A�����f,K���W³t,��v�_��j��:���S�R�x>m�KE�5���n�5�
I����.��_lI����Xؘ�Ö��x�ti�꧅�\r�tr�x�&�w����Aʚ�-T7��{��<�?�׵6����jD�\��,�W��jyِBj,,�4�R�8��ߗѓɺ�7좘Qhv���_�̊m�V�[�O���(\D��gv�Z&��H����jU��;���e1D�
ZXH����s[����-��f%8�>���թ`׃
�e{`�Z }�wKO��g빉e�"Ԛ�ɮ�9���e�#�R:�e蓳ۤEb`��Dht�������y$�/�ߢ��j��P�d^�7ܖ 
�^�Ż��P��/.�a�Z�DQ"I\��;����z	��}
����բ�Ih%&�����4:e��>E	fԁ+j��w �__o���'�nks��C�M�ש��yK�bo���;���&\m��I�}���,Kڹ��ɩh�O���0��"	|Q�nfu���>�B��Kӵ�
�}��h[�k�Δ�x�P�tpa���P)"6��+��	I�"r��Wb��{���CM���� ��V�W*df�R���H~�O�y�̓\�Vn�;|��c�tx���ó�X�jbҥ� 3�~�d��ݛ�LvRR%���ka��_X���NfO/d�bK�������͡e��i+�}���0s[8���BL8'�[b���_�w�����pVc���C\7��b����x�;��A�/{�<\/�����``o{�d���T�P�'���G̍���]�hl���$`!�Iy���9�|#�S��*�����;wF��1�-1z����L2�ؽ�;�
�ɂ���>5�{(m�����6�#���r��7�b9'8�@���`�P���������n������A�"��sb����4~��S<R�C�B�Kq�$�TR:E��zVR�1�|��������"P�.�P�5lJ�G6�D����ެ#7�$�3Yƛ���HO�n��EY�s]�Tҗ����g��"�D�n��.�X1h��\�Q���@"�;������e�+'����:�!s,p ��^8a�u���e���0�~ڠBQ�{��R�x��'?#�pyd��
��FF'9��y�i�o(�y���6��%#��ͪL���W�Z~eC2t&`�s�__�j1rߏ3H�����.�x�̷�[��2 ��&��񮍨I�?�<�̻.u�Q`zo��Z��q3L}e�[U�&Z^/K]�*���l��"�����NU�=*��u�[�n-��[c�*rmFL�߁��{�C�{ ����qC��!i	�(��v�z���y[JѺ;�y����1W�!)zF -)�Vi���5:f��#~2��͛���.J)��2�K�
���?<��f�;�:�<�R[�>���cP��h}�dlu��)#������S��3�3x=E�I4��̕;�h(���Z�=�ب��O�p�Z�|.i��U�i;I����H9o��� �K��Wdx���	d��+��TԔ~�]����&�t��;Qb�R�[;�t���
�ak��1�pf��TQ8Z��N��`;�ʜfe��^��j�0�v�U�pA�:芗ȹWm��|{>��x/�C�;�I%���z��ޚ:6�]X��#}���݄���ˉ۪��&l%?�Hf��u�� R�ݽ��E�ԤyP�t$�WpK�z�C���4�Ν�	 j�͛�(&�'r�K!E�b�S�
 ��рv�^/�s��������.�G9V!�V�fX���r���x�!��[{�'��e�$h���Lzj����s�%�@�� o"����j@��,�<��[�st�R�Bg׼������d��J�܎@��~�f
�k2����5�C5GH�y�Ԏ��[]
q𵋈Z�ԧ*��J/��l��WJ������%���?�Rh��ꮠZ���5x=�zᪿ��pXF)����[�Q����7�� ��Yf�a �;h��<3�Sa3��@2������`�Z�d��o~;�L�2x\�M�3������(�0�f�X���Β&����>����u���6|ka)��	��?�:��39�0�
`��0�m}-���0�g��I��rQ�*����려K��Y�A�9�/�$�8�x��e��46c���Oq$�t!8�$y� ��-q�3M�mmv��j�ֆKmG�������¯	"�	}�I�8_Oδ��o��\q��L���i%6?�%���U��~���6�m��� �3H@��
۶}<�X��c��J�(U�'���|D�5��櫣,tZY�e�@�A���:g}f��!4��d]�?����cPqX	��B�.C-��ZJ-���������7�GR\��+DO�:�J��җ�e���ס����/h{m{�9��ۏ�Fͥ�R6獡q���ف����N8T�jF�a���:�sW���E-@VGBNT) �S����;�r�T@)y��5��m5PD_+��Ah�gbr9���P��>�t�D?���=a4�
�.[�b7	2A�>��J$���y�+ȭ��" �:�s<6��FSv��k~N3�����}r���g-�e� 5o��$a<��/F�}H�y���kE�X�w+V���/������O�I��Bљ�#ǡ����i��p�����-������ޚTٵ ��S���pyP�t��K1���C�钴ү��LA���A��4#�$�os��U ��®keI[�7*sÒ� W�*�H)ƻa*Fv�����=���<t_ ١���Y��n�V`-�̹�� W)��\S�,�U�0M����3�0�J��W|��H�hV�u`aT��*k9{�}��b���\x6�1���6ÊS�bUH�x�эe���LO,!���kjph��ˠ����Z�Z���/�+Ҟ.��>�+�����܈O�\1�n䓞���6�wKF�b����@�$6(=y.k�i���X���
mn�H����a�?��
��|��^a�� ر������s��S3_���o&.��#����n�	jJrܝ�jNwN���VVc�~v�Bρ��c�J}6�qGC\�1��:��ݠx`�4�<i?Nfҹ~�H��X�@��A[�T��x]P�ԣb#�J�c0��9HUO��cգ=���2)��=K�6{�K�BW��w��:<�������
�R���~�b�*����A�U��_� j��My(���ّ0
�Ĩ�ep�g��.�O�������uH(�ZH�tw 7���˔B��{a}��s��y��Mٳ_���k|r��¯-}�Ȋ�N��?�^T�.�L���#�T�*��j�Q�B6�7ڎ������@��7L}�G��kDg����l[6$S�n\� ���}x$ ��v�k��}��O}p�E莏J	�Ӂ�]�=�_����_���<���#�W�0H��}�|ѳzǼf��-��"D�[���H�wl�l��xu���� �%��ݑS ���_`��ȝ)�jΧg�׏ w�{g��Z�d�˦�(���A��d���"*C����b����?^��=����*��z�0�6w~�>M�Ⱥ���ى��C�qrQU)e�����d�Mnr��n�$����I�)��ze�g��8�*+���\S���8���Y���=��^d�����z#���$5����R`4���9���R��l8�LurYq��7�.��+�^������X��M�XH�����'z�5'�̏*1ff�> ����3�1�����&1��S�H�;��(����-DF���➄�-s?�}�� �oF�}V��U��.,Z��JKADQU����K�	]'�9���A���ҝ�1�n$;��Bn���|uy��%�����B�w����X��H�d�$�(oy|�z�?uJ=�d�r�ˌ5:ܢ�'�i�.�98�0@�9
�I�a{�R=�?%�Fϰ��cw������Qv����0�_�'��*����F�����[�]��p����is6�O��4�$%� �Ϯ]����A�E��*~xcs! �ͺn��ph��&���v	�,�j���] $�a��j�j����%�9K�z��.q��Q��+�p���2ԒVl���U����e�1�e�3]0.e��T��]�<c�V��!���F.�' c0u!��N���2Ę���#����R����7JZ�ٹE��q�L�	�'։�H�&P���v�󯔳9y��v�m5�C2�Z��>�Hè2�ʖg�����	��_<>}��E�G����{I�rel9 #��3����cK�wv{%n�hp�y6"E�cf{�)���~75� �q�J2*��]x�H�%uؐ7�c r��_���2ge��w�?r������R���dZ=k7��R̒��\E��j*�}<��r�f<��w��&�����"���O�Q،h?�#1��*�x�2�^�ėN�+VX���}c����<�v̈́��q�U�C&���5cWs��b�0P��T�`��l����,��ڣ@w1F�M����������\������d%b�j����dbv圭�N6�V\��tc����M��V���3O�37�\f��5��~�T�QU�<��B�&z[{\�����*��7$�bm(��
ph�q��Ӯ�9��lr2�����ǫ���m�l>�P-|م�g������?�+�|��ͥ����a���MqG�E���W{笘��"��1�O�x�sn���`�T̉�IM�h�s��߬����k�VHz�}|��a�`��&ª���f���!+�r��4�k��n������/��~�{��U{��G"�6|T֍f��~� ��E��3�>���2GS	����"t����՝�R�L˞z���K-����t>�TQ�uq�)��zS�o��C�]��M�q���I��@�۪�>���#��ޒs�Nϣ�Ʀ$X
�`;ެX.F����n�5�������EE�D�a*�Y�g>m#<�)�X�ηL�h�}�*�0qn1o�+�+J�Z�u�&��>�SLTBû��I��1HSh��X{��3���;�9���8g���b�7���.���S)Z�^딦�)����i�'+�H�c��L�u�QǦ|��8�w�G`{�(7<7���/b{*N2��ݒ*/����l�Bd��4��+�� 篱���3q�b1	�U�!�/n;��!s]�z ����<	;�\����D+2/�G�`\�H��/��B@)&<I�RC�	�>W��vxn� s�H���]G�)>�p�T�%*,u��3���P^���Z!^�����%��j�ww��?��jV�vO���Ӯ����D��(`:� �烗��$���	D,��3�hy�o�I�7��`:D��Ux�����8-�7m�i1�l�aO4[?�5�L��ko�^�5/���<�d��!l֖cw+T�5����XQ�r�@*����P� �S�]ܤV���܆5<>��wF����;�,�N����,bN��'o�VS��?�zg���-��T�F�?X��p0KC8����j0���GD�h��G3���?���qq>w��{g%�'�{2��cU������j�#��t��4�dW:�Of��,��b��"j���W�&��ځϝ�5~��K!$��^�Q�U��t>󁟩��r��'�\�D^k��S�*K%<R���������%���@C"�y��cLp��m�XEv|N�����i��z�+nwi�,`fN6����7HŚ⭢����A5�Р�[�����v�\��t4�z&U�hg�LtP��s�,���ו��j{_q��^\ˠ'#�ŕ5x5���/�[��t-]s�j@�Q&�(��~������x�{��E�6��^��kGL�/�H3�.sY@�i*�e��JC�����-�iQ��6]M>�O\3�vԪ1kYvN��s@$������-4n*�$G;��	wPټ爼g"��f_塌��Ŀ���8E�i8��QEҹ�%y�[�%��l���FL0�����TFz+ᇼ6����2x���,��<49ɵJ�J�e�_�Kyc�w
�kc�ȴ`0����t�	K|i���2
K����2�/t�?���.#��B?�\0Sg#8�@�1z����"I�`��T���u?��K~1y�f�#<��y#.��������,ەx���M8I�>iF1�������O�h���x	��}���7Ⱥ�P*��j��P^��0�������g���N��)�&kK)-����aq�Wr"n:����YSO�s�.�f��mr��q�9�LW�ƿV5<��f3�v��Bw�G��ܝ�W��I2�������(�uJx��- x �R���&�Y��Gѭ�_]�cl������F�_A�������6��UBq��A|�H�ȇ���<JG�S�>�o9�q�
�9��T��5�"ZY�o�l�t�-#�C!�Y|�N�n�>��!U��y�*����������؃�yɦ6Y�ȷj˯K�jF�Jq։jE�I��qsvNlE��F�XNG��͝��hy@٢�@!)CJ@k{i��(�Z��,�w;ЇDC�)�T��ǣ��.	r�'��Y�Nt�*�A�IP#�����O{^������M0��UH�⻏;���+���3HH/���kɣ�{�XB��g��'�a����/A��m�@�3���>W��FϜ�8��Pƌ�� H��!���)�	ߴb�m|��ۤ>�$�����`�����k�N'Shyda�6ʆ��y� ��:�Sw��"������;8:�;�����=��6�K�q��m�a���+�(�L�hݗ7@F�e�u������^�Z}�ck�K�=�.2��sL���C6�D�w���п�+�[L�J[\%_�!,�΄�g^�o�I,�d���l���z<��M4����T����!f�������V�Zf�U����@L��ȋj�E,��s�Zo`�G�v�#皮�VE�=�Ek�. �����X38�%��(}R�ib�~VӇ�`o���R��}dҊ!�á-E��G4�H����Q={��e(�Љsj�g���L��=Q�SG�em�D&��o���z�S@6.^��b�N|�咃�T��t��V=�4-s.�9��Wl�:�S ]�2�v�����~f|0����k͕Z���}TqS�&��>���ޣ@�E�Wr;�ѕ*h��
�b	���PW�}p�M�LW�Q��o�4�n���9%g����	$��ѦXҫ����8�R�90H�Z��uI*q	3�y$c�?-��@�����\	@t��W���/�D*�����u��@A����p��Hec�Yin2(�HeXg����|�L�_���Mb�S��-j����ǹM�[�3���]��3e���{�K����xۇ�ޤ���ͬ%(��4���
���@|Ҧz�S�J���I=��	*k�ܶ��"��l9�ۢƇ�Cz�����4����
��G��b��8U��
��$њ[(ˢ
�|��S1nS�A)u�yA?Y�Hv�������x?qV5�_�744�'cE.�zP9���n��`�ۿ�A�
@2(wG�8��	�)���:� h��1��&Ʉ����A8�~���N^�Hxb\u���`� ��\�����w17X3mb�znˉ(̤����R�:Q_�K$�'�į���*^�%K�9Uמ�iuT6���Ĉ�&Y2�T*4~!��j�rJ'�XK��;�aU��ܕ�踱�c���=>w��-=C�t���࢖���0��cM�]�Q�d2���1Js����ը��涆�Sv؋���ɸh`�	�fW����oh�]�E�����-�"����zT���×_�M��nu	>����?�֝��Q���r�$x���{,�[幋�Y�Һ�3�]+֑����Y�ni�M��
$s�Rzcf��};m^i�7������vQ$����0��/���K�Z���}�r��P���P L���U�ҷ
��1�fVNH[:Ld��gq���QD��%�\@	&�;������λ?*k:�6�Ly�D�d�-��B>Ʈj�iGZn�S�m���VF��+<r:�4�.t(�9�[�Iz�E`�J�y_�í1@��g��U��!C����ac�,�.[��&ѣ�!e���l�_/#��8�������rK�Hs�+x�z"�����8��e��>��t����(௪	�[*�za�>��2���-ҐM���[��G�ʵ��[��?��5�W|�;z�Z}rO�[�\�#+{M�Yq��ҋ?��{F�w���=�4W\-�C����q"b��	T�Z����g�1�����Xm��6���a	�G��E/�ҵ��[d1ϯy�ˆ�IC4@�G�`�K&v�y�.�<�h�:�M�D@ٜrP'����x�І�l`�1u�jx�B4UNL�7(F�/�����av+9�l�W87h��cl�M��1|�^0*�=����#��i��xܪ��?����n��jb-Eq�o���\U�[� �W������7���u��\��H�[�E�%Ȍ	�pT>�+�b��)�^q�!��O�i��|J�UF�ź���P�N�Y���1��+��-�),�A7Aۆ�(����3;��ڟ�塤��s#@�0��:+aaO~i%��h
���	�^b4���G!s�;�<M������qi}Oʴ�m�X%�NX6���T�-��f�(�4��w�,��$|A�­gD�����ƺA۠H��E�Q�m�MIړ  ԣ�y"v���V� d�ȵ&C���Z�"�qT� <3ތ5$�� e����kG��L�Eg�QR���*��Ҹ��y]���%�s�UYz��� ��?1*3�Z��a�Zt�Wj��.VVq�䩼���bW��6��HBn�f3�'����	�i�nT!�q��T5ε��*6D�����;I�>:H��[�C�dNj�fl�N[�S��sh�ncvU;���(R���Õ��d���2QN~�����\���=�'ڇ-$k �$oA�ƶ��K�ve�6���Ҍ��G>���G�3�6���������q��k/'��I���F��>�L�:��hO��dE�ؙǌ8%��`噅�\S�� �kl��d�_�ĵ�%����hL����cE�����XEfw{��F<��h�7��ad�3�߻v���h�(�>����m�O����Dt��fӊ|A�'�JF��@^�,/p�'|��tF>�al?p	DJC>"mR��!�ې
�v]�?#k�=4�T��0ه�`�kھ�wEq�g��'_[z^�Յv�t(l/��JI�Q�����O\٩�q�}8���^�*�nw�?F}�8�7]�x~�� P�.H�(Y�T='f�=�Cb����^�AP~q�h9p��'��AW=��b���v���W�y�Z;	oX7y�v`gGg_8E_cn@psv#�Fza�B�r�{�6��)g�y�8�"���)�1oV���r�!��^�V��rl�,s D
P~N*R��Q�
�]�8�6|>�Z�L4W���K}�h���
j��H�������@op6
�y �/IN$�4�c��+4��Eo~�T��q(�Q��?KW��s�R�o��9���hOE����������'��}c��K���\Pg���I�#��Oa��y���Z^���F��S�dqu�^Cַ>��^�~����Խыd����������9�5�S}��J+T�4F�Kt���S�>囈J�e �X$r�6��-���;�� ���{�Q�����30>�H��e�G׮����(�~\��m�F��9�20�L��9�8C�#� ���|G�[����!�r�A؎0 c��d^���oP�����U!�,���fەo9K-�H���Љ�뚽�8+�����\�)�"I[s>ѕ�E����~�D��p�	����7�m����8�)�N��7}Gv>g���Γ��s���|���{�N�3���A%��Ç�C�������JɂU�%} ��Uj0�������u�ds~����a�b������m|��v�����=ρ�*7IR4yQ���ێ"�h�6�f�M^�T�1T�K���m�a;�#%x#e�'	�q] m��)�@�o&-��@�?�mE�<Xގ����`�gM��� ǜ��Qv�/\=�G��FB�T.����Id��㟆L���j� ���w�G���UHi2?0��1��
����s#�<��j#k���<G�ʸ���9�`��v�KHkK������H&��g�P�s���c���dL����=�${eXi�n����� �:W��`��	F��i�S~�I�\ӊ$�����h�"�XMct��iB�"�v����/�vG�X�8��;�\��ȇ<��V˲�݉7]��!5�wC6�1�۴�f���\E����l(d�G4 T�|{HALw�,�z���1��{>�#�`��4�,�Hl��
���,l+��W�;��P%3ԓ�DU��!,��t����xQ�DaĤ��Q=����w��s'�@^.�l��/p
�[b��xZ��t �c��#2�d�ִ��;�Y�z��+GMW�\��~M2ԩ��}�hA�����_Xt�}NS��U�pԄ�5�U�h ��\vOS���׫���Ze�;�~��ҽ����/qv��C��)SW]��c��s9��{ltU�v���}I�S��@��)馄���l%R`m�B�m"�_ӨS�PE�U3�N�!��JQN�璻�I�f[�t�Y�Qm�#@�^�����i�m.T�l�ƞ��Y������ؓޅ�#V\�&���w-hu،wF���d��f��+���"�OV�#���p�Q����/��|�>��G���(j7��RyM�m.Nj�.��n$��1�~tl�Y�C���%�K9C�X�37#�L�~�7�u?�Ri
|� v��1q��g������C����D�2���gEų��Pɝ��4q?�
m��6�#��R�QG��Ht\֎2�c� �~�s�
�ݱ[����b1�eyРJ��4���+�> {����$��3�n��e�"�ڸ?_J<�u �:�(Ux�m�֮�x�&i����kwG(K��(�̮����9���XfS�W�a� +3kbN&!�<�t���PC�xD���"����hc_�~�.�a:Rʆ�	�};a�`�U%�1�0��I{����D����ƈ&�oy�<Q-NwV�a��h��9!T��\L3s�2j�:���e���l�⡅$�0~�f-*'x�#':�v�jx��e�͑��)0�9�n���I��Y�͎RO=�>r����1mM3��k��$��	�?Q�R���O-WT���8WU�]�s"%/*7̩�@�Ͱ6WL	��7:�oJ/�l��h�Ǳ��t��p�+�l����Z�f?����b���?B��V���Xl�2`��a-�pn]�-�iQ!�E�������-�x/wɃx���0��r�����o-.��r�M��y��<^�ԓ����u�f��<M0bS`,y'cz�2a�����ZU�,�8It�˔=�W�ch�d~I��3?��|�i�|��|������4���������dFH�ԯ�-�?'�F�Rƛ\<Z�
�٬ ����{�:m״e�,�ؘVؒ����<f���s�����}2�Q悾.�W���6��	�Z:�RG����bB� �x����ԃ��@n����3V�Ѕ��i��(T�������8I��U�bZ�ꔇŻ�=�D́�Єs��_X��qX��B\�GW	a%v��N�s���)~R���k���>gJ��{��<�|���տwj���]���)0s@$�u�z+o�Sû"kz����d�l��:W�Q��o���T(>���԰,5@����������M��j�=��#R u����UV<$�M���b����LT	[�&�q+<p� �q[�5�#yw�� U�i��̬�_���܀�x��?�n���yӀG��%ݱ���^�)���㾇�T�ΛM�j��*,��(�P��c��=�{I�q*��J3`��G^2*�C
��WH�=����D%2%0������[�6n�L�vv���$�!������nR1yQ7���v��C#���"�nx��F���d�ۢ��^�w=�2S/N�<���Q�aY�.v���нs*X��Q��.��PAL�8몥Sj���_!�c.O�g�h�`����x��!*ޜ�|��.Sx��F7�TA[�7�gv���b�k�%�k�]�%0�ȝ�^��-/�����Z���dM"<=cc4�i��ь1Bꢶ�rh��2o�����I�H�&�����%$�ǭo����)���.q��Jr�MA�6mj��~fF�佉�V�L:����v�n9>eua�`�$������Ǒ��5��"�H�Gq�N!M���=*�Ha�e1k�p�n�s�<�S�K?z�Rk�=�C�q���y��{!�nFK� A���� �?"q�4���W��}�j� ,��RN�A�@-遀�`�3L��X���6�wc���[i�4�������\��q�bh��e��72�2�@6W,o2��A"�.��<��?[�����Ϗ)�*\�/A��33��h,fդ跑z���x�o�J_ь�Ӌ�A�L��ߢ���J
�d"dE$�|��8BJ��7E��hΫ־�*4	����T̙x�R��ǥ�_ic���:p�u�Iy����mӑz��R%G����G��s�Ξ��ڪ�]���v֔nֶ۠UjbNx�X���Hv�Rך������r�I�F���F�r"ٗ�t�6��ܴ���b֩���!-�"���X��ʚ�g����7�H`�n�S�2!�l��C���W��+n;��������H��E����}�|37��Hj��#B2r�TѭK�duA�
��敼�>��x�v���׆���^6�7\G�A	a�GF�[�4�44�] V���H��\��ks=�=`���ʍP�RrF/�uo�۠�62�`���n�h��>!��*П�c�3k��(��b��xt�~z�Ǳ̌�`e}�v@_.$l��rA>�ߕM�X�V�F��=�~x����
��u�3[{����.6Q�B�o�l��=|�(�A���R��^M��� ���Z���ySJ��e�
4� �����)�7r��,��4ӿ�b�#���-�ZH�PˁHp���rx������>���-����\��`����;Xm�%c����:-�F<���y���4���ˋ4�����|�6�`'\��cr�쯎��U��8L��)ʾL��>U7�3,�f�KSΰ��vŬm�X��P1���"�ևUqB@I���p��q�\_�غ�oHԢ�Qr '��۱jz�3��+ޥ5p�Ȍ�4�ܩE]2S�������Q�����"�N�e$�&^ϐvC���y��O����:��
{��3��r�j�6�Պr#�;=Ѓ�/��D[���g��۸֬#pvm ��3G烙Qs^���M-�klw����{x��V?cz�.h'P�4�(̠�!HV���a	�����zR�&��'t���~�!�䲱��o�p�������˺>y��t��9�c��9�E�H"���ư��� ���z*�-�4�8���
�p���=u�3�.�6��رF+�����t���e�ճh,���HP�����l�<��n:a�������q�kF��@^s�B���[%AE�c1Ҙ0\a_q�&%���N{������-��&":���n�L�(��2�$wΒ��>c�8h5%R�[f�C����E���W��Rp)�$����i����L�+y�����2�0��b������3���O�C4�'�C�Q9����ɱAK0�O>�h?�t�?]�RR�j�*�{fqb,bK�IU����9G
�EOL�9Wkg��ѣWa^=カ?�KLD���Hc4��CCz��%�tª:�U�\�E���\��u���a*�u�B*��.�C��v`h^��g昀��S�5'~�÷���F\�h��a@a���-�zG�����M�U|�P�ª9_¦�c�Z�͒�rtƙK5Ti;��o�9��N�(�Cn�vk@��L�Лv{���qz����р�E?����!�pl��܉SƔwg�0Ę���P5Lck�(:(�k��_�T$���x���)ʇ�*oɛ"�B�����ٲ�Qȩ7)�h��U	E��!>�����N<7_�w͋�-�`��?u-���|H�X
<�eqW�JxN{�f$@��1�
o  ���� *��G��Jj��<8��
���������`w2���F��ON�O���t�W���Υ���s�0:�ni�D��Nx�?����r��,G�xק�~ �f`"9����)R���Z�C�<r���aN[�#�z>i�<i#�rV�˽���%*, �`�>PJ�'Rs�W���g��v� �<��v�y�p�pN�tk�+�ڊ��X�t��c��Md�(���̔,��E��@7�9:��~ٶ��24�!���i%��%��)�l��9�_���tX~@F����J?�"&FIQ�u$���G���0�8�]_��O^M����x�	��E? x��:c7���Q4���o"��"_�l$0��Bf���Z�oG��)� ���[�Y�~a��9�^$�.��l-7%��q���>��I��jEi��b�*��ݜ+�j1<ԫrL/����h���zN?�P;#4�g�!�����x�����h�D"ׂi,KF�4:���ªH�P��]`�4���������WJO����q�?�CE����iR�������I�La�$���=1Tw�I!k�A��r�_Ԧ�l�=\�ܘL�P;��g����p�E��w_�T/�Ir~�'wz��ֳͦ]��&~�<����M�oP3�s���>Ѫ�u�Ɂ�F4�:��=�Z�l&�g6���6�M
|��:��bo������ۀj�
'����~Z7����^���v���C�Ί���t���)3l.vD�#�F_RtĨ�$��G�dY��M���(:�]���Ou(=������lMy����¹7?7i�?ɴ��>�LH{��u�*%���OW(
�%��/k3�`W���i�����5�`ک�v
�g)��ä��8��W�)K�P^"~[�c?�����B �1����g�S�JVъB�������2�7�l�:6f�dP�x�qwz>i�7csZ���,�+���m.�����~���f�0\���u9�Z�҄c�4�k����r�}ܭ��hO�H�!1�B0 y��U���5W��xs�+�� ���7_WjLs=�i���qz��uU�m��Wc1��r-�M]J9����/��!Kl)�Bw�3�\��	+�@�Mx�1�@��M+i11�0�Mf�,��:%R�	�_ ��ڪtr(IT� ���b�������ܗ�?��c�Ob���3>�b�S5����?B�r7�4�� t<�:%��ꫢx�@eIud�,�[���;���s�_&jM=V|*Eɍ���f��ָB��Wʰ�R@�&�?\�Dg�u�.l���+���>����^:$L�[z���~P쑞ڐ5�!���X�w�s�{�v{a�Ta1�u���Q��P��D�q�]>9�	���e��#D���	�S rqMiV�]���۩�!�h�͍ͳ�������e}�ۖ�ݭv�"7$K���:v'�b��������	�
�,wg`������?�n:Lf�T�S�Κh&���a���Pa�����Z��N^���������q--�p�V�`"N�|�����kBsd^��Z7�zl�~90�Z��j9��n��p�-!�!�L�i��t�;�<|')��놂$?d[�w��F�,^�-M��cHya	2�aB�_�Ebtf�����j:�����9�N���'��� d�)=%e�w���M�o]LjzՕ�V��i��H���v��ZEk!�A�.(�~_���ګɫfT���F`o"��&�"�F�H�x§�p6@AO�N�!�͙�yQ�Hi.r����b��'��r# Ҝ��e�����۔&'�iI��X��c�3Re����vmȒ���9:�?+92��c4�(����(��[{-�a��L�tΌ���⨯ݙ� ���*�Ndv��������]��#�3N�"���PZ&`�$7�a��} (Q���*��v;��g�%u�KY��>6Y��X�o�
�a�.Kv��B��n�'��'�2�5��q������̯f�&�l���[���?�nO�R1�>��фK
��d�r20.�KR�X�$���6���~��]���b�����w�9M��Ԙl6��vN,Căq	���3;�!�3����oK�����OE$�g�M���3m�G�ZA��Go;�v���r�iTZh�2�x�勀��
��.���v�����4`K���w�JQj�
��K�-!�a?⎁��7�����[o�o~ӅG�2�s7��7���)��M�b���-`RӁ����q��L���-���T"o�����w�
��1l��a�Q�5W����'ĺx�B�<��3;:*�!�16_O�yIP��>�i,|_,�z>��2
�B��^'�{5IqM�CvQ�z�y?M@�7ߟ
&�/��%8!l�O�^ӫ*��Cb"�rUi2���ڼ��������4xu�U����,�G34�VxSY�O��,�B84���qױ���LA��n��{qCx�r�I�{�j*�U��ݝt�n�� d��jq�Ju���KeC��VX���i�9��l�2�,�.��w�+�����Y؊���ڝ`��yJ�XD+�+��x�̾�r��]���K,.��!��u6���y�un�Mү=_���(��`+�Wd'��(�����F#�F�����he!U�[l8���Є��j���>��X�VM�%�:/5�H6ǸH�ه��<�g�z���0_�<�p�w#�Ą��%�û-��l}ņ��@=�����-� �S���i���L�h[�Q���A���-7کę��W��S���(f'oگ���o�Lz�[�-9ߔ|]��_�#C��j8J�h��j�$�L������*[�	��{��qu.�`�j��c=��J28	b8��W2C�m��l�ص|����ށ�5�:WE�r٧��750���N���!2I_=�L��M&�pV6�u3f����h!����_9N�2�w�HǢ��o�Dtxsh������(��a�Q��xlؿd���s-Є!�������FR9ӭ.mD�!�OO��OE�mq�l>�
X����'�d��ʱ�y���g��Nh眆�o9�5��y2�8���;Ғ�ԁ��$��|P���Pn�8��E]��ɓ\T=r�Y�0�z�6��������D��E��!}]�P�$�qi��ω��~��O3A�e�/���P<j]'tG�p������}��ے%���hHfV�OC�ϬҎ�Ϳπ���X�C��$H2��
؊�S$���:>�v�ߺ2��W�Qϓ⑗����c���#�ؤЬ8�'"/{���~�xy�T��?�}�Lw�̗FǴ��Q�h�ݚ�5�hߚ0�Z⒜�m�I�������zۛu�U
L=q��	:o�]�����ܾ�DmQ\;6�nӉ1gV4;"��t�$�8�-�0odP�<�_x��X���[M�����).w�vs�sӼ�=�)(�r�dT�� ���#RX{F֛)��`ї��K��P�c��J	a�=��W����먔�1���&����	���3)�oZ�K��F��k��8u�����c��J
�%��ª��w!�Q��H�4��J.ȊKԌu�EkD�����3�r�(C���a�f��Lyi����]+��{�%�)���w��T�_��J��ײ���6/�T�U�_m�[�2��5|�1�¾��q~�'E@�j��IƮ�Tށ�^�$�����pc��_ĻFY=,W�a��m�6;�������rF����B���:�s�Y����m��>�qU��& @��~���ҏ�u�瓙7�q�&/k_�	OM=���̼�z"��e�~ޔ����,������&$'ͨ��S��Sv4�i^�1���$�I�~}��?enR6����xk-ߨ�g�&a�`P�<����^��'"/~�l&!vnKn��=G�DlKt�yw�k�G��Im�U��T2-�LY���_�йm�"LcL=����޷4��uO��5č��pa�S�C��?/�kJ\�GY�0�k/o~��m:���j����#��(�Xa/�Ra��ʣ��JÕM�H��
A���ԉ8��W�뉧��L�G:G+�5������TB�]8�V�O
J�Qڇ�����i�\�+��[�#q6�u��*Ǖ2?�Fl��8�÷�'B$b��h�.n���;�����3�����1Fw,�����N�u񏐓����y�b��:����^#Z����N�R�̼�M�|�HcEL�|'��Hi*ﻲ%�����9��/���T�
s�cm~���)z�*pͭ� fJw!^P��,����j���w��
��U�T�����g���3�MF�TXrc�9/s��0>���@��~v�Ydڥ4#O�DeNYq�S"`%b�=2KI����3� 9�����Ǥ$3�>&����lV5����桕oG'�C*i+Up��8	�@�$P�D0����J�cqŮtDټX܋�Mp��v6�nx�9��$�H�0)�/A�c!�ګ�S ӓ��n��ڏ�������k��p]�0�Z"1|�i�V�T��������"��7����f���*p��G��+~��$�AjccSI3�k
�_��Ǒb����(S��>Ѽg�����K֎:w�
�^=9>x��(]�1��um/�y���+��kB���MKX�WH��|{�=)��R[�\@�=�_WJ�k�������zP}��Z=�L��;��8�6ٱ�g�P��8A,6
�`�u�z���#����D?���tcrY�e;}�,�mʙ}
��t�~�tR���,�LU�?���_�V�>��o����6]"���/�$����!����!K�|�J69Y5,�Nfr���3�D.���,�7���?�I��?��y��X����9{�<�tQ1ϵq=<�:O�-��Oj�o�d�w��|7�;'`�y�H[���f��j�8X��;���&�@�uzT,Ϋ�Jrs��"m�>3ɨ�w�׳�4��f�ts�\�B�=�9�ݐ��dk_С�Ǡ�C�p,���S1�G�ὲ.�j!m�6�C��N�V ]Cp��E����F*HsSe5}]�����*w��v!6���e��pF���F��V��2J�˅`td&Z�%�z��:9� \T2j@*�\Q--�M�:[
�d|n�l1w(G�>���L~�m(���'K��R)���X?"�@Zcn�,���僽2��
�[��U�:9�}�ng��2������Ԫ�wSHTO���e	�{{:{���Wo��2����g��ٹ}��$V�cV�H#�����@,��kG�|�4�?���b�F:ͷ��񲨑�`iR�g5q]O�F�9��+ƋV�xź)�\���u}u�d�+�>م$�GSXD4U��#uĀ,�DM�mwI����^R��5#����v(8^_��0ڎ�!/(�ʷ�~�!� ���٣�\"���$q]K�Ãwu�e��
 �� MhՒЏS��ꣿ6�E��A��UL�e�.׀І�Y�kbqJBI4��P�3���S� ����7?�i��ӏ���S��}�k�]�kAJ}:��	g< ������F�@$��d��`�Gv�3Z��m$IfUze�[�7�xo�&
�4�33��/� i?G�Y���\.��	�pbS[��Q:�0}������/�yF\�>]�o$�������"��1��{$�<�#M��*L�X hu�����E bj�P��T$��U�ʪ�7rW:�]��RvXf"U�`qǵ] �^Z�; ֣���pUReB`�e�n��[���X#O������.�W]D�W��Hy�>ʐ��oaw�a$S�� K�Evh9l")1��x,r�� 6-k@*J.���Ѹ�M�����������J�2�qp<�<�{��'�3_܏2���?I��`���<���4S�Z(#�}�����#G0g�=|�ɾ���r�F��sg��PF[Q6p#�
�@�����D;W�e�����s�� �FX#Z=� `o����?g
����D�}�~�z�����>T��П����9�J���J�\����0�j���V�I�Vd���N&���*OS-��6)��K>�ր5����cH~�?�sVX�=�}2���¨�a�Q�}_K�GG@f�J'AmLA-���B�[,����0q\4�
8r�4�.�{�;h�����דf��� )�k����Ӟ�Sz�ox��
�k�<t@�k~��N������7��&��z��s�����v�wm�K��Χ��6�R�Y u>�r��H�_VW��C��i��*������<:T23e4�[��ߛg|�)������槰$IP5%8��k_d��s	����Q8�m�d6��A��ʳYK6��ڄ�P�I^�&�|(s~=O�竔(�[����^�SB���r¨QsD�9��Mp 8�=��~,ͪZ^ה�=��e�ß��Ҡ5&����o���a�e���\���aW��}��/7��!a��U��yOop�-������_a���������ӜF�@�4Ҁ�LEr!T-���>�
�a�"YP3����ؚe��VC�hL�F@;��{�_$k�B�ɟ������j�l�Og1�y��-;�
�� ||FH�h��ܷ����-0��e�!m�H7|$K���O�~.?��^�R2'=NP�^<$���G����s��z��g��M�c0�ݥ��#4"Ո4;���q-�)��Z��v����3.��_��9.ۆ]=O�ή��&Ͼ�02he���ϧ�W��vhʵ�E���|[�����<y�_c{�̝0O�l���Վ4#�!��#�����a�,���+�>m\�3����t.��(���Q�d�����D2G�"�+$���˾�d���
�3Z�K� �����������U���V=r�:�^��Hv�����8��za��T�6�����|+��&��(B�5h�!dfI-@�,��bI��ݰ�%�����"�dZ��u�s�%�*�j���y�ى����f�����h5� 5��,������B�n�J��_�Pv�k�C��.��5>��Ҟ-C���蝁d�[��A�Ψ;/P$b^�����ρI@���,!�Ɔ���T�ܮ���,ag~N1Uw7_�d��p��۶�B�[��;�u�l4�kĚ|aB|�͋��ڇQ�A��� V�[�a׻U^��c�D�L���Ï�Mc�ulr�i�7v�R\�G�ć�Iûqz�o.t�����!2����\&��c��Ě �`#@^�3}��k���Y�sU��Y����ڣ'�e��SAmie<�	c���>ö��QYd«�'����s2�C<_��c<|XBd�<�vw>�e4\tQ��Ò�G��omK�oE��h�<�d�=��9/2:���tD=��HY��+�iݠ$:$�ώ:>��5�f��dڭ�ف���Ц�aʑa#k��3@�ю��|#'�B���� �;�Ă��
��~��D�mF��I��
 �["�$�̱N��@nI�B�7��[l�x�ޛj}�=Cߪw���LE��`�����v'8Ѻ�^�@y6��+�١�Wr�<��I�jPz�i�:�6�����]�N�s��X��8$e	���&�
�t�������!�2�}�M�R�}͉���8�>�7P�s�?W���%���q5}�/��iVI�
k���m�|`I���? ɬpS'^�i���F���}�*�ۏ�K��u�v��j�4�����z��������w(A+0f�-```Q�^�0�`pIڌ)��	!߿��ˤ���|;��/��s��h�@����&a'�S�^<a�Y�:3tT~�S<��i��*j�7� C&�߶�����`^x��f$�:	�}�t{���N���g�]M���{O��;|;߀-B�66}`<�j����6�\	LQ·6-��G�F��t�gB�ͪ�o����)o�:kx,�xH�wm�~m���>ٓnTo�&_E२\	A��@���R��mO�3\3O�8,3.u�U�mx��R+��A�Y�~Ȍ/=�оv��Ͽ�܌r���S���DG_�sl{�Qơ�O��9�jy9��=O5�E|8�
I�r�ih�XA�z�x�D��S'��
U���[T�J�L;�o�YRݨTGF5�-Pa%+G4]O�(Y<��B&��#8����]��ؗ�5w���-nm�_���B��v��1�S���5ɯ~r%W~��+P<>/��O����Ke`~ɪ���8�B�*W(�.d��d'��0���|��r$]�*,��H���fT��;*�}�Ι�{_�fX���	�j�fh�������I�3)6��yn^�/d���r&���)H��I�}d겺�42'EA|x�M��L�h���i�N*k%R�_B;$	++����&�¦��;*��ϹoAw]�(�]�xi�{�f����ӄ]��Dk�-APF�[x?�4$Ͷ�P����-te����wk����\��~��ŌL!�nu�jbz��,��Al�IN��v��ז� Ӏ23����
>:j:�azv$&o?�4�el@��Y��ŝy��y��β�D���{�'6o0�b��r:k��]oaÛKf:a7�_B��}�������MRp$��*96�qW��q�{mR�AT
Z7Ya@�$S�tv)�Mܢs10�XT��4�L����"�N��V��i �A�@Y��@���Y��wHbpxk[J�Jг��_�F�7N��s'���f� gLG7(�7��X0��;�0%F�u�����g��5c�~4�ĝ�#��w.�"���Do8����;T�f-7�Pč&��/���L	�UI~:/6��R,���` ����b�^�(홖k����AA�h�d�4�5��E�CF��{16���*�n��Y�Z��-��7AGީ'�)z-����@&h��W%p^IJ��a��{��=�7�$�S��j^H��f��Ⱪ�v#{s!]��i��KuT����<�ĸ%�C�-VV
;L�AO<h���Y��o懗C��X:�ۆ ���3�ޗy.� �吓:����ڣl �^a̩�X@�D�Z�tw��q�8�q�#�6���,%�޹����H��>�D���5��Z����kB/3��,���!�-��Ê�+L�O�AN�}~N�����ߏ;N�K�7Lj:��?Q��ࣹ3h{i�Y4�G����܎���&�.�C�@��ښ��G]KQ'QFdeK��J���hB�g�g@"	N9�-��2��U-�8{�@���$\��v���Ų.a���#c%�����v.�'�r���Yj������Odi����6�F��� �2%���L�V�^����%��r�hE@��v��ءwX5�����
zS��؉蛠�n����Bs����*>�׽�}ˤ���x���J�0���ا)<T^YI��*�.���8��ͭ���^��^���)������i/���<�Eu�u��Ec2#'ڰ��*�?�.krp���G7��6	������v[��w�,�&Tq	Ր ���4fR�#p]&��Ow{fw����!f:�Gd�?�ec��.��ڱǴ��y ��WK\F�	Z�L]9����<���fC'�X �P�<�����Cyv��f���w+�u�?8�^���	+��g�L��*�����R���F�H�[ '���6�%��|B��`�=ء�"l������^Ŗ��:z�gN�x��A�pa(s�����d4ɘ��MA��S�$ZjuS��:l�@���{4�:��h�5LuU�2���k�/�K��
�O;��ۣQd��p�q�) ���~1%�3�"�֏�75&�]Q����W�˚���ڢxhvo��e[DD�J4����٬��MGl�S���,t�:,���Y'����"iמICK�j�>��_�6�����6��\'��%]\f���#@�qM)H|��Dv�2<�	M���1�+�dĢ%~�\���\n���w�IȮ.�M��z���/���<�N��<w�J�����b�\�-�4���/���2��~(�,��?,��Y��C�� mRP�H�ee�^���V� o7YX4Qa*2����C;7�oֆ�O|U���Տ2�R6S\����3A1�J�Q:��V�/��!r �v2�5���XԄf�$ZI���|�k��[J��>�Fԇ:n��Έ���Bgm������fM��z����K���Z~_m,R��-(������������rc����L@.�MJ�r��T�']{���]H�9$o�Gu`��+!���|�K�R��W������z7�o�d盗4|z���@sE���P�`���apпb]����E���:�_?�S��"�<�.u�� vʳxߎ�����qx���o$4���8��TSIb���KC)qt�ȸ����7��A�����8a+&Em��:У�']m�T�+�	^���S��C7�I��GɗJ�	�[Z�h����ȭ����f�Nsf�%�.����뮝L��%+P��C^ǷB�zg�V�{�A�AbG��dB��o��E�E��y��	�P���G��YJ_����wϴw��P���r�J��G����
$��*Z���v��6y�yCp�6�Bf$j�V`}�>���G��t����յ���s¶#���?�$��J�%=�Ԡ��G���B����Y�"����{�<Pf�BAG`}�H?^��D�ﶩ�,��m)d�q��U�i6��fH���	�ʲ���pq���I���v?�x���B�P�q.s�0��%`��c�����G����MzvfA1�wS/q�+.]��F'wF�^�W�����я��K|U�(�Psx���V=�EwI��2��dS���O����IR���	�gT��'Ǉ�>Q�I_F\ɉ�
TQ��HS�0�JQ��ѷ�A6(X��晻f^>]P�cc�\z�<�FY�S�1㣚OM&HShU�vq�K�;=޵�Zcl�,��[�p[=�Q���
���^�+�B�nH��/��M�N����?0U2�'(W]�M���е�A��5���o���`�(=U�|�{>��v�qYP=ՠ蓚�o���\߯2`c_b%�֟9Q�U��1�T����ٹA1��V y����;����_X�?@nmx�>��Q�;�eD�f�y�F�5�D��q'��VZ���*��Cj����
Nl*1�������w�~ie��Nu�S��oMq��_7��O>	������}y�'�:M`�p�$iDv�J`�a W;��o,���	C9���hZ�x�rٛs�lv�C�!�� �h��r0��Z5���A���ga�٠�;f�/�ʐ�<�����9W"Y�hO�핲zQf\�J2aQ��$���A����p��c5������D��p]>nD�<6ci���t�M��WuE���k �o�{�\�z�1v�9�e��IRA9����M�H��ʈ
/�S��P���d�"������^�Q�ۮ���_���6bGP�9��LEnr�N��D�1�j�@��XIC,p<թOC�B�LQD_A@@:������G�Xq�x�����,�$�y����H�u�HD+�0�b��g^j�R?����5(]<��t����e���TT疯�M|��eq�۵� �X����u?�|�W�T��{����7��t��`�<���nWN��~eJ�|�`�W����p��3F�)�c^4a�qMϙx�s;ZQ��~V=���s�}�ٰpϗ������1�o+>�Z�8�ȪpG���w�q�1���J�FR�aj�t7��eիORn�
;����B��95�^��!m���rp^�@��8�D//ݑb�s����A��Ċp�+*e/qV#=�c���>�1�N�g��>:��*��H�.��B*R�����Kb}�1]yK�w]<xO:]E�3�x
7O�Зǁ���iU`;�7��c'u>O%�nYj���G�Ua�0�2VfAP��=�?�50�`(����X�c��S�:	س���q���������!�*j���! _N����
�~�rGL:&�u�1Y���x�B���lY�����'J�'
(M�\@n�`O��u)������`;�Ml+\zt�vP��6A5�F�e \��9��� �γ�`���аg�F��/�b�,�q~�Ս*�׏�xh'Bf�;�]��_�h&��6��CߜA��$��.n�qlWغ�1@ A!F䕣C�Kz�Qe���jߚ9;[%��:��:]��Z���o��)b��[�
�ߦh�\���p��D?L'γ˙�����v9�:�fZ�߉Õz��*p��έ��*ek��s,y
C�ݾq`J��V{^��H��nq)�3����Gt���9����Gռ	����=�e�w1�웑�!7���Gd�h4m^�j��ͫ�ʵ�n�<�_�s���� �_tVF�L�}O������p�M��"eo����n��7f�N*0�X<q�$��[�A1�fzQͯ4���� �E�u����ҁK�-U-A��~A� ?�2��	��E6�Q�W�p=��2� ���<s}Z������1KhnL�����?����L��Կ�\��Hi�����̳����l�H��no� l9��}��SY��f�<h����.c�|'�2Sw3'�w�.���is&O��9�q0��\�ٵ;���j�W!K7\�K�;���t��b�g�|��/"k�t�� %��2���IHZ�xZ9䤒�t�ZA���TΙ_hTbUИ3pW$\SԹ�^�v ��2����>ч��Dث�r�2�)]����t�Lne,�� �[@TMb��Cϝ^|�����C�W"�r�^&Rxu�b~�������-�yf5����]"{�����	�4$��.c�S'��&�T�9��ۥ����ϕ��2zQ&��y�*��Hc�9QL��YI�����x��r*�����vi@CY@O-C:|�*��6�vH��m���pl�FE�ZxM�I��ƃmi{:�<5�>�5�h���*R���q����ՙ!$�e�XL��:����9���y_�-/�G���y��\����^ee��i@I��$���aK_sW�L?	�cW-��^	�*l}���Ka�2ؓ�@_��"�mug����v%���dH��W�I�M����|Դ�9EoF�[^�r@;n�������]�¼��*�^8�NǞ`:�����N�!�Mԇ͜C.A���(�k�ķP��U[Ӕ%��^���#���\��ݑ���#�*�7M�\���#�;L�b���`Ś�q��<���}��i/��n�y�l��Rp��Z��3�ab*��#�u`�_����{�k�����:��b������֕ �XL#I���{j࡙B�1�#4����UlPh0�;��o�XITu`�ۏq%(�+(�k�u��1�T�
�P����	:[�&cܽ
_)J�u�+	��"���6��z%]�.t`hXY� X����a���]e��!���Su'��C���B�x�4O�Ý�����S��f�I�o;?]��t^*����W3��0q�H�0���
�%�P����gQD�R�`@������ivK��Md��Y�ke�
��.�6���C;G��;0o��ᕺ����n�%�H���(0�!�k�ɀ5�F���!�q��̤(���
������D�j��w� &+B�1�N�3?Nܠ��S]�:�߼�Q
J�s�[���:��С�%��JJ�h��fR硺y\$!h�W$�ϫI��bv��h
 *�gb�eT�+d�U_ubn���k&��@�����~0��@/�����S{��] �Ky�̇��l��*���Y	�W�j�|�D�LDOA���6�׈6�CN]+�ȡ�����u�=T������78�趇%�p�0�F�ڷ �n>�?3򙁇֎���$�߲�}\�yeY��f�S�dx*����f���+;�h��"/h�C� c+����;����uNC_x!�h�����F�����
Q�F��<�N��/?��]�?<9fX}'.�_* ƠI��&����;�8����xj�([bBՅ5�`4��)A��B����s�+V�D��(��%!~����7��)Ѿ�X3c�N�'_��e13��ߵ����͸ϲ�ꓛ �M���^�˗�N�쐭ru(R��1��ٶB�g	[	Ju��z��@$��bO��@��#Sj��`[5g��u���$�r����f�5��\�}�Z����B&�pOJj��TkL��o���Kf؋��>a����WϮ1������8�`��sV�L}f���V�Q�<j�FBp�Ig]���0�ҫ�id��nR�
;meU%Cez�4��{C�Hq�e��(���*`�ѕ�G��p��4ɭ�s���l�k�zX7ك�b�S�<G�"K�?�����2Q����|�Z[��!2��th2��
�GN����#CM/�����������j������ف��>gvD���.
�}�����A{���.d{�Z�u�[K�`�zU��baB����Z�C/�vGv�ర�^w��͌��b�Ԃ1A���kK`�ɋp�3�57/(������/?ݢ�+�8 �X�&msC��-��X���gc��3��[=������w�*�IC dt�ZQ�*�I^�Y��ڲb�C��=
D�����H���S,�lE�������A�ߜ����U�H��!�;�i�	��L��K���Q�1�s�R�^  �$rH�@����8}#rv��KO��8}I�P���h�(6���� L���	2ȡ�)�vԆ��n�G��-u[\��)~�@���Ǉ�p.�����"!��l��Hh���}�Mr +���q?��#�o^��R�G��MA��# QՊ�h�P?�a1+�m��}�� #�"��ݦ(�O&�^ʽ ֺ���k����!
�T��R}�01s̶�׌�}��A��B��"i@������d��.����4d�a�]�(�FPC�Q�Γ��u30�i����?����&���S�����N'�l���5h�7V�$�-F+X�ǹ�5=�ؓ���"��6������iw�z�]!Ҟׁ%Fj�{nL�{���ڶ5"�Q�7�&�}�
�FV�:��8�3��fF�����ϙV�_݄�\m�)�6.��Wr����lU�	-���k̘F%Ώ�EL�<�O�1B��9璸���t�z����i���e�/n��k�&'@��o�s�+��5T����-�D�
���{,��a�D.Wg����`?��߰i�9�Ŗ7�&C���",Q7?F���v>�'��>�Gu)�S,�RГ���T��D��f&Z��������T�:;�({�ӟN��j[Fǌ�b�U��,qZ������L����3!�Q�#��:��(r�C�??����B�aRZ�?��<]��:u`΋P|�N8f�	m����p� ��8�A�b�m�����<��6u=�MM\��b���%l�!�� .oA���oW����֤�`�~�?9�D25I�Q�c��%y 8K�
�|m�rZ)�q�"Ǵ����vk��$Hr��B�7��yI���'٠���эKLG��"�mҴ�����29�i6���~T��EpC!t:P�xY��}�\�Bg|�bK�5�9� ����Ry��$�ގ�k���H�D�9��0Yq�
���m�������L��G==7<R0+�\����8�6�#��-���pM���,�abRi���Z�>(5���9^̚W�&�������7� 8���3���K��b���S��� ���+��}�8t�Q�K�o��t�,���fd���3��8�`�˩��Ó�w[����]�@���wn`�T��ɩ�FӮ��� 3�+�D=�|�����_��]��=���r˂_2B��r�vjxW)]�0�ꊠn�~�P�TBi� ��|�~I]H�F��*פ��m��J���f�[�ɍ_@,^��r�uP�K�a@ �3ߣ��#�h��:#�V��u�(��ƨDJ���%�����ʙ$�1lGtmx �u	�.C: ���ث&9����v����0/�b�F-�!I�n8>Y�cΰMc?/6/�Jaʬ%=D��v��?Ě|ڈoҟ>#K�1}�Rt⎛�����q�m��}g1Z��[�D(7I��J �����Jr�W�	��:g�rU���V�o�?����x2��vѸ?�-���Ѫ�9l��հ�(hNN����K�.7��]h���p���	Y`��n��0�A�;i.�Yc���{�+�B�:�6i�9"���h*��ۧ��q�堁�h2>�e<K*VW�2+}2�'|Ʈ��]�2�8�p��fV����������T�]��
���f%��+8d���Y�>I�� ��<x)���|ߴy�������a;���WB~M �Q���c�xf�>����UZ���<����������N����.;�խs�e���e;���}n�kجe�V���*K��� ���p�_��yeX�8�^%9=���6oەE�;F�Մ�s⌇��`��������tto��֦��	]B��:���(R\�(�Vd4�zn%q�&3u��x|���D����e&J��_��#�)�P���-YX��k.�7���SI\�;[���⛘ٷ"�iBW�?a\#���"�A����m�Q���?ڳ����"��~ԕʾWY࿼P�JQ1��� ��
N�P��JPZ�yU���_�'ۏ������J2
M�Yߤ�j�|1�
ܹ�Gr\2*c~���l�)`�"�ZkT?&WT�,vd���w>=��t}��8�1��CyB�A�� Ovy�zwӛ ��<���
�|��2�<���췟 `p�꼆���\�fcL�y;>�tEv�3X�`�Yḁ�{�Xw��u٭A��/Xj����gC�Ί!2e�{�ֱ���W�K�)4Mb�lm�5 �K�������mN�|���?+m	�E�#��뚼(T�6UJ��e<������N��Y�2�>�����TG����lCM�����2L�������^��E��y��0#��\rD�,D֗"��pfrk򊸝�X��J���"%@��[E0�g�6Ѫ�1c��+���%�	����4 �VK6�%G��%cy�ø����,�S���&>jt_ �B�|B����wp���nH��w��j3��*̃5�a!�}d�,�2�:�W����m�ǒ »e�ȅߣ�k�v`ܮ%��'�YP��h�d�����Լ;e�2�2�'$F�{w��of�S���~�9�D +��D���~��.̎w���o��Q��6�(0W��ơ|�[�����d����iH��t�|8��i�;O�ew�ܑqC�I�V#�iW�K���'L����eb�t���갅� ��֎ֈ�G,��U�sS7���7a��(����nQ ��Hh6��;dE?��ش���ѸM{�Z�Vj�����m�ҿA��5Tz�Ab��*�[���A*W�׊K���\�������K�Dp�F���DTp��^`�S00�D�](^�=�q{��)~#R��,�������ХQ�d;���,/}��À_������y~/��.�a��^����a?��>Ǆ��4��4�a��1d���1c񀸽��e`J��h� ��F��Δ�a.> �ū��^�5�oۦՀ)4��_3K���@݉;Љ/P의)�3�d�bVh�6�9(͞}�3W�;#�oֆuq�y�+�c?����ߵ�"UMd#u�����>���*wꝞ�����H�5ZʛW!�7�ď�K�A�&nT��#��0��>�J��G��j�ԼK��r]ɐ'���9����\�?H�����ң�y�Z>r�«U��HZ��x��?Kc�Ŕ�D��vDZ�"��8����T�^�pDN�/�bٍ�$�[(%��N���9�h\(�o�!:��t��k+Ƹ�G�o�q���*9�����H�z�ͦ�2��P��^^�I�^�K��:���۶s��SR�g:�(��I���4�J��u�p�R/��O�fk�c�*%糮���������c�7WS\��p��K�������cB��>%�X�f|@Z��&���N'���y�G�s�l ,¡)�%�	��Ɠc=E�h���O�V�;ʖ�Tk�$_��+".�,C�&u��� ���SF)Fo�M�_6˪XU�!I��Y�us5L��Y?<��í�45#O[]'�9��:��&��(2>��~�/�+=�����|���T ϣ?�Fՙ��/(�^vt���=���ڄ�ղa��K��� B��M��}g=�5D�_ހ��y����݂~���4ב�yں(�Y����D��X�rW��j�6ϣ��#�m��%ӡ��U�rfeO��#�*�w��&�S��0�XًC7C��F؟8�#A)4^Fg
�}�<���f��������L�H�R�O������l��"�O��NzVzg:o����:#��I S0S�BS���T���*?:���}�j6Ҽξh!@J�'5�S�	g-�m�)��v�r���.��1�&^�{	���6ۦ���
��x~nsTB�Z'��
haqV�O�1�4���˕%u��i�`Uܓ'Ҵ�������b潚�Z�@��/�ۢ�.���-����U�6��e!^g_"��;-��,cn��'���S`�6����w�q��\$pY�nx�R�Yz�#Fլ��h�
:�i'Q�CoR%y3��E�:5����y��g�k��@��Dq��{ڤ8,<�k���z|���an�>ۮ��Gq��f(߶D�I��pn�s��L�� ����Z$��� �����|g2G�~y��O�q���ǩ�5�2��z�"c��h��	]�Z����cj3]���B�o�p�������c���"pwjXah�!}����E�:�
ER����%�`wP<ȫ����ٶ��L���:r@��6dXҧ��]��~��gQ?H���c��;q�"Ņi����蒥Xa3�>_�q1pZ��5>���9�F���fF,S�ݠЛ��O�$\&7�w�>?�5,N!�}�q�%+�ܻ�(nRK�-���X�[������x�Ck1�Y�8V�7���e�%	��)��j�
�n��R�2�;k-�Q�x�B�B�<깞|#��% �h#c��|��ش�^:dNő�Y�k*l��Q������j�fFO1"o��n]LMٳ� ��D>g;�Uֵ]�� o����L�^#s�	��P�d����3��]�}9��,�5�L�4I Z����Ec����R�=oc&U9Ɋ����י��[�R����)��d�v��+��LG�����p?D�G�0W�Ʋ�04�����lq���4�ձ���z����1!��YDu�����?};�j�`��ʹ' ���J��9� �ݧ�X� A,�5o��iV�ξ��Ğ�η7�P}	Ż��?�8�\��[!EC,���'�I�'���R��U� }w��9��6p�#�p���2	�/ᵶ{��GNǠ4ӊ#O�s|� ��54��-����rnζ^�s{�9ʩTM3�����f�w󢢏�HP��j��I_e���9f��,�=�O_���y��
c�N�F4ck��o/��'<K��=:���re��UP�����`�o�t��Sh�8�tq�X�*	ǒ2�|�뵦�;Bt���Dw�WR�u�(r�h�	��� �����3"�O����>�:�� 3��]H�4AH�S|*��p�g�Ew������v��sE�8qn�NZ��?��:�X�����u��$^�,����#Mp�ҥe�'��
�{�B��FtH��].-�7�Dbύa�?p��&���-��{]�u�!3��@#����Jd)rC����vK��X ۴�3���U��Z^:�.KK�]W!�U���� ��	�����A4���3a��g�t���8Z�/>���2����>���ؗ&5�( Y�r�� �.]��H��.L�+�� :Z�Ţ�@ŷ�!��ш�n�1_A��
�;H����<�:à�}����#��,�a-�R�
�*D�X�B���
TેLHZ��ePPU̩X��!%���&��_����w�q��YC�R*�<'�-+,����3�N}mJ��G|��co� ��B�eE�魗:3*�5���s G�:!��׬�{�ɡ"��M:��ѡ���x��u�q��P��@U����0���<�Y0��I��'f�N�	%k�}e���Gk����a�Ekk{O�6��L���V�y��Io��1�*������ђ��A��oi�%���^��YL��x�ߡ�5 ��V>��<~�S�d[���c�U��j��C�C?��� 1'�.�Ũ�~Q�����T˰[Kk�q{�T�QA�p�S�mD���{u���&��>�s�&��;�f�ҧFo[�
�(`�z׆MU���aW��x���,vF,A�L�!�_���+�&��OB7�(��0��<]��3F�oܜ�?Y �!n+�z�pI�Gz��^���8�ි��ȣ�Ȇ$� ���|�.����B@)����8�j&m�/��Ta�q�aY�J߾΃Jh1y0�?�ɥ���}h��z{at&o�o�-`���/ЅR������&v�}��f�>��<�H�vݲj�L`S޽�c���u/5}�m���~
�u�.&�~aAж��`�����6d�a��}���������:��C�j1L��-X?_wz}�ܚ�)��ũ{êA�r�e��B[��;J����X!G��
3�����GX�~
�3��Q|���^����|�+c]U�x��1�\��u?��Hi��M�qg���Yr�� JD�6/�Hʂ�L2�_te�W�Gюwy��Z9����b�k����).-���T3��O��'/�b4��ώ0b�7T'fL�f?P,U�����~�~�>,=A��Ā���%���iǼ�(3�mo��'�F��*����q�dRQ��HSb$�ం�yy1*�-���	�9L�_TFCG����v���J\��Ar��e�S��G�ۧ�ol#��׷�&���4$�"����=��҉���Jdenܱ�WE��1�H��E9O�<���B,����R�:3������XBuge�㰷���:!GrѨ���$�YB�S�R?��t����[_� �F�:�@֝����+�$�d`ߒ�+�6�g�RbO +v����e�8*�����]]�;�%`4�Rߴ��MO$���LD�}��'+ry��=�܋{=n_�J��_
q�?(#�Ƌ;�N�kA��DWמҡ�9��ؓo ����p�n��h�/����V��2���ÉŤ�\�fqA��󻬮~	�Rxʪ)�y�9�>5�+-/�w�E�W�����߽��|�x�[��Vbt�ܑ����=��6�f]�>���R��q�%\b"�6`��0~����ꩮ~)yDB^��@%��]��La�������j�Ǝ'��w��w��Ś�����Az��rǼ�=j�!	>�d��L!0�/�cU?��=.ғ�BK;z&���M��v�o]�]�X�b6������r`=B�rG4�p_N�:���`w���t� ���ʱo�@ڲF��o�bo���!
�h��a�`�Kğ0��$�9]��Ey6o��;��-� �?��K��0J�BF�vE>A� -�,�B�3x��4�­AA-v��d.�F��&�:� a���f���c���N{�kg�Tu:H�Kg�tgN>v��fmsT{�+��4����.��k�a���5p��Muz���n:�fۜ�AQ)�ƫ���Xj-�r��ׄ)���Ih����jez��(i�"$kܝ6�����S^4���+��B� (�\�7�[����nͱ��G�����X�/>wOhWlr� �.榯� �p��55�a�Fr�������1CO|P�jc��&�X0z@O�V ��KUh��AФCo���bF} �܋�,���d�  �ԣwl Pn`D�M]Eb���3�,>�b�B�'P�����Yc-;�I�DA���*�����~�y�)EDsF��O�.�F"��$�dQ�:q0�_�e�fr!�l����^W���N
������͞#x-�6�m�� �u˒h`&n�oX�@�����[��h w[��/�R��U�Ÿ���@=�5ME����Ĝ���V��?��I�h7��`m��x���R��������;���s|q���*�.@M�*$~���qdd?9l?B����@%�	��rԂ�4����c�8��Z�t-���`z���9?��U{�.��*����7�ڕ��30#�������G}8�ߥ�p�J?�/�|��Eg�����j��Rx���)�AN���t=��TC6
���x��})�C�:H��k�x�����5�`?�O�&d����z��@N������Wl��0�ԢFB��^�M��ծ��O�4r�<�!�J�R����`(�Qɔ���f�����lVʁ�����5������E.0�ėf��n<<*8Lq��L%��8s�NO�{�CR[�����g"9#WƢ�hC��mR��D��o A,�P�<�HCI�OM�eoPD92v7Pu��a��p�!>R�OK/���^8���9e�4de�سt�=�i1���_�Gu��d0̭|� YV�w��Z�����`�i�-�T�l��&�ƕ	�X��	���+�h	����HzEs�q�ک���i���O�� ��ߕ��*��'ȫe��rz#W��%3�G4�vW�����࿭5��H����7���"��[E�)�)��7�~B���[�$-�T���s8>d��:xc�6*�"J$�+�ʭ�P��GKC���|���� �cat�7t��A��}��˾�jO,&�2����.r8��I4g���4�᫡�k�a,O�����;��0�ɂ�D�ĥ�2;2<���W���=qCt����rV}�����+Sz%�Æ��oͼD_6���-�}r�o�q:<& l,�A�'�Y9������c�*����7{��.O�?�K�r�����'q�J���(L<��g9pA��91�V�V����,S�J.��O�����B��Ժ1(��2�n��zd�[�po% ���`xGO�_%�&�,P�q��}��eʚ�d�����d��>#S�^t\hJ�8!p
�L���q<͛Ps�N�/Ծ�:��ɕ�/��7M_=�=��d�#^��a�(TR_TZ�w�/aƞ�O{��� �I/q���X#��.6']��S��8gڹ(�v�&��mA�Bδ�M�$�WN.Z<��bn ��+ˎ�ȲJ�d��U�	��t"��!�����6z��q�r�09���39�k�~I�[<�k���=��q�t��^t������lJ�M��jG��L?��H�:�������OΕj`�{��?�#�8Y��Uhr�Ǫ�9�����!���0�޸~)�g!u���DχdΣ�k9
1����ǂ����dKz�MI8�����~g��lO����0�����?^z޼:�AN��#9ӗ���yo$|�S)���Ļ!�m�X�$�c������R5z��R)G��6���`L\-�waoKl�H���R��秼`M����1򾘙Ҫd(�a�OY_�Ug�cPo��l��qV=��ѧLImm��N��������.�3��T���&# ���xW>Y]�M#{}��P!hM<��p}����� �_���|��/���������pu�����u%�10�/[��½04��?{Hse� �fXLc�	��cM�/��^e��j��m�x!��.���X8�~��~��y��0��C5pj�B�H"C65�����}��f�ka���)�����\4���E�M�
v�!������g@Ձ_tkA5$2�J��tC��zu�_�U�=�$lu��ڑ9
^�&.e���+��4�f�a_�y��n���_��B�I�.W��o���ȩ��F;wv���U�]�%��
ҹ2�j"��2�aMV�nv�
>N�s���M�8?7�}e��M�+it���ah��@'�<�}�}��S*O�&|��a����v�7F�=,��T<̳:־�U��3u�V��w�2Y���@��Ru�=Z�)1X\K���x�R�x;ڹ�e�I�![h���S{H��	�������7��9���k�~C^�q�j\�骶ő��f�+h!�xO#1�����LM3�+y*N�1-K'[ZjϮ�}�E�h�2?���
���o�OC+e�N��Mnj$�
j�wM����V�`l��u�k�N�#���E��F���Y��`RA/�ch�l���[c�b\�K�o��WH/�r#����&^��7�LH�t��=��zLMK,9/e���xn?�}�p9Vsܝ�`�I�(�wOCӬ1lUF�Q�Hh�>�_�	��)����'��V�.�è]5f����Vn���vg-^�B��A͓����u��р��b1�|X� �&]�z��œz�.BX<�ϑ���eu�hr�����z�hh�/y~�s�Q�F�\}�W�/�%- ��a�V��^�xpQ׺�U��:vϡ �T�&�@�'����euֿ�9A���_e�Xؔ�[(��Y��t��y��{��p��Ix�zP����f�\0���7��|�>7ۖ��5�r{VN��>a��_�����0��d@W�o��;�N�É2�hJ�
���=-�����*~�1�C3����Ez�^��yV��(�[e$�Ӑ� �:4Ҭ=��x�����f��whca32xQ�����GP(�e��h��c<Ta_� �Qy	�79�$�$(:�y��7B�����������Ε���7�0��Ŋ\��GvO:W�0������ť�q9�Ӡ&����sK���>H�!m^�]	jj3`u���_�e&Ӆ⑒Aʛ�_(�f��%�ov"
?�X7�aZ7�q��[l��/�g���pc@��Ѥ<5���M�%��}|�D��(�Au�=�45�6`θ��J����}F\u�[�;� B�P��:q�rҋ����[aG�����L&�Ý�0 ���}�vx�x��c�>r��A��4��"������[�)j�8M��ލ@�Ԯd}������<^��m�cak|'����*����e�!����|�0���l��lX,_�^kE��7�������q�������$��,B.7w<�]{�4v��.C%�����.Vٮ��3�'a���t��3/��+�<�d}kopz9��9^��X6�eP��? Ӛj1������Ȉ�
M�qX��a����VmÏ!�I�?�F�Gy�7%��ѧ�U�V��]?��䮗9����^��'�ӏ9)S��Cb��v��������&ȷ7�_U���&�mPXET}_>��C@H5��i�ԶR��)��^�"Њg��6π|h��_Z)t���6ZtQ���?x��������V��~ƽ���z�O��� �>4�<g9�m;c��fu�8�hՒ�

�?Zm��O��Ⱦ�ӟ���d�7i��9�k�O����f~��9ݐ�g��>�Aƴ�D�2$��ͼҋT˒	o��珪�y6�ꁼ	Y۽'�������*T>��.<x��n�)�&�ڂ��'��d�P�y$x�4�%y�;'KF`��٥�L�/�i�g����$�����c�vOv[���,�b"�i�kk�y
���͏0�3�W��w��Ӄ�e�W������wcemvA��E�8���i��2T��I���iZX���J�O*�P��|���PiA 3���D �,�:�]?�ċ/���!L��Xσ���Q�1@n{��r裏�AM�k3!,a �u�]�TH==�b�P,�U���f����D��-������,w�:���+'��V~���>��T�1�\���gUЪ�5�<���$�T���ia�Z9�s?�U+!�K\�������k�+��I�ď4�����x�M_1�����qڹ������m��/K�4���$чl0Q�D�0��)��LmV���	��~q�ej���~��n��MG�4�oN�p!� ��U�`�����c֚_W�{�Kz�Ӡ�	����
l�_��`!4�V�[ɠk�V;�'e��E�3[��x�o�ܻ(�x�H4`�%b�?]�F��Wy@�|�@���J��(2=�p�!�Aj�g�moY�����|��m9��Q�V3��� j¥�}�$�Z�=�7��e���pa�*��jt��r*��bȏc`�?��hR0  ~i��=�!~R\�0����U�Y!�Ϋ�Jir���G�5A�ѹՆ!ZG��	�V�Vá�C�ŐN��U_�ԍn��g�-Q��rI�	�҆7��Qh�6ڬ!��= ���%9�L��)\�;.�>$�Td7�����2����xV���mž)Fԏ�RQ����o:�^�ʗ/#@���OX��ӝ�ک�5�����r�ſC��q8'UHч�;��f�yY���8#��q^�����&a����B�\�����
�bnL��ܘރ�O�-�h���c������J�t@g�����]P���֙�@Y��sM��r��w�&j���d'p�t��t
ώ�����t�澖	�QesTO�ަ���'5>>�� �/�=���n����`E��H1 YϰVmb�gf��G������(����0����򁣤Oj�N@.o���.0`*��Y�1ħR��!��B�����J!i!*��	x��MU5���;_<�o�H[�b����^K4�ؿ0%�������j�&&�]��K�Ix��o#�#���@'�08����f�rk+|@po@1��@y���ޙ��N��r0=I���v(v^����O#a� �^��},֕E|p��}Af�x�:,��j��2Z��:�յ�&���ʷ<�lD��S'�Ahw����F����J�jN����i�(��X$�P�<��Ɠf�5uN���HZ�No��!(�~�a�-�A���} n.���ϣl$�u6|����]cW��2`˾%?Pv9���f�>-sp���T/Ha������H-��H�p��ɪ�m��ߔ�dVP����Hl�p��х�܃k/z�ʦ������DTIσ�u��i ���?M�STnhħ�-�Q�X"0K~�$��L!�飴&�F�d��킩���?Ƃ��Z� �|��Ktx%������&?}����jT-H�B �ѷq�J�`$���'��дÿ�r\̴>{v=|e�}�%s������
������i���������1u�m�v2�j�Bsp��P���U�;���0�O��&`�'��ţ�������SQ�%�z@���|�˓&�,L��憳K�*%���z��<����ɩi:�#��l��>�ΐ赣�����\�QT'�@W�bȫ��
�r�5����4���	��+xu=s5�NEi��p������MJm��j�L%%λ�	����@���Ug �䆵�2��#y��=;5$1�Fh{x*�8��h����rv[ܢ��V��O�c� q��-9> D���tVܷH�Owld
I*6ފ��帞�1jp�_��3��N�� W��
�3��n/����+pn���'(���^��
���jh�=�"/�f�l0*7-"��(ۯ5}\�ű[��	
\�b�:*�����������������x���g��~����n��;̷�ȿeN��$����F�Z_V	 7����
���UrU�k�B��k�n�!��A��dQ�a܋J]AQrc���L詷yɵ	��W.e̵f�B�ʗ)=����k�Ǜ�R��5���P>u(a6�u����n������R !��k}�S:�����-ᦜs�ژ�~��!�^���o��Db�����XK�c�B��D���+[�0a�^�u4i}����*��4KE4��'"�f��s��)�Y��R�>��+�8��ŋ(�-?�`����b�e���D�$'-	��b�c�nR/�3����7-�*߂�K�)��og�a-H���q���q��`�\�̾��[�׏�~l��O�{k"�c������;o_X9�w�e�La��
�)xA��k����V��:ӫ۩��T�`/$�Ny��t��5�
��|�l��c'T�K��/���8�?�1�����M��8�x34�22.b��8Өm��`|Mr�@�l�~H#+H7>�b�ϰ>&a�[���ǈ�|R������^#���:ҥ��ƭ]���?3��>%�s�UB�^�)4�����UXS��n���o4�˘%t缡������e_4�������r%�O8��؎�W�x!GI���h���T���`Ik�4�j����Ѥ��%q�`��;~������t��͍��Ȳ̼0���-&̖R������l��J�q��d��QJ����-�"D�%�5F�+�I��QY�Ơ�)ъ�#%��J�	��-d�M{M�Ó��.�CH6����@���Cw(͍�kپ���Hz��X^�	�`��o!���_{O��f0d ӷ4�#�}R7��H�"�W&�LJ���ҡ�9Gk5�Lv1�7c�'��@��2�;����$L�5���*>
A�^�`a��{�� uT��5��8@z��l�"��X�m�m���ڟ���
�d��1Q1A#�����w�^�b�p�+�a"kP��w|���(mmoc�	D	a=�F
 �yb��a�&i([�J6H�J1Ky/�:�'H+��$��/W�@�s Q�ޭ!����x1~},�!�i��pO�Ƕ߄H`q�Z���kۊ�tCj�L��Z��~e˘`��W�CY�My�q9����0K���41�X3�z#�@�(�L:Z#���������J�Y���ᏡZD��6{�w��A=���w�Bf��}�4!��p8Ym�39���oacmC�?af�z�$���q����އ��� ��5���׶���%�ɰ��&�u�	��{y��C.����v��W�c�,�� ���	c�l��\gt�a����� �N��p�=���Z�}xId3�J3ш��$�h��cN>vE�
��xhg^WE���p�� g ������L��t���;�'�0/�6�۱;������ޠ1Z�V
cf�ي��i7�%15�p8a߸��_���C2𜷽��^�2^���.ӕ�Jz��c�ֲ�X���҈��R����IC�i�C>�]�BC�"3l�����-h�i7B���b��֎�/�%��k�;/�S;y�{�O��wuoO���[7�K�.����O��������m�Ire�A�j�'����L�;���.�OB@(p�h1�krX�t�D�=�B*�t�;���5�L�.�R_�����������U�͌����)��;c��(��ؒ�D�-�-{�h�������<����1�&�Dш$E����N�����/*��"��uw�#�SB9F��݀�L�V5�n��`R�I�#��^N̳�w��(��t�
�����B�ОwU�ㆃ"L���j	+�(v�W��>����s^=��@���Q��Aʀ������$�Vۘ�l����M�%ֹo�m;ߟБ=HP1�r�Z}ڜ/?W}X��J��ߞ�����d�~/��!�T�E J�뻯�|�+�k��R��e�;�˷֓�S��:Q��M�4U��/ﲂ�4e�>�j����ދX[`ʭG+����,��:���?�Pm���`$c��L���p�"�벰�N��Y�R>'۸�TNA�bni�8�P�X������%����k�G��|u�d|h�m�r͈N`�ߢ�P�����ޮY�R�����i={ˎ��}�r�%�o|�����m����Ty٤o���Z�D��;ċs�FlR)2�{�S���ϭ�"���ѵ����bԿBX�m-EW�)�l{[6����gx�W�9�-��ɉ�i}��>�HDA�"*_G��Jj��#��{�P�Η_I�޼Y�6��vU!����^i&�8�0�zI���8n��N�D�I�5�̩�J(���:IN��n���3��B�	�K~B��|ܿP[M�>|���V*ީȲ߮����ʹ`%�(A��!()kC�v���g���)9͚L���?�	��Ҋ��+�"�|���Q�xl�1��l&���V�\ �aC���E	�<�΍EGÊ�Lvq�3<s�psK����uao�JBx��s�>��i	]�"��w�OS�P�iu�?8̱ܘ#K�b�X���L7B:�k7J�@J�9�4�eX�2-����5�?$ב�#��#�";W"���<:���m��޼yĹ_�2a��P�iX�nV�k�l�!P A�ޒ�ME��<��\�M���,�a��?zt�ě{"�r� xd"�m�5*�U�v��{Z��vM�S�P��%	2P���J�D{�y�^Iv�(���Y�QG��f�S�ɉ�K Y�<T�_��׃���N��'6���b��M�w�j=٧�qm����$�4\Ab�Rv�gp��iX��q�L@KX?FNv�I�2���i�MӉ�5AO�������rb�\ޯ��;�e�i6� o޾)H'�3Ԧ��lYf)��&^�f��Ķė�����{��/�^�$��H��Z��KnW@eQ���=e�*!�bO��{ �;�ԗw.K~V��WT�l>�����g�g+cZb�n7�wx��ݿA�Q1Pl��B	9X�$˪>"�1,�KW#�.�mE�} N�|��Y�<�qõP�MvEl]	���i0Xj_�ض�Y��������#k�(�O].��X���y2AՆJ�f>5iW�p�����A:4�]��^Y�F����I��d�@~��l�W0Y����'~������~��)W��
f�#r?a��ҭNU].���v@���ݽ]34��0X_ư�>�jY@q+��G��}l��6�3�gtu�o����Z�m��dܛ�Z^O�^���p���+���Q?��>o`�q�����r0^�(�[��Q.�_��S�_�eONЁ;����n�n����-����{?��^����l��Φ��v��&�@e�B�K���kK���Ƨk=�T	4rT8,��BB��
	��u��B�h}Dg�{�֪ح���M/��n=���&�����(��G��-YWk����|�Rg�N��' ƑAS̅*YS�z,?�TIMC��	7�G6+��7t�͐8"�w�����C�7���~TH����x k~�P��m-���
�f������'$�a@WΏh�֭�0j'��&<x��9�|���Pa%<kߏZ��K���EQ�C'L�0���U,	���p�I/��8`��`���	�%�(����3�\\��[�'K{�gӭ�A�.���Mm�.�-� HX騽)�?&�BhH��x>Vrt�Ӎ�;�vON��Y�H@ӢD^��4���O#c��L:�i�E��S�v�;\�+���۔�#�R��+�~�N �Z�]ӧr��a�ŭ��߲��t�,H�[�fDQ	��ùRV(ޞZ���Á��,@^n��tt*���j��P���jZ}�TK+og�)�k�;=�E��b�i縭��uW2+*���!����w�h2?B��u���!�+����7�9.��pP4�)��ƈZʢJ�V>U��?b�p��l��6����9۝αO0�@h�:�ÉȾo~�Ι���c��XW]۽���xS�P�v�sa�~x�5Te�}��	�LMGGM�:ңQ�Z�f������7����ဴ:܁��i��@dI�ՀP�t�>�z� ��]��P� hrҁ!\_KR���E�p���
<{�s����M��ž�$B���y�8"=�Op����]3����3�$�	��&�0#�ח��K�����BZM�̗A������}<� 	t�%<5�$s�oG��U�#v�#ԑ�^��������Y�7���0١�fE�F��4��x���Zn��KV���@�X3m�4��� G
^�،�|�
��Gխ�����$��䩱f��LCYdnrV��=Z`�D���J��|g3E��[�$�Y�L�w`n3n���E��Жa�:UE>�m�؀��[a�����#����Ŧ��LHidU���Q�ϐ�L�Q�B�N�����h]�#;{_i�q�pJ֖�&q��cn��yQ�?C�������/�~w?��z5�*}�	�
��+���`G9|���?��l�O�|YRG���4)����'cc��������4�"�Yӄs�|�IxB�t�e��it��
U���"���*�޳!W�"4� �y�$#��d��o�"��I>��~�y��(}d��s��e�����zܠ��Ҳ���ͽo��yz��z�=%әa�7��|R�ׂV��[��xN�D96B����r���*�訛]O���Mg���/�<�5�(#�;�w��7v�l���ZL��q��� ���mj0��$�Gy��/�h�l����Mf|����^YL2���<����p�W���;r~��T�h�|[��}X<Y`*��u3x�<&�a���vb��W"g��&8:�Zy�%GO]łbFS3�S��5�J(uD��R��= �l�EK�i*�(�k�w�8o�E��n���Ԋ��#8�1EN@�E��D���t�׳�ä�蓼�jp�Тd5_�ٮc�#��n���O����6��뾜�#
m�M�l�:p���`�::�!�����,��:�R�@R�*��7�-��0#���*��H
zd[t}F��b?x|�"�{���U$��-��?(�1{-*�Bs�cM6�>�0�����X��&n�ԏB�~~����Rj��x$���`P��`���*g��.?�I��:$� �&g2݇��o��-z��1���']�)��C���@���̅���hl�ϣ�DWs�S�ʛ�d8-
yN�v�7_���e�z��2�wʷP`��
�t
|B�6�/�s�a�q�:B��Gj�B��*�_!���N::�������n	vuS��&�>>�|1�@�z������-P4\M딸�̫�tju/i�x������F6��*���W����T���ɑ|���lY�eoT3e�
��1��ca�V�VS�xiDs�}�{�"񞏧%�@M�a�:�T̥��x��"5!֩T#���+�2�Զ]���:�Ǽ6����o-��/鈼�b�{'T1�I��;r�4Ia�q)�;7�y�T3'��zԻ�k���>Y>ų��ٷ�$���}v�P��2}�x+mZ	a� �.9�Mgٷxg��	��*������͆�=p`'���a��+iiG<��2ho~Q86[�����|���YM0��:�a����?���+[S��U.����� 'pѝ�K�I4a����6�5v�yQx(��sd���C���I4�����
k Das^A!o1��������;6�N̢�]c*D�O��ރY�n�sM����8��/W[Dh�G���(	��C�4 x�z0�m���H@=�\�Ĥ0�.�{	r<ۊ�y.�yוJ��)W9E�^�8mIq5�M9�cw�|TxP����H!�9�N�u�Jϣ���Y�2T^8���m�D�Ur�u���9�����F'�1_� !+Ʃ=3���l[F�a���A�"�*t�\G՛�&�'��j&3��F�4<���.}�Qt�W���Z��42�f%a㔋w���+q�Ab�� Z�M��
��(W����Q���3�0��q2��P*�t�yb�Gn-h'�}�(�.< ��;anc&ǧ�B6[����6��?��C0^n(�T\�&S/K�[	p�w<����:�q��B�m�l{�ck=��"hғ*)V�G����|��-����dh6�3��X�P�KȒ�+J�eE����O-�i�@��/��y�z;` ���q �/`�Yd⩜sǼP�
.ڇ���̮A�oGWK�e�������3;0cI�N#��Ԇ8H۪�G/�v|g�S�#�Ehd���z���"�۩�W��ED�sp�H��܉��9���5��QT̓�rI�и*�?u���/F)K�s���܌�������|6=�� ='A����\3Ҽ8�?_v�����7 ٚ?��Q/�ct��8�"ZQ'#�(;�a���^�|�!Xc�<0�9��uЙҭ��u�zi2�V�y[5 z-��=�R�S�Ң�{��l.�i9��˜�>�	)
�$��y)����Y����x��G�i���h���UQԮ��������8���>vv�R8�i�K햯�5��x-�	|�YbB�˻5R�{���%��!	��C�ن����X랡1n3��&�i���@���C������܌YV��q��y��Eޥ������I�(���W	�R���b��m�]���1;}��������i��Y�r|p�k�Lou�H-I�[~��Z��B�d�͑n�-Z�i�l&h"��(�"_1���i��o|162�dεR(��O���Vm�`C�i"�5�*�8�:�e�i��^H��E�EA���q�Z!5_y� ��4J�Kn_����D>i҆���>�_�Z&;4��=����l�����=.Y�#zڒ�AE�d�5��2.*�)��+�MZ��A��	���
<��kTѥn@�e��V�L�7)P������L�.��&�Q<�v�Tגq�N�T8�JF����
)�;~�nR��S��,��*E�&��ԆZ�nM^��Fs������dMq6���}���"T�OB�����.��ZME��{*/�n)��`��f6RA�b�)TsN::��~�%4<�y��)�1��g�!����y}a׻��7��0tpZ�^�#pg<Y�|)(=���z�w|�L)U�k܈N�N������4����3�E̸���4y�.y�e&��8 , �|X����p�Eu��!s+;�bYI|�"`b�]^Tչ��\މd��#F8T���Ik-�8��V��)�p�x��j�M�3��i�] J�)���	L���Al]����k��Z3����e����$�ʹK������#��B,h��GM�5A�Ƨ�A"�?���oM�����z��@�Ț<�L'�Xq�yKω��]�Q����r3�D�Xm��9��4�t<P�������@]E}�[�]���;?H���.��,X�!�7u[��B`l�;μ8Uƣ%Le:�&e��N��ӫOB_o>xگ"��
����6�ܥ���MI��%���}��Mڎ�ƕ�����b}Vޔ���"�Ƴ>�D'm����E�D�Wq^�<<��������v?�5c+QL�2�Z���rޥz���~^�3�4�>s��"�����tW�X�Ӫ��h||���@��A�:�烣9?R�[��{U;� ���	'qQ�}H����>�,@�)��r$�� �a<��_&+��<������:�{1`��J�3�Mq+�v����Y�z�:Ƽt{t؍�'W^��\t��)X�#s�°b^|{��kM��$����,�Tx����+�nY���B�)���}"�|�����I�$y�<�`ڊ��7uH���+�w����6,�4٢��%B<�azf��CnI���8�´���F$$)�i�r�o�$��G�x֧��q	�$��H~��
I�\���ȻG���@�;;-eR��L^��ۤw�����1H�@�	�-\�I�����o���0��K�^�o�c\�%:�,�;"�iLX�Z�&xUt�e�@ys2Z,�Q�� ���x��ee���,09@���������yW�U(>�'_�A�)#��<Є[;��g�Y9<� ы�N�*�����R�AqS����~���S΋�Fq�l6��e�=��*� SLq!����Wc���j�2��|����&�8�H����-"��h�*����?��ǁk.f��aaZ��?e~��m ��Ҹ^��l�9`$���������;A�s�;"+ 4՞�(l��c��/���a�r(�/*o_�ZM�U���Y�.H1{�&Ǔv���ѵ�����3x��%��V6?ֶ/�)����kШIFKF���QI���lJ�����p!���ef�QjQ뿜�&��ێ	�A��`�~��`5���C�V8��t�p��E�!���f�j�
ȱz���6�K�n���O��A��3e�LH��+�$D(1�)pr0Q�>O�����Ι*��e�Xf�Q>��b�g�G��f˷3���.k�\�{���9�E���\�3A���:(��i-e��1i����<�t�p�ǖ��y�{�yrk9V����e����Ca8�K�|y�@'c��B��kKPp �{�@g+n�X�#9C3JS��b_dy�v���\�}�IV�.�ho$�q��-�)>�*��6A-[7y�Y�����rKP��_5.�9�o�ס���R�/X���O�RH���7kF����O�2�B�	O1��5��]	�������7b�M��r_?ڸW�t�+O]\��y!X�_>C�.�n:28mo:��ĥ��%���`�[&	4���
��f��єa
�N}�m���t��=MP$/u}��qa���U�|;�]e��s��#�4�����"���U\Ēv.I����K�V�9��_��SV����P6H��u_������?��r�Z�.6�jIͿ;����1�$ؘ.F�N��?-��V���Ên/��`��'�޳]��L��9�;vm����6Q��L�����M�vr��L��[�Zrǀ������Y8�4m甒?�|�p�������C�[��.���E�:�$1�F=t�1t�5cT��C.7���_���U���N>)�g�c���!����d#�HK���f�iԸ>y�/�J��F��_b��V�4��F�F�#}R�����ӵ���{��S��ݭ|�����9(J��^엾M�̹p[��0�rbfh��G
�e#�ƌ�J��YH��k+�Y' �U��(�=2��W����Fe�.����b$P��� �9C�<�]4r!ey��D�o���@n��FJ�W,�c�),�&��{�Ma9�N�6	�6��կ�6��߷�s'���,��_�����^/�[e2vaҗ!J:���hm�]��U��ˁ4��ĕ𽞵s�����)+܅tN�f���P<�V� H��Qy���s��B�W�zv�=����=H�{*�?n�u&��e�"�6�֬c�"A=�]Sdi7��J���sxQ���F�yI��� ��Rx�E%����D�B:@�aت�18$��0Jx�+"�Z�G�I��1�o���pT�Z����Y�����?^c�mH�?,�VM��ttdx����KH�o��B��J��A���c����&��F�y������W�u�&z��q}�����ݭ�v�
4�u��y����M��?��-�
��=�М̔��=��i�G�+��qA}��
-\�ɦ��R?�qJ�So�ܺ���2�rj ��z*-�}���w�lS<M�c�6d$��T�F�C����άG�$�s��,�������1|�d��b��*�"\�ə�6��<��8v\�����)/�W�)è]71�(��>j��"��1(D�F��w.ժ����D�U�@ik���"3̯�%S�� ﺇ\�|�+��vʛGD{5O6�'�jNP��?ʃ1�jO��:<o�U��1G瞰��'0����/#�I�����S�U�
��4�kX	��D��Hq���N&���*��f��41�tE^�0�������Ivƽ�U����2U�ا7��ʃ�k��?C�,6O�/9$��ŒL�8B;̭{�B|�7��?���e�0��b����ݐ���/L�OQq�����W`M���q�_ݲ���*������D�t��=y�?<����r��\�1��mgǒ.p�~�Xb4��Q=���l�1�
B.��P
�W	$+���lt�D����nV�r3������%�\�)���qpm�� $���g0a�S��R�m{��LWFmƾx�/�m��%��*?,�O!��#):cS�i�{�:�r�h�(��d[v�ֳ�y؄=[� U�n�0�b�͹��N+CP$ƒDh�#�M��@Tަ����vL_X<��H
p��D���p���
 ���;���zZ�K�5�1����k��D֖�.��7�*@Ǝ�yB|S��A`#	�3�1��&�0Ա$�aa�,.(���*��K�c��ź�HmzC�V��?F3+n@U��Ig�4{�]@EcF@�4faF0��GH�0�D�u]X�z��C[9���+m�Bsq����x��2��.<T:-�� �f����a)fR#p�F�SXj��ʱ�	e�g��<Q�~~��K�CV�j/HJ�c���ː3lۙ_zaE6r��di����p�8�b����왆BM��Rd8c�nFLԍ
O�;T`�+��3wҟ?��~Jږ�ƐO%��`&�@ɏ��LI��rF��z+j�ܜ��[�SA�֠�� _�D�j�k&��ǽ�}����tAm޽x����@�.����s��or+Ha�Xd����۰W��(�*�*�2 ��0Q��8l_�Z�E����������'4�}!',,���F���mu�Hq�W��ӷr�ϫ#����x@P]���]h�f�K��υ��̺t�"y?oY#���C�m���¶[�н��)�+�� V��e
��V̍�V\�.]��'��Qm��6ތ.�ޠ?�Z���w�U����f.��d���Nv�&���S�����4'b�w��}�%��da�TEG�aP���Ao{���Z��y$��Q�����yy>����z���8>t���$I\���7K�w"���}PyB�:���D���ʰ�)�W�x�p��q�ۻ�>�d��D�$��/!��:A�#(����v=��mj�?�t��
R�-��$��a�M�^��aF��-��Y%8z�I"3����рd2dkw0a���[/v#S��@��	����:С�L�aa��A�h��@ep{C3�̋HNڗ?�N)�w����)[��ᱮ�b��J��@���h�vr5��O�;d��тՕ|��t��sF��k�Iwf��B��"$����@!��C0Ԕ��+Ͻʧ;19�Gy�	�f� e���q?�|Uܺw� -#.��f�w�wb�����+�)E����:9T6'$	�)Bn����*Z���/ ��?�9��~�1S�!�l�����]ZZ��:j����P�Ecc-vɜ���5u�$.��"��'m�T��L�M��,�ф�?.�Př�
8*����^ޟ�-�h9��ļs�2��0b��1�I߲��P���s�hI����P��+�\AV�7��F���o�c�fh�U��kDM3(-����:��}M]Y�L�9�Vr-�Iw��!f��ɷ���y��4l�,E�J~U~�����r9n�%�I'��;]�Ė��Y)�-Q�N�4&��^{�����A�F��]ƾ�w�,��}���	{ڏ	��� u�Bڲ�d1�0�b}3^䢶>��*�Χ��<���I�S������b4/GVn��gB��	�,7�<�� �|�baTQ���l�&��Ǡ�KtS���
�C�%=�/3�T�z�.7t�sjMjK����W	Q�I����gm�c�s�� "��~�6A����B�"��s�?j�KS���?Цl���A߰�)l{��
�'�(��4zyv�X�:��{�����&���b.h������T�/�(t�
x�w�"���5�4Z�eg��ۥ���t�c��yv��3�8�ʴ���)Rb|D�jrv5��������aC����B�2��Έl�LA�(�<��i������ �"���{y(���� ��E%L��
	Y�\
�*h�{ų�������u�$zp-�P���y����Ȩ0 �y�swt0�����\��ecgerW5fs�!ǄRob�9�8x��;��?�mO�h���D8��	UhO�_�N<��	�S8�����3��Lm7�,?��-AnL�d��7!�V�b�������"��e
~
G��hJ�W0H+U�4�|�=m���{���Ϭz�2C��}�ߊ,|���[R�՞�q�����ny0�LcW�!3�4F'��4U��b��0��A��ޤ�˯��ޗ��ޤ,�D��~\���y��}+*È�|��7B<=ghx��s0���Y�����̠
L���{S�#�x���/��Ǽ���J|�����SL^m�kj@|�+���	���*8�u����(dfX���}���ث�`�!sߴ(�z`ٜz�W�C*ED�e�I�f�sJ�������γ:�؊1��d�k*&Lݽk�N4�ϛ�d��NrT%��/, q����{����@����R;6H��B�?�m���z���7�]��ޣ�v1q��ц�ֱdh�3X���J�ᘚꄡ �\��x�I��JLb����Fn�p���t�-�m�]�ט��(R�8�m�y&[��3�����+��²x�2M�;���6��f�� ���k/T�k7m5�Bt�yy�����������A�sO�����!�6���^�ӽ��?���#�
4go�C(]fя?�xW�Ǝ���6�Дi�\��x�����'U�{�0��&QwEj�FR��wU�����)�t��:�1�ȳ�7%3��5�h�����v���8��(N��ms?�Z����[uz��>��[�S��r#��G���c���8_ozG���Y$�\9\o*����=��T�=�f������UE��.r�vU[�c��t�VL�uZ����:?/���b��T��B�L[6Z��_�|�1����P
 �	���/���#���+�&Ǹ�A���]����J���$�����+~�K��<�!��t>���	1��Y��P?Ѩ�BB/	a�ʞl����+(�p�L�T ���LC���r��Sk3���&&v>R^����PH`Yf���z�oq^I�0��>1G�_��Q���҃\͑��[��|�T�!��7!Hn&��3���t`ѥO|�$uv��l{�q'�^�fn�$K��c��5����D�n~��yhYBR��<�9��¨�82��HD���I��q�+��m)�����\Yu#,��R9r'ٔ��z�Q�r���YY��ߊ	Ѿ�J�-0~�9
j������f�/���zG^�ƹ���B�E�j�~�"yW�i��(X+��1��]pl�ʺ��w�:P�g%�	mzKk�� �xY;
���#0�!a��3̆��M�@�h�k�S�}c�Z�N�;����`$4
gJ��&&���}����1;}*k}  d���g@�]�������c������t�b@c��R�K�<�����u�GA������m�*y�����0�����s�j"8�3���"h]QQ���Q����[���Y��l��D���i��4W���)��Ε�I,0B��F��\.�?#a�����Z��f��D"Yuu�C������w��U2�1O}d��+���b���1��|<��l�TH�=|s��F�_ilo��v�u�iH�R|�S�-�f���<$K�А���X���y�J�s��V�����}�ڨ��Qd�:j��b��<n�&q�W�'��SyҬ��Qbi��6��x+�),x��涞�"��
9G�C������E�D��[�\%�sңNYo��l�~�[\G뼈�8�*f�����Pr�P1&�6�ă@d�Q����m�׀<�AsȞ�>I*ڭ-�t��`Kr�z	���`�j���5~�׽'��L��f����;�d�*=t,	�G�#�J��/6I�m���a/�&�����X�����)��oW�3�ck�M��[�6w���ۄ~�:�j��� ���0z6�ww|��(�H�P7.6��~1�|ӓ��=��Wbo�t\w+D^�����䲺M$�]�[�\�\Od����q�Iϣ��+"f����{�׆�t��(�q�1������y��������0Ox#ɡ� i�>}Ԋl�Z��M���T�˨ws:��T�?����mR����9�M;@��7��+¤��ז{rh�E/�ַȆ�1~��]��U�Y�VB<�^���T Nj�В0�AXGn�,FV1
�v�{v� *=ȗ����})f�U
3ȕ/���i/Y�]��Ӣ�柤�\�[q8Ȟ�%�/$��a�EE�߃pHAR2�} sNq���Y�ߐ�Ʈ/�]n�hU���S{+�����c)�zCeί����oFZ����yQu��[�SB�A ��~볰��|A9�,���vZ��N�qߑ��Ⱥg��ǰ*-÷
e˭�7���ߒ69 (��f�`���d�"I��[�<�ӎ
��c��� n=�o:�kV�&~B���6iGa��[ 9�@9���q^�w��^�k�N6���Đ��������j���^v�ה�Ok���௱`=$ ��hÂ��ݛX�Kս�;����B!�Lc}O�ߟ�=�@���h�4� �gZ?#%f�T�:��f��	7�������T��G�CU��b|y��D�}DF��|�|����W����!Z���1x2��+��@A�(��_-H���%�=7�:yx�%��^3�w�b�t�3=���ӫ�,~Qh	�H2ik�ۂ���q�`��5�r�e�6�n�"�se�z�xG:O��� ��k{���#vK�2�,�%:���7>	�	6ܯL�jjleqBA�9f�ښF:|��|������G�В<ew�'��m��O��#->P3�ͤmt��ƫ����\�%�Vh���X'��̻#�M_;�	/}������R��B��%g��W[=do�Z���r�u���aPz��e�Ln���8���9+c�,5-Q�ML}�AKM����џ�bTR�&� �%Z%�5��4r!?�of�)�[Ӫ\�Ǧ)]r��x3,�1�! ���nz��U4��٤-9K�n�l"�� ��`f���M(�塵��1�ik�
I�K�1�;� �ҵ�������̶�W�b��'��ьN��׈��2C�<^�:�	�R��;Z���E��7���t�VC�nc
�I��TLN�K�ϧ~j{��������7"a���6�����DU�� }"�Ye��j�hER(dy0Z�� *��"+���s݋�˕��	E,A�S}Tg��H]�|�������׫�YCCp���Dq_�I����B�EN!��ߋ�V��4o���d�WY;A��JY��/Q8aDBw��`S]A��zt�D��ݫ��@C�+a�j���t�i�Pŉ?t>ĺ�, -�80~S^���,Ě{5~���Gѷ%�_^�I���<�|�Xw�v��O�*�����Rr��ZdDR��r�W�{�S��뛴�x}C�ς/��.yr�p(�݃��_���/c�YX��+����02h����xq�o�b)��2�����(��y�k@l������%%E�q�S�[ŷ���C�M��4�r�|V��i�L|�L	4������f�-7R���س;�k7�\������o�!��օ�B'��P=k`m]��]��d�RJ`i��0�~���rdPW�1*'>�bA�d�c�Ư�w@�$J��5%�`<x5��U$�$��*,�Z��oO�`B��6�|�Y ٦��Et�f�̲�߮��w"1P�a��)iF�U�B,�sN�;��V�ˍ٧;\���è���:G8��D��7>�F�ן�RL}�93�W�D����5X�ۼo^�Z��˼�v�_�殛h'ɞ�Mx����Q��:g�����;������ݞb$�� 󡡭8L�!�7���Ɖ)��į����6 M%x9|6b�hL�.�U|s�����9��І4�^�z�禝���R�j _��I[�@�J�_�PvuqȎ�<#��O���p�2�J��󯼗F��NX��D��>�;pX��(f���
)�J��q&\����2�P�@�6J�����p��S���$��<K:���&�to ��OL�3���ɘ�y(-�w
I�%vV���{��m4aK�<�Ɗ}H��wn�w�-��A��
m���XE7�*�[=?�h���i�I�o�N�@*���̃1:Oӏ8��+2���6K������5l�J X��
�TP2��K|�[n%�L�	�+��/5	��p��NF��q��3�%D�M��� �9KNT���<�6E�ؖ%��o���1d�{��H�G�w�=�+��T�������~S�C�!��]f��[��d1�I+��g�Ѣ��#ID7 �H<h �ʦY`Wwj�����T����sH�ð�8C4B���:�iydo$r�2�3k�)���������j���.{�)���\0��@��g��FMs
�9%��������r�4��<F��f��v��ʘr���1h,�	p4�%��v��Mr�\)��)�f���<����*2Tݯ)���0�i���W����M#D7̈����BV�*2[����/������K���a��E����Wb��I�%Rr�N�(��r\ �fa�W4����zKV�T��0�Ɓ��D�6/WQ�-�pJ���Z��'z;;#�s2!K(uݿ'��^@�\߈ �#����G�u�ה4�V��hy\^MV��⤙KT����i:�C����&F��=[���G�`C@��H�ל/[��\z��ղ��f��0���>n�}�������P(?����XU��c{�md5ߚ�P �Ư�պ�G[0~,ҩ�_��GXO��@i��m(��:H�:���t���FyMEE��%�P)�0S�U��e9�	���D���El,����-��8��
L������d��4��?VÈ.���#+��:��9�%�����_@�i���O{Q���d�y!�U�|�=g�L�e�`ɜ�����`h~sj�t����l=^�3���[G�M���>a���߳(w-��Y�����c�VUv�����:^��PZcN�e�^� F�	d�	���_���`�א��!dTd���ݢ��dC���R����ŋ6��kb&�n��p���yLgrO<_ֺ>̺q��vԑ�fj���E�6�E��_���$��hXܟ���-QV�J�����T|�a���[tww�'g�&3%g���DĢ��(�/!��d%s0i�0j�Ȥv3l>��>B�]���������Q�Y��>^�ݜ0ק�J��-e*M�8������o&�U��$������1�W����NՈ�"�ӑ��)������0��ɑ3��*%�Cz1�8�E*ぬ�(�&|пQ�!�N�A\�Oƺ7J���G��:�`$)��(�v��9?�@��<�@ ��RT�������v���r�t3l*�Mg���V����s�}�����Ȳ��?�Qt�Ӄ��3�y����?���%]�XI�>wEA&���-%�Ǻf�p9J(O�����{Xy���԰K~:���	�v��9)P��[R�A��@�=�� r	<���o)1�(�1�.�J���W+�y|%3(=B��Ğs�a���vF��\�T�X�`�}
�?�o��ez�vD)P]8��,xJ �X��P,T[�z>�tI\5f�E�۲0ZTI\�i�|�D�x�_<�������嬎��R5�
��*��ڈ2D��m���`��&#����m�E=q���(��\Ya��QG�% ��'H�ۆ���Dڂi�J��c�*�%�p���ү횉#��k�r�O.�A�;���1�:T`�
��8�v�}���ы$6�d�B�=��^2.��*�
2f�*ۈR�&Vϣ ��h��]2���F?�f��
��*9A����x���m6�\���GB�!�1�t�MK"���XRvS�t>G��#��\S��`	�� "�d��l���k}�9���o#�8����i���꼖bY�x�Ӝ]��C����㳛I����q�h���$���-��.�TDT�#���'�4	J.�xЏ���������� �S�����>��9�$��&����$R2�����:�8c��2ĊE���_ ���wL$Պ�}3�oŶv[ίB:N�Zi�Y&h���b*ћo�`�d5N��9O`�Zw�D>�d'���C|�e]c��e��m��"�8\<|Sq�oz�֦���lWj���������=6�XfB�����g����\H|J��h&Q_�����X�v���Հv>�q�!�dNPuq�J،#|��x"�h�Њ�N�KzO��X�A�ԁ���/�ۨ�XrbQD<�Ѽu��
�=5p�D�o�q�(�]��g�	��]��-�{0���%�PP�׍J��`�j)�V9�Oҡhe9����a^u���m۹`��V�#^�U��x>Z��aU��`�kRj9~I��r��D��ﱚi#�{Ԑjƅɐ�b[6���9@�F�w�ч�͚��^K����
m�֨�l�_s�L�-�~1��f����e~�O)�����%�=�<��*0Ub�����kt�<,%�з���\b_o o%��c葿�]���q�* n�9��ܱ�:��?q�[�_g��,n8^(z���e��ΌE/hk68B3.��N���[ˇ�qY���~����a�O�Jh��`�"�%��4�B&�W9�e�%�ĸLx��m�A�Ri�[.�[��R��˛�wY�հb
�g>`�rz��L�&������_��q�X�D10�il�"��OeSƳϮv�n+��R�A���//Q��[�3�
�c��h�D�(�G"�7_�I�dT{�@|(����x�׽I� ��^D�ucr%�ԇx�q�������hH�C��d�J٤w̽�Å����[q,L����J1������ee���a�z�%I`�%B��aN��p�~��ʲ0B��n�$�-�D����B�-;e��N�Q���v�V8�l�[D+��`Z��4Oe��m�u��mc���Ř�ʑ{�$�1�1�����H�#e �1��΂Um�����o��jϛ]�R69"��D�+���hU�)�v$M�ieB�W7L��'Z�S7A��y��0t ��*陀~ȵ�8�؋&(����t�@K*�vZ9�a<D���XDg՘ko��BD_���~k%���YK��Sa/Z��$�רZ��h�X�
t`���IB��P��$i�]�>6�Nf���nƣ��H1w`!A?���C�)�V%�q|���ܩq�=c㠱�J��S,_c�����[a<�{����Ν������x^C�V�huN�=�'?C,q�
䜝�J�Š|��,iY/]$�-l'�g�c�45����u�B
���1�4���e�_B�'�s��z죎����/����>ٵ�8�х�eI�L1���0�$T�n�J�LX�d�[���=���۟=�4�MO��L�dM|��nŶ� ��v�|��c��k"�[a�Ƴ5�z(���X��+�����d50�o	�X؏-�/b{	=p���V���Y��`<�nA,axא/�j�ڍ>��;�%R�eaN��K�ޅ;i��v���`Y�y~�Ud8�R�;��$[�xi��`�N��*�ާas>���nQSП��^!,P�C��y��<41A�p�0|�|�	D�?�[2��,C2�j����pBiI2��:,W����#_{�����aŹ^�L5�z�v�����/4�1��M��?Q4#��}��2ͮ*�v̏�QX%á���P���6�������C<��H]ĝ��"T� ���_��e���#�����ܒ��Ԟ��r�Ǣo�<v=��"��UI�U낭���hM�|I�/��oċz���t4Nl�8<;;~Ce���.���rz��T:��2���|�g�}�2<OMTWD��W��P���k�nPnپ��֬sz���@�xE�*BU�V�v����F*��M	r��;Hd�B��8����p���قC��pƍ7C�_����+,х����h���_��
;���Gzy�3������,`�(Q�54&Hg���H�G�-�� ��(5���ԍv�A�Ɏ��n�$XkGê;�F���v1˨�R#��Wc���}��F�cg%Ķ�3��
|�;" ���3Ȝ�u
jO޶��y��8��i�)�,�v��zb4�%���zF��E7����6���b<��O'�����Q{�i y�rX0XtG�ϊ�AހY0�H7nW��GP��b�s����1(`����i��K���=���M�1���fts#RW|_��L�nKF��-���h���B�|_q��7}�|�Du�1(Bq�=���Dy�E�E�[��bU�['�Ʈ/ެ�1�dQM�z�ڜ�$�r�90�~b��ˁ\ 䱞��	�$��y5�% ���C/�ڇ����!���4ë�+�"�.׈+[���]p�#K�[��g� �0�$�f!���M5z���}�ˎ=�CP�W��~�w��/�5�@(����t17h�.5��k�)��/��X2;��//��U�.����Es�o"K�@*P�'�/TQ��R���Y(/��z���
��웊eM�ɶ���@�H�!_ݝ������������˕SÄ7Gf6a=x��R��kN=l��q�=}P�3�~�bj���/$ɷ��F�H���uݳ�_F\i�V�O|� 6���3Q�@���¸$��R�F؟X��ʪv�դ�U�2�V�`���{گFM��)�zw#���p��ȅ��!ۭf�G�K��6�(���²v����O�o��V}��c^G�ۭ�@Xq����Q�u��.J�$��vs~�$�[?����,E���,!x��El����Bh�� G�{���K�
�b���uE$]���\�<_�47u�1�����P�6��]��[��Qm
tLj <C�Ӿ_N"�Zm�*Y+S�)�)q�v�뢿�Ye'p�'
��&Yi,�nQ��>���ᶉ>�F��0�.�eTT�	.��������ܒkW���	n:�4����ڭb@�k*�/:����gdHH_I3���Y�J�Z�3�,�;��겷�W�8� ���$���I�Dڮ�I��p}�<�7�l,�Wp`���b�Җ[�:J(Cˣ�r�ʸ<��T��ᩮ��a'��j��w������IP�'X��w����5P������9F¢l���E�	��c���&�˅�֤/\�70�n�J���~G5�d�T��]/�@�,�?�F���{?�]Rđ�Y�2��.�7��BɃH�Tl��Z�d� �w`��TV�/�L~炳'-`�Q̹&"�Ƶ �MG�7u�^X�Z֓�?|���EI���Ӫ���[�RE�D��	&�.P,%z|u�+Fmo�^%�D�D]���;nn����}g��mz��p����P��\_8��2dk� і����?���mv���G:h3	F*<X��ƁfLm�IU�B���Y9�'�>�w�#�|Ƈ��AO�ѾUgn����>aʣ�l��O�;�Vm�;�e�v���@NW�P)�sG�m��Yw���N<��B'L��W��+3Y����&S��G���s�������iCA+��b��>�1��r�&wK���3���"��W��a�Zy����z�>�2�)G��=[s7�Q�	-��W���}��/�`ͱl�R������]������#�ʯ4��h�4�0��H25��F8�]�#��Q�̭4�����B��*�#Ԓ��O.<\T���&�]��	��+�1���R��:�9ߤ���0I�y �?:/@��X"�r�e����T����B�;��.ơ�r�Z�^=T��z�~,�����q��|rf(b�\ ��� e�8�y�MZ�%��n7;Jp�?EX Qa&j�,N��2���5t<�e�vs�T��A��2d@�3(��5�9S�Dڨýx|H���9�R�L�19W����D+=����c��i�l�܍�Ҟ9G$�;�Jvg�_��F�[��B6�u(��|
'�9���
�ެJ="ύ5lrh�$�ֲ����,�t���dj�i憿x���K8e