-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zy6dUSEe93fgs7AnMyedgWM2dTA+kBgxtKwNxnUkJWIs3ycrJPztYIW2FHLFQaGVc6kRzZuByiOb
/X4dRVbExndYHF5GYFSlg4QGHPXuebgfT/cY6/ycGUYk58PwpbX07GtGgpiCt0CWDOHQZAzlTDkI
DMvf2tdpBXVK4+SUk+wqkRaS1TBZ43mwkophrcUNJAennjoqkCbduK/oE5hdzD3y+IVFOAXOA1cP
3rhTM4bg1HUuuD2tvfFF6dgXx6025MfIpCec4OZ1GcTqgCFLKHNouSNGlJx6efBzrDfmMUlVA1V0
qiFCO/sX8KHngTujGA8uTXaZOJv1/YpOPBVy4g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9744)
`protect data_block
o50nCPtAdBaQKBktT0xfrW+xV2tIFdKVuLUmenmojvRtGJqa29TMEJ+1+8deulAnG434KpQrm7Dl
hHIutS4P6UwBHP8SbCDsnuQTbtmivQiYISuaX4+a0sf6QGBuYDfFOSSIDi7NvKQcm7FEHZj9rHB2
vRU1DL11XADA9Nk7TDF5tVrM6cDbqcuG2TEm4mhi/l5jZ3Dr+yAnk6X4Vmt4U6eAP7ZU6COZavJ6
SGExolbSNVk4vvx1SrtHNZpqNN4dlRy9YpjwJObBsHifdNrqV3uXmHJQOuprRTwP/oj8BGujnZJw
orn4K2cP2FPvm+22ekoEQ4VLbLyMcTXiM1LFFSdjsbRL6vnAV4Cw+WObT6nSSPY14cQo2pfU5ULk
i/mf5T5jN9neB6b/5bwpMkGbYidUEs8RRIGmIm4UblSj5867fTk7IxzhheynvQ6TJf+AmliBzVjU
fapSLiNBCDRPF/biYtrIJTIgvDrwSTe96gENdmAYV2sdF38PczLkKBNcfhKBfrccsvRnOrGXK3F9
dKAsQGxmN2vaq8Lkpi4QV7USRXX58PDZuc0oa66PRbLVRmdH6bbl85tCd64WO98Fzd65OgXIHPVf
thpn97Vjaa5nEXIws/lmsIxci0FX1T4RRm1MDiaka0g3IRiDrmK8J5hbYSALleewBG7eYE+rWfwT
sYUzZmnJT0Ww+K2e1nOlf34agZnGaRJKT49wKbInV7oMClCe7CEiPkCXU3liz0NBLRVtxugpM/q4
udS4fpQssNGxk+bTHT7wKEORolbY2hd+KxBNK1TSADMGOMfWXMTCIA+dsLXF7/NFL/dyzL24AAu6
WjjkxuXrIIb3KI8bSvjlltsGuNlwcTe7N02bFTsLa+MJQwGFFg1vLgFGGudBl9CYsJ4hGUTPLwOi
2q/Wtb7HvvBqeKC+6BVv+8Nzl3w1L/jJESXuf8+cB6scN12n5uvYZgMxMlu81lFHNhiiBgkGJC1Q
l+/+T6NL9sEOBcjp4Yr2Q+3nWgxKbhrYJ6TMXuD6/oOYJIX99vkomdSQh5cTnHpinaEsJy1t28ji
whYBFhb9BKoKucO5GuBdDIAz9SJXjF4i0RT2poPOj7MyjcPW9i+P8LC57D8swjRp01NGLsO0mgFS
nKnD1KXgL2o/KVg9CaH2FbPvNXNPct/3L5YHO7XW07v03qXqQORROqnZ3NFuV/M7o5x5wGyUYoA8
43KD+8KeCePyHorLOdgkqLqjzcmeVwJInoG4MeUeVJphiyJslwNZDm05gzqWcRBjTYbNWu73B2yA
tHW1+KwamuZCAZGZK+o+DrJt+BVDStiadyUkdY+7KLV3ZY/Dk6pXki1cxH4QF+/sTQimxNv7ayly
36voU9AcGdoZtp1x0APHAbrClQVpef7b0itu8ebJEpmIO03CWftXi3yaDKXZVpvgNHz8d787q5ah
ZDXUQ0LfHWIJKeCcZtFAtQ1eW+5s7v/Zx6YYwNqqrkWFBJ4qgMpJrwI5/k/yf5VA2WLrRzhNyPhF
v0LbkMEVR+AREcOQOMXnEfccj3DQM/MF2V6kZERFSD5Y3iRmgxBwX6LttYuAWoa4BPAl6/lgXtrK
CaNvZkyGLsi1Lp5eBo3DFCxR0a05Bbz/jnX/LLU2d0Bfon523FmXZYjAFJOZ93VaoSWyonKY2SpV
LuGVJnYGexnTNbLZChG3GBnXgq6K6yTzyd11Iwj4UGcSuFJoj5gXa7MSGmnkv5YLjEKvP12+Ar6h
2ZwcI8hQVhTGDMOfQ4WC1cEnRJSahMjILD9j7eL1zPvPbW8EBTioOO+ie9F20XKAVuP0cxD43W3F
ralprXkkNYeYNy1amEm/c3+cFiwv0gOVa6N8J+fsEsHmRNdf+I4HMT9VIxx3Q2hbamu2s6E2XRwB
XzwXFdgLDStfOTrkBpax/Mbw0qb7Wl4fWgbz65J2kuocOEFkxpGG26VFEC7PutZ7Fzjj4eS2Bx56
vyXzUDSeWoDrIUW3TlbFDUBNrBFlQULKLBcRgNYRY7h839x9rsHSpM2VGbZvU9X3yB8fGL7YZJ0e
Oq1xXXhpHKsqThghMcxlgGzLrYKW9TZp+MR0cRTMX7H9G15mpjEx4NJCUyRFIys8hYrWdQyEJEty
Ja38Y0XcE9N/6slMiH5dn1f8UB+1vXKPSRHO9VKtBEmoMcK1/TYP3xfORmTlQlGvDGQofSC8tZaJ
9pKQiqyT6yFPzDnzY9Zeq9UXXzPhEU/j6nYhRy5FH/EK7Wjp5tkhJObx4k9+UwkZNA04uar3igM6
vOZf1tWTqf/HOYCUy4IIdxaDeKCdCEMhaAZHUx7VUAQsZ0Zs/JwXx7ZDKV1vDYkCozeUdZvf1L9V
+5jzVHdklCu4SirtaASQIOY8wxl5TBoyjMyN+GjxuRiaLpXpqGJYBy2YMVbS0Jm7TNnUliJRmMnt
lX1GFY921ADsjGVPM2HD6bbQDTrrf5iQioHuo+IbABj3Y1HvXTgR0cTGLsNxfarSdhj/SN26yagj
M7n7B1ruYW1oV1xYsgTDBBon6IgQ+/4myYS/bGvUfivcwJDnyTdbyJ9Dg9yZp7HE+c6H8871EkEf
Kgrh+O6kHpE2JiGEM0Bzw2iswrxfDPASSVhEVAvjIZzzwWplaLIjWRnNyyj0dOdHENusJ5nQf/6K
Wu9yj324fbh8qehMFHTY+6CN4uLLwOfQ1AoVPRH7artWaoRrNd6VS1tlGzzF5OLBxeZ+6JY2Lo5m
nHpwl3aExM1PbW/DsHIWT8OfzuRNdZszP1XF+k7wb4vZLen7OVQg54U4eBHcCpqyrsRADYQUVm4f
hI3CE1Q356mWX4HCod0yYW6EeNzk9fpqP8mP6eutl/i701BQI4ARl039Nkc+anz+Kfda1iPLzYLJ
CJT3CSZ/TYyX4c0Ayx/LHHtgOYJWcLbvP8pnKXnhIlRqTi+94z6w6OKI4QIq3L0WG8Tf29gzN/2y
tfUDRR7Gzks3DYBHFJn2XGeHSUrK1FMplXcpVW+/9otUXoVjEFMr/5pUqOgvfUxFFaso4hZ5IKI8
XYxf6FAAFTPaYjb7vSXJSIa+S/11suEt3VnHE8/TaGoQxBKrl3N8IUIrvWSNvC9SJNX4pwG7CYh7
ILoT5RftnxVHI8nJOtB/IOfbX2DqWCZu+xjD9w6QwR1oijea4UjUJFn4TxjPXn1Ca7BIcQ6kpxkk
V3pJkWdkK2AqBpyySmHlYKgrxAG81kOjYEJnmH1WYGCVCaQQ3ezbhu++aCeYDmlhAzx2jlWc2KqS
Mz40WKc+HyJHVaYoRJn6py0cpX6ilLyVHIA0l2ckGKG3qhCL4rmyRjsmCiuO/v0C+x8+Bq3BqiQ2
NF9Yi3iHhtPioxf+drRutLCmwtAFPFPMm8o3kFK4NHeowPNxOKmyLL/9u8LbIriy/+8V8GkqOkTx
WRiHJ7IqQwNE3igQqYztmS67NuI37iLfTQPbc+J9BWJBlKzdEWDG5G8pojofE4h+8Cz3dgePA1Oe
L5rN44mSM2yWEF65WJjp8O8OJSlCXVqovpAWXTxQkFKzj9SrV3wtCl6AS2RMiZ1q/W+gYjOUFLJW
FsquKx7OB/OOLWDxAuon4P4Ksjowpd1fzJq4O3kvN/BSZSwNLsfo3YP2f5nXV2c+rgi69tKTVvIY
VlsGSRZYVc1G3EMoDdJ4qpg6i8Zijf2u0eYfW7pZKVQcK4fpp8jnR47MpH1PVxs1pWuapEC492gq
JRzMHei8EWTGS/x+G/wUnMa4K4eGwt+XSU3Q0twSZPY/+kwV1Yshuz/x12GjDgoHCn7bu4pwp8n/
YYTsRrKwvwR6HHqB7qefo7IQlK1UwDmd+n/vHlC/jZPL/Vs3kh6f4pBBCDETjnnqazYfppWDIikz
SoArYxpwRGLGuMBgkvArDii9JxRQQfBwOkVGA8jHvQobnuOniJnbZ2EqJpZEKd+3oUlePGk3ilYO
jtYb2G2tahTYCAov3oWiDb+/ovOK5EvEEpdBQIUN0a6hT6RtVODCfFOIoy084zvb1ImryFV6juA2
di+tuCEq2/ZTapcNdABQsa1thLFc5/hvi/K9XHzRC87wjs8dEwyHhK1anp3G9u9TWjVlvxoCRW2i
yCIophv6FlzQnYnR+Oq73BmKj0NlbCvsu9rQL9Y6gNnbrXQIzbiReOI/O+c/vJWjxSMsdjwa4YLR
oxjPIM0OwTwL2QfIsLJvv0LFhUE/qUiR3eLQjQQZXXEVhG9YQJrG4GKQp2nSpMIow4Zknyvvivqe
vU97GcvhG6WgBPt0ZTKDmdbIuh7LR7utGYEsVDOOcHchWuT6iG8VzZRzYALZd0uXAGha0FS3YLSh
spaXhL1k19lca3kxO13CnjculFrT13ziphTpJgwopHzkup54NXrhoRvIm7jvX8hfTgDhvyqHaHJP
XYtHe4UY5s1BXZCOXXE9LnVZ9ABmfXuN0qyVjhatT7awElqYTKEvrTYHiccK+3B35D5uP4eabhql
iGEYmxXWGCs4UevhtWgOzGvPJ0QTAU8Qpm6kNQ13qFiFibo59g9DDOb9M7Y29YcRl02oFmb5b8xZ
rUcKSU33VUHZzRwKcUHcQq/89DDJfgAWlYlay+Go44+BtQwgjnajIPLD36uC/tG+/TWYxmugoEB3
jiXGmWKTl2sGfIf6YqI/QyR5BeRKndlx+D6Nxgew1sWG//TFJdd53y3QVuUF91oZldexexIVyfxZ
G7/TyRRE80e7giiKhq22TnHyVd4d10r180nDQWnOE10fu9JB15E6CP8YrkIi4GfGS3IhdPk+VWJ/
B/E5QLhmOfq6Ioeqv6KEWFr019jqpnMv/aLIwpTlLs5SLbfPkW3qrW6LCykjnfCimWKW45V7uCaP
XRLQqjngUEcofLVKvt9dEJZsb4PWJ2eXjWNP2N3DPCp6BhZEqsaeh1ll97pnDt/N9Fv/zaM21LUd
OgoielI0HiF5732ad1QMM65pRrLf79jJADaW5D952vVm08nlm+G/eC8+Nq1bTpB1abpCICTHItj/
1E7BznwTXOz/NgbjlaL7oO9mpDLtR5VuCQY0PnL3oDxGiRUgtm5Uf5Ab3ZegYgHVp1jRFzLwBQe4
NNqgibxO+ahvBPu0G2TctXgD2oeMnFoHVackcJiWTnj3/ryNPfzva1+f8WL7w2DzSbeUDMJmZTqr
7OTs0JG848KgchCeo4Eu9DJ7En1V03QzkXOJZim64JT2DMCto8/ce04W2OpS82Z0+SiMZP8tYxC5
/EXXVSE6sYXfKzTTIBw+2TLLJx2clTQFA2KnixXq2XyaUEo4nMB2B1EuYSpfspqKubExkFi43NED
WzeWroeDvxXsehEAqgl4I4W399dnedOQ6UbJAz2tNCrxhIbt6WiY8Mj1feIZ3TJApjU+SYfOieww
5zG952ldEPMXv1LlST4DWTACyj0N6AIUF8OFtpWu0PIjlVr6cGBoyZ6APxv+GmFm550Oi2U650DR
OVAxNYNJZnSrnQzCxOSvLVDUwA0RnFGIYtdmyMqDRCPwcyZ3x/fLKWwB63a2NSRqsRygnNTU3QGg
+kz0Te1j7QOOXFoXmBXQ+wKytKa4GXZ9Nsv+mCMV4uDklr5xzhdJxZ1lEZbm2NXTJkUcel1J6Os2
cX5tQVZAO39mKb9DMvX6Sh8EWniABZwA+QwFGwnhBOj+kR8gjVZWxJoafUs6CKOHXYfvV1N/cBtv
RL2PRQKEJApvI1GsrpUBqMBd7QOubYr/PicQMQbgtrifI/lMvkXtpxUD2PQ/O++Lp8XQRaeMrzPV
JgEo2IrVzBtKBrRWriiomXN2HCFZMoYm3NZNxwanB6xFVUAoObBPNNrSN5TQl8VNKVpI146okN7W
VAzqQCtzUyUgZZ4VuZEQu4SGxoO/zQzOOYAr7kSbghXFhlbcWCHHy4ly4MuyvOBk8hD6KUNk9qMI
i6VlnK4ouAPIW2pPRZxPRPTAbUheoCcn9JR7q9a/40iZCxl3qYrI9Sh/+46g6sWjXhbj2A7+XhfY
/qUd8H7DwUmvOqkuYG4Y45Rfi1+5XDVGwYshBEJSt4y2D2FbGnBPvL9i8GLL+ZfrogZ9fiZIPNKt
uSBFF0CBP1uN/dM7twRrYbz1WjaiCL9lMeURRPjCOlv2YAfGf+EXkukR52qDr9TAa1FhspE/KmJd
yXsrrO2C61ukPWRL40uD6v9rMxHmtb7P8Ao9oLzFCknw++8nYOVPvR3pmRzurptuulopsS2D8tdy
1olWfamzKlZ2yss9yomckAwNVD8GZfNs2Bk4k/v8GSmh9SjGhIB/aT72cIX/N/brNHVwfJcKn2Q4
6CdRxujYBlxTgCap72LEdfY5Z97ypXrBxylC4SG3NsDWZZ9BK2unEsys0HhGaBJdeSX9JrIqKhT2
WdfLaLo1f2sMoUV3tn43toCsFM4xGZeLDVxhlcRTdHod0r5/nD/c85bGeGGpiBb9OHz+MjR/vHWa
MxpS7LATozDFn3UF+NbW2U+jBBskYCvSwzwwBAsBtPyHROoV/QyGMFTahA1zvxNWNG57YndpCWDh
16RcxIxcvLsLiXCoZmAPCraEWTh96FgKH3oMtJaJmyEoh4vGI4oqpSXpoWxGEL+J5mMMvmxnwej2
yPTdEWs4XRvrOHidjCbiBNYOg6jBvxILFRm0mYCHBGc4A64I09BBWc6iPcfxhEpEdjeEUH3lxQ0D
ZXjTiwEahUP70Gc9zzFneA6asRvMMTmi+D0oVj3TgNx6txS2quUn26XITVo3y10jNsOimrYexsj1
R/u4mE9ik0xeir1AX19c1GJgOkqTMXoYsgNDQGRtcG/OvjaVGETjApPnaa2fYyEl6PoKyCw/V1Ra
mQ3nm6Zq4fXAgExEmpkbteKcbXdb7PnUlbPCazsw4pg2eW5pOZaUqMwJ3C+qHKMSMLRZx7C/FuVq
wuJwEi3GrlWKM96dC4A+OAe7kOEha6uGLk3eXwZmvQj7UsxKPvWM/VhKxYQ1qOpJ0JWPTDyZ2nNL
yBTEOUZvy81HyJIOYw74mh5J6VDhONauqyM0AEbgLEeNBhwPraiLv2DJZfjHWXzDRmSfm7KoiWn2
QRCPL/lVru0iOBkZPE+HQn+Pw+BsUp1rzds9fyAf81bbOG1Pe5F1+F36lg7qsg4CVI67JlRjP0vS
Nh2d+xUJkhq4Z5P+sE5Um3txEN4QiDXDNYj6bpOnlPhRhXvKSFXc7HRUxL4HDpPsS4ooVvaVkRWO
QzEDPjuzqhHSW+W6i3feNz2IVQo24z1cT4O/yKRx94JVVM5orM9xhtA4QF1Rkz+viG/Hf1/9lZWv
ruHJ4oZE31Egj6YsPMZNjeZocD+UI97eA1oj/NCKv0nJkPbcHk1v6Tf55LqMBsc8F1/FE8NoHGp8
mV6kP2Ol8rZVST5Cd7CdaGtM+6Y0LxepUlH9l+MwvJQUQa64mqxN09Q7LRsJ1gOF+xQIpxHiq7wx
P5kj2jqKOzjmeouAwigv3o59YO1j5fawo++kmQF4of6z8iFOWCF+C/8nq0hde5781wp0Fb51ijoA
YQoulEdpsvEC1XonB4QvfSkOCqIn7uNFs9mwX/7Rgc82TSgK3GR0r7AabSprSdDGJumCNUOydUPR
Q7HZCk6UfI5FVDri/86LUJxQnBZzQYTGxGfhP6fKXFYVtJGwQ3673eXCmRmyDPUdvvgXH/AX3K6C
dl/psrlnGwVAAOR9vwMSHadynkz2jaEh26+n2ebTq5hKDUfplm1aUAAiP1sELVJtwdKrs+9/9n9b
5h1naqsbFoHxwSqYcniPqh/DYTLrSSsAbm+aoqAt0sjt24VWNV/bcksjL70Wi6mqg9ZFKNd0D5I5
fVX+OakI/ZOJb60nyR653TO01CAzW5jjf9C/RIBUUgo1iPT+DD+LT3eseMeUlPNdlftVfBA1OJfM
U4lHaJm7ui3y/o855n6lLeurj+NpqsINDAnpSpaPWR/0/LMNoxbSUjHLkKQpKnqhyhKzOH9YrdX5
aNveea10o5m5YKJDopU2lp+KzScbYegi35yflM1//CEFf7b7DSXAfr/XHO18aLhNCaR/we4NxapO
WfB8Wbet27SYzUawPj2RofaE9pq991ibPMNBqsu3EFn8p63J6BwMRiRbmm8BDoLkgyrpg6ew+Ta4
Uds1h6erYbyYuwIckhWsUUb1M544iLSE2u/mZtbxQQjdqiKxh2nyU8Exb5EYFu88i2JS53ACPU6X
D3nzzxAqqvApBAtSgIgLIpQEKGD/5NiQKVDJuNK8wkfrZFGxAa/bxwWc90HSPiP+dSzeNR2LGyaw
LYNDS2G2Afg7QUmD5qyHKAg6iBXUZkzC5+ITY1+mPXcKjl/TLz/6UjGGSf008KiW0/tDJ1Xjt+6/
25vqMlfpoPRHM0Qy7cxoa5E0ErPGoRE48NEIZo6ZaD5fvyUlcFfEG+E2MqieWRBAAoiV0qKgJD6w
+e0R7pZw7r3bn30cRmlBjw+Z+QVYUJ4gbYT5k1RcagFiSFMG3Re6+Nqq36K29iuVKP5IgiQA/0l0
oHr8wV18LvT04EOHtNU4cQEoLgKobHh9BqQbk7caLWZn16lyF/GWXWNkqVyGe96UJzWkiZvtird9
1fsULouaFsPyrQWg6dT8AFNSzUb2/1q7gXk6U7YMvuXYKlnX4sf9Uy0qOgt9TSqXlFKaFDohF5pu
KGTc2ayBLxb11VqZlFpWOkv51hzXaCklAn1ppAbyV1+IXssXHjM0IyfkMX0fZhO0JOnTQdIRqbzC
/e7jiy3ei97Swbo/Jgp5hwHaTSwxJQQsYICdQ6Vd9dEIwB2ZC7W0t2KqBAB3uAzuhxpEjVPHz2dP
NBlgQ5R9HgdebBZg5idXo3/ONHYEA43uX2aFn91+PQyqOASQFe2yggksKMq+2nVi/XGzan8nTqEA
S1UXj5hKANpfYfkTmXKfvRstoqdpiEpH86d7GClO7rH31j4thit4f5iMUiikxKytttVkpE5mURmx
ZxpH7Y4wfteAy9Ib1ldzm/Yeg5YIH1G2wb0UZcodw3Bg88RuagTC391XvvA78ZgmDYa5gsWcBm/B
vMS7wOMJnOIPaz2XiN3Dyu+gU3gl4P4fnxZJVLMKj2tmMC0V75rbnWOAALVwBxSH9oIcnQ0TojdJ
FW9E5xD7ZxhwHIzjWq8U7zjfz8uh+rbTFDMnOwce2Z1oOGBtfUL7c7WXDfMRV5mgZaRUWPhAGp2H
omTRVkg1WTwTJ9dyTu1MVvWgW/rjzS42rBJ9An2OxuzjylGoOaX1pfLpP0SipNtPPRahfkdFqDYI
NGShaysxmUR06GfZgVLZac7D4PwX0yzhQ3lks+WhVVf8SU1kC2QJ6fYfCIUt8YV4qE/V8IL8iJrI
Rtr3MOOVRC5iljAnpjnBNSLPpBdA5bLh4JI+hHlgNtO9z+zlJy8+ODRUzaZg2ppS5/3CTXd4kIu6
3VzipoDW2Seadda12KV5NfsveaKCWofD16tsicFbej8vS5uwp+N0qdEOp7X2ZrXSTckLRL287TqB
drCNoXzqLRp/HcwUckecCEX+LJega1HiVD56qq387sHGG8nNpI8rxDR3a3Q5eGtIKysiEpiCnbWy
iHj+h/JteFAzYM8uX6/jLNjwWynXUWd1kABOGjRDM/m1QvWxZ0PEcOkDNDW8SvoaD6IaIoJeBOSs
8WSLogJSiN4IwW+7L766+ZBgteikp8Up1RBD7Z3wbyzyXBk0YCAE7+T6ZjiWanegg+ABWOsrvhK1
IEpPsQgL0jW5OarYMbglAAxXJffWB/jDeZpWSe0yUNgLYCRloFzIymAUb0eSxbESWd43j14/RehZ
GEgYA71eXXspLSvJq2EL7pT1JoTy5cLCG0iumLrcVsSdCKENtphVfLqpJCO1Nw/hvo3puscUXVnz
qJ2CjgOA2axU5yKO6IH5SCM+U78Oa7PPzRxo6+MTGFFRk/d1kXxlGsULhXRlobYuOJg16cBun5f9
91P0qhylQpokWHM7k09tJIL2SfvJ/olg1eD/KH2zgOL91a/1EhJQuijsKXEWydMDoWsiDTnre8Qq
J6vTPtMFWP0DUQ5HhG8V7tXWUVb6JPqj4C5GWNY8bXbHoCOm9fjoZl7eGyxRQ27mQF7KBXsCSn//
TXzE7MU0tkMSYI4dfKxzJq8W1+132V8xBLhhl76/t2Pakxu/h2ffAbBlC5Ilx43x6sZP7108EIZo
ae1G2gswYND8sfCJCRhJiJp7ahJoRYVleJFIRsix93dfjYBHpSBA0tTj1SeAmYEnP2q41vM2pCuv
e0rHHSVKwtSUFMSWx5lM6GjinSbfWCRr57ilSeD0hY9wFJ/VtxykX84QWwP9XIWhLVgf9htzw1jl
Kn42MwUqA23l2GfZWsJJT1UmOWG7zSXbCi+tSYNHcqktZrgdJXk5hF+Ac8LKq5q5fTNpGa15Ry9R
oUwFpZ3IBHj/Ua+UwjOKmZ7YoY3L4k3+pKWwOJ41CWnPHaEGpVXxHhJMR/QGZIbDghPNnkd3Lvx+
WHxFYohI8eY05gNcCFmhaLZT3opDAs1adYVLJ5zFDxpDSxhTX87umZaK9Mc36OI0PmcSBrvvI+K+
wRsCr7AoEulk0hXIeqo9HOSK7q8IHs8HHnG5VWITR2TnV3Uj6wB9AFzmVISWNL0rfyPzJAXsKmGU
StAMw/Q3Nq2l59HJX5yFEksAyfpkHzIoyTuxnjwGTaR90Qc19JSUnRmKLwBjrHK7TcB/lKC6wtgn
MVcw5rh9Ocr8g41vO3xMxHF2yJiCXGO7gMcXLLitea9mdhkTS6j2XR0aEZM75WSfdieReBb088d4
y/O23N3q9zXKvylAJV10MPad+djX6qVAwXifJrDn6VbdkspqWW3oGqNSvYfgNs7s5EojMfIb3nfP
i0Q4BQJP2gXTiEMxzyp1NHQ1DntYPQUQsT/tnhlYktQOHfI0VJfVbiVKIXqfcGufokfR2BJzrkk9
b2esT3T6mmd0YqihcufzyUpiq8aX1oiOSjcuQOWDSfVXjagEylUYdZXc5isuridg/MX85fUPRDnI
HnldUn2chaN/RKAVDX59qRaKpxkbZtg2wZ9zhYwe6xGGCJ1pa4oLxjMHogB1QzTwA5XTmb9qKCun
MSXLyvuXydLYWFh7BpmYWUk+eQFzRNFkjvrRcFHdcBGntVArfN7q/HpyJcfIq3U7/pprcB95W3TT
Svnk0qOnOblNqp98IZ+ngKnUJ9F3Qc/i6cx5/ae5Dk1LGuWE06u42XdCDowYGW0lp68KnEsV6xXo
ynF0ZkadWszScb5IAbbaEGIHq/sgHM1/naHOlHBIgAvmYQUrgbAT1/ztApogsZTAZxa16WsqROs4
bGg7wTWYumbvI/LLn5lnWYqJAv7BONeDlzM91nR0DiWF494SqYL5I81FrQs7NWWgUL/bv60BVoOf
j7DPL/jGt9J2ynX7qLdHliQtRNtd6jTdzDxThZvDHOddHjvrqE/8aSV8re1o+6YmDjm4ulPavb/u
MavoxGLW7tcDZsfrdvB8dnIG1ZvDo0nBE8sif30LRmX4H2/V7CM6z5xuN7K+lNSRb9cNdxdoLNWF
ffm4kjAzJCWC3QDVLd8tfO8syFq8yT17Zp/MdKWxBoLJruwcLDorx5o27pVhQ7xTbUTGICtbQOov
Tb+GvpvmNpP2tWsS3Gf0rzMFJdY8DNLGCntFLFU6IQayv1hTxrxfVeb06RDbtzFO9MkdLuQTLQxe
dK+GI6HIIQ7QegM1kXofd487jUHQ5q1yfeXRArkWzopmTQ9aUybAFF3P8IKEk0gr4tCQEppm5xc4
sPmiUeFfetuvrCwvPMwFVITrgxMlafvZWFPrggnKVUtO48T/n+tg4K7Q71Wm+lgJEIeDfrufHsG3
3tcpc6IOowjtMSG9f+YeA+Z5JB+WBU0SMQw3udToFRl354CDNpm76pbgnWywRSIQCaco6ZI4ncGl
+vhgQq2il2XNJSApZ6AVQDqJjpGfy8M4ktqDfYJDtEsfOfLIu/lAyQaIe6WEgitsgh2/SYZKkbHB
+eNUKv4VV5llsXjiugTmSjBWXPG2GmvczyJDCC0OKqlfkxe+PzJCXDKbXdiY+ZCzWeL29lnhq/hr
UKvhsVFl9hWTs/wBPzjkvNFQZKDz9CjxVt60/YDGbf+LLcAh6dmLHHlLNT1HGJJHeYk91riKSngt
J0fxhF1kmupAm/V7NEUlguXe4li6oUGPfcpVS8hCxOCP5MQW+C+b+smcvXAKEv7qQpK/ahjnYLGp
9okW0XrT3VntBerXqsZNXfoITXCEFyAo45tkkDTxLGQfPbn+OLN41JP2Ij/QDVUnEHllKq/5Pgd9
I5YuquC7InmPww/YDVEyd8ItcrV7gHODj0vZfXHu2fIWech3ZRH5n8A2U7Bo0+VjUNnT4IY1FSpu
gp4fbcjktK/FpUzTyNBK7QA2LUPEZbAPuX9JIdYYskRv1YK44iIt3S1h8nJmCUKuYBECESh5iOSu
oxAQcv1qACn069eGf5tajDc7R6x9M6OsK7hXeidt4bRUld+pAIXivgoINKx+b9vpATHC4O6HDDfX
lMsHHjrWrFH11OxEghXqEdIaWhkSTcx8q7u/Q/NCOiac7rQISaA3Gejt/FGvi2CLdTuyyZIjpOHH
tCtZ72pI0ObeCqRaS9bU1YOCvUY3Q1oyUO9+EtT2Rez08jj7wAfhGZVpSCLj7VwbaoaOSXWuoU6/
4I1UfbM8nbnGMdpcbT3+jxh3LPkROA+V5i2APIyuRcvsIRs50mq4pztJmShtNsPwcc3BZbXfJfCf
icx/4BAUZVqqCTy2olcPmVZ9gd6i4SjxihutjQz0PjWM9PEXFljoV2j+Si1KUTd1k2OJScRlN8bp
B1s3tQCNX8/WE3o7gX8WLxFdE/46ELVZJm/HXXiiAI9YaOn9gGMOumcyA198CWeOwaiRU9gEkZIm
dvM+Z/AddfI9kawqOcFyRGTCT+sbhsFkDC0Bi05L/53BdYt3BkQkO3ZriQzX5ew9mINN1FCJ
`protect end_protected
