-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
V8w/OMmvpWJAlceoG9K0wDjwq2VffMlHMK74rW/afBDyG1ml+hwLgufs4HiUl/pq1R/ju+ukOfk5
9hSDKFmdmyrggQGw39v6QHMd33+UAUSuKyvcLxwyLnLwPkIW+2j6SYRMLA1CeQKJevpUaciEXt7g
/yqcykGySVYrNG6S2aBqNnPiuZF8uundZlLyJ9vk0AOYlZZLZEivUjBs1HHPeBmEWcOMpGmbH0iz
mZ2BF9JycPTpy79hON+JZBfL4I9qmCGY3wtLUwuZhcKiBVtM8/x9QS/Q9m5oj2zmJba57VL/jFRt
rCuAR8dlc8ObiN/DDMttOFyOpKu8fyBY07acHQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
W0CDa8eDWWCiCn+pGr1i+0CC8TeSbfvb8TckVLFz6JA7Xqt8DTH+oC5chSvvrUY1Bb+f0ghGsctu
DWX1fXWQf/dtuOtJJP6z22KpKc9Fdhnqf80IPdRwgxxD6ws2kxE3mOtThX4zRFbg7B/Jom2nIxTq
0Ciit0DNlFlle1YidM+b0wMpK2i/ZEpk3CaZHA+0kkaxUqmRLu3V3afP/rZECLOFstGrUJjW0Ozi
ZGFPH/84EsLllrGLFG99rxHYwd+1wbFFDNn1nF65zjgjO5SUNJiE3S8MBa8uC5tyBHryRrI7UxUz
uBur844DsyKReUL4XDURwTKU8cV7OdfsRyT/G+uJ2kRFDmX3h0pDRDroI3uUApvWBCsVKigCbg8Y
UObR7c+NPEuyPmnXPBthK5Dcd0Ljr6gI+kucyGDh456e009kKbr03EtSHT0ynR0hVWaWBV64cbGx
eYB8LyS/gaA4fALgbSjZ/eXypqeEMEHf+c9YxbkwzedrLnVB1U45GRVugeGxICz6+mkDri24gvdP
hSb6E+EAs8pqgM3K5RLqd4/9kSttFXkBfASGgYm7YhN4tn9+opIjxGlcikqnmMFTPlD9Zny51ga/
Gveitrdlpxs9mMJVwT0ImZca+dsTXb7sJrjn3u+zJwBK80UUasyyAzgyEfNBJ90KOuKWpHC+nQkk
pTxO9kgakYyG3L6vpjNbiCeQQnb7fqsLCwjFoEC1cbyfR55khhJetNAHNP8idDjqrJp3o8mQPS9f
yp9ekt8vXOiFm34aS4StJfK9gDVi+a+cYCls5wyzEkcQQD/8QPjshML7dlPkyZQYgiZiw4h2IaHN
Lpx1EmnV+h52TEiWWs9YC58gBq6z7vbXYiNLLBsCTOWxgI8ba8mEVHxAPjH3pIq64rWjd3RrQiHw
NTgDtmAWq9YnE6p7Z5K3mjzbSZQR0z3TgXSXlFgICqTffi9jCl1UP5ZGbmpcYSzWUdXjNa0Z3FsV
rruUSKMTElbm87t3w3PbbJWhqYqKv9lFDYSG3BzdbPgdSqzyBzs601Ff1lHJaky44Phl3PCnpA88
DPV6tFldd15OycB5YG+IbOIEicsqw36cSwkPgLw2DPdtTjEnVvlXasfolLmgnSvsfBz8L5JCrNbC
0N83JTetFG7qmv/U3Y9EpCt67dphbCKWD+Ep8cILSDFghmPXz2gYR7Si2QBz4P6/qybBSEk7CrZj
1+Evy5a5Z5GUxq2yMulgeB8Q2H2NkJ5fpMg/uuNa2b+HxE55zSzk8BffW4GHczj2ILK6SbdTLT5b
OxczdeseNPrTxHud/n0ca/3Xe1nIvl/7jRxMM/C3k2HbgyGXTZwFfiT6P5zo3gYBsijZI3XClKj1
ZIDDUPsBWc17Vl1IPK8RdGifi/B3jx9xmZlcgHYzyKIH2z+mFEMNVf08UaEuIUz/lstd1Vln7+1r
UXRmNO+Z2CHZrxDHr75QBE1dTO8F1Cq+PlnpvefoyoSPkBDPaK/nSs4AXfNyiEHiInyVHvV3ltan
ukyJnEvAJy9U9uKYMQUmGnasEw427mqOjPX0O6zr9abqCNS1/byU0FVyBzPIWqR1diQeOmFGltGg
ktEBktGdSyC+1uT3oJkL9mAhQoPac2x1h+FeIn8ooVT5ds9L/jnf4/IJcxsb+4uD/EPjlg20lhe+
pxYXPVrJgh1KPI3R99vtR7R/GkI1OgY4AkunR8q4aoAQlMnI7mXQGivycsjySszroD85aPHy9t3Z
Ljf1rLfzAz7YLzg2Y6MAB5xSTDMUtv1tDUorwQZMWsKJUQz8jX+ixq4c3aOA4Z/ptLz2LmREkxwb
qFE4n2Vfg1qSK42JgRxW/FghR861T7wi8lDopGfXvmRVLMAbIYmC67f648f6R5+raJvphWaKY2Ik
M7OscCqa9vwX0zt6RG/iT1cGgUAqR/IQ7JLIfqbCWQoc4gAgH47+FApL5SmvFVz2DRS3HnmMrOVn
eSl+mVMnslfoF5snrD9tt6CcA7ghYrHjWwF1v6T9cbn8Ijzv87Fj+lvfzXaHw0utk0MC+rIWh6da
eeBOvneA0BmWyUD+tBMOzLMuk1bAjlbX9C0+n0j07NLX5a3IAVoZokjwBgeT+OhdzTZgbLzISoB5
5cCX5kHEukyNyXW+dmoJbZOV2ejb58J/RfcDWbFUIJ2FO0pwOUpWybR3PRMm7lgTbdVT6Boj6gi7
G0KY+kgboHh0twIlvyZxjvpWemwa+knr717lqmu4AdcImb/TCEzLXVQgdIcjkNBBtgJR2lF+XKXm
9n1yicjJODLm+hP5W+gFfe70Mf+dLKoODHLLfWzvcX4ZaZBq6Ii+1GdChfqxWlw5Tr7nH+MwcPzj
on93gQ2b663agR6r46DOc8XRV3oiOt/wEx2Vm2xtH8rvtSIuExJuXCugoWkV/pcuC2i17hfGDHey
WozoJq5iEMsByxnwLsIDSoyVyYi9/ReWpbibKf2/gwdcugctU3XXUjPr/YpEO5RypYJ8xJVG8VqI
OqdiJlDlJ6fYjnVIaEsu4b+7aXi2Z2KOXHEpNJj9L4V4UjRYWyiG7lYmSRdNBUlYMIHWk7iIlU0x
WBG+cxmt+EtqOvZk171CBmuEuLoiEIfD1xD8rpDFcTfFZyQe9/qWwDcX6DQb+ezJKmyCWH/H6DSL
0D9Mw6vljGey6/XuWYnN9kEf1KSfSrcGDhW5JdRgI3o9o3TZx74/VR7BOxuLE7eBh+5nchp07Xhi
JuO5FURW89+Ma/rQ5o7aj+mDkFUuGgxSn6GtNeJw8blI/RL7DoiWhYzETIy7hCC2WIhSiICjxpnu
Nz7fSIW8BZejI/o0LDrhKu6SFHdBvLSN+SlrX1DQr17bT5Zeo45TQH8vdH7E2Pf99zb0QXY1qmoS
kxLuq5NqA85ATJ+xk4dfPEglyrNL7b8WHjUo5G2kNyonN6KFpzOh3iYw9IC6zqhAg+chLHoWOq9W
r4ejCWSLivwrciiblBIF6Y8K4lpq+d7PO1DR0wOSXfEZR9Eh5GQOdHcQDMdHvvAL9dNlBUCZyh1J
hNcR2gYkjhdOkQSk6EFUQZFTVaqFcqiXWb9lLxn5lnyWnZOg4rUKCcSGYWBFwLTY6CLxXItRleMj
58r0+UmXq2gROK6nyZbHZH+BCVR/nqMh6uCatVOg3FSIhCgXGSJPEZzuMK17f9+4Chq2ghvlEwTD
kudczwxSMJfwOqX/o8mN6zan3VDR8VDckfF1Afn0QIFTtlwI+Egc5+ZNHgBvrhf8GSeOUL+h8Z+3
IImiJZE2gX7qNxxoJt6uCxr7uHNPZOWOViHZt4Kr/9d8jzOWgd4204lYn07BauPGWG3ZhbCRAUk4
Immhy/TLp1v5HBF4bYBEe6kve3xhIHN2K82fanlqTIwu/o1KDG0kJ255waZ8skgAGIyDKUhtHlnn
sXW4QbVTSYsX417+sU6fdpjY6c8ZNyOoJPRKkPl6LNMZZ5jU08ZU6KGcMEBrSO4/maYSYHquPbMJ
XN3zHPTkGMdbVJPGx0B0hTEtjZ8BvmI/GSAc5ZLYLpDnESjYXRX8syFKM8SdkdFc1/6EKYZK+tDz
sl2xO4BKYVScSG4944runUf2dPTjWellUrj+zUWtTSH8ZQuvbDeDmFJy+RVqYF60zOZG3U+R9N3+
ffiEjiWY1zWPPEx3RvsK3fTb2V/cF9liw6vhuqp8ojKYYALRYZBTEz3fUg1d3i1/RBvEDED/p5xN
V4GzPE+AB0npwJ+3ePsFzH9vsbHWuWpo/+ZjzvGnT9zkx7Y3qTTl8S///kZRze9lrYhZtiiWpaNM
9Ckkp22jS71O0YFGVILx8ZBucNstcJ/jYu5sW9mCGhS/kRgSegrJAlfAOUImZziOnXQ+DNUk/86V
aBoPaJx8846jjipXsAxy8NGyL3u6xyz8GAYaVl15f6kSRsS4acPvvNWwsR3CWoVdj2gnks3Gp15B
PwPdXduDgxyI9/l/qzDRhDMFlj0m7SX21kEGp+7m5/VyfjimsFh4VWCvu5Ig7KNodZBbUBugkWDk
GDygtF82d5H62LyhFLC3IH3vGU03Vc5dOurUs0E6pwaNjN5fehrWu/0eRCksPBf/IesQUeAJ0fbX
qmdjzyhXEd5w45e/VSqe+ffYxVK2gzcTTASXkIce7BKSdi35wxA7lAOHmcyUL2sq2cbGsoChDaag
3GXSB+QpVOfeaFJF6w6flCF/jJhZaKez/YqbypnTOGa8CLa7AoBtV2SLJ1cuNDjhJTQbd97skuZE
+j92+aySHxQhoAyMG1rWaoxdcsSEK2+Dfwq2N+4B+VHQHxHe2EiI7l2GkToBs5+3NhGdkfGqkyED
wW1C41jSApprtsMSli8W+BxorNnqSxQ/Ux9VzOBi8UndbPGpUze4oM5/DC6JLFn3fY3IiaLBhHXf
KrfJyvjHddprQ4EpdwDapGZjw1V+VU07QyRRR04mH81mgiwZBml62PsxuVt4ivAELc4BIP4+6Vkq
wAPUnf00N0T4q07OjLXPZAV7f/Gg7GtVexX690MyYMj8icU0gSo+MiMd/oGjqlGeEIZFSnVzje8B
W2BH+ky3UPmVLTcUPFP5QzjnjmNQ/v/feUONqmpl5tMpykwlKYADtPMjqVMF6mQeJRwaQY8VlZ9d
zwJPzEMKkuRGkucFVGumkCtAxYCyB588t58kCiPu6BTFiHhezC8uBezeOtheUQ/XBFvkK/2jObTq
rOMZhKbHRM/qoYpEAosUhpR2Ycj3wfvcVLmE1NArJJqj4lRvscpAIYVJxJQyP3V8nH+Yy2pKV00n
Oj29PZSJB8f68Nu3Tgyk7ei04/9kw3YrR4FtkC7RPeHJ0ZQ+55rsKTuoKgh33IrrzF/iA85Bk4zk
TXnAFsD4vyktq9rebZnOIzm0OWamuJ7SZQVugkYJvHTtcKLBm9s1AHzUxcyL2ErLGLnA7voQtCSg
vaTOQmkpU7xrPcZotOOvSTkO5Ag3adKI3BbIv+AzknEStXT61PIbfpVxf+s8kNT1iSxqOLczsHJb
VGSeC18JptG8T+stsUfuxH8vBE65L3+f7VZPPagkgKw3G6ALgSa/dUge8pu/UVJdqXQ98+BQYXDj
fQ2cCMiMTSdzIGxMZ3UI2+lvoiKuQCaloBtTzr8ni0Kpk46Xvru78/vw5pK4bKIoeUl1I6V7ofxD
uGxXEItaSydW9knGLsjMMijhrxbTxKHIb1QrDHtwp/sqvevORp+f4hE9VwJbyR8Tb2sSXoP/Xf2U
ZRsMnu6XTsAOMRoMfUbDpokDdyw+llFPKGyBDEWyzXmkM16rP0BThRuNrnA9+kMOvdFIZVFgjDO2
BEu6o+70kC2pvV/yov94UCAmyKwE/zC+NeGQ+UyNxeGgleHu7tn3sX0DbKh7RXBz/aMtlcDqrjGG
9pE2gnPcV6HsOS1fq+W9cVT/VgilmvuHyPBT1lcnhgAe4uzADyWGb0D3qcNBkLBxWR6glqjec3m8
xIkwdSTUx3oAYNWsgiSFuG3uretjwxzXIvzjfz9mq29Mz2LtZ4lJba5zvpfpjjRD66VprpZjHlnJ
3xSSlbKrZc4fpeqt5gOb3U4QIZ2780CVVXkG0bws60jFG0y9VtmdmXa/0PnfzxewZASB0A0I0LvD
zSUZcn9q0zltEVfVEquWb1En4GPcnGovVpFB/G+ywUTZhWE/7N7s8d5DMmUpUh4zxW+XBeTuB3gk
kyfSd2e8eQxAujbhy/7bdzMN0JAvchQV7fLFieAsLtBZVlEwgdKUGFnpyxpoHvlFjKA6xibasOpg
58FRnUKzufMWoWBzWj4yDHnCxd9lCdh1JNIaGIQRA4SH5KqGmdVYQazJnBVwgw/iHBlxNt78QhUc
543Pn8Wyx5Me3z2HZb9slX5ymqJntBjS3H/0FJLhTOGIeC+s15/stC8rgTIllVgeVTJj7EDtZRZ3
HRgjwC4XzDkd8nofw5PyT4kGDVZ9u7FDbDoOPxH8XEJNqnjt9sZI3XgvLhL6FcgikyBZaj/Yn6Wa
X+PBeK1zcfYfjjBP1EF0qKdTJXmOBPrA5k1H87xh+YpTZxDWMf13+1Fsa/lyl/hcqJ3iNb96bpSq
7HI8e4HuRBt3X6VhV9NFVC26lKeh3YRt1xl889cj9ie+pPo9FmRJXsWhap61PtR2WNaXCJ8SSvxh
BJlQojv7uagvcpzqqpTi1D1BzjzVm7XWpMxxoPhzYXhn7b6sr4/hyDXzs5o8DGZ4xW2qf/Ehfmho
txXYIw/OX4kuFt89Ctqca6TtFJZ2ICvQeE4zjxI97W/lhgWa9ZpBTUnh+0bNjpULhezku4+J76RT
0sqBCkQnfQ4JWb3PCiyKuTr2DYU1b7iEHZWwpJCvIuSF93/ycYhlmOxsppSQiaKJRYXNpc5TUOt4
SQWLVZpUqsmAVMyzTUVBLMkEnXPjGcISQegGYcLr+fczhEzIYPqw5VfpNaaOFSf6DTAFdGIcFxzx
6Uv123TeluQlO0+IWYzqwH/hsTrbYhdif0iBOi2iX/2vluA2iomcYHatAXtBBiC237i0XrPeI91Z
4yfoagIQqDuwFeMP4AlNENoohru6vU7dzirzXf2i5ki4x20XaDeUucSM1JnmfZ0tHwe0JXUtW2Lw
gTg+c8qMKuFrpUNKoroyvd/6Pq2wbqlc8hTvYvFK6sicrOPCRDOgOKoedz1LgIbZaGJh4nL4to/R
6G05ojNlBk3BymFxfbbEbbn+RMrdQ9RTJXaKtxXETKEW/Ld4S4mbpQrcPFRYCuyidzs/v9TnwEeH
06iZtr9ExYnyCFZPc6U3mBDoMLdigl14tOUo3teI2YKEG+xg8dvDeZ394CtHIfe4AZBGt6ZARblg
TlUVawofM5OI5YVmqwv81u0syLL7u/ABDg8eIaFMEekfq8Se2aalNREj+jmuHzGIgspJWOxm0hl3
4XIJgtMnPRNI/k16Hg9Wt8LTNYQmzvui6w7IyBudj7gHHFWPB7cShgUtRby4qMapI6E/q5uQdmnk
BerjlsSE/Tucx98f039tKPrrPScHsDvbkicg1wltosv+d+ug/tR57oZVBBFOK6+3nG/CflNNkovR
Iawv2FFRwhqbplzkJ2fMXe/jFKwuS0/ph7NuUtRVpJWFsKjkoflGHhmFyv9i9RhV6NINYxeDEefV
sEZm6qKdcYalvBp0YOjfFHIrYyeFkeY6SRaPQfuVUxh5M12+WC3H2F4OAjdUPlJ+pd1jRNeAvMFS
hbNrTd3A90a+4RO6rWYqJD9vZxI1sRMSmTo/ID6uAtUiPPFDodUFqqPY3Fb7L8jv1UoxGR6f1Z9r
PHBE/n3PNdgHVunRKUqNfdw3udBm93/ey1gNL2O14hYq5cy1++DrXW/SfS8r5glhMJ9SQAK3RqDj
h5JMQ6ktDxdV717djSM2qTUP8wkbVm9eMomV2j/n+OgSnK43iarB5xAGfsRrMw1aHwfFtzImZddi
RcTaew2K+t4mZy9gxf04d3bOzsyN3gYi2+UpHlFuc/XSzlnMr3u2wqF6h7aQCLxkKqe8Kleo7SJJ
vwoJXgiIs3//lHc8tiCXcfx7NbWQaKC6FZnGpk/peQp9vTGGP6Nsi1qnYv79UY2oQUmLzssnxczE
VP4ys/tniUoKVGulXMHDoSzghKzdMFkKTtiGFqk9kknz68gyHJTLndRjaNxsRjvAJQ+0tL9YlAZE
VE/DSC68iVCmirsDNGlIC3L6Vagu3ryx+D82NvufKi4Gy+FYr14KYCSEzqg2zg8LtexEXqu7OSvS
SCrI9epYDrGfKM74+fsw3wSTiJgVwHp15ZACC2fmmTrj5jhHuzTZA2xxvMuqjPCF6cv0V2+Mngpg
IGqCC4nAqWD3tM2IwKuV9zpocuDn+ChzXV52x2H8fZXjLVMvLzx1SVpecrBEMK6d2FbpubPi+kae
C0va5kUczBWu2sLCsFnprDk6sK1lb6jG1uuHBJi64BAMsWi2Qe6WYlFokTVIhOZnVqMfFdugGsgD
oJ8a36BxRqfO4MNJArIflH0SkoDvlB+AAXn51wdb6DIJflSnWZRyLONAy9oYVhifvjEflVwMZWja
H6/rOFyCTf90wZ0dfRPnLJ4FPn+nEJ1QTpTE21BlsfcpwgIQ4vXzRv0ge6qzRil0q9gBnqbZi6AA
i6xyNPeMMCIqsGoq/bzeoFMo69q+J64YH/yHi+1jYjxOGUqS1w8LCabcygyVuQIPntjKGRq1EepK
ErXnC55s94dXYSBXh0i8eAWc2ADG1b22ymKFTnsM2MYOij4S+7TA3MakWsmtv0XNYNes9zW34M2M
80lGU44Htw0/yVcc2ynph+mM80NlMyLrskKMvmI11Oy80qeuFUuV+Tn9v+gLb20BfPRa2T3YdWWU
dTdboNDxYI/lctiiG65IHnDrljTd08XohiDC37Rg5ncbQfWN8H42QVbfs8DDb0zy+M1BNTL0yBAt
g9VnlL3FLpdZj/GZF/sL2ONR98KCmrScstFUWhiJv21fuHENapGb28aVA4iSoX81y5MN+LsLxKz8
mnyVvK8FcmES9/2OQNZC9WcCkpmLbPDkP7elMGMJ9ZrerE9Znl1kwrWQMoeqbRkGw0B+oUmIuDYF
Flufz3x9e3OgM5+x+39K6dn+yt5Ia5KktmacXhVRDdoBiai7v7O4ewK0Zn4MC3HT70hglx3D0Jyk
tRJFqGblhmu90YRLZb8253Rf97NbsZ5eurDo7jzimRgB5W3DfHmzSDAc9Cz9RCVlnzHxuLwirblL
fTfqH6AYzjVI2hsFLE6D6DCVhgXtaCUs0f+dcwCudZ6aI150/iC5JY6aQuDft68/IWalgyw9kG9e
1JPAWsrFax8JRq09e2gskMSuZTXIGRlGXEpdnYPaWyLg7yx6R+QbPZq5eBVAFjjVbzDIGVZTS38O
kFAAlfvuyONcUMI3zpAlT3c1AxN1g0djfX94Qs5RczdjGDC1jMTapfW5A0rN3mNCyfKoyBnqupki
UZPwysrNr71bWLv/j/uiYwYqFS6pTssYfVd90wW1kjfZAVZ/S4muWFLGDWi2fK3CYy5+uGfFPauo
lYaQLxFhznEjt7DMdaMypb5W/RyRoW0Qy6puzW1k3/iLcvOKunVppoxlRx12zC0ejzhnLBr7QQLR
A7iYXFhj3gLptJrCJ8C1Ov3UhjgwQb+InQjSXpVnY8Xg3aoOX1/1MLztlwFLPuOo4AHLmwmyQnjr
LpwoaQj+94a3eO9zI05vyK/Iqkki6ZQEw86pvTWZ29xUkuv8d23kkf94m3Xh7dpHNrtyB3CVLrpz
RsTaSMRsulwO16C6lakTeP6mZnDn2XbCvY4Bz0G2xYyTaSrxi/Pvn2tMiZrEYrrUulOepWi3KkHs
RLoue7wXN0Vw73iyuluYb+WDvAX6TNhIUioh6suD09nWEUOS4qa5pAVQAMkl8eV/yibgIbXs2NWz
A7oqFNvJYsqGywh4/ock4vI7IrB+JW+5WIQW8mtbpJQIfaXzqks/GHPWag/qmxyIycdoq7Z6Z6N6
AoKYRTzkiQhfCFt7xUj8vzLLsaFDszgwnnpEhbohYnpHFv+p9Hj0ISGDcl11ErWZUtsxtSHAHS9n
AXUrt+32dbmU9d6EH4XHRL4g9rYlyHjBaXWXizLtwjpZe3Wc1escq2tBxPYYoysrEbw/n01/Uplw
fRSYi1Mme64+4dOqVO3mTV8ZnVAmhsvjwF/9yTzQUB4s84/7CjkX7AH3c+rFkYeee2qY4a4cFfKR
rnwPRr8avV/Bm29wuAD9HHWVrC0lZJek6K8lHSfoQxshzDlMaQDUZZZlP3e3awBT1ja9a496VcY5
jrBEz6l836jRmpeKdujTPrdjQVjbNGeLc1vq6BGukofbgZNkxQbFca+6UkNzlJAfJbRKqWFPpH8W
3Z0TWPXkV2wWZjrtid/m2Ps4sU5dwgYxhb0mbySa5FIFSRCq8MhRAxj4psV5VvlMnzKsSHVpEpby
6fPZxXIDCGHGFX5U4wf3/gHYqNoClox4gR49BqdlSEQqLiSeDqU1dLwcJ2tw5O0yZWsyWJGnXhNN
fnJeiPaMltTAXvxwtV3KisZLqVE3FI15FnjQjOe+eK1zOb2y0KQ3gn+IpNdKripHISuSyaEAjRV7
aIteGzcrZ/tnl5vAyaUj7WCA668iSrz0yk0tTaOJqRpMP2Bn3ZALRLR910qVDA+eH37IdSjLAURx
fzHFcVgeVP1LlmONGvTYopP9buXU1C2Zbv0M4MWh3g6YRCzo8zkNn4VJDZOiXsb58qwkFOg5LC+j
CPQPdIilUrAai5roUeEG/JRdtop//2llQx+I+lFVxf2Kwq9P8yEg6etYpMHmwwU47wsYe6q7Jr0C
zhHvnfRhu/FP3QHtSM398PqaolUVSrzyk+ByXK+rHRh0FNj9KOJCeWwjowJTg5r7YykBwEFxH30b
rmxoc87JEj1Lhf3W0MEkJzChN4Jo3AB1X/LSaz3oLHWxcPGsAO0/bpK3XvRdl8RE4UR8zkjpxAy8
k2LYUbYSSIYo0dxjVcHRDHZFx7n1/Q+4caAD0RCIYK4GOnmT3WFit4VXZGbKxmpyidm9GwEDdoXz
FFbu50UJPiuCPH+1u+N7TCha7vkPlrBqXARKskyBHkmvYTngB2SZJXfsoZLFnc43jp1TSGX+n82x
zGEGmlh5j0vYSGK6kxzbnfmQYs4GmuFgJ+zSbrW5PBptYUDAFue5GIQouaIS65Vp4dIH99GecrzD
fd8RLAueBI39o+uxsJETaRO2CJLTRzoy91YiWb/op2S0MBfxZSLA2wWKcD+hwFUOH4axjeVlqlkB
Io3paXWzZSRmLRw74C5+ggkp9WH8KNGtKak67ykegHtLlOGLVyEiLaTglzS6f+cAccOPxdgmXr0g
wYr9tmApWlS9RAFm2TWiE4LCrqPiMeZ5BGueh6DUMpo3DJBJ8pnrB9zt45fEd0pd8T5vldSjbv9s
YzXMYYPCLgu7Ko89hzcaP2ifmV+8ER/JVIaelo28AtCtleAqTN4mwV6J0dmd2j34LVIqcsjh+Qew
xlmO+BFTGUBYm9n62MKihYVWywA+vtPT7lw+HmFfRmcBjgjeJP6rvel2++HA+3di3+oia7/vkFL1
zqBza1LL8ypysX0sY7zvA4uQ1eae68lbkLH6rI6JozmO7EevjvOB+pg0+exk3EzeMYacRMpWyc5S
OY2VDr7XVb4ih4pHjupG11BOIzKfezQD6jATsf2UKfru9lI/Qp5TpP8mhSt31kIgGhiyp0tI+tYK
g5NFtlEqd31hkXiwY0lSHBiMXerPwC+7W/6GJF9nAckSClK8iiPqRgDz79wyJrtegC6/DN9og/xX
2Oghzz3DHVaogsuIwJ0/gCJCo3ELGQ0BFD4DpbYThatUbI89ociR+JNO9lytsmWfmWgZwLg1BRhD
RiDVhF+i4kCJdVKh2d6uL7Adg9kTRuf2YKjajNE+dCBIdE5pCwv0+nKD9xyWJNntXap1BL28DjI6
TmtSQbNRgWuR2ytiEhpLGhZkBMRfe0F/YIJ56YHfLUm5c+Gxzd41PI4532WwpYeEbG2OlE4e9fiC
kvCN3gWvk/+B88ppUC2n8BCj0DYQGnjdB7mHFXOsNMoQGZpOhXlavBfCCrT3EUJr8SZtp+/W030a
hpv7+G6p8H/2/d9Lf2sqhEm8Sq9W/BjSKlosc1rK1ZFfjivY4AySRFIDa6AMLYGM1zVuvles5aoh
MlxL+COH5jkn9bdK/JjWN1KnJ/lU3PpU5wylSP+057K+RCmtJ5c4yMLrHrCilgS/P8kV6cG89gow
gxId0953rTKSNvqhuZp9OfgBxOCuZqacKiht11qrAbJFYcRjhNC2Yk8koDE39bcw2+/XyZRPHMom
EZGIfhZEz1kuJOTuho/dUsJRs+lkj5Gt8NJ/tgi8sT1yj5/vWyJ7iga4nfc8H5Jefa9u7iY1Mna9
d3GkX7/FALGcOpNpg56DP9OPabeep7/sUTmW5l5H7mUDC1OJ9i4s2UUZPMMz+/eDMnGs6cKjnd0J
a5RWuxfGkFtISq+0uH6+3SNKnb/SJK0X/Y++gxTxs0y8gMR969lMH8zaWxdtUpQZ0GLKyJpJSe/4
hv5XHm8yBufmvJe0DvFmM3ZTW/+UxSmEoCkPcZgSmVJrVWzbmhzpFmvQpmSfD+sa2cH9VZKELQIL
uWUxjO/hNJRXhYeXZwiF0u3Nbo0gP0jHLkIsBeFgzeeGZx6C8dQSq7JQnMAETE5VPD5yT7MbNo8T
TKQiSc4mdScd8mKHSITUDTD45DKslS/kaKumu1ri7N6/Triu4p621RCzEhOKHKexl1dvTd0EMK2G
1jDrUKYfzGxmQ00fd4wGcetuTVHjGl939QY9BKk1LlY8qOEHW/CiInBO2c0CKmJOQeOG+6GQOaZs
+QQlBmHYBSU2yTDYX8joYVvRFpZp7e9YF16bEWyoC0nr938E0J6e+iD/DGzWvVaHwiqQrrzJIdwK
RNyNMlOJI+rFQPLnU7LlJ5iGk4DpDAEkg13otxqNyoAAFs5uqOpqeQBqlkmnU/VSdGyeBbChaCeH
kLoVzg27JOg/umpDdyOUdAM0CYSme/Mzz12S8s6hPvsTxwNQpbHV3UkJ47MF2CY2n4ZLeB0g4xxo
gYeN3uLC/zYWwJvtPqxOk8nF+mBHwnLkDtP8OC/jWEYLGfHQIU7EwQvvK6IPgbxPiWPBJRxZAFIH
NVs0OSAUbxLR3nTxl7PRgabv3bt5hkXcCCojSYgyExugC0UztIMYpmXWpD2WSUtryQnPmjHLbGfL
IvWwvQxM2JqOmvsfi3Vavc3v0CpM64eCe1CRAO2xwHNyy2387ewLU6xIJZalfDMtnq1E4uyzXIRH
YgsZfMfAy37Kk8Cn3hqI2eXAMCRZlG0ICpfL+uVr/3V9i14wIct66Pau8NYQIrA9CKJjIoL6h6PG
vK9qmLiE5A9JM0QrdG/Pp3NE0Ocj0MnHhsCMUvXhIPDGrw2sZFZcFlePpwwW2wICHLFMRQP7zHz0
jtF8sVauQW7tvmZKfqcNW3Derflyyk6JOuXZXCsDfemx7dHSgxyCmN+of3zkA++OWyhztmYfIEaa
USTo3Rt197pR8wrTU95yPIp+uH8BEobtcnsd3hC/ZMLPfR1+BNoNQgklMcvnpFaUFID9lTArybYC
uuiZszzo9tCJL0k8PcTb8BTBVakEU5xVpr9sixWWqBAD4Iyj1MiRjDiBpv5lA3jMEhPNTTnasGES
2N8PVImRgwDRcmWeP6ELyt8P8XPZEdfl7dD7VQ4UmJFH5GOEKe+Nnav3JZMNzV61zOaLKhRWgur2
3fZQSQ2QJ/YLpl5EhMimHZRsg4Qr5IQWUwwOhTAyqxiKz1ujjDpSW5HqMNsQPPZqsV4BO/UHysbS
b5Pv9wYUXpilQTfAVCHeEcWIPCsmzsoU1029bHnXJiKiYqapP4MtdDQrQkRMQ6UTI0w+u9oTadDU
nEC86rEjjN8gF1dSErFUQP9bzKhU3vJBURIzMvxj53wIU+DCHoV3b1ATgjVOz1jXZ83OnESjlJCy
446gd8e6pfXDE5MSH9MOaMV9k6jj8qY7xDuPKt6Ommj1HOdMSE1G7EOSjgohAr/Psv2xuLL8vrh+
X1J5gKdI8CV3336Ksv7IusT4TwLWfq3Uvpk/+nbxgtNVpylTxOU5aP0WV51T0z85lJw1pbk4OSMh
g6vPn4+h6RrLgt1I9piquqOUc30xVGdJWNaLt/NHlpVMLiZNnFkDwB1oM5kceCv0vyLAv4pTPHcY
CW3f8CUSz4Pmc8g8ZLCrf+d85ZR9WyKOt3FJcZ4jWC9haN+h5WXiCc7LHNbuh6MlD70SDSoiW3Nv
XJ5tEAUJlZAPZYdGvO5ubGGU1zp8hchjEMvKbZUbMiPkzi5CppWWCInjNO5PkS3ETTgOqeqNzSUQ
Nraw1VCdQhx1nn54Apa5yjEXCy86e/4KZ22a4R6S61tFKucFmFQ3e1NZ6ou30G2ObWPpdauRtHjO
aMwSPFDO0TaivArqgVeAn+T+A017HGniJ6OAA8WQfPFndkYq+PmpAkme13Du9zvj3jZSLwS47CCb
yd/Vu81Bdas594UWUKDAwfSmp5ZaX30e/H3QZS+7EgEOKtiDPdBsyXNjrg3XOmhGsqJztryYMJ4S
BqN5rQjm6N790LDsQYCiU7RA7mzAgpkhfol9rDD2hAsDXYj0fLQOmr+HOLD//MWzP3kLXA8YvGBC
pHAl7phV7TqcBsyKb0HXFnYH8itAUWEqlsECJ7XDU7Jz4C2mKQDiLSJI+XDcte2WLxHVdQgkDUlx
oPFYEJOKbCW/gTjDICbHlIL95UH6o7jVYzHfMqVTWjJL8TqLcPXByx70rW1v1SqHfKhPIKtQ82iI
ZUg70onxcnMo/7Vdb/ltpt4tT4lMFTVYZpYtnIEl2sGcJU3PdKvGkvp69kv9roBz4JYMF1HHruau
2P3tYOvkon6l8aQ79zKviZ5goAtXbKVNYJL0VaFtarWytvKoTvnhN1JQUErBaEmqE60GkY19jO5E
udSJNbyCvjjUCapkQSmKGQ7NPEHRUroYBwtnrTUaoyWlhhhWnBSEGNTTeQqOO/324AcTaSU+aGW/
rGOVqswZqGk0UMSrVk7Kz6OiDfy06O+9pbsTchUFRESeQkNu72c5vwfRsL6BU8JTMvpTlxyMyDCG
zqSkGecrG7jO0deXklp46qKylJel5BW52JrceoMeulF4LrqgPZgP/eoOHYQpKMd9ukCqHBlMpofy
V/FTIgVMwJmrtG31LCIM3pPL+rkWMgYewI016e1SPMJqCKCXfnihNCaRX9PU0BJiJES95Z3m7hEa
Q89p+9qeZD0JbsoNtIRQ8AYa3wcI7c89/RFiPqtOUj0o4EPN0g8T2HSkYishZ5rybzKfRAELtzBE
WpRjNJJHDm15hndgmL08FdAqXjKsuJkFDgwm5TA0OVfqftVJYVswNU1bHzbsNLaZpr1zUse0vCe1
w5COWnKQJBci2/gemFiQ/zRJjRwoUMQF78W73evgPBdVooTxdVMsR7r2cQUsY2dpk/wMTF6q0MI8
CmeRyRvcXKBwZZqbMLxhXJ5HUYW7zF9FqsDeRSM4073SJ7zfPfcjbBB4X0Oyw4JpA4OdXq9S8qab
CoZSwdIhz4AtEJMulLH8RQi9Iqsjva1M4/50xJ+GKvRFZunCr1EONns7x8xpE/o2/8NjD9GAN/DV
heTyP5gI3qbE72+f560xNu/Ex2xR1DP8MlEXHMTEWLEf6Tbqu7S0bkHC8MhsvvtxITzY3fUgVxwl
qE3CReVRnaVgwpnVoRJDpPnN3vG0jvU+EHwoqimumSCxE3FZJ4bgNPLnxq7v9nTCvE+YZQFCqcgJ
NghUN69UbqYFyiBzAKzPAZaeL20jNvHNq+L+Gk1v9n1rKhIE8KPfcfv/wDUSCevDPXEKg/rFpmj4
RiEUSBkXV6+vBGFvmNPLVYFpNb++JPHSVVdGU0MzWCWnvzcSF89t29JWMpnl32Ptq+G/i+sH5qaO
/XImiybKhv+qOAyOK3tYPXyC/aH4gZrMYgdp3ODUQLmwPQNEzLymjbkRkm0+MZMrtoGjNdBKUpIo
TY926YnrtDSLQXdBrx/daOh7QPh+z/FsF026iFp9jE9vqt43J4g2wIGuPvypqkTTu0NPEQi6yZn4
7dpHKorfoSTlGSYxNFl53VpGXl5JKJ2l++nKRFC63La6LcsamaORGWk7rUZSjxOc9KQa7EfS1Iuu
03RF39R0aX+GSfP75+m6hIDcdWzYbgq/Vd9QrgGZV9FHZD+uR3WzZ2xNSeZ3mmq3QShwsT3Jm9Jm
VtUioamGiQou4F+MXL6ofpG27tpTv8RGyrPess3onjsNPMs54cK1PToS++WA2TCBxlSwao7gsrt4
neyRpgwvrCsvPlHCIYsyF045QzbXy7dfo2aCgI1gXqi3hefbib3+iKmZEJ6kieXSlANlJs8vAveM
FRK7FHn6HtMM220VxOnMwpVQDqkZjHDG3AgztRww6rx4hVO6XK6Wcv3Jkz84PIWkfYuWQPMDSlJs
SA6Dbl61hekSzWmdnU1vY52HcHmcYbE9fmRMBhvDmWU1ogCVAC4b4WN9RBCmGkWo0HRMc6RI3Bnc
d0q1kfD3mtUa6V6cV0L8tMQn6zVGAOUh2LPLoO5FHe+BK0dBZEsBVdUexne/2uXXb/NTrolfviUF
R9r8htI+Bx1zk+fhCGN/hJrDVxtbR8tzN8bkn0npQVPtUvOTzgMqpiXfAS0CEYe/fNTc54SzXJtD
64c7QsOVzu+KJKaR4dPp8HJz6yGkDj1p6pT7r90Lih53o61ADJOEf+Tzgt3m9qgqD9L4P5xrG8KR
JN/qONR2mQOQCoZ/lIWRjisFNACggPwSh8Yjfd2B3NVIMBXSqqB/H1GhhRo+8GiZ90ZbjFhAlY8y
Oz+KoxuHUNWWjRye8LJkf4bj4Vxd4Z+MZKJWjqRwCLhmIBvPugd1G9GnzRL8lzhN8hkzztEA1cSv
l7CY4qewc0rjjWehwL8G2B8YvRmdsoaAyJRCUSV7YcoTiH/GTXDYBtNoRLmr0lzKtFXOu66Ue4+g
pC1+GPWc+YVszP/nlaRTlfx7ri5+c1mtO7HEyIV7xZu/oJsiLG6t9seETnC0Lw0t0Q/3e1SQ3Rni
RY50A7vQyrc/OK+mSEtXNdTXLUxIU5oS8gpSPaXhzD+iCM+pgF7k0KfBm3mBpxhAVIvgK3XdPVfp
t1Y2Cv0yiuy9s5DmRUQOb+Ac7aIB4+u9AxXROKbkerG8F+sjpMmkARYY5YNeDiZV4aWvlvmyyARf
XgeCOyAh1M/SKO+HP6LH07ubgIiBQYuAB553Qup25fJXSPshNBk9PkFfOTWIKuPJEgb9aRanzC4C
6Xpq9byvoGinubJ0f+mO2+QSx3H55o51rpFjWYW5SS8D6WHYu0J68lImce1pveoD5vhSych3HqBT
W2n9t104Q7KzEWZdssBjjG7BJ4rBBxU53x+sGocdzj8WoLGJVpfHOWeJHQrrG5jrsXAe/fQ+yLf2
+n9KMDwlGbs+ywuHqCwcIy4P9CdHlJ5y70KW5LQfQ1qKl/z6l44q+TDJLfBYv7eMFxsCFdCQ8FZo
87v5B6nXEW/y0P4jJBU/PKL9WIHL/qido9zU8pqoDuLzgKKEtB8HLi6WiTa1bAEbIKmzEjR5nvI4
UCcnaPbSuKJJpPyXFH0OB9kDJMogYJnMhBKul6NYqQVhdHh8wcAp/Md/cME1Hjw7S3awDAprPWAZ
ZBX+AsDp6Lj+M3zkr8A+/LzwB9QbNcBMkzfU70bfnoLSfR9INLQinNovhTVkTPDc7/wl4vUcSVjv
P16l+W1mhNyFypk/1vwfig3B3pdX+vQcMLCHB6mheJj+KyT9NDr6EMczXqi5bPRYXZXIO3zybaLD
cLJgYFR8qIp64QtVyIfz5eaI/GhZVotigdNq6imOKPAx4rJuap/JkTZWPR0siX1Sz/ZJmGYkpwBm
F4jU98zvDK5S/71/E0O4MMQbDyJLUvjS1mtjGkkflk1KkmzI9tNEdOxJxpaOubH35jzRTXCnnNfq
fWwr8Xs9dzEoPjusf7h6fmO2anVGTx55ztdCCvSAfAkRnYK4CYlvvGO4B3BmeL/vYTnpGUpPXUgL
Pxdx8hOW1sf8vwN4eSl2RJAA17xidSqWUje7IcKE/QGee3p1JwFrIwL3aJRk57wGwBLPDrBCrfO9
FhYaYq3qXOJC4EFaulI6OXU8YYmWjz/MJ96TTCKCqHOZLNNMWr5LTxfVQ5s/vAeBM+8r4S65lTSz
jLS9Ij0ayR9jhIAOPN0EWw2a3anJCgROdlqq8O2BUqAqBa0N17L68USnO+U34QDPxbRVVD+DKQ/Y
aPqN6IyJhAqZg3tsG6lD7Nb/L+roTLUVF/bDq9EwcTqqtMrMbv+CmDR7jNGORhlQhdzh0wngvi2p
TGpcIghb+tz0zFxayQUaoyWPS+mTB5Bkrj4ABIcllYJsr/CAVyW0YVem2rLxQYnV2t54aSu5sLEd
+j321J14uLH5SPtHN285gj/A+VbgDYKOp1AkBYHtrbas/rVdK4M/KF2H060W516D8LyZQ6R0z38p
79sPSvjwtzQdezwPbsBDU/7w3P74hQPzbe4yOKf3hXr2VT1M8lh7ldGevP8kVgsx/xUPYEgtWxd4
xyH9HgNl1DikxVK98+aPqy+qYYV+qr2Bi6tzfU14jK4TYH2CS5Qk5FHJWp7ouMxH8bLFUpYdtSdw
pVzB8vGm04i78EM0v2vU0UPg9IzQFq/YoSOBi+NzYZuNE000P7TRbZhM+5KRyuBUeyZZm1EvwonH
2tY9YmztxiwfRqY7fyMf9T6+UiNuiBmOiVUNs3s54prVdmnkJZ8phH6EBKR2Xma3Tis5T7sksf5a
d1YRfCF9lRNaBAX+u2GDY4LedHWwAygkperue/mFp3KxlHIAhHczCU59uc4FOvJmyEKcXKECPW5x
Od3NJrdptAFQqLZn2zCE73n+6VN2e2tnNT8NVC/yXS5EJjdeXmI40p0HFO21BKCNUHDRV/b88bY0
1GoKcXBaLY2sa9oD2En5igkyMO7l4y8aNBQGCJ7gn00f6wrgW5f3QWOSf3DUjM/4uuU6/l17NnNU
KgoIjgMgpRkkLnCczq1rjO5oycnaWoNvVyX1RH9ZOYn02WFSrla+J82809BH2yf3Q6YoF0zSKRmh
a5XlCCv5B3nj/6ITr+W+x2vwQqjsdiXw5Bi8xEwvhihbjz0su/GMMulJScX1j1C/f7MfKzyv25od
yFY6sWmXx7z3bun57K/zFjX5j5je8MnzXJV3/07pqdlhC600KRl/m20of423LZyhUKIVicU204n9
ZCCejRqTp75giaia9T4jhKswdXiAT3KzlrMg4nHujj/lnYU5LiGS/i1rn7y+iE6DCi3bWlKe4sys
X3N329aMz7blDNsnnBHSP5fSyNG/NwUtpNt/zJImAyBbtJgUKoQEcNrc0vB4BSfFT8liSZ7ok1Zg
i4GDNRo417jg2NZRUxL7KewuYVE6jlbt54+kM/GoffZ+OSmuzi28LcoqoR+Bdp1cPyKtYl4hUTPr
KufYsdC4yw0ddpBgZr9F15Ttl7cRZtBlVkKVjx8mTRknsIIQgzAWBhdwfEZIowNjaDcKg+o1s5Z8
ZQ+tjYbVqq7AR7ulyxdetsEe957url85nF6TouO/nPF4aeL2P5/6XhhtR8qCYMl/Sy7HSDQXC3+/
tUSBRMg5nCm4RIiW1Ofrf/qJOYFiKXZjM0MIK2hiXI9xkyToSIGAs+HmZK27dbtKIHTrFxBttBcH
XZlCVgtWgE6iJzvsUwtT337xrPlIvj0OnyPX/w6QRPBpMwFfesN3jbf+rFpXaJQpHJdkcGMGiLQ0
Fie+QQP1Tj0VkY4wf1y8IAUlpLoX4BMaomT8VcHPqj8Ttv3CcFUWz6xpNaO3Q03lkYkF3/MIgM9O
l7U3fak6/2QXVBXvJ49/E7dt4YLKUwtDs2WjEifCMZwmimsP31VAh1J8/8YBPlOJVmkDPvy6lmid
efJORMAGakhoTww+lzjuovWeKw4Qc3biN/rCoQg5SRIdbLh1PFIpWjHVtBpKb2Xse8Dv8poi77nJ
mrorE2huOdICe3hC433qIanvoCy+RK0XE9RZ/Vms8C+uixxVnQRL3xSc0HCcqjwTc4Ids8s9vfht
j0GyzQ1oLoLK1nF2qfj36tqlUqw9OsXK/UOPUE3NtIpQMb5w10c3p92KenGb5OzCa7++50/z/kZv
Wz4fxwC/MVe1nnUTIL43AofPAK3FgavtId48Ap7nXMviMOiryXzCy3VinliUGSi0XYRfMKzUPguP
S/n8++fRlpfqHkQ5lbn/6Fpz5808fmOyOr4ULJTrFKXdExyHZ8n4f2SnFIwBYTcC7gpLtJp7AKUc
OByM53Lc+8WejxsDDnm0x2RTDSJgJNtRMsGDgmzNjAVR6cyzaUGeJGrtyj48HuefUxSa/1//wVVQ
NeYnFe7ruApg21vI0QYQqqm5sJyAA9Vd8SpzktOh78+LVaZoUjxdmB8K0ntLrdGQs0r3NbmAMWWX
D+u8BLTKKURhy7jcSJfsBMV7VLX/Sq45JmAV80IGkmVAtMujr2kK6D35GTiiE0BGUS8+8dq++R0Q
0KbXy9+MNSLCQAxC0zSOl3ZpiON/3o7n4P+Lcf8efdb1gg1piXDEkaLQ3n7aIXs/5YRYRQ/Nnc1w
/gfUsI8VmyfFQNSHT/etqN6MG3wgH+eB4IT+WF0FISfIl2ZOGAf29wDlFBkHo2z53YyPrciMyUV5
iymuqF49bcke93alfuln8PytYW/zpUJFCVMzggbIh3n9sgFPYWksqaclfA35d8xxtfDLlxU00Gt8
Iva0kJolzI5URJv0QNxDdmsswKsKJYEs1QaUmUXJDjvq6LpO9S4/wW1eoFDSqINjOI5/jd7umdMV
/qgJS1PY3Nmcu1+rK/DelszRJP9yRlNCrTNcDKA/zR4TRlbw0eAMJPd5h94O5DmMzunHvuFrWDZM
i9i+DHAj6QTBrTrpN7dZIE5VZohBIOt0junEf7mtGOfq/h/MpW5g6PyqCK/a/VucvtemVrzN7NNe
GY2v0AhidKrUuZzkCqW4ajKu66HYPpWwSSJSlAiR+4IhpW/HxcQQZAzglhNbJiqNUyzOhpOYbXde
tcHcP+NdXzEg7gCjWknRdcVxk6x3LEqJY328/qVzNh/HHxsMi7xCcknzUGEvcGUXGFXXBdPFF6Hx
jIT5FJYoPT4IAxN8qNunWOKXeqhGIIYTkfziBAp0LyWBlBaoR+3/CM4/IGvXfXMQknVdEeVO/bUY
ccDPanXMfWCNUZo3YUPyZqzbTjDsqwUXscM4e9rUG/1iRrItJfR0mJ8ww+ttqVlnUXBQT8Hiuvfc
16XLbWOX2jdrL6L7cruLoFI5qf8To6PFZpyOEL7jIPM0CoZ9dg/1AHWTZuNY6TycD1DY/1a3LH78
Fj/NoPYP7bM7ptmiuwdNCuH+EGT78+X2JuaGS93oZqBBtgjWcMQRopqCmgU/BXuLSre2uyp8xkna
byBF0HlAuG+E2vO2bqSJIm3Xr3EM5SE25g/+JzawgJuEgf5NvZ6+OJa3txIGoU74r3w+/+WOZFvM
Pwkdw7S1ei2V8ip2qIrJQAZp6VYVsWQrLpfcmiI1NG1Z2dajMiBtWT8FZCg4qtCFJwNH8Z2uPTq4
MRSJNcN6VL0L/MOKRDyS+xqy1ODuuFPtLeUnEKgO/MWybzovNINoOvH9MRIxM7JTA+hHnQcULVYA
Yp+7CeAG0G5sw0Py1Vs6JJ5GCYe5DvFm7yo5yJvK7GMgQ6u2ZuQpyySZPOAtz7+EwjThRSztKHRN
XOHRXdtoRlx+jfgzNhcL+szLNwTAW8YtFwcQ1sh4/xLDi6hMEsCijay2a7u3ZNXq65s6zDP7zmM7
en0RJ76a2zZ5HA0Ctf0HOPFfYmpdzHqUNm9LMNySrrxeKXH92n6XgiZp2ZpFFihlDYPcgYSBZy26
legdDIQ7f2Lmi1aMdlYiCj0WMHm/ltmsIZnpaV7dHqf0DSUKAVLrVeNzsbwURQa0qRqmt4TLEgWF
Jqf69F5VX73peSDlflpUcGfim1IFJViubcFhTwHqYiPW9WfzdA5KtUtCq62JMbuacX4lYN8sYJRG
7vWmib5eu9eJCdG+mcTuu4GhGlyHLZKafTglwIWI9CK42sddj8zrjitAj08q4izB8sfsjSv+Y3o8
e/6riE05uN6b5V/Q44eU3iNYNUcxrO0yUDapOEEke5/+UVXJrPQTtAkibu399tIna7WAQD9DELM2
o9NtTGOtdRSxltLY5Ua0acFOhpnMhf3DYzxxDr+rMy5oCw2zizCULGps4Qt6xuC31WCA89UxvHUf
COu6z3C53VyYPNBWo/D4t1W7+lEF1R+jczMpNh7L8Zz3Q62EAXrcwkd/LzNh77VKUpYxytbUYXod
CYdF4Y1lMa2ImD5kk/AilZnItQgwpa0Za6b3PaAYHj6DXclGE0KHruIK/XAmkTsR82TF+bG4D6VK
OyS2HboG5rXlARYF3RQ9iN782rYiJkUmXom3yVHHJWajFWurHbWQqVwD0YXdhNcdT4r4k33C5omR
G75sdFTFfxWQHLisg1vLdawNpoyav5lvJtISDqNQSVBHbpA9qiLz7cgO4n6d/3Os8/Vx67UWHiBN
SRrJzhr5FiIR4WfH/18uNd99+WYDc/e485Jjqzt/YMzlAq1n0QOzLv9/PCEoj7B3QCMZT19w2/4u
fOAdKZ8KpxMba0kyMk2T094Yq8RGKgjs1NOJcVrwk8k2/OyWIlwWrV/41SXMCKlelvmPvS7/wN3R
BxG8vsqLoKA3beY5ScrQer5FcP5BsE2oxRv3zrx4jl7D0t9aJmxrH8D+PM04lwaEu5AednrAPs1j
YceMDULNLJkPDngVes4ehbAQZ6nm22m+wpRgtjQjHB/PbeTx23viEBGk6W7gvhNNwQbksEHGkUUB
hiwGGpBamvtyWA2sITmlHaRaocE8sEyAN3Tmucc/szWJc60yv2Nq/g4r96a4qWv9ZIWg2M1Q/ycw
Tmw1sGhcgAmNGlMGPc0w6bpQJ0l2TtIxc46lp+MbBTJgMAvN/00JWTBxbwhu/caGN/xbTSCWSa0b
OHC4OXfPC+K9N7a51IPN0qsZos2R9JzFj9IDbf30to8tyCsnu7ntPhLvo0EVNFdfee7XnoYKScud
1m1vB9PtcJ/d4/lO3ZAo8ohf7WzQnV99F6KKlIU4NASfi9Tjqqv+s32RAQligKu75Vfb1fMgMXj1
Kmin4kQzHEk5Uv9v/jB0Jh9Avb1E47DWc5Z0aHPr0w4MmRAQzqkvW4HPYg41XlG2B0Seyzghfjj2
k0qKT1A9iwWGM5j5GilGp3um3akyukV9ATxB6shUeSIJq0PHJDSQpywQvHGditeI8ThoTOmxfNtf
dE/oaaS7Ln4+Cuf535T8aD3dpXd2NDX48VRSpF0S7H1sdusfPrO5U5fvSs5OPXQk8R/UJuP4gbUI
0DUgv3AotJI8AyR12WI0mKQB3OJHxJmvFyRQwdRFC0LPxOFqg/fLzQEv2nJMEcJczK8SmWC8rEmr
vDiNRbqCU4+ccOLesCCWodEZXdayMiFW7yPa4WJhN+7akWrX0lULqShJ/N8Qi+n1cMpROz7ovC5G
lCl2hg3gmBgJKgfIxDYCppwJO2IzdGsdiA2uXGgCvwaK2yzpiiJwNZ8HfamSKTryif1q+j8YYoUW
SKUr1uR3W+eJ7IPut1YzayCijyogP2fzB5WlSeWZfQNgFA9NTn7InK70VYmWenR26pKD6ElbYpSd
ZPeAqtKeChU2gCTJ01zDHOdC1uVFuUKwrDxeEJWVU4GHL9DxrjL2QAEyn8UogIyk1tcR695vxaWB
37P6jAPlVJwtTRFc2otECAoHuStcpSeoMg/FXIciusFsmIa2vJ4o9b9UJ3Irjx5+C6Bsn10d2SXc
rNOpQHDb1EXwKw7tn+w5fwZaMQ9KquPGBRaOd/tFOWwqxe75xN5ZqDEYlu4sOXzmZqjrQjHn9xMy
xwhU7rgo7k13BkRDy5ECKLMm402jkfjZIxhZ60jZQBLyRSoBbWMExzPa1UtMo222iH3pKeARhW9T
oafoBbQsV7tuzEnFY3OKobPQp5709VPV7oV+wBqMPHGOCLuxLSYU1rmU4AAoMNxPt1zrmAX4nfod
kRpTTEjp/hoecstr4y1NZ2IjcEDO+9X/Ratm2D+timOTzF/dCCec1tJxRR/wZqLWjkH1kDCRoRDG
1fA9y2ikKEcCCrBQvjB5kFpH3gbWZp6LAJ4rMKLT266VFjNXkCJW99Ju4XflbuCelpH8HQSSmjD5
3vzfXNr+xL6aWCQhKvGNRkWIsoihahkoSQbxvJb7E891gz+rWXwMHvEqC2l0B2op4DsAxQdVH3ht
Klu9tbH9Awo5mKa+P+a76tkgMo/rH0sJTqpDxJYYDiC3/UlH+KLmOwY5ZQlbvCpQVfAwVm4A2UBz
6oCxESqRqG8VbeQZMC0K6zLEKtqe8F4Id2PdKnjpGOnKqQ38fLgZq86d3nkLABu3vnf5qwDzi/9m
FOZlQklFqtKQ8qchpYSyHrcXP7woZAtXd7aqZWCtlAClFqcBOdbF3uK+ZnJiEpH6Lvlt/O09/GX8
oznCWS6R+jKD/oClf5anJCiwRBPdZyF4AoWuBW9+xtXiblLgG/fbpeNqo45I+DfhAiJcr0lTaoPM
NeGH8A6Gn68Ei8VVkDB/+Wd5LrweaP4uZ1Pnl21krpyu3QNZpz5vdTMd1hIi9xC/4XkaTeUN/old
AbW7Qm9uBuaKywmpsF+5oORu2DEqWA04MW09JvCEOeojMts4YiA+UVddeQCcClTI6hKstzuWBrAC
h0Oz7K6ig0MjewaVzdHAQ+Libbtiih4B875m8dT3slVtfnx4x9A4VJVxhQOdaL+vGm++jBb22m07
ded7w7mUFS7zDnsBlflmQc1G2XoWdEMu05ZajJvFr6Lp+agc0ie/Mf7V6JoOzitBm6jLU/AvS/3i
b6uZKMpLRRBOSOsgbPM+c+33eWJfJ+FTSAT/FUa1Cbx/DmZ2d1/w9gv3OaFFihT5Wu8bJakv3Hhr
q+dhVHMMZj8cPFLHBFhsrcehX+DM9eWel5uzLUauuM6++UzsTwGmKZjCEr1CWe4guQAV4zGfuJtf
n3giYyaDmfusgwt+XQiPdM2bzklsZacZUWZCHUBLypo7VwcWRtDILPalcRz8fXwBW/UjeZczGmcG
D69ZMffOq1AHb6SV0JpBPqLPIVd3ct59duIQTGDZovjeYg/ohDzs8ZwwXvGyG/iYqiaDFQJ4i1EV
LG5y20EOy2XN2Wgfd3654ShWNxleTydE8Lryge5R8+DEW4i/KMvcrW4XAmcR+t9hvFOIyW9Lvztp
mpt5SfqNfdtCb5RKcOZwd6Q+S48NkIIEFeZWozCFJCMyhuJkGdqfUs8DedpwFF6Y9rXeAFmUmKr1
+oSEGn7fMy+tfWJoXfxdT4FFsX1PcfHjkdhBP4aXQ728adptDAkqFSdRfYK3qP4k79D0UyX8pAfV
ofFByBxzFU8Mwdqt/Vo+Nv+6reE86x+YTcHadMnxS0CJF+TMKkSaBTj3KZluVhJ7YqkRV2znxx6E
P2rU73j57Z+fJe+a1cLRnazHrAOnpLqEmpSZSwIwWcWj77e2YVMjmuaU7VTI00pikaXRTPZEYW+A
iDaYbaR84eVGBM/IqbeTCTivFCFE++TMzh7cObwDjnywnO9OA6BXNdR2kc8c4X7qSqQeqfJDZG5/
Hpyb67RLDmZlxkjSrBE5rm/JsttOKBcoyAEahzWRVYYUQdSxeZWtx7LxvKexC9loYMi0p2y/zlWB
cwLC5Cfh5yzG1Pe2T/xED5unMorcMiK5rISKUx9kJx0Z88pdv92MDna0zDa655yOiMYTz1xUgUYk
x30tSOXhd0pqib6vySaAnL/mK/yJCA/Wva62WAFPhRZMRrNQAVSrcfldqSRCO/LSpoMwSaKNsu/T
+6cIhbAu57TX8V6UDHK9ehT1AhKzcGznJrCvnL2mBbTFUfznWp4JNTWgq9Z98jiv6iaEj7VudGoI
slBQjwXl/cw56jAgjDU66OxoegwG2Y7OfuI1hJgxjL1s2TYdGuZsSF8RZODtFo6azMGoKIIzorJy
ZORB/cKEWousiaMrGaoCpCzTn4nJ9mvcNgf+gvmxCxCe2T6C8U5L5CciDutkgsMmVuDixvPCnand
XEWV36WXA4sYI0O526Vr8ZGcwSi7pYfiK5+/WN8QB4riF4TU4QtsorHhYjX3yp0cERWGQwJZ1zWi
kJPxQKFnFKmduzJJWGrY+0e5szrRjUvoJ/otmZQVP89d6oDn6pRoZ1yedHx9OYwui+vAq35QI3GR
dimmN6mug4NJD8BxA0bXx4YYo4ifMpgGgaHwW4WSHESqABROU3EkC5QKxsru86zg5DnEOQNFOTdG
JdUUtdTpqj1mUY4M2vOsypwAbTBUoaMUohsm9Hus1Lq2ieQ4pzzDfF6TFO5AHsz5YSjXU/GVtHB1
VKCEEFPy5KlprMQjZUn/Fwww3wFQy9XgiZ7aJVKc1TxkJ5/Q1pF5GwP0gFIBisPyczDpoJJKvIde
y7kMP1XoxDwZpZn51mo3F9fLg8TakqvuPsLPtgtvys88W5puVeBGB8+BX7ECiKa/SfxUkn28+oYV
FM3DESEANWjDQUNm1t6YbOt5of6yjqcaiJJsCATIcGv/Z0VBYg3EVDgP/3ZhD2LhoZOCziDOxL9u
OeVQy9jviLWerWH8Wp/q3smFbTlaaEWite1kPzzS/d9dz6OqYOfYBJERaAY6VjL2uZ1eYHPe5UQ5
VkTxGu90930r8oCRdNO5TCilzVFV+9G1G5booXbaBGLr53szTYJCOON/i5wuby+Yp6SmLtQaGSpx
mBqHAlhRflQyB9fHhXbkQz18rDlELmZacDuCu9SAiG+qJSrMi4Xw1CFcgoo649hLryvtXTX4nmWT
w2z0LEEmPD6t5CYX2OO1b9OkJcha464n9w6nOVDnltjVHxQ/SJ8K24DGTARCT7UjGqSs5u8uCFLT
78pFDi28IN32+XcQg9LQP7lvKkzoeQSap3sbIbu8bsTNbqtcqkBrKlM84ErYMD8x97tYugvRUhrP
iwwTp3cG0Kztlw7EQX4LA6aNVffeWJHtNhHmFpMSNTsTxLi+Xn1Ir5J69+v7Xdn/JC5wu9e8GPkY
WA96935w7EhKqMMB7I66h8P25ceAcgtptorYr5bxURUuTpX7DKbB6uX+fUQafj+0rCnyAHybnNjb
31XU42Oqn1EUJJQM7JfqC+iM7YSdnq7FbqLZi5y1KYAOgKXbttlEP0unebpHqn0enHy2jpx20WAD
Trx3SBr2u/HdQ/2FWvbaSgJI1bF2cdJHVLwKzNVotjr+uObtegIXWiILawG9OqZ8VWHeHzTf/qOX
b9IVfRskVpC1Awt/GONBfA0di1TUB3rjrrkZEIfeVhhNv1v6PtPer5fL6Li13ZuDGXwtXtW7ei+A
wRReP4BrZ2MxuQZ2JBKr48rwdByA7sYkPqQq4xV9/rzZRyRBlyOeGuBMccIYAwWhwqlf3YnuMKT0
ER7yMRlaL1cKHWsoPx9uSTDdsi4g9gcDh2FUn8wkzYuIvkcp0iI4Lye22nKzOc/fkoS6acTYK9ln
hvYc595DeQTIepVdwLFNPXYfmS19Lcz+aZIK07OLjPHf4qOLcrwo+7Q3tE8MvpaV58g20ZGeXZRs
N9AZIgQRChIp9TAgUjrL67sVAj4kH7scxR1SzVWzQOu6vAtDx4w1pSxLJSN/lfZ9AiPlkcc8Qs8m
9OEndfYf2J95zkcrqUQpF34VZYAWVFc5IFo1siwIjKJQ3NvZo3QhZ2a7vA4ZOWaGnmVK9wTbQF6/
Xp1cyM17peURyIxii0qySu/cedcWyMy10EHx6rAJaQQOe9341vvCrj9TECs1Wi9E9XLMdpwVAlFi
X3hVMiOC1WXG92C9G33gPXOYwNkgiOtARVrnBFrtUgRMcEDGcAuse3gH/Q+fWuN1I3/Kh0L/Xrye
j9HIWpLzFNZHmUdVdovqIcb2p11GY7ItVzSfBxL65THvJF6o1jkiQXQt7KTB3WBixSzRGc9dNLCJ
k6hZusENZyTfASPA9ID/XWNUrvvoNI1qv/MfPtsSH6Jt2tGz/MPojll0WIbwDUT/uSvYzlbLDy+9
yQo9SlpySDi00kkIGRRAa3PGSRUpAS3P78tqwQbwGg/Uwt43thcH5U/LwOFcx4mX2YAwbTDzrAQb
MszERyv2qrqxzjMZJ6+UM1CGJuNp5j9JcI9DeEIiczcNUbf/0XX3EQn/KW6boRvsoMN8HMd3IX6L
u0lVgSVJgfVOVeN2wiNFly14gk4aR6B97mF84V+yaQ1JiA1IjveP1N5chxDd9Yeebz8no71gewJP
sWcxsK3UBJsLSiuaDy3OB4esmPxYyjv7OgygatNRhhXrbPoq/WLUMxag4KomjRv5UcvnhChSlYFm
RetcZmHfUdkSff0jOjvLriJHWT4wFXxMV4SkoKedf9ZBNj3B3qwDqXESQ6h1bTZTtMeV1evH79kB
0Msy+nA5uISUkj0xQWdZ/R3niJW1PaV67kzU8dHl/pI5Ck2MbAxij9/AEIcuV9Q0/S5e4ihTkQER
cwh7x2Mh5DvRuRNOMRiwwmKpcA9gJNBpx5Oy1WkoA60h/kIShxlu99U1di2GFahgYi2KQDOosawI
f2A8fxUVCVXrIN1B6xlM1Ia4dQo7OnJNUfh15095sLpf/KdQJzFTX7GiBDJqld119BBPTZoFkvwL
tgPVzn+Jxq5JeX1HOFzuQzVrv/YQYMQDXsYi9vea5V01VRIR6qoexrHwu9Xu8h4ku/lSyUMdPv+D
NB6un7KrXfMMPpwfaPAJ/uRxtOyI0BUJIyiKfMuwoB8hEpfyQk/mCnNd08csZvlu2D8sqQ+V6g7/
PhL7PSOXIXK1P8tBiwLyUMQf5U8hu+1rggUXhiuC/5mK1iinRpo6zrFgyGj2wBvZHrGs8r+6GsBN
Lilcp8W/XpEvl9+k/523dE3wn9N3Xz2Kukbcxus7bhN9DuYNTwUAcS77bq4cqJ3w+5405w+R5rB+
A2kGZZ80IBh9QgG+H0mNZVM9GBSDyW7xTkAryxCUsqpLEYjBewaGhhZW2z1GTUfPAcR1HHSFd+cm
d3vY5NW7sBwsAOB9HvcGUR2yPnJTa8M/e1nb+LAbvsm/uoxvsJl9LxEStsg7EWP0WSdSqMn33kGp
BM60xlAYCZoxal4nw2j6dCa4RuvxkX5X3T1bW/nIbpdzxc1DXJiQ4XIjcf0vKSFSZa6Zd1VVNK7T
7yxo4AIbfmycHp4o3YiAC1DP4cqJg9+r5LOjen1FSiQ0oDB0Dh+ZDBglguOCC7oUJteN0lV5tf5E
UwvBSrVKIJVSnH6+OC4m9ocY8dAzB4jZHmdWEEt5jL9q0QKkl7Go3/49QFZTSmDelb2rEODKAALC
P9PxAr6gXYm5JIjuClToh50VN+cZqzLIpD8wa7XNLZDyzZU5Q/Ew/azgPHS1MS0fiGWbQMt/M8En
ENntmda2XNOyGkfF1vtveE2KHIQRW/IJeWvPGHdFPuTW9bINB4wqAX8vxSHrWv2qMGJ0Na7zkK6P
C5Ricg7nHdFGuFcWzbLHTCdFstBqXKCLquRDf7DjZfeN+LUg+aFbU20bZkMgjtQupsA7HnXvp9En
hDOjMOYnDknr2JBNV6RXmwsZF0s73B/oBgzQGeDzNBLeZsTr0VLt/8pIOquIPGxtaIf7fj67syQ3
jD+BsjMJ5zrijE2ru2n/3TmJb5DNHtYb0LzMAI9RMutWBxUNmM0xtL2QIIYIH0kVuYgb6EWZRX0U
7seRT+gt3z1ptwMd8sspx709IVVfEvDBUbrDc4P8Mb54e+O7IBqZXpbCb78pRRudV6e2MFQ8XxmR
cSyY7R8yeHwLYbYbEkF2uVRnEBB9DQj5YSv9UunXmMBIwVp37ewoOU7PRG7fFeU85xyqzAMY/TXZ
b0MpPQxeG5+4pzQdK50hnJSqTXEWBEnp2iQKPA1DGoLti1L9oJQjQWpGgW1/w+1DkpREnAW1wSIN
stdTbMfU7Un+eERrIaKQynVXYW9V2J6sco0uWc71QV/USROenBWqOvgucY674d6Df6mRqQ/VKsKJ
Hi2ntjaWLOcnziaR6SR5NJafPmhm+JjINLjP6u/Jt/iktlteCaOqCY1XDAtgt//XI5bcbGq/SV84
rWYVqTE3+fOctM6At8fSxQ31+NrHhgrRiBKiwxu4ML5j3ZWzwhGJKsJnbj6a4NgSd98eMvwh/xRu
dMlLD7OmHWpF0GBvB0UCH7UIvO2mN+uJO6AwCcQQhDJhzx7N7neB8pW91GlL0lOTunzVJspkXhfz
BJujaAVR3j76IKcPuO2PZkPBdhFSAZUYq4U4bUwuwTAFZ7Q0lXfNi0g66MEk8hWN1SC8PQA59m8T
NLQXv995M5x2QkhlNqGiR6rO58v1HUdcqCCSGOwPl6Ff+9/OlJZvK0ZVTWX5N7QYGHgd3Uk6+suJ
96jzFFCm0SDGEeWXLik0T/gl/mvj3cgyDN2C0Qk3S76+IqpgYUZBi0GVLhIWw2E9mbf6ViYt6f+p
mVIYYPQWPXq3rAjiuVb9QwsA1sCLlmkWem7zrMEJMbqpyZExfMqx5todojyynjWcOyzoOUUTi6kR
x5b1B/VJlCmMrHAvVMaVod1WvqDkZ9mvfV3mUkQ0tVnNRG1iuxobTvbmhfBCBfZ7v2TADT9KTIIy
24SlB1tgRpp2C/qJ6Qb6jXIkc3h8Aa3lYs5lUKq1xowi1bQUfxGHEkGuc49JBVxqvcKe2b2+TWp1
rtom2Wpv01An2WDWwD3LwhOadWEmq33pN3Ww4+g+o5p/YCo4+E9hPEsJ3OQB+7RdAKvEzcJbtlPW
n33OW/M2/+eJ24bYqGzqK8JR7FMpxBKcwRyRWNsv/KPji7GzJ5WulG591N7r0VhgZ0psFKwI0oeI
x5R6p3u8D+rLOwtCJDI0SIbkciT6cuaPH4aG1OeCBGD7I8c8DW4BBvhqtBE3psfxELusNeqHz8Wi
d8KDPHG6XaOXj/d8CWKTxJzho0JE27+JXGiWeHcPAaU0kaIj0OB0lVAs67fYDGxN0oZdLUL5sDUZ
o79KiZP3ZO3mImXr7FwGe8ksQYBcdFznD4QASIc6yP9+eRnmNhqoJgSw20Q5XWMnG+Y7DmDr9JDK
maESdsfk0+kNM+2HzuD0ai7aUnm7VAUfEUtC9uTfqx1WYfckEIuKqLiqDZRciu2ptT9RTdJcDq6K
C4gBMu35YvxwV8ddYkJICjPKI3lzJ/dFZ/smtm+iAwz9xAhOrL+RhqdpUkw4SXaGN/FY4eZ1KXeb
gcWLxgX/zjhmrjpCQjYp18E9WtrkL+vcb4Y6qclqJsp/5UTYY9U3YL+PNNAvcYNxVdqdT43RpeEk
e7Mo908K+eFf8lBOpfEp7TlvyGPVkN5B0NlMgavd7NbN6llpB17fNikGfznTdT/84vYh8xEGUOao
zfYMMJEO2Epk75rjlpjk7QQ9oRN+h6HXFZ/+9gvtZ89e5UdyiD7GnLplBxam68TDkszTKSMRvv/q
vXMcLFoIcJGRXM5V1jsr+pJWbM0Kgy4V92pHYo+qPAOKzWHk2iQS0jx/Uxoa98aBEup196OH/9Xl
heGDed2kNvp+gLRIxjChC6VObux6lcbxHDbrZz2qAGo3zAeK9lVGpKorsomDuc8+BUZ5I/35gy5u
SGAm3YWSSuOBwZ9XcS1eFJZS2+7pRjrz34/LlHrqCdOs427XrE3l9qhWZf36UfwW+Qphoa2KNnUH
oGSKKuUuCs6tKyLX+5Yk3E2LT75Waz7olRP9M0mw/xc/MEOEuxiCvEZkHkvIwgLisdXSXs4vtxpo
wLCatsPIdaco+VGSw2a8oAjRwXJNEs6ArRgaAYcuuQAjfI3gfqjQrlMcaOb0wyvbNoPjFPX7lQ77
qxLqoZXgOZDCr2o8/XQkmAnNqKRqBcYT83Xi8TQ5Ye/+VLn4Su0io+Q5Hir6WQqRFUs3lmUnKUUi
nH+qVssAoEVwSssQ/sVZ3t9BInbzC4eDbT40r6T5cL8nvLPQJMkMFoGVPVNYJSNxz+YfB5WbUbzm
6Xt5QaNLOTZa4BgGEo1yaA084Iy0GUCaVfJcvty9sAzDALD01f7/HsG3PRtdkgeoNelxmS7tKS+j
zEJ3FifRrR7WvcZIJtOGhCWeN5UJQv8/dHzhFQSRi9ne+gO1Ha9KjobJ/+y49QQorRTDI4HKHKaQ
3N0u0c5CRhEdIxTaeG7Ejx/b6p2Ey3tsCaZyhXZJ/oPpht9DzBoO1vhI9F2Of7V7W9aHTt3z1MYw
28+AHWR2vpBtj7bmZdUiTmyYpO/3UVusWUzr5eAzn0OHaOWZktrU3okO+YI7pt6Ffs7nVyoJmeVb
UolVIwEMx+HNxfub+QXdCB7X89+0pU0gz0q1Yck1O8u/sqXIwm7buk5xs/T+Q9RfMfUkl9odE2c7
f8Ofa/kagpVx9GwDmHFSV/oe82eeEUZFh7EtvB4l8KVKJuDcWxLzKa41Dse12H5pxs3GNKUp3AD0
tLuxG3cvcR0buMOgqD68fUwC9h8HT1qkJIF4hSzWtJXaQgF+bbcVV3wNy4EpdyPHnuE80i8bPwgh
MPNUFSfInnw5pp/L/s+1jHTuwMfDQBmkVlvX40HBYClNm0J+gIsPOYbcRoiGVJfIL0r6dl5uqNrC
+hHqzTbt4aQoXRKFQu2qPewg02dzpMf8JstpBvb9S9hJUxTjtYLvvLKcxDOe9Xp5WaqGsekNUh5f
Nk+z2N6dH8joAEcGV1ffNn61/2BT23wjUAS2NRHWzSOguy7ggxe72sr60NL4PmN4lhANaSniRNwZ
2hG1zS4AGMQHFGX1ssP/clYt/8CPN9+4Psi4px0BQDRyVh/OGKer3ysl9GH0oI8ELUJ4Z73To8dU
X73oPeK0Nfy2RCjM0Vj1aGmlvOlHUyhdsJBE2U9h7S0kBFDvA128EV5QzyL0XjG5LQ5BYog+4iI1
aC1vj+LAzn7Vp8mnnd96pW36H5Jore8G5EJe2lAylKsrei1MARQXsNHcujKlK7NVLKeMgmjkRMpQ
LrI8sWVPl47YvJ72c6wU9Y//OfS9BNS73PfxDK5JEl0DQmA45GS/HcD6Y324FJc85d5LjVEXmsIp
sn3virfWa+87vJ8M0nQHJdqeONu0kCOlRRXIsk/726Hs2Y6BNgu6ptjleUaGcPnM/7oooXP0mRvu
RfcT2ZtPkCcDebqBDK2dNH1DCWm9RxmMo7WJQW4/dzFxvUEFJX7AeYTabMuVlwgHgxPGPW14UbvX
o005XPPwPT0Q3Pblun07INIz4/DqkFw/mHtBKV51XkFcmPifFd+D1sFOosDlosMbaoZPOqcsSo9x
tUpPtHlzc0MFwmhuQ/5WphEemWpf34/Ynt254JoWzaIv96t0YAuUsfCYPh63pzxRMQk0vWLcyQBj
Kltp/W3bond6tuHilkx/Q7SPLgU9Wt8hAuTHX2ztwBmkkZOPNrMLqv8fv3+ghQkc8T098Jss2rBn
hpHJviet4mDTbzfH7aHNKkeN+XrMlBQYSFcPdL0YbKfGFR51vtY+Ly9DPYok+9gDs3Ke3VkFrSjf
lIJH8Cy80mAXzMpZSVzxmbO6NVwCliwECeY9ywxGrFPzHCCEQSHiPZJQhvtWoGQY7++PF4By18LE
Arbj/TkBpv5wIWpWOvHB95xOiZhzjrEmaokF7nJq+8mpaCAjwTs3yH0NrBamA5EfgOwgstfernGU
ikE2+K2F16nlfkVAO10g9xEHQdpBZHvSfo05sCD/FEl3Lib9oV4UouclAUpLuEkkFRSJR8RZEo30
0hZsAbE65FsZs+dBRSHGQv6UIP+dVMOYWWf9sobfZuxnur+Ag8O4HHf+LxIvGPlFVYl0c5PByvyT
1bVbcdB/IvCFaPvHfPRhkXPqriek6WHGiD4/ynJEOl6ACMV0wXVdtSIgsuSiYxfz2ObUh160zrQw
CCMcktyOp7faoq86wY/j7n0dMG6skn4w94p+goCoLAGgiw33Gnbg94FLgfxbEd1MIpafYQJ1e/ud
ayZiMWt4W5/ankaD2WBY7+xeps0Fq8ysJR5EWCdLAS+ZEQTwaTF+p75U/9Zjfib41V0X7yc8iUfj
6VdBHuxVb3vvbL1V/0iZI3nhB25CCzMet5fsVosrKxKreVxcJdH6d60FN7diBqjUb5lEqEjwS7ec
3rrThnr0mX/3G2aAIwo8PQ5eVsK+d4QxtfXl5Otxwdpw+Lf6dCndWaNFZcPHJRp9aIp6ECv1TvkZ
kTnIXhXbN/X5QWmAxPscA6l/B7POsfezbIsX94Lo2cSVgHc4KAQk/L+n9vW2iFGmZ4Mh8K4U/Q93
/50SiUGSmyQNeIrntdyoCsLh9WAcQ/PFQdFmAzMVyDHdsy87Tf172DaSX8Fl+mUffOCh66XOA+/2
jGQ6Pcqk0WIR5dyGOjeISrE7ZajfRq1WAm4FEH3HykJuTENJkFGuZLT24RehR8aVfTPgt4O0CaRk
KfE5jPkBM/t6TJ2+i6hyl77ichSqiFkl96+y8k2IKSTaIIEhDIf+11thABS8z1UmIYLazozl0jVM
R2oCx+tU+B+6odikaUBywtxu+Z6D6l3su3bw6v5JmBruch9VJ0udA9ZHOEHjWc6F5vk7AFwUJU6U
fJKReCne5+I0esdz5ND1DzX5Tq+C5hldSyt+dxppO0Y2fX3sm0nZXYcSA9s+ewYaptAnMWji62ZJ
2+tY4IAFHZciLgWLE/wad7cARKVMJdiGa4We2NbL+d4Pd+I5bUSpfJKOMF2FRq4s26jnBXDLxGTY
RNZq1XTxlKSAtsFdWpTMASePk5q1g2+T8qsKh1P/hbWqMDrgWTrILQLbzQDjCYjcMahPqyhZVQuC
qMJPfg+kzpfjxKgal+HkF9tvWeKtWoPNezqHx2w8ABB2LIWzBGVVf2QqCRCG3GUxsQJ8MQxle8ZG
ePTNsBBkMPFJKzTpiorb6EFWCanJ8vTWT29GLO1QAO5RQkDEKBe1pODj0GD7fPdMnxt3IsAfjSZ2
uz4Zylm+3BK5ehjyFgsWnjbG/7GI4OhHGpIgESr+bJyGZ0ewvbDJmwwx0zZxGJ5J7jOuRRzblL7K
AZty3itpXrScFlXybCKQSthokHUHpg9Jn64rbaN553WvlvavL+iRxKGD0+9nNwO4RNvM4FL+IhFb
I5E3xDOKOUIolHvZjuQS4A4wqBlBQDxhfur7HUzofkM0cLhnI7PkcTP7ZNAF+Ox+hWnPKklKlMuQ
/wAr71NazGYkcfg03QkVrodSPXMewjsZ1LhvlmZLsjwjGxcUUZkI5EFgL1YKtYSM6hi0XvgGFMaV
lWSxCKvFC/uZM0YsjXaLkWoMJm/mW8XOLMGxfFS/cR/ElrAztrDJRu1nucMNjlzCOKn1O/y6lv0F
UzkbYZj8lhATAHxwvv1dyvGx9ojBvNt1kAyVNA3KKkxmx13hHlAeJ6VllBEuH03jzVX6zyeU5f7H
HulwofLRAjCIauP+cMVsvqTe96iWL3NU3UIZpg9hJbHkh03p6Fqnh7VOEYLz0jVmVvelOx1zKXkJ
XDLRWfqRJfZpXT/J5Jgbqv3hFqJqWO0I6gE6mbT9C7kLNBr1yUsK/doIP9EKRPv0TNFB14ThghsU
GF27Rn6TZw6wCjuG6NSKxOgTDhsnIvPMdXU6PUvS/USIwO6Ei6f8yC3iG3cVt4yw/EFRoy0FevlO
yB3U+qyGfQuCAFXKk8XsmWny16e5b4mHtR3n9zOF6CANn4sUbfUa9NAHq/znc/wvjadR9LvUwJRA
5ZyVv1TSnaP9yPHnNZmJeIp6BE/aRoJk8LQfSaiyhr7UbxaoiU5zXzyFjAvYBAlS7Yc2vxm+4mS3
o3c3KBvLdgI9Qf4w+lZx56+9FWMxpHlqlbmSESTZeKbPRqzy5V6qkaWycaERKwaGzKT3n6qWLQeX
wN9cNBMfWTHAQLL/RB3uQfO7LeiCfvkFy49MbUgKpvvaXXdkETAjiMyj1OzpnHhnvDYLsyj0UbmD
nqvYsApkuTBuaFObI0PYhbiMYJolmzDi3ZDEj9YZm53jlHBT5Sks5FN1kbe+NnOJYUPC+O3FGeQF
k76uQz5NFLp2MEuKwCj5Xc20KU01JN91u+aW6nOCBx1Tf0s6in0+niwkbO72/vBXv6Qt8zYEwoXd
s3ENTWmrhel+NhOf3nurIO+K/TPw1Sggj35Bg8ZtBuTSsktJoidGe534oDqjgDzYYj9iAhCkeMaf
QkPTZabP85uHBDFF1pta+gV1VTX4bv1yaS+rgXpekjwjhXmNp6Ii5RP9Zkp8qgMev0LVgO6eX8M6
EzykBOo4SNeoXglFVZL9p0Qx+ydOcaAQx50aumX97Na+P36dXfpORTT8QWss6OJB9o4ad1MG30KD
OUNQFUPOIX1mAIw6gKyA+/zZ5eHQsWSzBizI3gQHpBk7Eyw8immSI3c5ad3iUJNdKOkNGwGhJeSo
+PY0DjG5gB7AfSy5KoHRtwM2BFa1sW2iXqKpT8sEBQN84uogrI9TiPUEXBci55xOfIvv6QZg/Y2Q
ZzcAre2dRNdd9EMV6LWSsSAplzSmeSs/oy0HF9Y0rc8K2606FeBdlEblHDtOxsPamHtGY6z7xGAG
u5KlV92MlGNzvAdETjzzVky7J4X4d3hsjkYfaJl5/VvmGAumgM6S48kNuvskXdlEpIBoXQI5I3nT
T2S2nRjFa1w/HOHwn2AeaUEZKMVb9tAMzLuQoMvamRYIuX+wlwHgeSK57pBaAWaSDG3Rr/GXWAT2
Ed/Jhjf+FZbcaksuXq6LqYpqfns0Y3rON8KssbVwIwFK11pgVhFf0bV7dVy0K98iRbOpJbwBu6dZ
DPPKO0hjxSC54/jfWGV6SXlIbFHEQc6bEimV8d0rcPqBbT6vZ0cJ0G0mru3djrxdQsEC5U6XPlz6
Qhrgtf/3DcjmsFWiCd1l4e/APVvYEmg6keQGmL7LvmmLb01sOB190GNlE4XGqCdJ3snEFq0qzdnv
aH2C8mrPC6QvizW3etjIWmst4LzGXsalo1MPwYF6736OE8njJZnlpIJPqmxsaQUolxMWk83UGXsk
FM77Naec5SEygM0xSY08w4deSj9qtYX4/OQmv2hR7W+zFoBCao1hfzxkb9GX7O05Ahk5AoMqrCF+
8B3EBvufUpuRqIyAyT3YldHfTIK/colIb9Jv0R0+mxYgTNxBEsqecyaTNmLM1H/1XcXZQd6kd9Ye
0RooJqmUw6MoWMvqtd7gPAJgMrFPiUFILHSD6jq2JS9VmzrRKhtkV2IuJBoXYMtrXbUxI37MpcGx
RMlHM7Oa/kZpX17c/SI8exJnwkm7zThSa4+PvxrHcHdBNZBTYCqkO5s1IGQph//a8QCOtmF9KVjQ
7IC1BcYGa9YHsuZyRpmiFECw2rVgc8pthPpgiYCIpE8S2SpJh+3R4rpf2CH4W6flCWMzPJWHNsgk
9NPAlBITx8LwDijcCDfqAtEFG+blfEbnHzgEBbni99iKB319KOxZQKGuF5SuJzPAqJIpiO2uhIpy
+ETKXFc3dvdyaEaFY3hcbrpGLXPvxcrHw8Zrxj7lOETBM4ztIzHQIvm2OPlhC38j3ksbCTT0AN9U
rUvRY6RVaBL2R/QPjirY/vNaJofUw0TJoE0sQQcsHi46Vd8UNvk4t+djXChB2OKoQaGH3b3T+QVi
fmWUwkbUN+hdNM2Z5j6O2a3OCJOGaqCY5NNVICpYJFQ19dNOqcbxefd+RvbBGcDPRNsxCe3D8NCd
L64+n8enUafDD61iDSW1IAtOABktGx8TsXWr4yREByR/ANDmAbPuz3MMb8Wbmu/CMrs6wsh5kKXh
DgCHgPqnZqBJEdWwki4IbEtYj9AeQrvHITWludLALq0plGEEK7D7vbDNvDG7Guf6dn2Wdn/WIMLc
x+azEVljNLCt3mGxfIc/wx5V0gAcpw49ixWAYdLFLvAza0ObDgfxR+PPz+r4XLNZFTmHohtFfnZa
f/Qw5uqiqlhuQGpCHW9vcfWeY6Fjaf9w6aMcPRRuNkFas8LrraDv3zUf8MXkKt2S1CBEVmbkZ4S7
x5tEPD+O7k1bmhp5kknlG3P5x3SfjJ45rbAiu+A8tLZ5zs+jm8mnsZ8YaLP/mCdUwxMTfjSzc4Dq
e5zRNWCMHPRD+oc/AAKJoLwg1vGPRCfNMc5eEZnf/TtjAlm3NkT+emn5t7gHVRLUgLcyWrmCgoUs
djcfMLT24iaKDUi/k8KbzA6U9pSLYADUQEx7eySyVvrFsC7U3bAA9bXPetFPlnB1KTjv/6Mp7IP6
gA1ZUpzC2t7T63cUCzoxbfnZteVJwkSmSccasTunkE3Mxvrf6DYPEvg9nZS+yE29UdBWpxLbfWsS
Z6njKBfraSjG2AQWxS9Rz/yStkLfJSx9frPpCEMyVvB6RNWwzeSzwfD8ivqvWEot3cHPT/y2lqfg
CXIFvn6+IuAilbIlc23VS1lMuVu3tUUh/PnWH1vndfbDPF8xbYitNeJaSY1tLbBXwjkUoJZHWYDo
f94w8+QQVa54DaUq/y7I3GMLxvbCDPFy9pKPZQc4ptbXmbkuz0WUJbyM/WPJFwO6Sa90HWu342Hg
gcGy8jJ1qHY07Wzz1Gv+Ngpk2WHMTjSUSc884ovfPTgO9VHBSA85d+Kd+F8S9jgDIVeQ1b0RjtzF
ibSbYL6Cxm3YYdXOJUvK3SYcy65b111XIr0S2AAFb4ILQP+in/8QuQgbxAkWd/ZJ7ka7tpG5IWnz
W10eZXk9I4Spkc5fxiBg7LyWoV4Wo+0mdC/Ymu8nO7m0cXNseqXLEyrFZf6ym0r7QSPqI9VfkDRG
5kBHej60433HAU7rOVjwXv1wl9wimLhmWMY7gdPBq/G5z8W+B5g/cjSyT8hWffbG9CbiE78tfnOv
GorxeP8FrtwjVCbBgljjP/1uveYOCG3ruFriZLsg6kD3jbbLaBmFN/cNxc4LOAMWwocUwt/3DSOO
t2H3b25nFqkGNuKCyWo4ze5IN/P1DCKVKFi6Won+JAWG8bBuRFnKCQ+Xgap6r17Z8HHNiMvihV7U
NmZ9BN8JdrHLNf2KPfTCO/8XFfuippNpOmsjW2U6Ben5S9vT5s3qdEmaS0V9U0kkhT8iGDbqvdaL
2rjcopVSZkbVPXrpPp1PNjxxB3MrOcoELkmlPQvYsbYhwIMPoDiDB7V4YCV9Q4j2jzn7hCyBupNG
/nUseco1j7XRY3GBZuCkb/KDNolO0ox4tLeaNCLiGFZmIrmyi+ku2/N1YxG6mggZIsoGXwsuMKQK
w1k0EaZXKXdpqDavD4GMXwm3Os8wvpfmFf1RvBLcMNsrigfnJwyUv6z5xQyN5U59IesQKNLngDNJ
tqazPV+mJvEIazrYgx1JjGxC44ZyRRQFbZBmKnJ/A5FbpaazFXs7Tvn0QQIzgw32+t2Qx14KAg+W
rQWfL3gGnvBrVNlogU6KKn3riJ9qyEJ2VUpql+75QH5SHBR5M9iPh3Z7e7iOQvqjojMrpbgSICGx
2DwwlGhEzrfd+QazjNyD/xPRWL+Xcdtjoq/gGwx54vLIHb3JsSmb/NtnZulxVJNA/grq7gZUdcVX
OFl+FY67CPC2DNXwi8ltMPQzVuPmLAKBLLYe8xDsSHh2gyUMRYWUPGyL7DbHQ4nPblgj+9zreso+
S0xXdh94NXA5nfpqfxDqND7pfwVuhUr8l7v0NzGvor6bzDxyZ4HHNUgxmxJcreOzbmvF2UhrpJm1
+jRbK8rai4c+tXQssuWVsLdX3PDCSzRylqFiXtBVnfgr4L4k1cgZAp3r71ss4gb4YZ8Ckl4Osz2o
L2OU7UJ6TIztXK9QBuWkQqZk8Us1YLlWdg05/M0JezkF/J/dI0BBDRsaR1PF9cOe28B5NrstQsm8
KO0YepPa3wLPeujXZ80PctCdNecfcxYDAZV0EmCAZDZNSK4C6iZtLAYzFW57s3YTWVzto9TgAHxC
9bS5j4J7cVqNIivgzIRMCqARh+cDcZOUuOy6MQ11Yfe1MyAWYTmO6me4UwgwAItZkWQCXP8YxguY
1/+2dfIcPdMynbMn7++Y+gZmcMY/LoU2XmIQukPlXn1Zb80KIvhuMrOctEwHAAyMySmZlT3gX1va
/uvbEUqiQolswvWuEEQt+6iPuh/LwZ6FzL/3cBN24KZEfg1ezJgJJfmuPyLDtRzJ4zZpD2q4r41f
RYDaKmc6/Y8qEsSHbmETy5AJQUNb8feulNrQ4iVqeEfGP7vgXJ+8J3zoi58F08cKQfi+6lktw6Ux
bCbU+Nsg6GKNbyyY1CqnVgtlkZSWzDUtV1u6T6BZvvSW3a7BPguX1x4VXnNVvPLT5Wx5KU7rd1W4
dCLN8OVTUlcI6DPrJDo4BFOXmaihT7SiVQpBNE6kehVeqqf2xEq6B/CkOJYBZWtLEosE/cPR6Aa6
Sd1qr+mjFINQioRunzOqzXUEn4KfYYMB88J/gnUro1lZPOw2asfVKB3uBYOxs62LdE6DbPwBy+8O
lU8BkDzalwk7QIkdBVaVn2+hC0ZtLWeSr9WAqN79+8Wry+IYOZhPPJuVo45JgGzogvOzFx0yx2R3
rvlSkUY5iFCzZUw6E4+7ADe+LsaNYAm0/RcDPunl+lyEYeVB840ODjqJoGqn94NXvFwDbA5cnplb
GCXgo6XrR0ibNwYTbaLMv8Y6wC4Ib7Hegp5Uu26e9EJmZENzWmykN10HSdDw9s1g5M3OHsBFoaQb
ARZo7Z2OZxguN0RoVhaBjFXDN8MN0IWtrptGpp+OSzYtA4fiSAtTgeAPC5L9HteWeJShfo3RnQbl
s1NGEXgoGMwSuG2ERFpBqG1iOH91A+F2JzwJN0j0zydM7HG6+ikrGs2rM2e/iGXhNUzAQkQdUL7A
PdsS9ub1aajgtUHhZqOzYhCfoeTsxbp3txPktNwRTr7vXNo84An6AhXF4lnuG4i8LZgDzqCPLg9c
x9jqzQYBV2ryzC+KmwlOq2zf7FWIxlbm3fDAPo5M+NuykCB22KDrroa+5nfEXMhBoB5uefQJSFlz
kxUbJwaoDCFQdlA5egjVA8u3jIhMHlvR0XbZr8J35Bf+lEltm8/AQ7Vahcc78rTaqWAfB+92bnL+
AyWl2Arw/5s6O2/jtSY3ct3Tb84nxzqPK7POqFRwT1dksN/7cfxLlWbJDUOb+aXSp+l+GJveEFO7
kJ8lMOOG6CiiJVHUVD9nZvA322OsuraREqABEnSjK1WODYKWJSg2md5k8zD74IxANQth2VEdCUMd
f3iZglNctA75LhVqNB8uv/OW+iKvkUCAMGSmpxuGWklu2i1Yo3ALRyyMSUD9NLuESI7GBNsCJ914
UcRyDh1YaWMVnyiZasggtW2NZdIoDTSQdlrhh9RMq1Z/oToJFlJhjT6g7nYL08c5lHX5wrOdkarM
FrWYigyTtjpINxu9Ey/YRPb91r01z7mC0qMKn2hjl5uPDGsUpcqRTkzJHUB9IqzUt4P4wCuFK8E/
hN6gY2TsC1i16xl8bc3olGo6rfwGLa75HQg042EF7u6OXEkowSIgwgCMtidfblxBMDEZU98W00wI
oZR7+27pxmL55k3TmYrTFLtquGKC42noHWowWWOjNrR5lTEQawtOFx/wHGE4xYDhsHmvRDN3XnKR
j1J06sJeZeeRY444avl3BkFCiTqNAfmys1DHkSVmbV/j3keuqPR6ihnRd/AB109sKkEInhF9ukl5
uSAhuH4NebjYwIhSkWHSZJrIoG9nKgd19CrasbaPgic1Xy8NvZNNjV+Hxo6eSAjv0wtM8s1UPkxI
m8+QYSCo1JItKjdN/RqKqnUQ3x0PAiYgLUcMS042Dy3+K7lhPQ5sh5nwLN4X/vL3PpUt/RamrZ/h
HTN9TpbAj4KLMsYGREGG0e/KnC9GdnjU9h56guheEc9Q8FFXy8XHyKGIw8dIjKwUk348+LNbR7rk
/GWh03huV7++p+33x3qDLZ+6Y3V2vjCyLfZqH+LA92Q7Gxe6Hk0seZnxEgfPvF55GqMDSHUieDX+
AmAY1iHAaMYbhpJzRLmvzrYQ59QTwxjWbxokf+ED53Jmdw14uyHKMOg6K8MecRQcUspEsrSdqxkB
bRrEs/LJwY5PxpZ5b2BsfFaXVHKl+B7SzxToGT7CYCO+22vIi7l/hwRnxdZGVlym/F22Zv3pUt8f
KM0nukgDhmyC7x3e8PoW4cmQWAxKT/fH7j3sC2DlHGBtTxmFdsWckLbK2beCzqhjC52qLtcrI+MU
TXuVIE/4IOaMQ7BGIcebp1AYEKFPAHGb2WJUzJJWqQGKejjSO2As7ZLMz642m4FHR+YLD63sTR/N
3PMZhB4MAvWoh2T5XHzLEDvRzFXu8brfUfE0n3WlorZ1iODBp/AW+/o/6vx4wJon8CfeiDFYC1jO
F6g9Z9VmabzUttezsf0cyyI7f2AuJAKDuaNJ9ubkU63QsWydSicQ6k7sGLvVCW7PLud4ZS+nUuiU
09NJNDN4WL5d+wdlbODR7sLikEcWzaIx4MF/HyCObTCTbEmSJXNtPIYY6fcCSAQe0cuysEHJTjrH
PLrQsGNysHpWeZuEgUt1A+VPLaeZ0Wmdo0nHtje8T+Q+cbty1YKb712hmfiCOnylo/rVbsg8sHZB
RjV75ApJRP80abA0tNDdqzW6diCmXJNkvOZWmPTQy9kw4bMKKel619zFK0Hyj1WoMeyaYa2t80HI
sMPneplnNgSCi3wxrVYdf5SKs1XHooQMcWPfIcU7L99xhC9so2WFZS5Vf/dc6STnz0z+ItgAz/Wi
WB3FXbCiy2KBUJjwm8rphpG5ylS0iUaxn1qgtpJ3rcZ8PtRppfbTBOCb+QKMMSZmd52GZUB9Sw3c
31inhKlfOnxJLaQi6Tmk5jyBvnz4gz1+3b8ASeMj7vt03G5Hteu2PB4EgJTdh+FVSxw6nwb5RTaJ
xDgBYHY3OGi7AhhNidM2pt5x3Pg7ICoa/cUVzYv5JYy+6QKstxZ0p7z7fuhxeoNNJK3McCGaLbvS
RxLoCy7onM95lPf6bIk7XyahY8IJ3SyJJ5GNB0aOJ0u4CqMuzEBUjLY8mHoIUGaJ+qHBRok1BAw8
rLhz/BWegUF0zLAKL3sP+dE8zCC0HxZU+agu/sE4255XsRPzlNoOOCJbmtE1gqBzZky0D5YagqDX
CrRFfS3zxXcBHGnJQtGYKQETwqL4X0fLKnIgvIYDHFhQW6+qdvLFUbzp7VmNtR9virXuuo/fh1Aq
qfcAr2gFiav7YxruCfv43qb3SHuC270KxqXEdE1V7l2Au9kA7ooxzXnjBBeArlmIC93OS/QfOQ2T
pE90jSobwlkAkQUCwAmUcwk9myIoUkd0jcnEJxDlLllXnykMAlHXqNpYAGDN+m6PcKGT6c5mNRZp
IIGkpcdXzHuwqLUL0q2p03YoH1F8eMtiLmli24CeNBKZOIWqQST1RDTr0wz8cZQGVYYxHnfWC7aB
7NaM+y96/4pO6hB2apC1vQnBKVMFJvAmXA19Jf9t5WpGWeZGp0f5U8ibb8+q3USbm9DVxg3k9RGM
EzxyE/EorSpbCEKZzwrmkwdWMKdUwoVba/q9kA/3XF1x0NSsn33gcCeXbbNZwxwzHuhwu2H5TTn6
cG3qP8ofCXNmezVcoxbP1t+wb7fcnqnN5gnIlIpr9M7F+xwCvIGiCZJUk4z3xf7e8zZdlMTw48vf
naUwNBVQf5vbo9NESioSyJQCKbG1unmzZpvmjIVM/6Y2gRvNmvOtPT2UG5LNMxJsPHV8r5HlZw73
Xm9lrUSWAZ5+6bgsxaP8eYJ3187a/w5c+n/LFKg2iaifojZPK3NipT6nnZ+E7w6DWxhn6/unNxeP
4u9/GFzhfnb1dArcdV05dd6qbl8kktaElRLo6tMbp+oxFEhBcCv+W2wlwJY2KtsS2TcmR5tFLvzM
TpyTMWpsG4Va2OA11mGyyjdia+oEScHfVhyNiK6qLUkrBr//Xinu+6bAoV+mmUgG/OoKqZRc2bQc
BOdLRrwTOzQInRfnf/OesMw32eo9JlEiWA1RFLR+CvAsYu26+U2hT+aOyGvJPJbwl0oTC66j5/As
zZLVJUN9OMjhJkuDX23ucVzRQviqOxO0+VOuL5RiySrIqSvzkdxbMTm7EutEscPSJzHHdlNH8YLV
fo9nasriEGVTPEysitaudLUi2XNvPe8HarRBIbGp083pM9FEI90iCvwZIgwsMo1CTdcR4J0lMq6n
XcjY/cEO2TLWa3mIQnc8j63feVlxcKTrmvXPbobZg7RCDkB1jG+DvfQqyG+6ccvjOvJ6x0EIBPWo
boZNsVVrGkXZFqR6YzykhKPbAit3UDBJ45ldKM/JXh+dfTJe+5qG7STekgQV28I85gbSYczSifBF
aQXEiNw9R5YN3fbPAqJL1253JtvXcxrORLhawF7jz4Xiq6b5TURdzj2rpPt9az51zVsTj6B0qOZQ
gcQfg0CKQBftFbWMxQDMeWMNgdWEwh/4h6ZG9S8mqn3FX5Gul/lgJ1kuoiMkwyvrjRLxjix5WowJ
auGbsLnm2dAVT/mXQWSypfiMPV86LGfbSNn5Y66OrtqdJQHV38DNGp3KyhXzxG0FcjjqZf26RL0T
SYTvXk4UqgskNlYfPfACY7a286CXedoqzmcwKZ448Ss4nZQzw8mOgOKhTdBjNr7odaKQ22Ne8TCP
tat8UVo3ZtdFxhbV2rCKrv5bHTIhDdrDvCxJqzvZcc8eMUYfiBoGiLuvlZhug/TEfC2ZeCneKcjp
hDIerpzBSkA6yD8/caQ/zw+9/QXrtO3e5tMCgHKYxoiE0dhJ2wcTvYN5gaEIYtGllfkYaGQo4eBd
U2OTEnrqHxWkcgqcXxp0hS8UAm5CrZIeTFNgsbWGvlD5hSm8n/d6YxWZwSAiRiNC5dJvSKNgoyyH
iKeAn3uUvAhyA0iLlQDL9CI4UJg5UWeP0qQm+wkfIKnVnlURbdi25K/t9sVXxtUzYQXSAZ+sfUDx
1qsQadvq1lSgnQEMYzib6Z/qbVFLh6WNaE0S5EKSdOAPpxzEaaUsUpnbp/Nf9PhrP9Iibs/8OWzH
L5SdgNeQT5TxKPVReP/FvwjZbQN/3R7LgtfcekstdL6BHz2JtyS8N0Atoj7/x9Hix3XQibzZsd+B
W5TTXKYnKruVWkGLhNXdF/X6ScWdjaXWSzBWVtiDzf48uStedRHvkrQUw3am4bMUltmCvffSZwkx
iVf0uxSFu60+LlVdOucVnKEFAbtdVSafNwSKn/9V4A3kQ1f3SXY9chGlvalgJEqYkVWmsUCmrC/k
QSXhh0s+YND0GHHrZ2mGU++FF82b3ZT0gsNqGs2G4QPy11B8RtJZeiRiJR2pQoCw0TXcnpaLwpVe
I+me/hM73uzpUw44x1NaQ7yiRhaAjrRNi41IyLz1OA9yOR6vnsWSwjwo4Abxr813hT3bgXVdoyYD
IrT6I/V/mU7Wx4LpLiZg7ZXgwguUmJ04hU5FWR20HBHPYFIJb4AamoXtOWPu2t7BSqRtT3OuTP5Y
yeF8uUebCNEBC2J+fjp0WbRbdoEgmzk/rHGP1V6OXv3vpNpOXW9LeDTlXjXgZKjKQHdOLt6ZxJ+u
jVVBq9kosb9yRDLEl6HFOpUMxdnXGcegsYkiM7X/Jlyi6oqvQg5CrPnp/ggnVXKtzeec+Zjh+3TM
lQr3KjMSpJspMKfcNUuDUiHXYOlKB6fPL9POeeqWsnh72a5ssuzXkiCT5RYQur9RAAhpYrfKZ3AI
ZCXTM6Dv7kIisu7Vjr278I1gUX9id2kUY+dTEvDZYrWFttCs6HRThddhacWVcx7jhIg5ir6mbrS8
K24dncqkBsQQDuLHg/1Mm3Y5Tg8Cp5d0rYNAjIB5dx+nwInDRJRUy/qzDC67kSGgkzfU9v9mWNP9
gj6DIxmUoOwCoAktK8SQSzqqI49YX7lNaSnpDp3C3l+ejkhyETWYo/OuWe4gj4ZHeee73nqI33oh
qDFN33q+0cadP458pnxU6suZb0Wsw412uyh4U+9NdeBP7NeQtAuBlgbPP34Wo0eyBNgDj8F5qrJG
9KSu1lovvi+Ez/UWuximFenEsnX4roxCKZ9Uaz3vJ2aLDjFLEtbooXfChc7l7Ge9D1wx0pSKykPM
MVEdnUtiygoblgxhhQJOpqte0DtQ+2OSUaHmO/6GvzuhqusaFUcsZHHt7yG4dll2EbwAC7YLiFIH
b4vX2JBxqfk0fA/3MNScMPIk5UZ7R73Xa4mVei4SYiUe2Qc4nE6uwCTIDgMWRO3pzNIa+Es7j3Zv
LlpUWTVsgz92ZBQsuwv5NGsXqeLtKTG4DrNygXGYXxouW0RK4D8nGAjm4VWnUH/a8RwdOhn0CWNp
/37/98He7vJxIqg0Tn7A5VQg6lQ6gyEejDZW94EqaDkMP5O5FVJpBUg2/K5KAcGP3PHxETolnMQz
9f9766iDNUZN85ugBeENU0RLSn/xlq8xB8Xuo8RmwQk0TbDUlY6LnoaaU25f9VOU57NIRFyrWqa2
J1soMKXmC4W3mSFW8rPNKbKLK59OiZ87j9lkGTNsldWdN3FId4/IlURKdF46JfN7Tckl+Dj0sk3/
w++t+iOUDa2n68X2hhyC5EYpsTTuXnCa2alz4Pft3qf9R8NNWaI+zxuyJVfoWrNL8YaOVc5QAJFR
7CShkFRt5duAzuZHxjEDVJ10eYyY6nKeTLquNlMQj5SCD80ny4wv5yom+DCWl25AA+7psWyh8eGW
Y0jm+wXLPHm9vYMWZ4smE2YVsTN5WZRBNMHocoNx5GsPc8UHVCFOuUAh5nvpiRSH1CJwgLbis3yr
h5yZBeVpHTgwVrESuVm7+Wz6RayKEGr3VOXXZpiuMmjxmhbE9tqkyfiDfJefsfxx56CAQbmvde95
JHkV+l8YvQGPqDN5q7Yj5KAk8CWoKk8hS/vPsGVEZKeKWDxagYbF6PVfoaYKMqQC+fxPA37a3JXK
U6FNm4mfrn++SyZdrXjVVc6QQTkQzx7qXt6w0OxF5i9E0Nsh06JQ+93jPbFTNRVAodjttCTYgAaZ
52gzCi7FzVwV7irYhZyJNYtHyzvSrE0njDVG4ICQXk/8T5D4Dsh6wKbEdarFuac9ALtLO86yRnt3
qmEJiZJDPZPG3ooEieLKMqH/GsHgCz4CQs4/t0sPPtZqKSySeY73Zk9CgBlGbYn81B2sHPlBR4Tt
kdBRKgMDyBcDPdqTm7UPNJ6f1RdFLt2xlFpQQPNQauJJTWUbEJsyWv/KxUu0TNsEZNha/RABPWLn
tR82RlXwXlJuipb8XCb7
`protect end_protected
