-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PZt0+IBchYTbBTbXO7H3Gb7IYbwmBc4qhSARq7hlkTfJ9cQ7Qe1z33hcjyt2qMpswih/rM4P5hpz
Gf7FUbux+f6/7j6s0qrusu+WaX01HjR+zbT9rzl5XsjbY7Yl+TOXlm87mCByKgfspz90mJGi6kl3
khPziZ/lQNYJWvOHc8A4BOxfW/PBl5GBpTElqqR+5X8E58aOgb6U4XJF3qorPlwsAmHiiPW5oOmj
j0xE7sy3ThMOtuPUWublzFk+kyY2ZPI9UzqrqvIpo6zYnq4IztysJrDZAztA/xHeEz6GCpBFsjyr
jSIO35NLO7YuLh5vlaN4464KlV2EwenjkuDq9A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35744)
`protect data_block
ES8FQeiC4GoEATGSheiXvsMYSH2za+Rxd/p/Z7r2a3A9WHB46eMcszlIjNttLWDAOyxEBP0gjYSW
iFdibUZjJIAbeclADuLg5+f0YjnQE4mxTNg6Gfnzcg0vKB5J+1oMiyq8nVqpYvy0RYOqvh9Ul2HF
IgUN4y0KdrYQiJ4I1EDESlOY1gFGj6gA9MuqcwxJ/04ut4l3lkZsduuPhIJDRmgHzVPWuRREziuZ
NEOvdfOUHqtmYf9N4k4de+TL5sTCZGSUpsrjHVstucYAGSFwj1NutuWCLJOzIAKiUqldFH0QQr3h
0pB10fqCqQ05ZjIYs78rIoXEV2sn2jImbKdcmeTOWw3dUmOb+MpO/Y9FJhGCDbZ1zDh/t3I4UwGr
VlRAUXhc/sfON9iV0UozRuDIEtyxD1WtQd4D8a5Tk/JGPNN6ECFzb4FqMSrPNLss99neDeu2F6TS
koF3Mgd0LCnMD47zqWqz5qjUC0Oiuz16kTNGnrIMIwZ8MjnRng4fdeSYZqULzuzNKBawa4k3wZBu
Nw8z75SuvDy6MjoNWCjnBeJw5Ygesw7dfiTRaPtWthwI7Kke/DRe+zlJ404Ucli/VaQiKpnDhF2X
UVpK3RB+n7Dt29uJxRQ7TW5KzB4XQaxNKiKUuelp6rXQzqobzTVLD3qthXl12rzskbDDDs0jbetW
txpaFdx41rzLOV7N9e+HUg32Olqg3j6kfsC/XbmbM9CayYtFQ2XJLtUwnaavW2e4WPukr0HlKCSz
rB35CXYeWJ6Wfar8b3hqPdlzvZDVD/u0xUf6bE55wDAvC5yQKLhwfgNrg6ZsqIeptp3E34NxpH5x
KZtqMZBN7VWAs5zrTzutB7FYBIVYu9vSLgyXtQSMfFXWGknvy0yntg7WtvK0Nh49ReB+gYq3/uYT
bu6lSQles4zISk7PbSQKIYUEveBbfienoS4Y0TbCuZX+vTgRVaOCowo2YpUSbqBcZQJSdUtuk3TQ
i2dN0+NgyMDBCpkCjqEj46uy/htGJaJrYRjX95L32xb9D+wOs5m70lAxg2icvh1+qNX5D9Lv6EBE
Ebn/EP/3ixD2FZYC9eFzmvj0PjUQofYwzj+LmZio185BR3OvSWl/LrCVFb4BPaCHOOznBHFkMsMv
BG1B9epFdCTfASgcHqOkkqRD15lZdFe054xdWB4rfDI/oJSHGI601kCMiHKBlOdabG0a5F4dzqMp
Mv/KxzhEa4lXZGFA5Qc+P7o+uDsf4wlI3OibC4G4nJO7UveGELrr/jg4T+GcR3lUUbCtLeDvcIST
J3mTCr5WDTtJ6di3gqP2pJhyo7mz0Pi4ri7hgGfrvzyBtp2wOV9nUE+dMZb8RnYYOh6NPg+fA47r
P0Ggf80JBwizyL0A47nfM1cqPYXwXtLiomnZTos3vFN5P4gisG1C4l2/EMSI07cC+Mlw5Zs+Vss0
LdJDVu//VoXELY8z7p9kJP4rGFWTATkBOb25t48Nuv3SQBBz+suss7UyjEz5Z0d2HYs9itxkpHt7
Y1ucolpKsbTBd0gokX2ioKtMoJtTPauzFyd9SBc0b4AtxX0sWgc+nWv++CwjnWmodfxTerjyKudN
1KKv7UuyXC6Ihjk1r/qeTHatbBY0Z9OrXWx63P/Oxf9JjDqTbUMkmKLmMaV6M3HspAXt5gneSyvA
fSrNKx0r5thzfxcuA1HLJLaWU+z2SwpW/tdS20fiJ/kCmW9X9RYWHqXy+KYIM2nK/twsZ8QXZi1U
0bQ8mpr/jUyQxLH6UD77VlcY517pkJEwY+OyZ/zbaK+k+VmEKxJuZh5WlC6JUNcVRYJCVCx1Mw61
0O9geaAIkP/mYLrb8+Jdfbsn4LEmCQ/+AdgBqdGV+QNes3N1O5XpgR/fViHWCgZfDYuFA16SQL8C
M1UCtamN3M0VuJv4lyvlP5+ND6OORS/LtEbufZAp0VRsoh4eyUzKEhF3OPDytUKm86ubDIxwhCuu
/XBkeB5KgkWvvHdko8CHdPwA6s0iZ4ZQwNgVl+5ksPejucJFSDmHMoqCxc2p6ncDKmH57y2lZOtW
c+0cYiZIZFyE2gw5j0oZ349pp1u1jJycSMFEhAvtWbDa7KIEbjjAObXJGSILJqFewy6hhvE3/zV+
Nb8yt963LxJJADdIzQaxP5ICOWkLC7xn+Qe/CFBsT8iCLYfcQxUTqd1EiEQ4cWxReBu+nAoS7eXa
0zhp+dKVLYF8chj7ZdOr5Xa6gyT2vXUgTNw5UXFoWaYXPeTGPImmNTKYOFAhNGHhUGwg+vmPSPn7
cmKf/W14r7PaOjwn+w+Uc8WPY1PY7QkqZEIH/LAj69my2qV6f3FktQBb+9nqRIFrSZ3fJ0Xy3IcS
I+KH9W5NuXHBKsXa9QB41kD6LHMKeb4BA15UhwLvKav1Gc6WzFmq+XLv4WXTafsIFhlvL02WMwpL
OB7snls6Ix4j0AHXLWzUgZll4PRk2BDw6+QIIWD9o2J4LedxMU9dJzDp3dJDrOa3ueldaqkbxbSP
adP6wFNkyUQppCO9ESx4NZbkqNy/SGtFvojX9H/VHLn/3nKioWySQ2h6kSgE4/1K4zYb0/lUMpQR
LUnI5dtoFXyT2HpTCJrykczizIf09hIQBbrpv0Qqbomv1MnHFH2uhV990Esv/Aja1Cgu5zWsK9jX
gjul1IFZyHhL+ru2svaX7EnLMupR3ct9MWRs/Mc3/NGs706bkw98aH7t6Z8q/ACxLv6C/yLfMAzf
gAoq+VXjOzOg1dgVsje3pEhw1nPXmm94YDaK324b/18nsr06ghYb+bjaW2doz+N2bEtDKzKCV2JV
k4Rgg8fsJHhK5369Bre2W/kCyMU/jPOMZcBAmUFN78BsC3hHEuxbxWAEiey26oq24BQPpQDYtm7J
SUHZrRmDmKXkkd2AFn6bNryA4T94CmCrymdCsnGFuNKEmWmMzW5/Qhb1WYZoaov6Jhl7mLfwwgJ/
Yv6eR5gejzGfRj5oSYRFmtZ8D2Z51XqI+FhA3VUIb+Gc4HtgJtL1srA8qOx7jAR3MlBh0Zt5gxCr
UX+TncTYM1ayTsUlhcNIQvBE2RzA/q84JxuooW77PUyIwoB59RzVOq9qCkik+tthAHnhntKObOeD
FUe2ATC+N57nXJYtDjEqEiM13vjgr8+Uc+sAl/nKV9W6a/qwzo3yw9csrC61JCwS2/DVbDf0A3QS
DbjRetFlo1cAqltkMCWprVaKVjpVwGX3rS0boTjNuXhmHyiDBa6iX6LbFl/vEcG0Owb05u42VWiV
Ticn7Vl88M5kmO/ggOA/StsaiOg8amUoRHwERPe7rrpQh02v9NBlbFB/7ZAV3/4ahHW6+OfPcvF/
0MX6oV8l3aAf58Ij61m8Rph/l0GObhluO3EzG9MFUeDLDNFvplxiJEB20OsMD05xZ+83/90OoHbw
yJECOgHsiukSL4uqq3T5+r5ODy+4//BxrE57Xl3iCPjKqvJofgpwajil7M0wiI20u5kgxNqDACYo
30jCfClWAakEBxm6uJ9MR4D/mZ0rNhFo1ToZ4pFniKpbfN4I5d0y3U1hqPB3t1FBhEYIBJjywmpi
aGJsiJ/ezFRX4cpHf5xPgQltyZRRjHIK74vGIpvEkd1ObT7P9IVITCy7848H+h765hbXyaRrpUnc
vKLnGEGJoD3oSDMoH7jHo5WCSAsqz/JrcXYC59njkpbpXUVpA0/NHTmrvL4YQNBMFobSv6YTNpuy
tzCNFX/B6prPyu5QLhm5Fc7Q8jPkKZEWlaJnHiZooLKthlAjuFaI45BRhPnnby77zQ1tGKUDi18S
P45ILZf7mECElNsy7zapWlExqg1jDZIMxpwZ9I1AvLH79eAPHueC9Jek2+GMwfjn48KGqQdwyzZO
CM0XuoJl+nAKr6lPagMmtCmMPPCLhE0WePCP/PMWVjtad60dyqZ8zDu5FczSY3YGyoXa0qJgY9yo
VW6WbhvCgyJQnqTdiMggkmMUE7XG5rac1we7PFgvgBVUVD4YmLZNj/8aPXtbmIEthE6qAWnR8Hq2
8xCmFOnaGSoNkJOrESblFpod9XnQRenxDjJWUtjTfQYD7BO/dmRzyV9EuNwjh0Ia3lXdeg7z1uQQ
RGo8dcLhkt2cgwt0Vhbsh+b+CTzxKWaMt1OmXVhhfXDvCl0Ypg9meKUxJCRv/dZqnUyg4toIgOv8
C8mOsZmlZp0IV3CD6hAWeGowoRGiAc54LdcgDBZtKhdSxI0GLLzLUuFZveCr4UuiAJANV93g4iNZ
syAiXtbrlJ5NTYhJxpk71UjnPVmEBXMXOO1hVqHSCRtbsvMF3yzyfPYGBQVutS3395QKKEd6eq59
IXk24WGtDXeCtx2HGyoeqon9eP1sLcgRq6wifeC+SHsIfzeKAn0PhEoJa9E/l+fF5NQSqEdYoRA1
J8oYHq1HxBKa3bDozkZlRhgSl/vxUm11+YiqTmaBA2hzl0XrjhEuPNGwIyr5pfUjZvYTtOmzx/v2
odXbgS3fbadfv4dYEO8EW7J+yxmWn/OIamBZ+Hsa5S1+ZsP+d+p06l3qQBGLFHL03cON3jaEM9Ot
6VxifL3zRxCkEhbt7dZWU5DDaP1ZEMtSJ5cfLhLNzyHO70MHdtawZw+HVmcpbFH1a4AzK8lYVrzX
PygbeQ8MThYlDj2GNmxpELnLpyE9jGYsDZP28sdVDyJeKCdR0TUCGR9rhQPfwtOfAqm7kPu4WHKo
e/WdPVHBmZtWgevnKJEMxosqVbsnv8yPPCH2d6zewvspFKk6nw00qADlNeSDcC2ry99h8dnY9c//
WZju1aCTuOFtMQftQHJ2aW2Y9CJCVZZJKd4A8nwTn9uy5ONxdTegR2qLXk0jwbOU8DTlTe6yYXc2
j8dAuhAhtxd7Bap7bCZSGDDcsM2TDcJQ8XzSVqlIPGK+VqwJU5PLWtvKP3ZtcsLDzWuH1s8m5c5D
WD1NX1bDev99yoQp8E5Je1NkucCFaRhQHiTuvVdKdO2jGAZKuHlZzQR/xNxrbCIM8S2nFey+RI3Z
PihvUE2UhN8yF+zonWwbSZzGmuyKdoB6k5qEcGi6oEaRqZEm5dl74Wm1ooJmsxvjPXGqikVTD2ex
7OmsO3ktdkQkvQU19s98Srah4O0KMuWD1mhRQsie3c8MqnIX1nCuCTnY9fxofPDcN4pWH7DeqEVR
CL8miOCcoNShqo7Uf6/M3N8R+d2T6M/1A+duDd6khEnds83SLJPkMf94M1JWVN/liGnWDUk7vTX7
Yr6MKXH6f9oRr4H3NO0DoQam1JecZBA3i6B9N6oHGy+8z+oQ0RAx2UkWxeWtrOj8A/RRt3/BrhQl
3LeT9QdMfAKBFRB51c5VafTKakkRLAqZxmPOxYSBUvuhH8x8kDoVyghQn3EEzOzHfeewRi70RK9Z
YUIeeLUPZ8G6ZMg/Bi5MIX0jdgnbIbjObSxYjjYB5wWA4PPQVdDON7j8tHTx1butEMF6tmNnJvoZ
lUz44/WfsTwlxQ1QBTbzhNk6JNVzL98KQAL+Dq0+thvKTPz/GGYBsJhNnySDMfG0iIqKclIJB5Ip
jV8mGrxLEn1ej9CFKY9Ewm9oSGCQBgunOaillFqcGKtxP//QH218bJvh3ZR/RFo+wrBOeDl7HbhU
hoOyED/QJp2kf6tlrHUjWIy5Be2ooA9YuJ1MQDRjOvVmXKRDRWAMfHbmRZUfHrSr+rtI94WqVrJV
z+vKu8LFmU4Z4FK+MGZ9G8VSPrmtYt0i0gmU46Of+OLhUqKHOAJvHkSi/aJu3UmUZAsMA64ZewUK
t45U3q4KzhW633IV05oxdVmveS7zB8b33lMcbhyl8B74ifGepi7o6l5c2e2BkR+rjb/XHr/NhGrM
dWLLlglgEBIRFDMCyB9MIXijy+2wW+3CMiuglfPZBLvqnw3yZwDElQa0T8jHvtl9V8mbeLU5BNHa
Oi/JTl7O68SnbfjGejZesmtC1HHzslDi12wywWnJnVMGnnYvtzvELXrXoOQpTfChunXddeJCC1Ds
oOTN4WGXcPV8FIg9CfL2G9iFLbCl7WGQO56505lEK5h6XliCa9jnq+3ro5sOFPtBNB0FJt6frpa2
/3C6sKyvgVWWMmUdNcdGYwQMAbjHu5Cab2p6K60s6HcrxXmBikPAsISHjDQJfqC3wAGGuH/MPwkt
Qk5hGSJGURkl/8Fl9hpcaWAuxAmuhQFQO8oZn8C3SjJzV6UgIlZ2B5L43zzOSwTyiDy+uYEdhppB
m7QeBf1DBi7bDrUJX1NeMeeyXGXw008Y0iZurXomMFB/d540gNHBDmoCAZ3W/WqfGuWyX7SxOgQt
VJDujHqyEoP/2YhM89flG54GoPPmxDKvo7zLj9/rsEbY6Gz8ZOzBjXCDhZmaKjtJql5gEkx1uQrY
27TK4FFAV1552UCxkRVCoJEV7VNGggWaehqVgVK+FlLWHfcO0wqj5q6nI3cG9THniQUK3uDfD7Ph
Rlhm3MYCSEiqpwSWlHe/8MhWQuHBEI7V+81xSg30tmFwhKlgJ9olvXhkReu2gTmiT8OuDc1wub7m
XZd44N+fmE+ueXfhZpN5cdyam9w+4DARcTV1EpO8yizlc4/WR2gvpVZ/9W1Mr7Uuaric48r9DQwX
JJBV3kRPMtZJdpvgw42BARqVXGxdhH8kMlrXdjqtCpeehPch5Zzk4mQCuBJZ0ti6pGgYvBtsGeOe
4cM/hZa5MIRhT2cYiuBYOc4q3soYGeoXRuyUoramF+avklU1Uno6mUSpSPS3cs8ClwGG1dkgBHlp
yKhvODiU3j/0FYADiwEWa4hw7piUT91lLbxtiGa1hTsyFV68q7jwNIUP5EgamPctnUe2h333E1qH
P1Z67aoLWvyTlVzWLM6C6ZcHJg/fHGhZFDMf4tpFAyCF8Jway8h8XYagpfsQRv72nTZTVUy5v6Sm
axir23wECA/N194fM+jsQVxysnce+dKZU23K57X3OlShF2htUS/ZGhlIrNkKA7L32im8MVJcgdWv
F9g/qVuMcw/m92kvkjAVPQUc0yu6hO4fdqlFQum2YMJWMzWgpy5Lu3SWGfpAKMNNmFqWRht8SIWF
YjmwavQp+fvkPT1ary/9W0usFJ0jzyRBaTHdl2qsoM0qWglFQaFdrya/5GrUhhv2v8O3OP9M/zuo
r91oyqEIM5l/fX/fi1D0i5pA2zDTr13MOmMnqFld+tbptmeVtQZjfK1DiYsW/5PacEz5+nMk8mJM
MQvhvmxcfKkJnPjVu8jf2rqlr6Z9OdYJcusk7MAdCYIakq3amYd0lIGHGRA9NZPYanyrxOgnX+Mv
ecilxX7mid97q23faR8gjqOK2C7M/XjQjN/9v1BpkXtI+dJ20DtDmfWwJtah7JIzbSAbQ0QBTZha
kQ/JmIcdCT3b/gUlAnWEflB6qBmpj8IBBM2bWjSa1WXfbVBYTqzleEruW5GCaeBUaZbftmLfbwVJ
wNwyLCXBy/5LZojfC55stXtKwdUkFwRONsGNpThI9+1MKMdjGrGCEJGmywqSQtdImVN5Bozv4a8g
Em2jSlfeu44+cGUqWpxB4eul0Cce28OZVDXbudhyqjTJakTtvH1/0K83EA4owjV8UArqeIE+X3zQ
pL4zYTbkAPj+/d11zu8L+qeodSP5bIFuh7TxAKBGlsjUYapifwTVvHetwGdCtaCKnAwvaeGBAuS+
PAE0Ys/Qgj2xjwlXtRic8M1X9CuVShU4nI5S4Bs8fAKmS/0+vjoWA/NDzfy8WMZZMA+smCO4wQpy
XBeju/0V2X4hH3qcGom614Y71Hu/dUmAQ8xe/Pu7NRSPk39SPCyh0s/F3zOtrE7qR2qHnD9vPe4k
sHVP2s9OVb0mhnYDJC1qOxcsQbebpJYXYvUmWAL3TW8ga8uvO/WeXzRlC9Uc44Y92Xcm7JUs4a/Q
MWXnuCIRg0WEb8XNLhm32gEICnP3pjqYE7HgZ6hCWpy6XW+/oXikcHkQXe5MDY3a8v4tCEif8gNE
wbjV/1sN2D4nAQeOiRV94yFxecNqaDno0MJY/UvGrUyc3TWSMMYsOLGRKW8nVQRjON8x7TDXSCV4
bqef7+eUi91J+BgMCj4pRp3ySYMEWbWXb3W6jwkFcbT8RPzS2uQepCaQewC6DFrfOIAin1M/o0Ae
LVPnHni6D0Nv/Z/62G8OgxN0ZU6AiQF5OMXRvj2B5IzdYgbI5h9/L21W2P0PLPoktGOyTUxQdps+
+FksNwzYcoYztUJ4ZRB2pUV99XN6Z+mY5L4XDxIilVzJ1lFJQv/5gTvCklSqyfX/AEGrdrfp4GZW
5jXdFlrV6n0byzW39DRI6nVOn1MGnyx9R56FNZgxe5HwvfpgFlKxZvgpev0ArPfaLN+ZDKXvakRR
ZSf775mB8EK/vgd/FG/2Vgnwmf3zeITXx9WxxllCHgzAKI17wowDL8UmFiuGYVZmkxs9JH1K5395
/D1HAgVxpmWIoDMTU6gKK4/TkDyekjvhyiYlAcmgsgSM0stDLmTwxss2b6WPFi43ZH/IRhffK7Fh
r1Hwhb7kg2MSxsUJSDf8uVFlQ08/COYRtCJt+KbQCNIBXz2eskYxQHT1CdbTeQD9LVL7aY4I3UpH
Z3CYCY+OYf1VxJQv3t6ZaNH3qwvtxST9F1ofdejbrXOMMOQNI4xbQlXhu8ylFjIdfWTprCepPtZt
7GPR2/Xcjon5NZTfnyyP1hQTTu+F8+qwlHrW+YsrRBE7SlGznOBQs4OiH0AIM/gQYGR0o01+W3vR
0z2QaYGIk+ww9WwFz/1FpO8evbTIpd0svZBRh/uWiObdKu7aJ91Fugd9JO/ulmnUq7U+h81tcvr7
7l70sDcbzUmyST88Ka6QSCS5H+9mnTKGjo6MIdbMlpQNScPawXFCHCLfYK9EBUeODEyD62cAmwQ/
LRkLD4JR7oDogE+g7PA53ULBFW9WKSF9H/pI79Vbpj4dFwN3F07cAdzbcPCnxy8p8CzXdYyKoYf0
i30zRcPR46OQolcf9KaKwaNhIa7xpkVXimFIlaM24Q+gG9eP0hjTzjkuOElN7r1o092aCYkllJ52
kfWMLahpwTf1/KquMHTlCXY/15bBY6kqaYKxZdyGIDYc4FU7x8Mp4LQi08zMicixGqBdAvkSJCSB
5UDzA65yV8OcMkek/T4HzPVBeEz4ch8HPmmzof6InP96J8WsrENlryfmXuCsspiqAb+9j0GkFtLm
qDT+aKmTF5XP29O8HufvbquS7QwYR9Qr5pDpBZklYJ5mmNtdpCuH6iZ+RCUdrv+c+Mzcu56AFVDC
u3fJH/t9PPo8UrFKiZ/dqGnUNugfWyVxuNpl0p/eKPmEQ3PEaX8JipBbQT74SPiVZMvZimNm457u
cwcjdUajgXO6nHDK7R8PVbjsH7AVunCKtOjX69z6MoK/WXBMRpXz6oMKkPrdMWjBq6FEgdJGZx0O
EkkXxmyWZeknAoe39K6WRzD9fz3G6cdZB703RMsQAXxkW8W6M48xXROLPJ7nZDS0DFjy8UYty7GA
l1pjsvR5di1mN7z4/su6PDEcpr3eDi5XfqNXwX2cYuzhzLI2ORZcuWwlJto3+T2uzSAKhfgYJfw7
hVn13liA0Rv+Ltdkd07XNXO3Obctv19c3+PrCkgNn5oXeJMpgJGoE2juPm389zDfBG5l4uoC4h6Y
LrHxM2W9JcLgldhlIP22oPWVQOwdgkNq6QN1J9rM0txrh65wQ79/gPBgpacjjtii47+TtPcJEUHL
a6DCItW1iblxzKvCuOfGsJ0nNHJnCDViT6JiEzt7wYVN+9Vx59dOD4hDOP90BxhkjR1UEACORyc1
CbLvpRYlBC+Rj9+9QFkT3IwqxmvO+M7A+QThJDjAm5A/wei711nnxDd3MFXMWJ/ew4Qx7d7IjTEZ
Z5K4xmaTa97V4RsB69Q0a1vXe9vtfs1qbEc0THPkAPsByEikuhWyzcpk3d1Jowok2vEgDUv6m7uL
OH+nB5mt71L4ckPGyxjFO5H65kWxGkVVbdyO7g/NddZVUsnH1mK+4+GjcykwV8lkCBcjH0v/ZlC/
CGxx+DRitJl45VnbN8pvShwfV6jZMfdKEs3hhbN9xvFW6V7UiRUMywK3mOaWZHDLBU3iMeIPu79S
ZkENPsFtnKYHH8UXwuw2vNkK1TwjQNHGEAN0YSA80XuFXXnrNCbGIlq22Mtd5ae/R7BN1b/I2Ger
aXoKSPJ4Zsr9V208xPqatlSEM5O7UQsNoCjKcYEGBJ1qRQIgnK5hhxYPKRLnVYHoZa7WV3AlJ7HB
rBkvCzVfqF1WlOcS2RKp71pypGhQpdvD6/yTiw0JlFtLz5EdXebGFjM7Nbv+e3qewDbvPlXI477V
ezavzncKCeiJMlbcIzAqqMZzF0rnErhZXOjzpX5McXFvzHiqJn3hCw8SjDydV+hsnzrgDBCrFH3F
OEj0SlDpngPYDWT6RlYcj09KhapMMXfWqn3LtbLmz1ayVf6F9FYa6p0ZnkwCvMqtvIHdkH+9IZHc
cCoM849lWOInYT4JLA9Nsq5e1s8e7L79ynjoOiBEWXT5ssWmDhK/BWCf2FCYm/MxPuEYVeXTuENH
2OZaHbGoRGur9d324XIFk5KHBIWwDltvRNRU8PSrmE7QhIvz9o0vbGvMr09JcqcKTYHwLiI5odQ7
vtIDSS6A/LVjNQMwSQdGuN0gufpqJJmMpD9JQB/lDmmaBsWo0E+9dYNxL2Bohmu2rhjPcnEXpelV
Q6N/ptnGJdtbuWBHLeWUKSDghtLQdQvm0r5tWEs8ksw9uMg4Yd4ap/MIFPYO0kRM3R3U6FVQsnaW
mVMZnh9N3HwIuIxNmlw3UjKinO6kRqW9EjyFbS/XOEfvzooGcohaQpFwOUP2uST7y9oFlXMmrMEE
GRDNieVnwjf9prXit9LZ3ZI0go+iDX1i3C4GbDIZjyqdQ+bgqW6z+4UN5ZWRGRXmIpZI48laX+Lp
3F5wqtZ9FNUQrD1Dg434WbRsACEhHpyhrz4/KZ6vodBxgo/R53IIFox/xItnw6ndNtHnt4q6syAc
naTygbZVjlWHnzf0KAPdl9ycow8uYmFDkYcy0BG5zZMSgKtolkIQUvrZNkiK9FAmfDboWvPLvcga
jCZVHXKi95M6pJJ33G81izwxXV21lID9rIbplpkhGG6/F+WSdLPaGfHhmjyKagN37gG9pYwMxk0T
GXNiQhaH8kIrbEvctvJ+6D0R6TQ2A5TpX1D2YhhxCUSJ8+IKKETHUd4RX+iqi5AtEb13zlF0S+A2
RckG2yBwAGd+6Bay+skA5AbDkosYNu+QseTrw7GtwNItHh/TNgdb2ayDpps8M0LAjo1/8LoW+9no
mub6hNvvKM1Xj3sY4evbBwA+q/ddqorlBdmWnskIg6e2OI44aX8tMevI7Atnbus0TiQFNyH2MSw9
BBr9/GUNwtet5QtyaplpokVFQdcuoR23l3MhmYqkBC0nN1nHyBkiW9i2mXycRvIQhBWoaSdOfMdk
EunyOjRJi5IoxqblH+ewl0TwPmEJJEygEWXseFoSL4OthwVwcqalasfNoxtCUOPawWvOF8FsY+Z+
CNAdgjYHtSFhJGo3vCf0eSul+OEP0EFwRpeQSMe+nkWZmG5DCedlLBykGPli7M7UGpYlamtvnNTN
Jsw0WHLIa1ceuh07bdAY3lLW5u6ctEg8TykvZrvNj+kWrJYznbcfX3oIBucnGWJ5Xajm7oP0ZL2b
ber9PwY93gV7JaNopgYus31XD80lcJyl7FRl7JgPXJZ6BnpEBQedDShx1JtMoaLn00KDwnqYgZCy
XH9aRaKLefU6cgqkYciAhx/HtZCSdxpYPMyOwpvsRzrtogoYRGo2huFfGnlLwxVEuFA9JNGEyPKq
IOE4JqW7jhjcn6zNIh8v71dryPw6W0b3TjQ5jg5LnqQKjvcwBVyIEGjCwMxK7w1iRZFWfQ/mco+w
DPcmTrMljiUFmnSuANcrAaa+ZA3qXGQDd2V1bDJgXolD95hmFqnHrzX337LCNAyyqqvFsx4pyf1p
mWVBjMciX7LbJezOHhDgj8+HzpB4DPm9H7/z3ZiwGIvzKPZ/KcRDfGW1wYPz/kl87fSBepAwZ9Re
wpEXjmYMJNSU03FJKcANI57rs+IQ/QF5me9LOAdwR3cg6G4DGI0Ro70eHYhMJNfUJDV+AsUgVuKb
s4mmjEIWffN6WvCEivqaIfaMa40BU0rJqmB4hhMegI1B6XLIA4cg+xzkd6XVjlCYJzGKrY2T0Wfj
q9OYyvSphrYScZuzA3aU6mWigX91VGxY7wuKFYPNQjYw+/3wEmWpJXSsl/BVUw9+/YJVOdXrp4Hi
73S9PBMoJX40DWI8J1cNVz4xdNaO3tmK2ez/HIGcc6Cewxu4RaXCgBPHe/6KrGWu3nW+vSI71ei6
7Ai7mj/dfJT+SD7rIsw457zFmY6Xb6l1u89i/GcrSDxeb/Ar2p9/mK6UMf+MOasKudqlQiFQj6h4
Uy9mN2mhYxNmYXGBT3jadWTD1wMJFX2CenZaZM2kraiN/Ao6pLT7zpAD2nBisVfaIF8cbKoiiR2n
sKSn6cAFpc3Z1mEZ/FAhOdrpQY19VXlwZ/OnM/IhATFBwt8I40l5IECduyrykG01QRnZ0ygmICNq
qIQB7cqBwhBTd5FCdiHn0jpgT5Kf99vOotvs31gdBGK5Uz3KJuto98a2gj9Wdgrb1qK8Qgc1pdlb
dBIg377B5k3fV/A1qDvySdT/QkO0jux+sfNb5BA3eo2ERYv6/hA2j+JKsYibrD6EEkuXstj3aSpH
R1bbBS5rHurIMdXLulRoH0S+Ul4WUUZDbB0Y5L4+u69e39b5RqUifkA1pG3OXENM+jTBiJKf/RIT
PrO4fbGPwK+aTTuY7++h9Ks+v7SizEWo4xaqmuKxRdkYrObVtTknL1joOvsXqWIT/OtXmFX14JdU
lycxDTV7oD6ZT/aLbcqFzwRchk9kc5BWklWFmxIGVKt3rqzZss85kQJPJaEpIK636CnW0gnc2H33
LUhb9GGMpkSmn6OS/lAfnoEb/xqWYwFXXp0loIn51XDX82WwX68d7YYetM6JMIBTJsMOO6V2KEFg
IRSUlOOAEm7WTYu1FAtd/iQFDitz+WZIwXEGwKiCR1jJwTkg0NZwOUmATOZJ00sXnScHxXc+L/Ix
5T5xvkJoqEKfETsMGsp7KIKVlC/BXO8/9MPjQ4kaSmgjD1fIA0PjgvK5cTXQ0KITmX1YEg9VfPB/
WvZmMq0EscdJKjw0C6AFDPaJfcCHFm9oUZHANX9NwYcqGY+c/2HZyXiNhsJjFWSiIi1dDy/UZMYx
wAO/wWmdndnQSpIN8soGylI2NMd7bs9YZiNcBoXDNBS17tim8o4UFy5ckGhAa6y1777gl07ZClZr
mbMQW1s7hjurEpeY4XmZcGQJg1kpUFy7/cwR1UX/AYoA+mizqUKsZE57L18x8Cgc+BzVavTSiTBm
B8fwm24atEt3TdaiFrbeY6/ohhHm3JtwkI8Ebxzn2TBatNTwDNeS4TjHm3gvRULLUJzvmsRjuLz9
5DhD6CoEsp4Jnpu5kQhohzl5jvgVqEoPPuP0n7a8VNumSct3W5YxUBf5y6cXvwGjgjP6Ry+EfXlk
R7ok+OqQKQ6RcQsYL9p1x1/EXQDz8nrpcNbfecPEMMqwfaL7EeAqX3akBFfPd+3ffMU3MSw1IAmJ
R2PyxaUzqDTKtZOrupdFCJBZmHZDV0y7+vZN3+f1UeB1Czpb2wUKK4AIMxzPWCJ2VpJ1OcSftdcH
7z+RNW0FBz2Wo07SvKT7oVRU9MOhwT4O2LJrMv9S/gDvorvY6LiXqs/RLnIfaQyf7nkAJPYictdf
nLhkL9NcRnE7d3s7ZjnBdepm2FlCBFVCLQfTrnA1VK8pzm6x6U4dcPj08K5Qhm6E4pVFcKl4eNGa
Q5TEspH7AEAlfBRIHdj4RPK9FKyPmkq/8H5TbXxS4kQ8YKGYwhdIdXYr+4XpgR3ZEsVe05yt6ZR1
vFn1qSqJisTFFEG+tL3OAAyR4t01yZXlpGtt2DkAsVp2BI4GnWYyjL8/2jLu/gWH8nFpbyoG/xOR
HZn/gD/KJZO5kHRm1b51CVmX8x3X4IVJHcea4IXHBvJOmQIuVe+STFmKrBka3Em7ens8DWgmG08v
/x5cESthgNdNyp+8iUdLd+6I7uchmzPoMYtIpDwdZt5ijFH7qc56JanYtAws5AKi1IpuMasqL8zT
S5GRyWQNWQNxieS8gtGI/U8rQKMaBBbusR4YuI3DzStQCtjeeq/18CIfyLQtOGQ69sCSdZgsBQhT
nDekXKnnb7u793KZg6Kt0EIn/zoJZbEm80uNRCbboXLaJOSQD4yw8V5Gz24KL3IE2of5T3+apXpd
5g/rbiokxWIGB8TcXsY5uvaz1O3dzalYDXe03nJCXnTwT+GASzVqgOmW5c21dTx/SOB4eR4OX8T0
LpEuJB5BOCkVh2Tw80ZIrDTDAAdeUhrYssQZ8I2jw6WwNUMOOxW/Fsqs4vE4T1hjV7YjA1giN5ux
iyyVPpABLFmxui9ROLHtpH2JSq53/CL+gcPjvf18r8rWLL9S4ZbVqKGT0SgfQTEaPOeR3VthXwcE
0qGxEd87UXxB2TTW2vOc31umV6V9XZ6gbEq+T3hbYqBJf8MyIYQ4jVkBxkcvmEqM/NvX6nq1Y6b6
wXHOCRUEWgUSyIqGoElZhHGW3Kp1rOKjxga+RU2BFs+xO2wgl1d6jphBjHWQq/140up7X9dFWAUz
zEQZmEPSaF6PfpFFEbpUgYYL06FEn8fjorLV93tXV1I2W0/5cRANdTdib02jbzxbnriY2qQxusF1
/uJlYQlDXENqtn715I4XpC2HF4llvN8SqCWMjEGP80ZhQi2xbFjXNFT+LvrF/JGZi9xMbUsPQwsw
YICv7638XPD/JGAUdAOLzlNENrLBo24llVB9C8tgq3iSrXbdRACrkyji0yzbzgNIqyu/PQgd9En6
asQhBs5yq5xhE1JHkyNJNVo7sqsLw4V2u2BVfZKHD9kKyxnKHs1XgYud+/6JjVpdklOq9K3CB6Fu
Dks2aXWSxf6rYmbc3RqpPsC7/TY0O3sPD0kfufmKoSM5RfhvKZ09636WQSSI5eRlowmozJzXG6Kp
7SyyhpAauxOryxOqP/E/PkdgOHBJq02fcgBVMHMjrfuxdwG5SzVHlR7Wd3iqq2F9Kw86bqdpEuWA
rgYktKI9zX3qevG9sgqhfQ/Buzu/rA5+8sMkupTxv2IsShkoJfObDxiqXyJeJ3Rznco8VfjZYVpw
rkppXoMcKsj0DzPPrHQfUt9QTPLBvSo4oc8BatTYr0ZX+lEKF2weqDbwz+Xt2e9J3+GLtI8AyR96
wMeHoTOJ/GEH99BrLE7H6b6I/zFKB35nRdy/XKsS2q4MNmAc0WFAM1cTcMN9jB8eYoSWU7IzkXSV
UmdlsyK59Yw4Dkjh1Ly1sOeE5k2VIxv9kZP6PQdG2v3BBXHF53ObnzxDoGftv/mjqpu4qWv9n6iy
dKgXwZNGbZX8mjpuFKxZBtU6UmWlLjyLr5mTehkbuPlMtlNEIj9EjDGp+nxZNImpPo6Spp+J3h3O
NUSLuAwbnaI0wDntMYjETVCIl0dEVZ+lepQr5cuYvNP1FSl3OWcVGlIkfLKnZpFfh3GIjx62Nqq1
QYk8YksCQ+GBcrFcSV6wRwl9BraJuUNuO/3VE1gjWwwJZHtvf8ZBxmEY+Yh9xvdYE3ZormuO9x1y
W61cBks+CIrsVQDd137q+BoDsn2y8b4+QPn1CFuMHQZuuD20xf2cCzjIB1CMlwLlCnEf+xz3m5Tk
GHk7E1H2jP/NBTN5RlidHxZpdFOR6fg5AsFtSFCjgviPJwGs9lxvevC4fv3S0CYQ8LqOkvWk1WLS
AIpZI1MV13ls3kZ3/cZhpxOIXQC1mPoGAJHm9CalOlBAGusuNUXJrkmR/BC9n4wwHMpxMIlaTATc
rM7PnxEqSTRCeY21ZTJ7afsAQKa4lE3K/21BqYQmTHzji8UqpZsVbhPeeL3cDdBCmOifYoCRznUd
7QGZRxZSdTGA7LXJyFznfd0ep4oj/szhvOL/Z48+ulxIwbcds4thaTKDJONB6G0OPaP7D/TAXTYC
R0JcZIcVLUDdZUwL2ZKrv3c7TfJq8EPH9hmlwgaseXt4GY5uaFrnNKgN6uOV5tTOisJ0snM4MX4q
W8Zg0TeWQCcpwrlDRMpQS+FDM68M9vFyvreq5MMjV1kBU0iQOHoC0TBFuFpkYM6xR2dU4fghYr1D
eVr4hgQ8gbINOyd2AQIi5HXxyXrqrM4pB+QbQbjdr4KwwHT/9NmSboksEePHmFMVyfYcsvMuiwFb
fZx+F9P9gVDSAkz8A9ErCf4bLmQSb6j2bqWIue0yiSZbch4l4neRZQmy7+S4a6dfOgklNXD7nVXo
Jom2l8WKyHC8zAv/uY0h68ByWYT8M0ZUk/LGbIlCan7D/6WYYAgVRq8D+pkl8ptaJmybg0BFF39M
fAwO7ViyDREfyIMoxliRTw8Mh9m0OfbL5gWCtljp+l4PfEqptbASsSRr8ciscEfLtzdKwxXXMWEC
LAm1ANYS4S3xoTVVRxMymH1SnmBNqKqI+W1FBo1zxuegGW7lWvqVF2MsyAoebVu2JtbNjdZ1mp99
mPYeE2cCuQB5BkAO0eP0J8wedsQSP7uaEGBNHWGgWwTGvUt551w4B/ugJKnezPkrjeR4A6LDikYk
1WTBhgfqBoDRUGzeMgTdP0ZmiY2ydfN9ITGIq3LTVlg580HB9l4RzPkTq4ya3wR87S4iR6CeZgdr
uDxhL4RU4ZMu4HYBEyBIcym4FZkKxInsjZzzXse31QXIdnR9I3GzGqDBYncWta/eRKswqscA+zQM
iNXhwRzqhNu5IpS8CVmR39BfQfTH0zWQblrcH1o8rbCOsgVU6ArLKMsOz7eR9y1o/Bf1GfpuOpGb
VeTBgmjKhSUBX6Im/a5C2RFQ6z4B9r2qxkXRGBGvPil2YI/P0kDyhM9uHREDB4fKHrNURpoXPUQe
Ku8HwFxeRDL490T1KbAkesMu1OVwhOqjox1et4Cix6InDnZSWZSAaTaxkXKMyIO9VXtY0l/PZnbr
29R/rj1CrZ/n3y1uVkPB4c78TCxoEUvFU5d6tWabCiJCq0SOT7m6DENZoU9lt511Pt6airGrhwx9
kr2pa/+DFVY9I6WE88Jg02pJqifvcp/TRoTB1D93EpegbV6gkh/iFhfd9kQoCRlwaN40/2hcsTEi
RwwVGJ3voTpstXsirmkjmJTxtNQYL4goMfqtuM3HjtjDpPF0g4vfBMNB5lr22i3KliYG5F6tS+ji
b1kePJmi45hiP3tmHSBq1MzthLLAhLlwExs8ANg9aW125jKdEWc/rXE1+/NxKPnZEoiTnMP8YVpA
a4wHXiGe5tZV6Rw744WZ3ouvb1c/3Xw0RZ/bpgv+nLyOa+I3piBob71HBs3RUjrlYni1datqNfxG
i+bpDwER8UMihMoZVUMoZ51+ZF/V3BGEz/l6In2LUXkGAIK0rfkW6O7L9lgke8RMEvD79FMnVBNl
M0tfbwPvnItBfd898r/hLgfJ0pkgWy0Iw4qlDeMzb3QpMyVaWvTgVI8LhtPf2u26FrpkNM1TAzlx
bGFkwatLP8mnup9HjUcJLSWC3tPlPIE7v52BFjo5wy8MUYmiXhi2t3B/bPEh9AjLgbYsBxMEWur4
1iWx6pVHB/uD0rIEK9S1w6e7oP2khG+Ohl+k4Us7re75TN/F2GjvXMq+cuDbZBGlXDMXA6o8SbzA
kkb/OPFIYU0kclQlf/Xzum04+CysvP4h7BKAU7PUqjDuC2WakQAaAZjATh/L5l+Qu652fWcNzaUG
giEXre1iYT1H4vuv0qOU9aSAHcWv7xJZpcd+SxCeZzdHi4LPlZHd5sMArTJIwvOmoNeBscD6Uaxv
Mi3DYGX77ydV7Bttr8/sk1ezMb9zO2BmSj0/zOZTniVP0QBUEeIvTCbxIWVaC0zKgdMLKhDFlEHJ
rbuiVS54dZZFW4mKn4zIXNOFMueYkO9cu0LCOxoJIYogu/PCfc8rDlBKRf8o5Rfqu1EjQ0RjO+x7
Xb/Fgkvc/r+5xEkvk4H6aQmLJQzKK3dP9nM0EDAWqawAhI84iaVWY0gdReIH2BSwaQ7hPzvzznMl
fMlsqkMrZmw2s3jECBL9ag3+bkoEqwkaM4R2gdy80OxUsONGwpuSvv4N4RpY3zGffiXl9mp9vK9G
aBaNuWkFEcokz044l0+RMqCJ0hocY9bzxGijQvqQz2a+AIApp4jZ8MMR2seS0zNSdP0bPTtko5yv
vMAvLEt/rOkUMNx2y98+2IaVenapVOK3JBnqKNvbj3DzRryhAzF0Ud+l8TyFHczlXTQ73VDgJSbc
v7ULLNOmaUkC3mXFS0a+rQxJakTJyIEun8o0CAZvCWH5nFPZl9degsdUphVQXX7jdga6ZDN9yGel
cbP2ljMPQBqcVVBNPYf+5fps0/1dmDA2O+e+yNXeyU6n8X28iWw6IMFbkKRjdur0BotrqKRYB4yZ
c5h/bYP031G1mATthneG0tgp7Nq2nq8GDuqRMWc3IHZR8J0g0jm8Raq2AdJTmBCNos7l4ZZczI3H
31RVCwCYxM9uG9dM8QvrtVRGTX45nQBHK3Z4diHpy+iBo6PLIgMd0fRz6YFXPeF3QS/kCoFwOOI1
qkrwIf1OVHNYvCTOq2ctDrEBRbzUb54j3V2xbOw0YxAcbRVh0enB7AcT5HZ4RHWNFjLAR4okdxu/
pDAElfBfGhNCHqm5mwudOXXz8FBmAP31dSgCCtGKQzyRPCDGoFWhZ4khrGecbw+FbuTPCGQyGcZy
gfi6OeR3WMytG4jFe1MMhboE+EGGrDW5ZHbP3TBaguO3ldvlJQWFsKPaNv31h2do8BK4gw3C1zZz
QHya1lD88zJdg9Iq3R8LfL2jN00pT9B6ITFPyjC61RCS9jaaA82MXIrVY+/gUhYPkIhDKGF0lsG1
/bsEEeTt8xZPu/C7heTCA1INV+jBntS7CMqCvk8z+VwURQSfMjH2HbSHNwsGxmmaFMMD9e8tTlmJ
ufUmlL9HiTs9FND700Zkik0M2RHnhIF5WUXgiK5fi+7zXVE2rnDz+TVIxeoALrtat5FhEy5BqIMm
/Uw5uaiCdTQQsLAQUpL6nc3bVY2sRZaC04luPI2dRxOYrEwkxunlRuNS6xs3BDybpMpbAxV4H1p3
bdiIy0gZrd8uZzcubaQGifhmMtsg5ivf6weq8podpWrihZk83ULQ0ahxAfkFb6QjwLErjkN4R470
m0yHXtDJeRBei1PhIb0OG3lKY2W6CJHpifCnZX63CNak639UdpLBVMe91JX1Kzlu5L6MOI4F/QP7
nt6XVfVjCGNkofbMXABKSbC3YUV6nC3MhTI/6M+KQ6cu/cIZxBLk1O3qS5pomqLuDGF/y5AT1Om8
ARsmZmCan0zeyXjQWuGAD0B+KMxQy1S56RKJcUL3lGJx5upjc3PIHidSds99TVRoBzF59EBmjhqL
rSycZXhU8GNMz7r1XwEv10p1musqQtKM9vmtLtBGNfXE6gzVVg4SxRWwJR1nPFncHIVo/8RjgI5A
Jef25RQ6gOCeHJXUVa2RpEV2FFjsFRKIiCOfgEjbwj+WDZZLYHY+skj5XgRNZkQ9ZgezJ1Rk5aw+
nvgyEmfIxPCjUwjvrplEvRMhnob3Pk7Z2yU+vRPa7Lxsy4W0/deXpj+upzALNsMDsAYssFoipVbj
VBq4mLutvXNBguqFDHF2jDy1+FuUZgP31y1shE2rMW8Q7fw5DXLUEvNDZK5X9xpPPqxj8mHOdeyn
Q1K+em+g1HyOoddSM+jRXQ2TgZNgGx6lbsT+9PJ+tBkX0R5kWwkc8yC+/18tZv54XVi2eOvH1JOe
YS7k780E/NKlO1BgrXg3mAQI0Zvr/rPcQIiL0Ivul/1NnO3DQA4x+WlE5hk/URqtixAId6dWKagj
LbdqP4Mu0K2AOWD26edHpWoSjNoib41QRx1TAuS6xXCA/j8Sw50AyF/4EMZmUJH1im/bfhx3rGd4
2jzOp15FtiK7nfHaEowYF0yRPWZVYFDYSRiKLvI0H8udXHMG7Plgj3hY1RI3gboUeuN34xo2BLf+
F0DcQLf/f3AFp63/+eEsI4gHyA9GXGK4vS2Dirjv11muTIr3YBSHa9XJlP8wNhervs/wUDpr/Yt1
/v5kmdceY62UTAMElakBEcYVhUTKmC3Vk8srcP2GjnIYIQYBP8Qc8SuBr5MzeLrCnLIJdl14b1/w
KKcViSFkh2QBgGBYz+VktIpcvjD6dqMtZZfxyHYaU6O9f40qrUCOjxiFledKrwUtidZVhkcrWwBU
bMIowY7PYQP3hfaVf3PMgW2jxUzm/ldCwiiDdLhLpIh8sfmytFo4WsFYRrBrA7LgUGTMo5OpxUTn
I/iWpTtxY+Bki2K/rWtS1J0acXEq6iQMeFJfIzqSJSY3nB/53arffq1cB/2ACEgTbmLphz7SsizF
zrt9X8RywnvMPGMG+VXCPoqHJmMxCJfpA2+zsS0MeGbKNUxr3FR4XmZSNpNm8pCH6bCr5bV6lx0n
dkVh4unBlnoS6TN1S7yv9NUu5wtWIfJvQe4suRELrdbG3d5wErvlHrdVMjokJy4FtbtbTQBP5JB6
fcvtYIE1Uu9zlV5G8xqBA1XfJKCoSqwQBtVvZJjOaWr7Or6pbca4QVEldSZsD2LgRSOQWrFk1YxN
99HhgvybedCssog1zKZ/vImninBrgGMX90o2poUea0hPiCGLMhQuH37NLTRr38zRssRZHIPR4Fs3
rKrzy9BThbIExedR0fBm+ApleMjA7BFyhOnje+SYwQETQQejAJL4nD5n0O+n6hFwLaMuqxtgFDfM
eE4AbO+ABfcuYosDtfnL18rXXa4FCdXSxxGnmxuuwMBy8W7CsINBjvAx/H1C+Bwzq4PJ7YTZ9J7y
or7kTiXIOyd6y6jaU/aDOlIlpkwSxDK1jlqCwurOan6ooDaZF7yTmBz2BZVTuKwRb2igKTBFl9fk
qP1wvUY/s8xBo5TKBlPKs6Roj+iXidBV3LPDX1r1MPUCyD2TpKWBIoCH1A/glwpA/tOn33ABdCM6
FvQIJzlrLqfIXCryQD2TqPDuCkXVkTFat8Fbly5uu31uMtG/1hlqsGWqQTpQX3I1thMeWSeM3Vni
3flMlZVLXYilgKKxUFKpxYhoNy51CpIAM/Rp+52Lp4HXya1JgpzUcGg/hck6rcKl0B2Dg5VrekGM
bN9DW1Mwa2gGn7ruapZ5mnEzMQfDYzvd16Gk1zYL6nyIhZq1YQFmKjg/S+ps9SKgtVoQSvdqGKA9
FCJ1ezY3k1ffrkbfirxdYf+Vuna9METQuaovlchpbDkiiHgT00NlQWHgxuKAniJekzsxOmfCIT+z
Qq178lAS5maVFdvDRlAeDdvFWrJR40pAiB4mK2j0dx86RTjrAWLR9LXHwVjvE1/5vyNLUiUpcHAj
2Hvz8ugGP0Bpq0/zWjWVi8nP/jjPmgERxuZQQq3FZMWSSFhLK6M86Nel1EPIBlwCRuaqklTWDTDp
Hi+uAzh3Qe2WneADo2MmsjtkZrOBsaIdDjJINwMa0j/jdxSgex/3YB97AxkwnBOEiRQ8+ULEz6E+
FQsUl13SG1E0av2YD/5cwRi/WKnwVk16penK/TguGJLl77bM7hXVeACRE+0blBIDUAljGoOEgIe1
iur7jBRsb5IWR+Sb6aLc0DTZ92/R1YLwYDrW+6DSQ5W68X1CK02dEvYxSIXYmj4pyMObVVQYijCB
ombnx0ciMKW1aEOzsdShg9yaeoA3yXVOyaBQXaXWDoOprg3WjdRBej6x8+d1EN5z1Ee1e6/KxC5M
XXvz7ssLUtYGWzzD2iQewmYu1Tz19HQJg5hTyqNjjF+vR3AdSu3qnWleFcdQ1COklPE2U7qViKnB
e+2gaqOZ6nDCQBPaiwACtGIafBk4KsIVF2mGChSWnZprrb7Xi/1m3JW6hIo/VAXv5cq2sUNblNoE
KikwS+0w/QslBhTa7kPqF6ABrYJwo/gDVC6ziPJFrIStQMGItyp4QlOdsyzF0JsKIExctd3HowIx
IpdYPoUYruK6EQZFAIZwVt2WQaxF2QDtJ0HtWZcbiQFXeETRtEt8UxtwhehvdJ64b5KBGi667ssT
XESAaS4kAwKKxFGqdcqAJvWHh38ymbd7Be1SN/fa+Cql2Zfsysg2XJzZmqB7uDIn+36mqQSJvwC2
EJO1mEUYhsGv0LvkqFTlvf23u9Seogp+frOV5jX27l3wFOPhguDFd4CWRm2hpB/CeipH+M/QcLtT
koApTsgR1/iEAyN7Bo9MnvDGjYcvWbHk47lAcw4lsFslJ73Qg79wRPAegWsWyrBdaDavy+3GB6+a
Qkwxe3ypbB3Ixuht++3ReHfjBZDzfQUPtm9OaqinOkpE3V8/sN1wW9dWf+/rDzhN6xaYt3vCHYBH
oSx7UnRik+cJPDvruzBfBvYL8XqUyGSkJI9IJy8bDG3AaoGNce5tcHYH41UVk8w9nvavNOHnw05g
fl96GZGomw7kqd7b/JrNKuY2uh3Rmt4iTDBg+FjWPIsD8apIvATagjbL7FP/vdbpN5enopeQvioe
cowmcXmdi0rsdTIjGagIuuwlSXUZC2gQ0L4dxbhDHruM+8YE5NfnQA5w1RdwetA7rSijwQaBBVHS
aqKRFh2NtZYGeCKORdnquaHZCG3aJMW2z4SMEBxg+II/3T/APWb0CorvHMwlKUgV9mLNuBGE/rj8
jMN1O8tUbR2jnD0SZ8V0wIvQjkJb4dvTEQ54xp0OZwfM77884bC4XDtLlz2g0wFTExG8qnBRuydG
dw+tzmD+m7/7ojN3033if2Fgeg22fN0zRd/l92uaDaXA8f6QiDKbU36a9UB4ETXeUcl0KqhLVoWV
ufStFbFb6MYWPl7SoB3XuwtrB/Ysn68wYCBE80QG31V1JWXiftADaGsz+OcvtErenqJVnA5LlABQ
O3hYYVtJ9MZOm0YIabgx+gDCybpQtLL9WE93mPNV+PXm9PyX36u6rvPoxXnoVW9Cyt+bCwfxst3Q
fX78XlR6Xx/QfgDUvzC7+9hgUeRU4COAczerF1Yd/xe6ytpoQgefNDQFB8g6JGOIZ7pXvYEAm5+V
ssEhoVITqZXntfIzMvteUtzwcXdAGokI0Mky4shDqe3XpGVPfDfQ+BIfNxYStjI0juv3yWd3/WCJ
qbUipC9nSs8+2UIWEzILDACWTKEDF+Y4YGiRUCtzhRzBT84DU8yt4D5GUKgPj13qeGIg7jr2I/SM
foHFqzENvNDM628gekYgmb38QCUsAjtgZ885/IJ/eqKqQy3rsJsD+Ri+ZO19q5MOBe+L3HdJAkcF
fh9VF9e32cQPH/tvVJj24zb84zdzhJjvQ0J1F6DRSReONU+e5tkd6deBjqYSyHjfsqGG2keYds/c
0RLwxjwmxmPg6/WiZAqSNG5qJHIg8vnlac1cssjekwzOiau/LjDvN/TnRveybWmP+ixRkzwjy/9u
ZLpFA47mlFMvTngjXyS0pzF0CzHzmGwYvPSn4UiJnz9MWab6FmBYe3Y24K+d7zC2nvreCLUVF23F
OvQjvZ8qOFVUODkhBEOFEjR8UZ1YfRjt3J5tWNa/GWvfG8XRSAskZaat+0IViQH2C2VOmK6kXyy0
QTl2Twi8AEXp6aanYqHYlUkmVB24/rftECFoPfqzgx0yPaeW3SbWNHBXoWAGIAqsUtTqgxUyPKEB
S7mMO3G1gpg0y03w6l3fbQroimS95btjhEh9COQwl/jOLFGgv7/Li8GpJt2SA/Fo2DLNwhM1FGzn
jlXvBUIv8cVtmZK0LNxkPtjuo+mP5uZWNgvu0vA14rwztG166sgwdjblXnBu1Cl61nepvSP8MI1N
FD9BcN8Mga1yxbSK1x8SXZlxW/E10/teBk86e7PaSDg9uClwxNS/VytE9IwV3tkqaSnX9agMTe65
WBWZE1bQJ1eKMHq9z9YUxnVAmJfKQD4bq0GmFCmpkMvuebbrdyCxRK71Fkcx1M3twxR9CBgMt4z7
u//E3i6lFVkgLYsnPOHbhLyuFg3Mqgqx9n5+rUCAJ31pCZ8JqjnfQggNLOBhGbGaPJY+2YWJOnTw
XowUZE/20zhQ6BiDjwq+T8cG9kpFj/oFu6Ec3BEenvx/xBg+sTF27e6wCKRDCQcqYhYZRxxke2Zf
zlJ2VLrHqK5QGeMj/Dl5lbxe4wzHZ+VV+rvekrmsObm6Ft5rgQlt9rVh3knYv4eYb6Wo7AghBjZ0
Q91P/P4guMzVx5ewCujhiLArCnvYGx5LydWDXYs6YamFoxdt4++p6JzV5nUzeuyN2LHxePJAL71v
oula5naLY9DfGrejImHl/bVvhCNtxh4dVAZTua14zcImCjemi+Ry/FS03BAlBIP5D7fes5O6g2LX
Qrubeu5jg3CmuZ2icsdT9AB+p/v6pCAEY7vkPWfa8rPqllo7jY1b2fIcZseUMixz4HMzrMni2r24
+KvVjAFxNwSEOEWhkykxxQrRSVzbQFbkE/IdcS9Iy9C//y+xXvjwwidVyox5S2ag9anz4mauEDNz
aPqBs8HTJaDUqGDVck2zAoH0IAVJ7ig21sHvf0mEhYouMDEJDtbUUpq20C0kiMcHir4bpO5Y/hLU
mCYCUOIjH1W+qByY7RlRjaUbVPjwrVcMc+xVciEpK4F23AXwCsuz6zTDzACsOnBnWoBoYxSBDHef
JIVwp1UnNuPYniJUo0nG4sNpm158rNH20BGWYU6xeyPt/GCAJkHsv0fg8gmF4wqRve9sYfs9Co67
h2iw8Riv3Y9YQNAHjOG/hBSMf5z8NqI98zsGNosCcyh6iGt4HQiWVaM2oqPjKzxGwZG76aBosT0I
/oUdMiWv241+pc5YqOAKL0JYsvSN1k4lQL6RXrdXQ/TU0b8s2SE3K+6ILmHyEn0tqvFo02w3k2DY
nQ1tejCZSrPcGIoS62prBzeOsXt4USiwXYB/9NBLSCCdhjcIdflgs/5l+cRrkIDhM6w6WnhrIwA+
eCKxtUTq+TP2IJl15iz7w7zpbLN7D+PKhLKJjoy+22NFp4lpZQFoTBbKRrUSNew1LQS09FJ0eSeE
3ZB9v2+uVxKmZFmBWNZK7DJVC7Z79dnLuAcEheZ11zew9g7aKdagPOBr865mBVXlk4fipMmlpQQo
PYHIs0JTXH9c2p00rFpv9DGgJru0yOfUTJkC7+hiiW2C9S32LrZzNKwCkzuRmOctx94qTMqdfwVE
Hu4Xwss46ZAqV0KrkZaf/fbqY17KB2ZJItWGWO13x4A09l1kr2KnYPhKYfnIVV2U4Mk8wHKAIioG
b8WTnTr7i9/jbIjYPvBlThZLhyEFGcIQUTBcyMZdANk2HggPq53exLrm4CedT0mPeqIExPkSBaQL
trZmVs90kPuJI9UugqYq7DDrPjueYyypq4/EPh0/LS/9kyfNV73gSt5YNA+f1SN7XNaiT2kGRGEQ
+541RMIloFJc0Q6LuneLYO0DKc9Xl9QAkpiismmeu2WmpLiTA2F3JSjxru3+65VuhegZaswLFBvX
nQU7iJ1i0YiaffLc/GeVmQkwTp5kBs/Ggar2y1DAuReP21vKzK1jKBYHugAO+liM4u5PtkjLl0OO
Vpn+rcEEHd6RYnydTZK6L9/vm9N2rK04TXbhDlLSaqSA7vNIFkQDwL3pk9OQ8K1VWKdj9KtqybI2
FnPzUUdRGA0tm2+xCTc9haY/bRagR5yLoi4dclNQYbnYX9SOi1lhRMJj+wgbyzIEPD+gdo07cm+c
lxKMa/AKUVDstBsG8E7MQB6JZH+2zGiHVMnBQ+hhtWAUj/hNq9broXKckaoy/NkPGNRYf0bi9qut
0Z4sHpYR1z5CEqLohSmCuuGmtMc8lS8A8mJ3xKsJMWz9HT6xep5VjHH3bCZkw/2xq0KUAPmI8J9G
zui7CHWhfIfaPaC6WRyr7o0KA+hEtKMqm8zFlU9Rjvsom9rHhgKbmJjqt8RCV1oLpQLLWFbEiNJK
BN+rq9uVzqJOx2KcgIa0SG2kw1DPDhjfuvqEYk9SgGeKv/ma9cXvq/nZ1sP/QECzzn2C4FWQHWJg
v8DL5g3kcU21EKUCwHuz2biwfC2TGc/cCFg7Q9DuP3GPERm3u9CmeFGheQHp4SMFPRArY55ViOBC
YE15B8a6jEUOhMEdyetVmJlYPDKshU2Jcj+z/G27w6yNndDorMv8haouo8TXUJ7CDym/fHSWff3S
EXgfeu7+4OOz+vY2RWeKYNpBItfzNIjCrwnXd96L6O2JWZPZGyHXXvttKWEKZEYrXXYE+Kf8yYQE
CLhaMHjPlsq08YljMcOC1PpIuj15+HWRGjnqzilUY4wkWy+7C6vlQ6i/DYUxTPyAGUw4qzzD5B51
0m+OAImSMl8wpBMtF5KiRQ1aj/TZHlxsb3UbaE3Rhm//poBaY14obaG+IBTgrmBzFBxopTVh6JCI
LPFJVSf8bvuhETkscGKt9xGkjRjhi/OffjR6nofb79txXgEQ/zGyj+ae6XtEqZxmgGnh+v6l/0Dc
S9/7d0f5C6or/R1kFnjPH72jyiTXFX86rJEVvLp3rsZQ9/EmJAmxlL0V1BuFM0T6L+OV83YZJL8q
R1UoaSSxs2PZtwWlsucaHAmqZ3E2/OqsF1BxI5aPgYB/KKqNO5RKXiNsAOvLvqPoGBEJbITAX65o
z7mg9ijzGtkwSZlDfZVHUnaiTaqVnwqFuaVOID0Zm2lIaCVCJmslD0ek75QqUS/wBoH2CwmJGbPn
aUMAZ6szVEdT62YwRPB1NDlT9N1yMKLRPEtanlmto9UQGIojhWDvjJw6I5gI94ACBNpt8GC9PbZI
wixXlXuuGm5V/dBEGym9xLSn6Y1emrw5YzQce7eJaLj5MQNFNO95bnCpLLisN27hegLrZZH7sRKg
rGmybjR7CIuigCfQ15vaORP7BqM5u4yhlkpnApv4cQWjlRhYuLOkgtC9u+6lbrjte4ufQCXaA+sR
qx1jYnB4OE7q2UeYGHaoTZVypj8PJEkYUtOFTwytLogAT3bAhuCBkjGgvyuLOBCLHT6BO6g/AmCV
v8RZItKOZSzP+QfL4QL/fdsl2LWsa7wIfbEoWVCrGFSfE5CFRD3gPJAqGU2ZsKAQkBF7oeHzQta5
RfD9AaAs2/UilR3B3OIU9mdbbfGj/r1dvU4pik0hc4z/pSr66RkYOmSHL9kdcGylaQBmAW2i/Hy7
5zPAo3Bf7W8XluGvS3Akr1+xqbYRySsnoK5ubKp2IR54Zh7IkeQ3l80TtLuZLsyZktewQpLINWBa
WD5pHJj8SzFV4EE2NsEMIISIOSrSyrtiTcTvmFQXWRwGDlNtYszVuQKYfoEyPMoKM4yvQgYJXSz/
xBKwEd2hZziRINTIokLXyZMy0zuej47FBqYbdTUWFD7OxckJHEYWqVHWkgIq9pISuNLczJdFWUYN
JIecpqziLL1uKMP7ZEsJnGcDnXM/4+fPYCvWKZpH2ihjikiZYm86+hg9fLjT2KJTsFPZjFM47xIq
ahr8kwMkXyyKlJmG4d0TPx0RN1VzS2MKEmBsU8SBtmjSsxWudy5cat2f8s7Am1LtfHyZD9/Yr/jZ
nMeQDURwAS6Scf2fjCzgQJsXX/xDlEPntVR/sIM7vly6Y+rceu01LK5QgqDtpEUiP1KpUPoYyw3m
hL8NW9kQDPH/NRMVY8QMBtqzr6S1+Rb2QSDsslRV7nCK3GwSkuRS6sIFsT1lqUXi3qGYInun99u4
e6im4/1iKq/QsXK82RYNOJ2/mZgS82Bj4P0g/7c1EzVBuM5wh3Bt9Lc81RHwrZ+C2TKg/3mUtp8r
qfiQ/xSFXrMfEKIQtPsCMonMnn3mphAXh2ruu5bS27S8uFaLgDpn6KxQiDJ5cRQG3F9tpJPAwMs1
CzorCjxxxnIHNYHiKHvqkdgmuISFmWt8hJ0qZuEEpRZuJTO9QmfkpHR/s2H+kCi+60Oyn7hY0Ztl
p+0Dv59eSn51xwADKLrMxOT48f+pQfEex56IagogFAgfqXbUaiNQLb7a4Ya7KzqMnZgh1lpfGZBp
joolQVyTOaW53VTh4oUuSOV0GCDPiatsn72y7robCR0hqUpJqdbqMqYf0XJD5usgQ1hGJXCw2v7M
3hH6jKbVfoQexo/D0FMoK0RVfDr93ePRgbq8q0W0FwLwS4xugbHg+paKbnFh4jEnH5HdHw0fyHMM
O8+oj6EU9JfwSPiLs26FIr16R149fFpupG9INiLYUwPAn4Phq1Ps7YoR0VdTHVfWehUWxEk6gdyZ
iqEFpn3gpkqWluhRkXR7beCgS4SQyTXzD1pACQZ6pobpX6ZRzP1xwwmF008FhsYqGq6GmAEUQBvp
q7GWeUsyzgnDapzjjY0gn2Qhemm+baKrDzrm+J2bGBeOeT5KWeelBCqOzjDpaFKMTE51g8cluWYu
OtmJmnexHn9sotmFoEMgdKNF1padMvzW8mAXAurTUst0OVoj8ta8OElovT1Y6zU0ZuzhUXOo9ImC
1cabn9nxEXpa8LrugeqaRpHh+HnywpfLrGx8Lhg0rhYArKYMzwc31Se6MTskNAhQwgaa92CPq2s/
eKnWmBvdhxpgx8RZHXtcgbNzHjZyTDn3ZBlDBdOvqmOkU4HSxlrna61x2S+GJ3dV/fQ5w9S2oN0x
b72uqwnKcPs6J+DVCwAePUnYaQcpoNROAOp4R6QR5vvKavQzgRh4UvyI3Q9YstQYy+CeZQjQUZ6U
+5J9QFkxKHZ7KhMsmrJjSR8RbEdRdugRzWbnO+lL2dP2HfYc+pxDZ9teZawWcM29uAcQ+4mVpHHf
G2C5L1edT0RnDRB19+GjkzAcRdBbmwgqmXRJxrT6xvrtfHXMqhCszywncCjYag5bQ+U4At9iXtil
N/24nwyNMIxdwriRqEZkB9exx7Ut+UuLzqQCsIYA0aWFb0WUglJ36PWw8DvlyGH9vNULONkc027l
/Xk4s2beL3Z0193+7OsQH4L1+sJ45k8u4lBkgtDGjpRhVAn3YY6xoqBB0mf/S+WdddlEjzmtpydC
WYQijDmcYy5ektjQzrQujthNGM+rPGLHn/dScdqeC9gYYUXF38/u1JWAaMYJKJsuKAYXDZUmlXJ8
TuCyfUq4ipET9DtYnIEVr/WgO9XXTsc6zMrS6TW8WXXDVcjpmUpV3jPggc1LDVSYXAF0JpMt4iJt
S9DqI3KiH1fxmyXTgKjs/b/QsgZ37L47YbKCMl7p4/b5BjXWKVVxawSobb28zSuZBEfL9yLWtDdw
1762jnejqL76q6OcpnXinBPW8XeEsFU3n0zTyDa7yQJRnzeisI0/ocO0f0Y7cLOpw9ITYi6MeNxC
KjtF1pFJgKM6QchrZWEslSsT3b07El+CsOeNsiF/1Cg6gTvgzfFfKYM1NB/3dBhoDL0DJSlqp4fY
6tnu4y3i8553p+D58C+ZFzw5aq0lmoQmad5TY8TuzA0tOQBNHgjxGYokxDNxjakD6NpmbsIiTn8G
MTMvl3CyLYZdBDSdsOTPS3siKcxEZ4COppcuNbNtDL+qNGn6kAHkoEsR6Gv8QuoXMEsmGZVgLWjq
D+YK7hYBnkaR2dYsW8Su2mLMDFYmJeZWzWX2OThZjvOpNnli3igKGu7QrtCJQTHrBGjKr7oIROru
r5PwsO/jau7vFJ0vNdt6p6JJvaIydQPucAUYPPGYfh1LigowX/6VU6YZNtOrG/cHDVJHzxRcloD/
KtPtXsBwH08iXieWKbY5NrdwEVjmOAHo7JLdVAReHT9QE+3d/p977cb+A1PxPsxmrYg1k5PantJA
fWt024rI2F32rqOypdrEDjf9epF9o/EUg6A32wHS4j8MiW8RdtluMF4u0u+TJRfctYs5YKqjfCYd
s36L92Lr4ZQJ0CGTHeY3/Owd0+YXdv9DyZYJ42fjl77zbZcb+ZhLjd5gyDwjfvibNjXpp+K1ZX3X
WPqadkpXXyhf0dxauTfg2TU35xEyHZ8/TLXS8nyIxM/bS7ls3YVCIWRLF+t2aLo+3QcneJnmLAkP
8w+2+nN2VyJL5D8FdCYsfSv/9KmnrEVmPQiXGEsGExdoTExrXzXwAxZCt/HVzMcweBiUG+Ykdn4E
Dl/Ic3WMiLQrIShIOn1LxeoPJbbfj4yB10IQ8s082Cf5/c5vIWC0yOV2M5x4ldudeRmtZzw/LETo
EDaszTxQh/lCB/XwBzYwvUHXLEjWL09JJZ+3gocnXGWymHzJnisE/4/2jBqBVjQUZ2N2D/PpcA0+
bbQEE1pk4ELIvdjuo0w013BKYBitgMuVf58yrEQFYpcA6KEpguJ1vYVf9QM0TEoNRS5X88LHSx6p
KPn64LLwwyC8+wf/C/tayxPVEqpUY60If6agWbCqS4/NsnMxo24uWvVTMyEKfFoOnHoqEUYQJAqM
0xHhYoB4U1mA/o3dGr0aIjFFscfj5azxywBP+qiivLoZrb4BEWN5WTHTz+rv8qVehTAsQrIJbLxf
2m8LHj5XJkFnnDGTmd6AgjlqAUFidmSeRcIA4MiUYJs6NvVF9WtGXAgDbtWyJAcjuO6Hqc8h+AWG
uC49RQNb/SPRTT0Vh51Mg6PZVY3fYqgW9kJbNlv7Fm9KxZ++w+55DbmjnThXipdZnP7GHFxoYu9O
cdRty0ike7zfvwHOY25fVUyvIAUg3PiU91T+EZ6VbN2CY4Kuk9raSxiEs8d/DGhinInPCY2ukMzi
rRyz6m+dVWVYinQcqANBoJ0sQCTvjcas0sm6rEltht0qtD+XIIkxyj5jRvo+cL7RZoreqUMO/oDN
S/OClrCWqz8kfspD7P10xBQf4dV7mPerg91Gz0qYlBIbOIW4eXOX5LLE7T7dVteaig2jUjFN2k1H
BXUrN7zajp6Wg8SHStVODkMYVD31dCdCaC0K7qi4YniqUVT1nTZVrvi7hqZNmCFz8HNdmaIN7QWY
8xo7ICBvWpqtVF5778MGl//0c5ybW4hHAxqFok3uIdmkj5y9c6vJPzsfep7SqprTWyhkvb+DUJ05
cem+cktJmZiva4Dw9jOltQiunFKdO/vC7cAV6jDWjvD4x4wiaYb/nieSEeUIrQlro21mVPJdLFlj
O/3VeNIRpDMIvWcyBpDjgEwOi12zLAlz2P+UpPZzfdgm+X2KEWC4smliaurztPLmQSbNoMnDrsMb
zFxitI128Jyx0SGCc5U6LgTYAjJoR41PcVuna2BL5jychVznyzYpWGMBUHY4SVE3rPX+SzSfKQ+h
tycyTeCK44JAo8S9+1eUPnOPlJch4AEpD+C+hYY9iy/rxmCyBfkMPCDfMEQGF9FtobVjh2fjWWbz
LqAhRfRvHbWEl4IYoThQE9JjKULGyZMaAUqAXI2+MQ381QySdbiqDdgjrDbC5AeMiNBkRVGmxhYJ
Dp8gRXV7zer6fLN8PrP0pGedhoW0Tg5CXtxNChA748BrSe3ugJMjMvU5ujtlyvmUDzNH0ek2pvyT
o0vcWBlzQRMt0Vk0hqnSh1L/FbMQ5786FGfelrxZ3S6m1F0NP6oYwIav3E3zxpzNee+f4kpyvy36
h2nAeGFA9pR7foo1w0BjpdlBnZqBKB1CkvCtsJwEGtrzJZb96QXaM8BlQYgdtnAnVr8tTrjyDOD0
3V376cIakUm2ESlwm4YEfVKUHZAxTZvNuaJCFTGLGUfdppYqCNPhiX789OIoW9d7pIxSADxY0A01
oL60P9o4gxT9CxKp04irlyPTD2I/6tiCxawSYOfeP/BWzY27R7O79nD+sLBxI1HXAVFDNF/WpDPT
Q5sh9+xkNhV4xZaXA+eCmViVK4oAu+nn95yUIWZJaO+LI6/d4kwQJk+jGCInAUfdiuiRmJxuTnCE
5K8UR8dizwt5CkwJUI2+D4IWUjtOVI66geiZSWdQgLpX9hNJw7tiCzcfrq0Oi21PTc0cHe4cIlFV
e6ylYpLWPE/fCqAtAFbF9tvdfvCZVN2kLiSYwG1+1sNiac401jBGEwN6XnS+YHnR/2vImTUvNGVb
c4b6zzLJETNpcx0NgVABtw3lqt0mXpaktFmzlso8uNEidkdYun38sFGSEbUDiRPAUIfMv1iiL1qf
tI0mPL4QWBcQA9KaYR6hhp1Cy2RryjdUdWLmHCqjvrRRG6jarWxjjsgmcBrQ7JdiSmsLYCRjPlsZ
1P0id3Z0+oMZh/vH9MpXJlScAWaqllEUOJlgaeDAwN6lhd4GCkhNCl81E87tH6P/dghtyK0J0ANo
bxYXP+79X9Grgk/Rhd1z5LDTZ1OAVkjEaPrqOQjfanonEqIMiE2O/wrm7CTB9V6TgZhWV+IiXYLm
oqcvuF1Tc2/KpkAdGNnM85FNv8PaMDnMXfJoV4Sl8m1T9/MFmcvFJ0sSViqQAaoauQoQz5eXcSlJ
JoJUyMGyIWGAi8Vk3OdFf7src5+D7jTMPXgUoCD+2nYlr4T0x4Tn7GcPqKhMP7LM170e382sIw3a
o7FFf5ub/LLgvqFt/rcaNhenaNOSg7LxZdI3i7B3bQ5ee/QWupdeHk7xU3oP+9JG1LBHZcQ56KHV
kH49qXBFzpb9g7RGU/MolMRtcuvaUddCR3GG2uXC+boeMaQXWgD/NBuWJyxfWmNbR6QfL1Ubel27
j4foYDd7nVx2xIV/YX/smsSy7tCI3fNf112dj+AECLrefPpoFxSyipel0EJuPaL9nwWLMfan7jJa
ObrYGQUpmD0rZnL943/bsYsUMVugj4ac/UPQFOXYdwemhqxPc5MZJGtuL60ozV1Y+EKw/iDxQFpl
3yYW5sjkhHOg1oamm5BXqqhgAndb3NNGoOSgGLqcBR+BLjL9BkhQfBhktSZJ0XukEqlZ4As4spZ+
tAep0cQ0O0mnMCfMaYIjTUN/Ph1niJuL9kP5BQYCGLJzzDdHzPb042Y+Pou/aqurKjfAyFsu5wVJ
vmUgchfFOvyBH2Q0E0iMzeOfhj6vmDZUq4fD0v4IBdX4H0r0FZlPftG8ueed6kiSefgHfPIx50ck
XdSdmkqi9C2LObUqlq8jqIAu6ebbQ+jhH6sYbKVpez0bVJve6NMq2NgVnB4wDGLRsn/N5ImtNkln
Zoy2/KORoOEbW9xrwPqCHHLu3dfRwssGUXRW4pvfHOwa9Z9aFZ/0ySHormcU/kVTc5Pe80rQkVlK
1u9E6OMx9fm3b4tcz+NTXdu7TnPraeABIr2GwpDudJqEKN4pcRMA4HuWYv6YDLL/ATwcp66Ydp4g
QP8ZWG88iVDxihFcrvACXxY+HAagkwoKeNV1oB2X7WrwKKPMvkbUtA1OTPHEyVzGg4r8PZrSZZxr
qiXdX6vGO6s7V7vsLD4cxNKGKSnDc7fXrS0jQbIyuQMtseEGRJkzlP7xJ5M9KHDKEM5z6VdcYAi/
oqrpEb6ogLG56RMnOl3RUoIbYU+Qv8gZ5QZzKGSHmx9j+7tUbHg6NlthZ8AvDdhvi5PdnqEKy3tz
lkcbI0nbz/i7hH0m6ncOQYYXxVGAWv2p04twynkzJgYp+ta4iANBI7WTsfPmyFzg9+IHt/cBsQD3
0xos5pP6J3wOZaKRc5LN18ps3weU+06H8ujPxCpfDb8IyAQkjIABLqO5B03+NKkXgrP1FcT3jLx6
1akky9xfrBK+D3+WsXVK5TdtdrZGY/ddfe0Gwgzky3CmYkTWhRQbqUb7CjQYiF59rhXqLxIBC4yD
OOx66gHUX37Kv+qUTTxG0y0pC+vlb/ztHBZZft6eOgj/hH68EA17ppBkDsFtJ7qtnPr7ibveJDWa
vASFhkHqXg0Pd980BdkuysGIK/geHf4Gd17WGzqaGUcHB8HeNPS/93M/AJCSVGnGwH6luPIwMM8t
IS87xQKfmr5vY9i78luskX2wx+wdFi605NJjb5F4GKKTSxAdBPhqwA3dZH3U013YnPMYo9dF2Cq9
2BKp5Pfc8sx2FUpNcPnyTNrNv/YW2nbapFZ4c6pV2uVZjyiem3kHbweMEaijgfR0ec2hYnEHHRik
72ie+DemRYRfo/OHtOsfGjY23e3ys6rAwB18EahBR5Pm7xvb+zbNfTLYszAp/0atWquN8hPEdasr
/pCpFgeuo95kE4qVHeQB3vQfIXn8IMeQ1tqZToK9kkkeSMyyrvtqULuozPiix1/FpbcmkW/WaU/Y
R7W39eBd2T1g1BcLbX7U3xTbicYscv3auowFpUWPhIUkYpjZYlev5tnBSgQN+oC/MuXuO9eh4wxv
25cmw2HgLx9QPA1wxl2krgA8UkkG/OL0OQpk4rw8AmDHzKCnPI0TwQhpQfq8CvCCXq2yWURMmXHP
LFLih35kcHadEZymPJPUU3hVmMC/wH34udr2KYY+xueC1yHA+pHQapllsbS25iNwUl7NsNG4jYB/
TUAh0ceoPLRY+dvWjSKpY4mWimnOD2XtJEQ9zZk/rMp5nK1LUTDZ66LJOcn0L9TeJlo1NXV+iNP6
PLd3fUietLxFANj+zt/PyCxXiD9UD0TKZQywemTkKsvYZo8zmYT3cAfS4kR9wbHfcvyI76cobDh2
mk77bYw4w08e1FHbWypXQNqKVWYnWv68k0NkrkYCeN3UHw77oK3AiMdW6IVGgkeDw9LdP5UK97gl
r1eDIh19zzxBEdPplZUNR0JaA5U0rT8O3hf+667wP+wIN0y5DJinagVGuLC2IZKjXyZJHEp3Sv7k
f5ivS8cW70Sz6eDmBv9VhaRuNOMJ21jwHgT+ZqdpiqbIStH6d9IstuWfjZ4M6t3Qdx80JHpy0XdP
EyiMx3BPB7DoaNj+38cLlysl0BBdri7/PmaWdeU3u8x9Kqsp3Lb0nZL7y8lUb1DSU2kHmR7QNusE
wkcXEKukgbEhmwIcyKJMLdJ2HAN0sOjEcbudnZSDL8rymUhSTnd5+Mn0OfnvHWqrCZO+1u+7QT5Y
2kut1YySI8f7L76IfaLybqZChV3A6lyokDeYZGuwN39qVuWHHUZD3TWXH6B8GBJ/t15kxif3hwXZ
js9xTIX98HWclq8h10GmQpdaP27eMR+xKWyiWg9e68eIcloKv9o+izS5gNmxfg3g1MWfsWuftdwy
YM5N3KPZJjLBHFfgYnPs6BhicUgerNIee4w+X91au4m1tOvPBomUC3uwx1SswdrFCgvZXVWDyYF9
ctA+O+NEfWhEhJQjcFViezPvhPNwPufjbXnAnkGaBmiSZbkm+LB/E3eNxIeMG+nLPwpnB5Am+eYz
P7tkAHE1UUfQE+S9lWuaZKcmnT/aVBZ9blKswHnKJj47LQaJdSwtFx5tYE2q7YoIPnq1nvR0tBWG
haqYnjWhrXEghl/Xol+FknZIi7soYeHxZZdYVtl5yA/ZuDAVzLCoG2eCc5b6QFaM680eK2wr1laM
yvBg0Vmyhzts72JCpaoHdVokF+hWL/zLkV0MHvz1TPH6PLy7uFvMJy6Gwa8VTaqsSrKtb3ECkAYt
K5/njoTxYhBh878dZS54txFOnEXq7onv/XnOJNh/sJLKPYQkH8jtmNnW2WamUWuzcWpjG9GQA9hi
nMsXxiPg6KS+DVxFE+vv/nx5ljSkUx4T0EgAoX7e+o5Bd1rn6ruHz3uNEEoCMf2a7Kh1SV/x45sE
Bxqoi2jzUpaKKM9SGPITkk4mtl8EE3V14ijji4DXVX8mRhEB8JxO5yoaMHQhR2V40/HGJ3T66AX3
S+UKyrkz0NgkWQPtUzOB5CNsUFT1h8qL4EA7YmISBgGE22EcyrqA1zN4dsKc7gqDFhMTw4RjGlc+
CoYgF2x4+OEwug7bWDmeX86lg98vfF3JG/iomTzkyisrb96d+v2MbgBk3zfzooWFP1QqHONXS6F7
Wriwt0Jpjow4loVjHf2IsbUoD8MIJHdHlyzjWhgicmown3C780syOIPIVL8jkNoCkr1WNgkEzFDQ
zZnAoj5fDDpd04xMt6lUG56sdghbIp+nc3+u6I0GzwPqXMflLLWqT6Lxo57wX0S7QI7agO5x1wLA
RUIfd1bpeisCOFJ8EVYrA4Mj1USDfi6Y6KZwu9EyNEQ0l1/OdTjzY/ZgTDGmal4onB/5r3WJvEu+
62KzCFtjuvmlSzOqm18t97Iz3xwSqebvOdMEO3HNvFsnEhevCi3XXb6TRoRa17qWk7YizzZRACd5
tZAIJ4nDU1n7tc1E/CcQCnaCfx0J/e87RMwjyXJXFjHdDs7SmTER56I6LKmpblIyLI2EKjSKC+/S
vUpOphNZJmkZ742zlcY9bKn9KnwkBbJa3nYmkCQxKv+CMwMVImHBrcLIvEn/8xxRjcPtSMKkZlmW
uXVoi3J7nMmPf1/x3NajpyL7PutO6KnLMnxGjGYrw9DzOP0V/AOcjeDSMnI7ctlBRdHFaLMPnWTA
58xW4jaZLBzNx2l87wHlZmc2vsD7f7kKhYbS4Iih3GHYK/5mUQIp+uSbRwyRwtGJsnkgiS1XAz5z
m5D24K1X8kSQvPssb2HATjbhUdLkfL4w4rRgAAiFZE3yNQwOXE2Ti+2evmK7T43H9A6e6+jBpA2b
FSr6D9uaoYGhmhB5uWxaOZqvyp1hkyqSHMMYHqsyZzV9v+dTOwxs8ZAK/nI5PUY3ltXa0IuVL9I4
SgtZhkLH3hCC8UOwcASxrc37kUuE44mypOmqaJMtfTKTHd5aQuf4Q9inTBNG9qvYxu13vIzTp7dI
qArJrqgggGzb6fHs6xaRXu55O3O6Nf7sBCUAsRtRQAVjHAOWluf/BYzHwAexVkiXMHh2I6MbP7bg
a0+SlV2NxKWvcEh9QPoopdLYPmoRlZC3fEZlYwYs7fbEQMwSgE4ihJKy5oB7e9BIueXCeN9xm/Yi
RPZJyp7MTDZbz6/KOR6wEsyzupaq1CY7dchSSeqTQKS4/8YRsHGuGdiBiCieEMLHFHRaYc4UPk/c
iKtGWcXaGgXrdQbAq+7fsdiKXshLx8AwAo1Z3jktdnDPViQ4osvRoJ94hPpVLcfbBMMZ+Rd44PWQ
oAbp7ev2b0R9VKDdwEvsmM8CNUQdGF5pGwX9bakQdO+P52WMAGQiYsVJrqg0PaR53ecnKFwzhdTe
xWug9I9eQihvcmX6f3EC625T0Vgz2FsZmObsBHJ/l3FEtkMG7ayyHEaFIgOQMyoNo0vG1qc/vd3r
0SGMwrO1xxnqtb9DS3G2Om6wdTAgqTVGgNb2fBqSN9aUDPZq59gsiM6CANFLRKA5VyUbKV2gZRq+
poF08NnP6d7DWm7j6/nhseTb2z2AIauFih4BYHgTEOfjNM/sfu12qcv4SZu86V+txa6b98kWK6ho
UxCnxMExQz8M35kmGofi6iXSa31eF9Wj1x1gy+LLkqFDNTAWzJetFfZ8YnmeYLFEL25LKjGc0jjT
tkAvvBcEjQ6+gfTDQmsb1M3sT8ezoPKEHu3breRuT1iC1N/rPzPvf3oD2PE7/teWBBKlrQcbFWp/
1fKmY1GzVVZXaioDCz4jYn3QVGQBU+8SZzzXh9nLPyUKhtZMoZhe0PAYR7HXa6y49KFOd/5hEhla
r1r2UrSVJ+8Yqih+LCXeQPOexNCKqyYOu7XiQLuaigKx/GBBn06vgg0BarcPwdFyT9myM3uBA2Qh
ylOOkMBAIvEynHVjLyT6hWpYxaXgwyTTrI01Xf5AgJVFaP6K1ksoy1jOdNvQWQlC/BgsnN8fp6YG
7k7i6GUAkn/AVJYDfz0UcnpMg/6J8rryqB+Uuc4wv9s8UFJ19DtpoEl1AByiksKYBkSjT6VO96ta
2XYhvEu7elhaAxAju913el5Oy2QVTR8Dodjb/ABPFTcLn50oQtLfc343xMq924rG/zeD21Vtb4wr
Uy6BxhERIgOeWEdbagkZVdwlFsqo/2310c9JvUUG5ShkNiGXI4h7JSKC0CJoc8K8hEmGySXa4yKR
vIosUjvfaYHtO7dJrBC+UH0cMep8/tCZqolzdjFladqm685686HaPr3u1fPgRMNREoO0xwhol5GU
Y6wgpIUxJLoWIMOD5j/j/pCTwpMTbtyVEDhnbBBFMGk+PwX92UUHLdqDvWkSFhdheGNqz68xRIe3
Y7XN8tj3bccM/iUT4q3MDSsImwOL+Jcu8uDtMqsu6cOnzrFxF9pa3+defOXoaRaeSM0F/5WSwGYt
1kwg95cANykMQnN36NzKSOUasSjmIFknwqLPWOGfssouMNpAn73ORU0+xNuMoDU83wjjMlLvgT/z
CanI3mdGa5guChc5o2XaETZtTuNzvr0/4YVdFbu6lKB1y8WQvVDDAqFlcsK5lbY8K/GEZOwLZsqz
4w3gcWdr1oZak0tB89iFtTxT3JIITGWKWftbzDgBEn+L9Si8TV1qt9W5nZQNHP9VAwxxdn0KnMxs
PShdGyWUe0YU04Kv8yiPNIwAo7aLQ5VaKa/fir4y7uzHHqkXKwrlNwNzd6YiT5f5pq++IBLzh5Ba
FNx2jguvply2xNOqmyqyUMILRnR+rOao7d3sxE0gcbZQwzSswXsTYmbuZj7hCkKyB3zpxVF3CfNs
8JAbzP40Ia1pPh1iIqtGsrSJBINvCzkEGHpwSbYm3knwXHxE9Gota5Fd6Q5WRd7L8dP7uXXFgwm9
k2/z1kJnMasbGuRCHMuuy1MRGZAChpSOSrsV9THcy+DlFVJum8Q/nbonAzilSlFbbTgoTjrc9yRn
UH0v+YN5+JvM47rJuOKmGTTAcGT/Xehqp+dOePl4esfgRDozlDkk/mC8qYjC6E8z3eEaB8gTdYat
bCXYf2HiXla1YJbfs81FmGXfZ3kOQPoqfMynySpK6MX6EL0eopIHSZIzhcBWZkkxG+YSozT6yl5M
phXeFZMkLb/S/LqlSdviJVEnQ6GA2UExtPzj3etV7KGq1dCY0hNdNHhQ9flvHaztWe++OnZ0ux8O
6NQ4EC9b1L8zIdD/A2+pwAyrGWzFlMZKIxhoDdfry4fIXs99Tl131s1EjXQBGnuZmgmIv+s0cc8h
PpJXnx7841pGhimo/qzB2V5+DsutFaU2jLHmrlwTUE0K2UTrbXl9lmlfFUEoGB3Y9vmIMlZXW+dl
nVCSLYG2rQvCqMwoGQViduAi2B5MboHRwCB6kgQX2JHPj83+8q9pKqUhvMCxQ0e2wMzeXUjZp748
b61LRPi9Y4Oq/cTUZDMSKcuutsCiM5UmtQgzJA1SgNuHXhA5/Svhwh1zbl0hIaRtBFvbnkduKSmR
KmsOpHRBjm9d6uCSdaDRzMLEzpqoVZfO+iP/bsatU4A05vhs3b7yRErqRXkTNv3MYoiQNR6gmzP2
O99kJou5JO4IHf230NdC+fDibGI+ryF7yr1rnjo67zteEToBTaPHlfancYT5WXsvkQi7IjE5sOgF
WClOc9+NKVZjsWHb7XR09aZnV2pMbnUqD0rNUYhqXcaHMLf/XKWcm9O1L6HcYW0vXUQ7KIh4p3eG
152crD/cfF9prwv0MCUPVYdTknHRGxvvWKwgzUj2Y6SPa8sr0rc/AbPZvMxxLmxeGy7uN556q92d
NR0Fh3fnAbaX0sLWbc1gyWvJhSplO1YlQwptuQoW6FnT99mdVklcwCQqxE6yA6R0VTi/AvYKgXL5
3LhqqlskyArxuaBPK02Y+U+9XjDnLHGyZojcz2xuXcHznzwk5QEeFz8Rj8CR/wl2bq7+naWSnn8T
nLbEg6DBskUhkT49OQbOaHYe0VvZw5E1XR1PZ62VX1GHeszRtBjxSTBcdZ0RW/wEA3uJH0OV3qMa
sfmUy1XQj+yAPPuKRG8CUXA89Xo2dJ8U29NVn3DI46PL/x3EpkyregUXQF1cyFxx7xqTRCJ1QCaH
JUcsoqNGyLiqDKF4AODAO2m2qgJK4zat3/r2Nl5OAekhqX4sLcu/LX0okl59l0YeRQOqmASdzRKn
SY/i+BJpI4J0qsfRqzO28ek1udF9FkCyGsTCuwdgjHYGh6HM37gglDcjl2F8fX8TUjBrRCjqpGRv
b7DIqaHoW1IhVJAdjI6h8h2x89dMttnsSNT1umbYoJYirURFbaHhErztmcjnxThDGMmnmDYGOMTt
NdYIvMB4GKYd5TaTHIrrtJS1JXv7TA7O3wzHkMu2+ip7cEY6C6rX3cSJAo44qK9Ae8h2FlAhoTAM
g+JWs0FiUxgwstHE75P8yJ5FzA0jNy5tacJd4LSzAeEj/020xUgx089EY+S0QCuH2v0pRInv5l3R
rNlV1Q3B9TVMiqEfEpVZ7noR62+IcoMKrTC2D5CwjhpZU6jhPHEqFoRQqw66c5HVHneMLDUO3drE
dVhwN1xrI7ES8hM1t8XJMKSWIIo9fxPBGjYKOG7yhLvz3Ziu3dTaGjcH2T8ZdMsF9VIsyOUOJvh2
zmPlK8PLnIN0kv0asL8L3JCU71T9i1bRjf+WcTWftGpL2yVPxWrfmzxVG18kVUIb5ACXffdkxar3
mtwKywObL+HTcGPPc7JqKJrzYt6YplxNQuuqEDjVQ4YHsEWb0lqotGRcV3xEKHchkAiQzQY/YAIk
WCw6Lc2bBdalJA/eVIIXblujaADhD9cpPrumQVRgb7aajoJKSdcRvZyZ2ypzbFdmnspZhP3xigzp
Gc8/CVqHZqobshDprz85D5EoABojN8Ip9cwvhKijuHooNBQ0x29j9fJ3RqUafL2g3BHqscnQrNyh
NrV1ORKAzdj9VLdYqyO+tjhF/WXxCad8AlbEVDuyQVCXZ+CxswPYUAcRRs1cCff63ZKtGYiSlWWp
yro1AXYN+Fcl2iqjIj7UYDF1bNa9SXCzUu6dqfwuk37zQk30u35cgGEJKoyK26FHXUZd5si4SAQx
xGXshFaKWY13843r+58vejf/NJhdPawnCzIxZih+jWjK7+fYQvznBA6TCq2p4+rzempNiGPOP0Uy
mrPTlx7z7H9huw1uicXPq48Drh3L3ZW+anY7ONhHl7BqduCjU9Zs8f//Fmecp+4T6Ai7EYrNnnrR
RKvATw+aRi95vW65IDfTKGem9BVHeBKgtp985x9pBNnCHX7JwZmll+/1ZPkzoSnGobjHpZ02xn03
nTkCB+a+d4MB1wcj9goWlS2VhMbp/Nb+ywLH7WEKqsW0ARfiKE/nvRfzn7HeUyvzmQ0OZAA3HhnE
PCAVtB4X6XPJRVnOtHMOMn5uZdVwGOzBF0XiL2idHTi33uMzpQZhHA/x98QbNCCoiT/zq8xCS4DF
nL8Vp5+CDeiVFZOHaO74ibZHIAZ8CKeCSo3v7ZQNallhiDVB9MX7iuOYSW8e2vnLnK3SNerlFdyi
NBTkLjGAIM3EJQaOYRNfqsrR5fx44a8KfvYg3TmWwI8x1SA8CNvkP8gX3LXEz/355zsnSrK0x6pA
sNJMQXJ3Zbk1sDwPpc5+sDbxrenmnd3+4ZnEqbstkOS1bPx0J2L+E4xrf7m36XnYI5/+wCasKBjr
YUcWoGOFm2AVJas+/X5cmdNgpoSC7sjk91uPa6w+Gxc4/YcvpC3Vg8CYuBGyj9eEVIQbhch135E+
LOgn5cl1lCK1UZ7rOPq2Xjvwmlv6b1mRx1im76lvKjQ1wBvPOTTBgU8JodpiW5CpCAz26JZ7sL9v
2ii5uWg+1A1itzxNW+1pRpdniqY0We2wAf86hieB89bu1iLoROEhjH9T5dY0IYxMaqz56XBoEcdH
8Hu4FQKOPbMXjvWyuDuA4ixa8bBTsw6nSHGAMObN321/gV+Ja3gbi5TxRafErqdh7L5+5Ht2Zath
u/DktmjQWK3iGugFcuWb0/tkkZiOpBd8pJGsPJvd0q9Rjs2vTtrSriEPfNYEW2BaT3tSmSjWKqVA
apxtSxppamJFGN21/sPD4YK16/vG9A+Apb82t/r2Pi1XTIyNIUJVt6Apn1QiJBGPrXgBe5YU/KVD
IZcmv1LNdHSbuZzqCFxHOBNfwLy3UNO+BXnSs2wx3DuLGXfZ2k9TCOGeahizITIbgA+aFB9yeFwp
FSHNWniux0I0O0b6zHtHcTIAi1/pxAwVS6V+SEHSSIU/FokYmarsVIOmYX71TuHU1xpgHZuHO2Cr
b8zXzAxHnZu/QmgLKJ02AUzkZVcbe8O5jBrrmcQxQVu1Wzh/cqhz/50q9pnae5n57xJHDeGeqAxg
joMM5L30kRGJha2adlLcRAMUyiye0UH0jeHJAbwY9CDvBXKJAsCgtHrJOXeTMMj808CC6GeSTrVA
+wBzIVhmZAuQbmobiHlhwFG7NH7OtfqTtHPiZcq71N1/L3HoyABLCd/HU4HuyMct7lEXqmE07GDf
w92NFG/2N+xzuOA+/OwSmFjZwgDq/NLYHS9FpcM4r21Bk9X/oS6OFbDqbndzZBr+mxgVqa7I49Io
W29oKnqfuAG4ct8uB7g6niV8ZhBGQO0X8GbkEpy+8bQDJOUAHDlwrIS4Wno2HdWJhUO9tuNzkq3s
Prc0ST/DiTzxQZdjUX0NL1zQ0yDVZckebtgW3bRoy8c4zckEsm98Vk/g6RUrd+oOZWyvG8IZhBhs
4wGRFfaLZ0clpFrJN5N4FsuISYjxw51oHpTCqDcdMEJHnQHOTHs0fHfXBauvIZdOAv0ddY7iz2Xs
64pT474JNYJtr/tIqjhLjFNejaBz1J+zKv5KFv9oRFj++KBwcBLHICa5hHShWj+p3CmAwgLiS21f
ahjDsctIgbw0tPmiQq7G7djQbcIHCTIena00NH9aH8fCQLlcHBs2rhjEYkh+QhPYexOdKWIpgfXW
zEH4AHp89HsXf9+7zXBENvnwswkyOwBhoKnpKXopU+/asIsCSlMztGKwDoknH8lsOhYSw/iFbyqu
Jcbz8U3peYz0ntf/+KCU8KreDyrjrnEK1ehxDTYObHUVmUlr5HoKIa4QLPQiZOdscKV7pZrDDAyn
lThyixZ3kTSa68SA9fW6Dco1M+VaTnocpp5e3gWMi9v6xarQq83RjuLHwxjXSogDfkYhuBdDAvbm
cbpkrRPUd9SzGxokcA35KkwOBwq/XsrWJ99XsbHJi7J0dPAXSIWq2wNNfjiiA6U4c7k4dCZeXkow
xjB4zyVDhjEzo7IU4kPnP/PowOQqtNWnTgsvyA2/Ndn21JyknN5P/IVTQwdaJKRAaght66Mn84rO
+LUgoUlpKHXiELiWvNELitCemN1+n9mQI23ren3HLDttDeZ4zBeG8Oz/JSg3PanOYhl4tS9JDBz3
ju4drrSmp3oPmA7sQ/xP3B4mp2X8n+2d5woqTnexuKO0Z70MFeDJs3vSyWaEjMqiqS7coS2o2tNn
CArjjBVEeClO4F9vNdVPiDdP9aZhO2sNXSei06hbcQIkbTa25V17q8f2GGr672km9JaSUPrY7zcb
rFru3JQprTXTlWvF83PdFZjuVWxtTY9S3LaFPaNdnSIGQUU+PxoZKqQg71xq+mK56p2DqNwVNGEK
r327mdzLxLgrP+o8YYbDuo1bkK7MJ9y2NEDY82gALU/bCnuS+t/ksxAwPAjQC4uhaN1XaStUld52
Yj/ubOu9Tj4FIltkPs7i0hD0k1BIjFhIh6lwXzinbhoNJsHcIrMjuxsjEPKc33rGaf4uF9eEacq9
t4h2pk5nJU+3Fq00dRiFTQVb/Me7EOJh9FaDztSjWggdz1Gs/kHsIB4Vok/0Un5MxjwaaBqF61bw
SoRKmme1/yRpmIL6GKFa9KaJo1ulCUqwyN74mDshhmBimmFLNswpojJzIqKnKymMOhSfZmgJh/Za
txTqiEUu+S+NwcyNc1l+cL8zfiY4hEZUFr8ZPy0edOVdL5PsFPwzbLovYpBUvB65SnTLGVUuFS7Z
VvdBUnZP/1tgHu30dDPyQkQg/lBCMJ87IS8HYJbQGccnkXmk/2wt5QPvQ++7qACfxK90TWhGCb+j
qjHFqp6ILqhstVbOj38RkE8e8XpGjS2kh61dHKsKCt+aAPenLAIxHp7oDXo9nAQ8oefwwNhJEe9K
Dwt5WjMgx7qzWkmZQJQNsdTaLAiciMf4YfDT0F/7llhVC9tW1y/BMH9+x44CyXMpQ/o7g3DG7YuY
bk3faC+ACS9eGyZfUqBrlF1hvsMFQPHACeB6P53FTGHMSKHw/kmKCsZu3Z5uTTY0McMDancYdnN7
ic5EFeIwPQIJTNeFrZNTRgzT4oeIWacWFtHmYK+/BFi7LBqJ2jGcT3wW5wn/bCxl2RfYzcnAO5kG
Hw5kjSSVgMPhb6rmzzg6YLzTrIbbAQ1fBH5lLfBhtbOQ6rBRkLQTHAN6ze3OZqmHDJELF2iNJ/Hi
TdYo/kFP4wrzCeQb6j0IXPUQNtxvTXxZ8eG3QGJ3CatRA+UrQK68mVd6jTETv3O+JpLztqWdn2Xl
bFBDUGTxZ5fevqo2v+2rEI5uqTe6lODStGRUABXAxmah9TIbbX40Sq0ZGvMsV40ig5C997aeD/X2
L5hZy9PiiuIfgfKg+Wzn022QroUFW0eIrz7G/G2F/K9jMwD+6BEBTj5iYUXXRthVv9LL6lRupIFM
4lKEprFoSbo66hYI/oEqZged+9HxM3sGrDtb+oiyJbQWmpzDqnwMeXcQgS5ZchBtiayY2zZxseeI
4cmOC5U06O2zUmSzcW1Bfpz+NKeRtKgE2ycc7iCw8SS65X3dcK5nv8szicj3IraIbHEJqgjb3+/d
vlRp0rpVrH2YVOPqLos6lpO+Eula3nslBx4LmjtONKkkCVl0/AYi5tt1ZIfm80Qj8nUh/thaNBf5
OPlhZrTF0w5zZcB1P/Aok86TUs99Wvp7dqtRmLV+WYlHjMgpk6cpifzmE42WrNe22BQ5Gas+70QH
RNR0DW/mgBaJr815ILb5rMpVSdJcHzXv3JIPCHNTwcMcxfmk8qa3oFe0zf0DanvaZdvd7D1rKuOm
XvBu+6emryoUTuDfqVjy1sR7yk7GoMfe/C7KSO5EAx5BxZOEnY/N4X3BGRhXXvtcdUwTC66faKtk
iIBUxFnJ/Mr6juBeDvaWr01j0ZyFy7bo1zioPgZd66MiFvrkkfZ7onSkD5prnRVrp6X+NAukYyg3
19Hi/w6iZ6ZhKzPDNl8NaO4cfQyQYenkbyjsNKTi3+L7u5F+MrmeLbeIHZ/6Pd4BrUl41LBa2hAb
/qk5Fvse+IiegbDLWX6VrR9e1IbPqvLACNsO9NyT2AB25KCkAHN910bfJLCzGJBGbjQHr6I6KLbf
ZhN/bhE1k4Va+g6Xeb442x00CeBW91Y0lsu84QP1IR16OtnYBfSCItUMZ+y8NeEpH8JJ8iny0hno
rf1yQVzX0KAgk3K4UjF/Tk2hJhZctiGy5aVnoeosULCEuXaDYer9rr2OlkYhDMOoV6mte9XH29bm
s7n9x7hioBbvpegYzOUY3AA1CYy86ZiqOWl4D+g4Wv7zRBZf3zNDZ7kOV6q6r5d9ysmU+cZTtMkf
jPP/dhKO99Rihsxn4mFLxakFvHEVUUhcm2Z+BGQW9dGyulBrubmnA4PNBjdCwECM40+cuPFQ9VBQ
XyK9hQfbVYTABV+nchNTHd77+Z/lKu9qT0sb0B0AdxGpoGYpKgfmFrulEqSp15YQkYyZF04t3uLo
3WLOccNeLduPeCdzPISAWoLCX1aY2Ggt0C7Natxp3craWgKMMJZ0BfK2gfXQoWhbtjO6GRswk196
tNb4e0JBS9TqKHwvIKUDKMc4+Lmxcsrn2i4b/5ZPxMZV8cecBMe9AabR2QDy+XC2zBWwAYvV9b0Y
tl4hzXl4tf5KUo8MDQBvDOSjcJXNbU+46KJolFY0SOwKY/4rLCyfDCVYFT/nAMEuhtetLlKZGA3h
lp9HXiVBpe3LBO49bV/QLbGmN2ysDKS6kp1g9xLwwx7jymLZnIFsj2cmwP5jiPiyyzS8HcSG8DhH
CE0uL4QeQLJ8hF8k6nZawG4v7PM67o47j1QzwmgZjnOlpEXMKl8FubAax1MdNNjHNDKRozXBWBWd
EOLhrn25OIsKWrjssTkg+Y9xDpaAcj9Ex5Sh2mvurFla7c+/Sg7F2rP1lhE0Qr3PPTkzp0Vld6Gq
KRiJY/fx+EQQRyfz6NJxYBvyPgnw2w1QVP2YgEXSvgcW31hJBY0l+C+KLsKTuYB0/PW7+GYyKNnY
mqQ1RluUTtyrJUUk06H2dLHzT53M3KwnlVpN3bHjuUR1iGWOJn0mA9IJ5XB638g9ZM5x6FTe3qCy
n4gRc4u16YoX11A3BV0ukDk91iTPElM/zx5BhtxJctHhLxpwSw4evysWdDOOd6le64GkxlHbk4dk
dq5pFZzaMBcp0JOV5guLXG2TpUgy42eS2ybkTcMWeq0v/Mef/BgV1QfE/ZeUMYDzrgO21icRck+r
6VH2wlnsV/hc+LZfSXjYIdaW4pxN7CAik0Qo/0Vdxw1v8udShnJshFlt429QL/LBaXmONK+Cfc74
aYvVYKs4IvqAOb6lNpJ1IY7rN9/DOcESvVqKsPsdBCOHpYKPZJ/I2fu79jIwofwsJBID45w1HU/A
/shLXfKI3n1rfBnFjXPEt2ku5cJ/Flgick4otzV/Az7QuYQ1LJzUj0BZ6dno4QLX3vp3MbtIieHN
4UR+fjinXUJ8QlS+rlMRwqrgK9qc8Yw8g5FwpNVrQb6uRQP86MBJ+XRL/zu8YgcUJTBM+G49Pfyj
p4tMtf0/UcOp87fWTV+pqeMjjqqizA7yxSqpMvuur1nnRLM60TYKpO28r2FqT3KJ00nQ9BspZ8F+
6cOMMlOruU/tC3bC7CqiADbv6Hi66OijATWR8vUh+Z77cvIwi2cDcLRXfkNcVlCD18KGStzW8R2c
zpOQ4kXasKzQDfX18qMPkNrc4pIbwnRUVMzE85p452SdPT5god+GuozPuMEq+SE+umWh30wMY2YA
mENVENpkqrqyJaY6V4H/c8H+d4r06/myDwz7Ej0YAt0PCehDQKST1tFXB8aYTu3jjpInJjUpmTgc
muElc2DoLxTHTdR2oT3xqGyY1DbesZqBfROtsAqxakD3tXixWuMGguUj2St9zoE6+sGpuYGw1DiN
7EWS30ir1WCxk1gTaeLFeLoaU1NGUgH9BpJ31ElHnrcpB49JLga8TGZqzv9xsLUAQM8LBVkAbYfk
jhm/jww06KoF7YC6OmIJ6BAjU28xud/5JDRkbeGyMOwQfVn2LsOs5043FMeE/L+KNU+bzfsenb+c
9ZgOUwK8uykZ0FkVw+MRR/ImZW2NKuAudSGXZ+XaYh9AzoPDPwX2GAtRKI8EduKAgdvSVquhV1vV
ihYa1mm7spuh/7d0LC5W1cf+MS4mv2PRhFru4WY5CGSnxHBl6XMyhx4TUwCYbqYDVZXU0sfEvf+M
dI8EvEb9JRSc4t6TSeFaEIQJTJADzk5WVYhcWiMgoOXeaK0Mnx8YFSI58ioCJfrSQoGYgIfhHakX
SlqKspIoRbeVdoxzTwcNJePuxp32cSdMJZ0V2GPQArfV5O6f+1j9oOfKBM/mtVe53ZTdB0uebfng
t7+yfz1xIpeMtrMuo6WLhDM58ivghz/dYo5FnlJ1bvfy9HWCp0rKeBK21/6OXWL8CGbwqh24QKQ/
YrHfXYHWDq1+RSak8gbs5W/+otkOcIa3Ze1vupo+TzZKoU9aifzKlrWvA0Q4bvqe5X1GpK6/grqg
mny9Cq5OdBsHNzBm9nDO740oPG5MdINPjYzGwmOxcEKybYhJ6FxLEtwme0Ih9b9oNy+OpZQ+0F8+
mDXgu44=
`protect end_protected
