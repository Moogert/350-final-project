-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ji4nx9VOZTi+U4g8LtJmrwMQ9ii5jHGnETJvjQpdVkihmf0aO5AKfv/eHNVHanRjKjZRjpPIDC+M
TrwqtLDb9YnM5z2+mob78bbWUE71hGbZx2f9B4xbtqImlaWguD637N/ZsfzgPNgrs+URNs3UUhyg
jXw0/dJ7ucJnwDzRstEgAdiAREfGxfHdKM/fQDD+x7ktP/REKAtiJx7V2xGfl4Ylrem6aYiSPBQ9
r0cpgKJksGBAVICr1rJS+d6cPy2N6j6Gs84LJw4xkAs9Iryh6t1Z6BGRQ6R+qntY7sBWP1TqwGJ7
7PEwgCUnRK/aSkPRDm1bXLtfYJe6vJ6ZNbtS3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
LQewsZ48u0lerc4BqnNLo15IzPyh7GqcqtGBYmT/QElwApnvt4hTWrmqAGmqq4LfC0uXVLOX/Rif
SLoe2ubjqBkZrpOumhbNt7cjSwyUCokto2kvba5N1pn+FSgpMtQ/+nWjF/29XIdx7lL1SINHUdO6
ufUzSnUFXZIjVqd6NNH6/AFaT8NdVSud4F+PYPkvsqb1krOqzmVTVs69oELFGKJQRPdEUfHWz8Rm
vnvA7v8ooaxsWf4wVTbpPFcx4Q9PpOZ6G4mEnN0t7Caee4a1ZCSNqUZMIWyINhaQkZ/edMg+i907
ipm37/eD9sfN9/qPpIaDXyr/96Y8Gk+4/PhUZdfXXSHrTtirzEVJyRju7LhbZZGNjRS3uG9yLjWx
lg56tiuO+RdbE3XXyNqyyXJLLZ0qngCvKx6gF4d206Gu3XY5jnRmiuNJ15RMsJFX11ai9HDqVqFL
RWoGv2KgTqQ2Bmp1L8Ip/7vAWTO8IqsTtZt/3nqIF/F1n3Ik8tzX6PCDYjbq/oK45WG4GU0r1JWt
H7fgLXj8Dh1U8gjLm0SFYGht1/ToBtPBmlcD4L+Tc8myJLCRxhEScz3uSIJztLvfvP+rxqeNcYRf
DU4ohL2dB/+8Afq4x6uHj4AV6DPCrgVFAxHhzQXrLSnIQBLS4gcJSogm5kLksfMQOMsa21/AKpS+
b09kl/Pi6hg8WCxXPhHli9cK8RUQ7Faj411/sPYWp84+BybPAVZ/GzXEx3fGiiyVLhH+wvkSwdQn
LOA0DOMRsxGR59kIorxyL8CIm0Egt6JPjKdO/BK9zolQ5/KXZnUYNIqlz+0wUrn2QEWItLJze3pK
xt5UU7o7JIE19bLQf/cg080UzUX4r1D+OgHGLVz08ZIbkW56iBKp+yv0XSheFmNB6kgp3G3CEjh2
ZJfhX+61ib8sUdGJ1kyBVR6f2H94VAp3Vj9Iiovfy+l8Ts/rpy8FM9Y3tI2BQoEcr8ThLBS95FSX
KDQSBiRmzg6Yth7V8Bt21VL2HnK90zlQZjBUVEZ/weFCHlhvit2Xwi0OLZf8M2KtA+ejQJ4iSquu
6MVumfnTh91U3HKkNkKzXvi/nQ9OylaDOIOJIbyrUmzA2lX2CH0yLRksUayvuH+MlK+RCVoz0srN
GscSwRmzQ2MDUXdCwGLgkrz5wK51v0Dtoaa0lkcA9QWCebNjMt3FnDmjJ0al/k3466/G01kgZcnB
mqjMNdtIMgqvgg4eJ9Z72g9UtSLkOXwaCSu6Bhskqt51gOE9EFdTwtPenjhQaAQLr0lnLNQsQvR5
AMfmdTtEele/pcPUXr/qY6+Sw2g8gyb2giRXmtObdmdhbci/DNAiBlGDVoBCxGl+aLQmACUGZnuz
DdjevYSAoBSYzRhw0KDfdvaqp6Bf3X/pV77dql/Z/kVfXEGmSHQU3eUwQ6bhhQqwpP4VkaOtiOBu
tdm/NxQerPV7oZbPPYi/G/R3be5Xp092+TBbBGXRkFpKSyvSTGb3/WmtIa1ns0+eO8Dy+JeiaDp8
4R0khMnvkR8o6ATpssbf/I24lWb4P9I9m6513xYK7RLXcewbiqFnp/tYdPd9bK5RBO8DhSSf5CL7
h3N0UXBA4/Zw6HdCVX77iRTsRT/ql9aLn/FlMRGErsgov5b5u6pCtUc9vWQjkqrfrHy98mPBDOab
cDMMgsgTNBpep2lwdRiXDjAp3j+CJ4MNDarIl69hqfQ4mAGH3ymPpA6cUZ4+GXNS0/jZo6ny7FuW
T3tMbHYZcNTaaeYNvamRbvxKL1l25wMplaREyrRMANdd8Hkq53qYhN8KNd9Ss9GxsOBOyj/ZLmNH
mispWAmQUv2O9DbWz2FycrDivLZqTMEYxo3l9yf5GZmCSMk6eJ8jXf6AxDJBUVtX6ipknWbktvK/
D2mu9X/sKC6Zdr5zTLoeQcUdDoE3Cgt8NThyy5wn4zBAWoXfgPRrs7XrcRxsLnB3TF1HjQuPy3iL
qRRB3g7Aos0sATP3uPD5ArANYVAA/L6cWfrTerzc+/AKuhm4S61ntt9PI2+KAK32TyfobEhrFwpM
zLo6yEWhFC9utjSNYzfWbOqvw+Zw/ny7D6lWJbG0gaPeyoSzEH9seeCmYz2fVVnlbhllNOMxzjZp
GHzXL3xLrNeXGcNvt93PLq87IIZ6uCEaICHBO7HWWP+lyTsSnjp2djyUyGIN9kl0aTC8v9T8lln3
p9xdpVr7F1Hh/QhyP+xm/URX0H347zUM7gCD2bAs0Ml8vL12+93wMwWvZP19ce1uqCijUjU+wKZn
eZAY3spgjDDMz2HnWJZKVvuY8Ze+zCjBXEInzty7Xzh/Oygs0I45z9oBHTikrCRNlLUd2wx4Yk6a
C+rdK7/luAAOEPnvoEkYGDwgmUrvSmZ7cAnq465Gj4aUhxJaKMZTmHNkIZPAH290rVdDMY86pA+2
HQ9eKj3KYYgHRvCTDCG1awhE2ADjviFW9xKzlD7YLlT+y1Fhf783AAl5YgmRk9dxnnWGkhWMn8Li
tvYpj3a+2kqYXq1Q7jCfUf39ehW5ZwMF0cDGIPOiyt1mvr8cFYOcbvpThfNRqAYsaEE1QUWAUuOa
5Eb/O9gdRC132yVA1gtyd92ULEPjAJSuWbFbS4IWEieopyyIDwOk2uzn/meN8jvAvJhHRifgwFG+
ta5BxSltRS7qyZIPv6zZ12IlW4kgung07gVT7WiHhpsVYsD0gL9QaqCS9GbBEVtTmXzHqq+ZYitB
DEoHw3F+mPo8dUET/OiAQWVIMqRmicLY4WqwKNd5WZn66kRA2v0veTdgDnQQ5hkjDkEIuiYjFRpu
gddn6yZ97Dw3U0H+0CHSvmsLxSvhaVDL+OPlMKyXKJQKrgtD8mmlNEOmdUsevLB6V7uwclopPxfY
k/syFLjgzVD9G0luTCj554uKKba/3ZpKWrUzOxwV7DVeCXAElW13eB93fMDGp0tCRn3roPt4vtol
3nSER8CoKl0hzMKldgpI5xKc5GINKI1MMbxl4Y5LPXC9g+Kfr3iflqAi8IPw2r4lS4J4enPfB7kH
AEPJWZ1u/KZygQO/j1wefYEGx8VAOOiGkxcMeXPWCD1wsGO5ZRPhYVq50Wu6B+oEZs2yTs2lBH8C
k3dOsQUZZyoGi3I8PncnT2xgAitASdlop9AL1fOH5Qh5RDewtqLwXuBkhTr0N2+Y9k5HQSc17Xmu
jsDwxb8l7i5jnQQ7IbKzLbk980L1gM7TX1ZxIpuSY481MJCzCrjmoHbzCWd1wVY8p3CP0Uo0R2gq
9dXN+A05yBxlu3RVrqRU0EitsvOrBbYt0ThsjZfHbfoQFucAEAgS8QGrfY65rJHssYNda1qmjqfs
SAgPcj/KetEtzZQEBwuMpRwW6FCH5xf8qfQyv4JttMPEj4g3AHabGlNTdC42JcQOCndwinEH8/tR
s2z6WQeqniv1i3dnLLdNsHGA/G+icUCgmKIkDbJ8RdOn8ooDbcLEIkT3Uz4Y4EWzxRky123ypK3K
OPKZA32gXNRa43w7HH6tuvBPPT6OTdHZFmEdxrahbiopMS6anU3ieKABy7HH84FMW/Oei7awL5YW
5rVofGR2KaVyGUIynxA8GDQ3xaX5Bcoy6wXHusgJgV5yHMRg5DESbO3GIk8wCl1vu2tOnl/jRhCU
rYtrEND29tnlZBxfYGblZG4AyNOTSPz0/O165pSswqnBXNoxal79uYkgBreBAR1a8cTBuJA5eEEt
jZAHE/xanE4pa79wO5/YvDhyZa/gSuRJup1WQHPRzp+ZsPlvlLp0X4kXuhIbgubBgVJqD3Ghma/Y
hc5sqaSmAPiGbReZypAQD2vRG2te4fKuS4U26Co0q5g+KXl3pQ5TWiISQj/GCvpevwQp/mJrP1j5
Neka1/YsK3TaYMSoHQ42zgqvA69/oq+8nx+VO8xMWtKt3SMe5v6IFqWZJ8AEXnTz9/hHGISaaLKE
RbeE/C0fYLLmGiF5btQ5eC8Ty45T6C3YX6SoeK+rhfidBw1i1BEopNX2/TO3hWmUvuTbjhxbJI7n
w6v7qGWZfs9RQ4CIbcAbvtyRQozar8RrrOlDanZpkinofJKNmWXCH8SKJLzhEUrJ0naTKJ10G+NN
eXvsa1jK2PaqTp+AkyYuzx46czifuUtzt6CrUd4D0uabK4dhj3tlU9IUA7BrsOYcZFw8OATk5hVx
SPxAisDOj1D4Ok0y3XDr7yuZAu9sJjKrtbGupti4+2U78ifmttBbmO1fKTycOXdu2JYmMN5Mb5+8
VU8lYpzg3iBzKPqqBWkJnZoK55wiExQqMPrASpNbMgbeCyIM+OolpZbrVY7SF6220/tD8i3ZpILt
/BekJcN/Zs84uz2lQingbAq6q84o6aDXWmhGQfdbnVfYHmBqzDaruqkC8w9dEOFfhi5VFzbSQGIS
zcj+HJFW7FDV2d5FHOvJwZ6ahDyB+avpq+HH4BwDmDKynvn22awFjoKn3eMd9jNUIbxBX3jX34Ka
+EClp2KoD3RhkPYM3sKeGyi3U2EKhjH+gXeptsEC0803zEKXeK32eroRVYbmm6NosQHTqdbal2G0
2v5S7zGonR82n+FlhM9Za7CfW5rKkKCEIhjugbQZoDs7EhGOBbsSWORnJYvZavNB3ivr1qGKvLxI
uAvEUWVOytulJ3nVVrbZuIb19E4ZemmkgbGcNBAWsDJNpoWv/hNGlFx/S4YC3jKpoOfJmIlr4xEA
+xqKP9JdOkCIQlm+6zjyfp7y1zrQbQ16QD6ZCnyO/mL2CyHQKgYS+5K3/iNSgHuivKA8u/CxJul+
7dlergRomBzL4nFAyax1u39gkR3ntWOWWVMI5iu+DwmKwKwJfHYP53tnYoGUv7gwaYYlUNaShQaW
rIjkNW+nXoBCqRIrQmnJN9UXa8YqvYMI/85OQz8CwLBM5zAb3f92GTToysKjWTMY0F/MBFpbMwqF
at1e1hrKq98IHP/iGMxpcrYIEsA6lbaB+FpJOu9k6gQgiwZDFRg2Bk0UBYml3fnXop+h2YYsrncS
jcNnxWz+rhRjPeLcZExG1VYyJLV8Jb3r2YhWdz+wyuk6KK9HJekWMkgePcflgeH7iailKxxvwfv+
2fqNrsn6N/9QHq3bRAD3Kt67D5cYQJ+X9udkInvEspm/ZYbgt8y24Irh1bOL8hPnSNldfhdTGetP
RClHSmEDEhqVFJS/dRPFav08byeDClRzRUMw4ZEQAvfI++QheG7ODjEIMWZCba3cpBGITY2gdMhb
CwA7DknY3xE2e6EevgGSSB0CP2PJ/iOtgnOHrbjupfg4+2cdD4yaav6qu1RvAXheGtGgu4VOo1r7
Wlnmcght1ylxdNnLHCcjuJrnwXuEmD+ksUiIWLSjVzfpc+xhqG36v9U+OVRIOauNwFOw8gCuTHp4
3hBCvwsOJrEdOXlQUlluhS+4ayvgW98r1fXomMoPZuIOVgtdiLzfxTq+9672ODSC9vLVXxbw4FBc
FliJfNJlA0ZiCPySngCAe/y+IGJ6L5rvIapJhUUd64jxKPzxkBWVWVSac7/rqGDKuGrGZhxEDNo+
bteYqkqsM8x9GffS+xnZmRHtWBSwS2fi+CaiqIFnSb6wLIUe3L8oZs9pMroxbfknOZHL4cbv03h4
7IPJ155l892LvTqTZ58rRtFG4xNnxIQ2CzQLztzgPNPd4hSNSszwYdnkz4lU1v207zG0LAXVtB++
KKnyrTntT/CQ8VKQcVWtRO0dnRpqJO6HwRZJxr/mc7REPR4zh1yyydTs4plGTuf8VDz5ZbS4yLwz
RDHGB9H6PnzBqq/5uyVHyGKQIgDwCPVsXadKkEoGKAsQ6xllSC7+xMyC+jsRmIbtxw/mo5CmMUln
iFQDg9UJXfXj1eF8N+s34qX6hK3rYqF3TyS66ppr+vMaXrrZ2STJQKMiuxFlWbNRJBMYy3LfJ0Lb
cGB4LPkAdPvTacqiGzky67kifDzu1Z8x+j5omYUL5yWkM4GEzX5E645WFDnQoR32rTvBvNa1+0vX
NpJvRJi4NYBV6YPOvZ42zQb1676kDneZRBhwJg6Ci4P1n18KhvvtojTbeAZNOiyLSnOpeGoqrcgw
VtiEoh+2wnWCtHfyaive7E7EaFT7QW8E/6VN8Dy0MCRANysxuiG3Q0fLDx5Dm5dWgHrvXimIzS+l
I8dNmJBjGoTLKIDIH72KFaqFpnLKrTpo3zv4E/kA87NThS8aE3XUiTY9dbj33btSTGsX7hT7+Gy4
84sQIGp18MusEiDkoQNF0MYcKsPNpxmIu7a4WfZ4vTwRF498E2WLG4FDhPC45U/aWJAs6ewHq0/z
kET2J3R8G0rL0bbqXr0bAjRknNP57zQB7UhZ50TOJXYb1ZAL+JWXuRkwDdzlBBckaTETsak8qHr5
ajEQXU/l+VjlDasslUIfZdqnfkrG0zsSv+GxfC4lf+cQ360ar7w9gp4KDqd8qsIUkTLMKnPECRSo
8N0d3HuhBaz/2j3X51yNNQIxlFCmQmDD9EUuy3/EC6hPLzxBTfDGvjIiC/YEaHTyGmn6wpYF8obX
P1JfEo3XDOW1W/sZLY5N6qLEnNZFx8nKq5rMYhDq4eSb+Cqw4ffQvo88HH3YT2ujOKsJbaMYRiBx
Lr7N6OkXb7ikbx6+QaJlCZ1f5icbUoBkt/HEX6++VihAAtrTi6rbWqdMBw8fh4pI62ZxnurpUrh8
QC3vPV3YDHkd1JpmYRlKcs7VFVmm0aYvG7EgyhjvFWplfEgL2P23LKkN7DQeVxZS+LcqlxJnlpo2
Q8nAgabi21a+SKIUupNFAMWvug3eidBVKvo2G6M2k3xGpAQJsUwf2LRpV/rfjYOfQSZ2doTNKGIC
FLdSFod65B3l++fZNmwNeY3lYyWmLcdKsn1IMdB8p6ln+D5j8SQ90TCCVq6fsa3vGarSt1dFiEr7
qScDP64RHlSZwngiHbIME3ziaUo6pZ2u6L3Us4euOK72Hf8xcA6Y51UNolADNvHIY1c4TtYDVeXC
KPnYyMOiwMunP8v8uX8oPSa0M2cvCQHV/Bn4pUAeXIxS3SN7JiAiLePlWtd+WSsADOSBUl6PNmcw
gpEOq1j85kVULAfoMuCmJdEbd5XdmgiViqv723CadqfaS2znMnilEcaf7/lNtplrEibciHbp3scU
jC4n9/y2F9Qt9FY2ClMoEB3exoZH1zpAVsRLBtXAD0cXuyDuPFwtE22Puz3aAPS7XY/Yd0GknXIB
KwmgoKMzGqYPTXYsrCxTXeVGuhz1FkejDtH51KTdD04Qq7fcmkNPxB4r0CLZ2dFWXqAKLd0Rn20B
ykFibsDriNJFz/J+PeagWBLV7W50dOHpN0PIkHmrLsMKUaNb99fLQ2CCn6Kx3f8gihNnmLmWY22w
S8uACp/HmQEPppoVr0+CcY1sso98oMJl28tgzhTPSvlth8WNZHcEQL3BHXXTgTLnw6s7O81NyuXo
MXLS31I9ZgBBXkvKH+Q/PbMe8WDil1UW9jJ4XpeSQX7mPbhrhXnrjDlNjxyAH/nwoWDOPaokyXhZ
LEFds2Ou2DDGxzx2PP6vrEXaPGF0lNpBwnebfvHjhZ07ypUzGQ1InhoMrpek1AENlge7AfR4D0AX
XmQ8mlFH8OjH9Jm6eMXrAd4zebDSuGXv46vR3Ia8BJ3DH2tC80Zj+IWjc4G6uKGPfAU+UY1VDGHy
ggVcIFdCMl/8/zcMBlsYZlekKyKJhVpoeOXNJCW3FLmKGde1ZpERU+B+NucWR7KHxjU/NioiNv0S
zB7XUookx2m/Mg==
`protect end_protected
