-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UEpMMzALaykER8D7bTqE5B45EOIdUY08BplS0xhlkA81nb73eUQUdnDrFPLNnlYaj96Hii7n4ufH
xGAtsgN/Ep/28UywEqGl0o8U/qP1u8TcH8ZS6O9fAPW2hO+7kDhYPsGeGI0/hwNoEvAhQ0lzBpnS
AR/W3QYQTWDo5CINa3Dl+RY77pF/inu9e0lSVxWybax3g8wtoTIunliuosZNJPAa1cRs0AAqo/zu
+HCF0PVPbbi2rWSTAob11gkhV4DfwUpDoGb3GDZJI4hUHp3796KHd41tZ4x8WN0eNC5dKhPIK1Ze
I292PjhMgKdGTWB5XEKbhlTCPEkNQ46R/gyygg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
xZ+8H6OMoqiDhMcGA4/yQfhxSRXYFCjhrFKjXFByM+pR4c9i4pq4F++q1Rcj5vekh+6cx5K+ykY2
MaUwomcQDFixbl+a+0P3jXltzfFuWletd6v4qur6FCfMmVEcgdqXwEkh1v8kuP8DuG1Mky7VouBA
dQgTPc01zsGRgCO4LSUDVkSfcOmQQI+b39rufNN5eIxFbfTGvKFPsNcZhkLRbbNvIosNuobhRo1s
idF8Y9G2amdtdVv+TRYN99A0K5OMGEIirb4qQSi+WWer8r98UChQwY8GMOP5A71BwjY1QDq+LtnA
PbhNI8NFvr5dI+mG/TELXvtIqfl7ugVLt84nYIFsySdDDBcakTMJIzySBf0nMXT7ha5Q5iO004fg
SwzzsiTHf05tIMBT9yl/mDllD05y1Vsi1/an4b9VjsRAKp3ySa8bpER8BaYppZ1Efq4Dncmer1Wv
Gtmv1UBjKNAvfFhK0QvCnh6RkMPeALenUB8dEZs9uFE5FCKp+WHgTNPj7E7QFSXLoKpKN1IPD0YZ
rijXBEzmAqh7g4onf0v7I44D1RaQx8N9vqq+x2Tj1yzpJ2npayV4xgHwn/MiHN38JarjfIV2YBrq
tsyW7CigQm2mLf2DmWPWQRUyOycsv4TOxWXGMjj5DZjiG7Ew9jzHdagiPZQfCZw5zdgIVGAXIONP
eJYEHtsQ3lsgdtl1QsIDGbQ73W/QUssOGTVLjH6J57CXIQWaoNx8vQ718jGw0sqxooIWDqhMfMmO
h/2WdmXy2iO/bj+KA9T5l9zyKjb3XRHjmWKTP+QpnRIwMQaiEFYyOrhv6E+0gimBkc7hzb74Z7Ot
lo6u5TIonPx6HRYzw+WiCGpvguUcDKYTsFCDoDZ7OjkBoCaZCw4tF3AQl/BJT1fSq/+zzZARD6FA
HoqHg2h+vjwaTvuXwOBkaN+yIjPTthOnigMCDNtUD85vRa+7hQiyiZnftE9O6OllmxpvaqfU1TtO
aDf7euixHdiueV1qQ3bTTTuva71xK8rp915Cas2qOGbETHg4+kmNGkd9/fzOXSzXwbK4cm2yt65s
NrsEQMDrTBc1v4JRi6tEMTqUN2eHVG1PnonAqRsYkIU8LcI0BWOqP1al4F0Ieu4QM5QNYod+2cs2
N9JbzBwuw1SIfIR/Ok3U0vclp+m2qAXO/tVpaUXIJLr/W3m5ZdI48JKpDZqymTfWSHr9wUGcKx8T
6xZAwQeXo+H5orYDfQjoLnaqQ3p1ot+KCNEGRfMKOfSLo6ng8P/v5QgQd55vybD8GbuGtv2O4lFU
a3IRCD08yT7iEvt/nEU15f22nZxMoU7RvKoljODDc5S4TtUInjlN69ix6jFV8oPrABjozpnH6cjF
bozE4e0VQtqPNZJAqdVyEUC4+J1VqrDH4tvdTaak7h6jQJrCXNnQpuqo/HAOd1MUUiiiwlLcbgT1
QyYSFRdu6mICdTf2CYmyRfNIpOf9jfRxfqKpJCAXUX8y0e3bnpVLbse7zEX3KafZ0ZmDuxDKJ9YP
6FrlMg57md3o7c0EqAS+sab6wKVoduITWiKvEMiLDHm1LBDu/r8491IoSvZklm+G4t7Tvc7SALDw
NeppqGF4eHJdArZhwYLhRWjE8u1HExwsIoG0DrxkloTnXJw0afXwXKtYA/aT5IWIiL3Wb0/SoUi+
DQBwNq1DJJOTSPtlxhPrRY8+NmtC40zymudDodyXdql7U4algXVuCDI07l6DTg8tzvO7fhKWOHYC
fTy50YfYpd91PJi3BOLgzeTLXaOxgDa8g1c2iPX6rkp58M7zVi5hsEBDv9hhl8OIZ41heE4PMf9A
W+MHoGhJGyFWGCTG0W1HYa6+z/iCzfNoYCi4wrD0BXd6e9Ugi9L1W6kTOrW06jxQhnqZjY8GX/Ob
k7OF0sXOTOBT/KczQVt2ZM4G7ucg/4/QTq4vq2nxcXKvHq41c9PDUgcyUJhpjTYVmFX4XOwatJOi
u2lNPFR1OUJoEUyH4k3zUb791KQCQAAv3lnw0fjE9MmxxBuZ1pQVaHo8DZRw6wpS+ghHbQC3TRuI
X3KU0yA2MxHLBwfSNQDlHUYOY31g6hHcr1wE9T6vnhLzUw+zkYn+/Y9PS4KCA5QpqwAqGIZpK/4E
btmkelom/xy+/yKylsJ8oHklmd1jjVnSvsTkrzwSpmQMYkosPaZCqaFEkuv27Ibn3p4E8JFKgmAq
v5TQ4Ly1m3SWH6kGl2d34O8mRKlnREREEzJBP4EDMewr9rE6xMLMbOa37/ginzQi1U0R4XGV/Kls
Tsk+eBS4Bhr4CZ02rrny3+2ucTp5hPwKJeBaHq+SPwlkUyp8LiUCy3mj/JNmxSxoPZU/XvzyiaMR
wLfy6OuXQ0D4R77Clk1qCti4lsgcZ/+jY6m7rw0kI3lTWFt+K6PeBRfibi3X1S/Bfqej20vLnT88
VAys1vznsZqYaZTfOxkS1oKerftormNyZUL3FXbnFTJ91CBbmQgQM3A3SZWAsSi5iPkZWhBPhelg
/e+wbv1u3/nQu8CAsfF3ZLC05tDV+bsVKJru6CrFiit9FvZVkgAqd7RbU0LTByn2RwXCAadDruuR
Gq9eMn7PlgJqSb9vnvo+DwsRa9F4GmLobMN35nProsz46VRAt5InVmIh42Mhp7GX0cWJjjZu/0pA
tCF+QhaSFCatW8m8de2x0L0dp7VgMAKydPxUKX+X6RlUpdW5aI3mWmH8d61tl7LHjDNUeD0CtR9B
Ol6h9ohAAJ1MEnQh5ZDrdNiu5Kw6QZXUChQ4UTHm0OGXcKvfJFO3wH+NaOp+2nHWSBibPmuwQegq
vErzJXUmJ2I/GL0lATEofdOpLDjRbGKzCd9l+VAT49ctvtT57UGAkrPoEmBofcoATAV6nxWWDXrP
JiO/NKxSlSsSDt4/uOJil2L3xPUioif2Z4KPsEWdGLL05zwNux1wrW1kkSrLaCD1zf8YVi4KFWj/
ItV2kQPe6+OtGtdJj47wNqGJF8klsYCuMEhxjkLZDM52VddqHZlKQON54LUjDgnhgwY03FMkTqhP
RB0Yb/O+CNxw2QhW143K0HTln/tPSDjR1ymTHI1siUoIENzVUrqSu/Bu6vyrfr+oT33xW1zUEgF+
aztbm1brPYxpkWO1zv4BURZbSsQLG7gkogTBRgy7iXKBJfpc67Y5nVrvzia/1SQU/dTkLG2y8ty6
eXoMHAwsZ9EAKYoPmxlxv9tQ9yijOBsYOIybu9Y2cYfotdfOGN4QoGpoWpR9xPzHhVtJB5KV23b2
4GpZrgjdxXINuvahjOxFGKkX/y5mUp2nRo6jwgNotCODzCosE+rCSizX+d1Ffb86/CtFFtwS+a1A
ZPukthzeKZWHl2d5XpzYS9x4Mm31cM/NiFbe68BrFbG14C11lLmXsWlI9JcMv3+RE8qFH3Jpt2IN
y9PmtlgqaeV/5gnLK0TUN6gPqZRihvEbZCcZNCoeL8UWKIYIyawrvd7dUokAxlsX3Gs94H6ndnP/
hMhCayU+EbafghLq3fcsPZ4vxY3iBQnTPBcYRroSy1RsXaG6lYYpvks2PPtKkQd4oSqbiSqgtAM0
hwFDY+RBf3X8OEO88etwNrrC4Uwl0giQT1bspMrTiR0snTpNdnk7UBEhq5SqcRNRhlpMfZMpLF7d
yK6ICI1REZl3F8sxtO6NzrDF17fbsQDxko6aMrznOhCj1GRBgX/UpMwps/HGNM9GUhpVmqeWCKQ2
AOXuXfy4q2ijhj6WZCRTDpuO3h8OaTKQnsupL+uFZ13jUrboEoIhEOJjz0HgAVPPA0G7/SCgq8Gd
Q2vi7x89CCQQIotmWrvRyXCDrYNhGcLPp+rnqLJhjH7p6k5QjhiVsgDjzJviNlS3Q69cipIlenOD
p900QSy81/orPitlVZ8iTvjCVV2t2TSPKyWP87vP9uIk9O6eJZjc5twtvHU7YBeo/r4qJMybwXp0
MIKBXfLiUu9ewvh9pbCekA72llk0nRrff1W8U0uYlbEn/dk88XxEsDO2/uoeWbBSnRomt/8CHZdP
vGHO8bInobH2e7vWcVJ+B5IgD5X3yaWZTJ89nmiE37uTYsGQcwnmWtAK5LsiG1fHIdBN88Yil8Ow
pQ2cs5cfL82Xqnk+CQnqAgcIADPRsimaSr9OsZRIDKQ5WxJv43lvWy8gsDGm+nnRVCJJ204BX+Cf
DP6zReozM84aWXM9MilFeQ+jVHPPh+z1NjJn2j9EVRXV9SL6/F6mbD+r1agDW0uF4dkflnXTn25z
N0zofhsTIDE2CNArzrcbjHYi2L1AUzmweVpdXt5I7fI/MKbbpUQSuRbJxEuwao5cmYivevg3Is+Q
tRYFxa3a8yqnI6j9uSCka7EH1KQfBzVMWtsGQ3vlNsdelsaDqPCHtJOUqGk/FCWcPL7Yiz1r5X1m
RDTO2Pczbz86bYNvEHN111xVh+MNonMtEjtwz3U7mr9FQSNT43lT8XII5BO+YfI4OWc2hd9qRtXg
AYkUYl5tlUaZhOi5rfCrU2QvvcxIxqimcYhtTKii979NRRaFdxul16m7OwAE46QKIDUCOA+GslFo
rNccsWqKfMntoMD0evgmn8/SSju075tXiN3RoHjeMlRdf5Zcj7JtY4Wv9nzziGjzvlXHJ9tXpYps
FxfGUvzF4Io+VOTUwedKhjTGdKdFuMMaLknJItt8gMDW/NURhFyHwumw553j0ul6SsDr2sj3H+d1
3zuZmoYHe+DZMrs9k2UKfQ72UU9VEnDRUvnpi2aa1gqMEbCMRzJjyCSjeyrKmDKCehOgHJ5CQ8mr
4LbFnKw6lrdExhS4MopwyHbQDGOqOG+9Kcyjv4+12wPSyKP0nh6uG/7vVxBl0xKEeyVdeey3xQit
5CvMIWVoQd1o6Wt/XligyNwMUrKCo0y66+1RonZNDDDXDnxk6Jtm+Dg4NzavPL4JHHO32tbGd6rg
Zwse2mAIddsc/gDLBwsapSsVRhjeEqpV6fJC73EUW0ga/n2DAvRtCmVtBX7/ICOjDFnzuI7k8wbe
eweGYqNHyeaqDrvHPI9Cu8r4Ee12xBg31/kZvMrFyGRVt3IgLaDOSPDgnYjtZDGZju3MubDaYDon
8rBgpRDlpgxnaMdCZsmnVjOmtDu4M41X4L8Yb+lJyCU4ETzs6eXAW5IsmX90bCsKVxyrImMxcfKu
eHuo/mmOPTU73bHH1VFxtWyQtqlvhBnMS8svBlFsiwTRpOWTYDh7Pi0qHvYmHZTRQKYVSAsPGjET
EpQh5Qk544c2K2DLD5l+ozds/K3aKHKs0li6/umPYeW4XwPS2ZFcQHrFrlBLi80XTGXBJdKw1gzt
gwIR6NXUD8DDG0JAlq6vVO9q8G+Vhwsf5k6Qno7McemyP6agzhG4oCBfUhM5c+HVh7zGbtTmMZXj
jT7O69wyf9UWob6vhKOTXPERPg57OBYLIBM9MBBSmrea2YUgvhlmM7gBOSmkL9uXyBgX2IRlQsX3
Tt5EKrd97j/SsXeojz/MAzk8aUorr0dO2fM8bP9F6PHa5HbEVEaRpTaGzH1J/C9WyzLPm2yTFAsu
+iu7Bd18eBIFNQKtqzBYYCPtXEC5i9B0xXAXuy41V7FmYqngNTd0Yh1t7PaJL7ZhjpKu5VA+m75X
PAeY6zI54Fk+TI1wKzO56O6J7ZhHEuBfBcGULfRFw56g459aspzSOAKMKJaBCvNt3o6pGE14yw+0
xhuWI3Js483LQmPIgqctx4zc4aumViudNxNoiS+7H2OhVKxjH9pNXkZdzMmd91P+GQ59geOSrpUb
9R4NS11u9VggSkE9yQUXXxZLxL9yRyNeY+ZPI1ErjGHgMRBJiW70ZSfRaR42PWLQS2yhS5fQLRnD
oLv2kDB0UAIqtJsYTpcGP+nd4Tlk/g6IGkzFyCePRYWni1U9wNWGv6J6kw3Nctk+KEgF6xGJAwuY
5TMTMwltPc3irfCbNip5NiooiFabPKx3HEwRV6htdLRa/lt5sFFD0/I5kM4cuMsu7+AfgdOC91Zc
SZ73UcMqjvaUJe9NQQdwIx74Uf4Y/ScEA/GLYgLdb78tCAx6BvK3izmvwFCTguBW0CvZra0oV3HQ
5KFP7YIFUm5H6pziQnvYk8LeX0K7n4p0iF5WdQvSi5oM2ZyYh0PuzA/FuBJG2pBjGtaqO+UfyBhI
dGrUuz4zhE4kfSiPzIt/c7PU0vjiMsy30h0mXm/sUDpI/zOwmY4UqUJLJ35EZUpcKgMFBUiLc6nw
2B1IH1PvogFo37IXFqA4aSDgR9NE63ESxQCjvbg8xzhPpL6tPkfHT2k3kc+VL1dlunbZgE7y91z9
jq1yM+hdErNX0uG8YobGgTfcVlgYX6VKNmYElaBfxg1umuUyugCrmeVQvJSolIzn2C3rm24iEPFv
DjTy+d+Z8Q2IM7q2pf4c72CiGh2BliRCHg7+1RpUQ5UYp8/fjUsc7kEC43jz4MyGNHMFKce06p1I
RKHhnhWSHnDBVKnqQuN8pAz1IkpUAud82ZmFDedtJe5DWk9OM0CrtDFkj7Y8HBh45xN+otmUUJ8N
NFcDYhW2s7sXK80lB8m5XY6jyzKr+GTFJIetPslg2NWDgJDLbwTRKiP1gUVek+LvlaZ3WVh4wQtM
pZ0DXeJzhtwbkeb4j9YIOBOkadsl8WjGQGfogh7VHiqwHLLnUlWQc7uNr1OL6CvoKshoAotmNT+9
bdGnl2G1dUTCeXn+qHUozFBmCmbLk68Ts8XQ8KOFrKMOlGB4GqU2ETEB5QVpvX9341wwhyhZeuOA
7Jfk8eAeXvC1RMtvinCw8JAH3sxxL/+hZ6PR9TU7u4dNkcR854GiZpkoUeQa1YtHdv4G33ucHwNB
T/ZCI3Jtbe2o77KXyfiv5xKRWsvecMdZIcomiezMaD96W2Pn/CqEgvW6j0ID8nbbT96xny2E6OWy
zTecfip9YQtkKJKhPRWquFSCBB4sdtjgjYSHEk5jAr/1FaFSuzox+krGmz9YvUTDdrzFF2JW3Em3
sSkOlOIAOeManIAmSNYqFFJhVCCw/8jm+V+vRMIoWLJfgxcXmha0IUT3WXgBvOB4p3lajH/a1Wnt
hE0/ejJDquf6KyduyiwFD9DaD2o6EGJJ4jcli58fSBZhz18xZfbjAbNeMr9JxgAxTrxz5wbVkLKe
svamSR7EAvVmGSH0uA0dzQ4bx2u+Sb1Slzf691nVHw/AUt7RFaCZtNofxdDE9fsWJSzHQvA1i2dd
BlRTMvorNTVIJsC8DzErGk8h6wViMeTkLlQ+EtffpVcFsGJAU7Ie542Ghl8Rm6+n3uvz/2RDak86
u8QVQ5b9q0oCUzUS7MmarceSP2pJjjuOlAqHmBYmYbiOiL7L0y2wrOZpumJQuoX2C+NqrarKzbB8
3pQvlxoRq2i7Q8UuiH/PABEHHe9ehRSInCZGGM/Gawe0of9fLBBSJuN3kz6sevnjwEuK/5clCWu0
eoifHEfkdoBqIA/0mXYyL1VrMBAiwshnoJ/KfcWCpbUt9C+cIMG/xyS6oJe+EuiuQ9KU71CTQ9iF
D0vpOkGKltOky2opN7+azlrNr9Er3C1pE8QX0XR5//K6jJuJ+2kDsL8/MWGeg/ldJ6HueXnwehUc
DcqUtsMLVUXEPGTP7W8qMDm0x17jTdW9Ax1NXkJ3vdOuJ+z+Fe6Amq2DYwW2MapRDqFOu5ysWHJk
VgYHz2QoWiWYzUdeNoghARDa4fHKL5PVWcbHoj2+hPyhNULRscik1hA5g1QMCVvwoIR4ujagbWz6
ks/p5EoTiiX4s75ZFQZZF1/rXxB1ikB+/lBCBpkXRuJ5CbMiHFMzti3ADgu8dmdWbBd/Goy9JToE
fPuYxozh4obae7etCAuQ6RySnOUHmmIaZ+RSWXITcWUbscdBx2Mmi1TSBz+LDtgJnorjUeMesoDF
FXa7Kf7YeSAIqOlrKRFn1vpQnNR8qa/dsQGI6SzbIz/B20kaWWGy1lZlxmrrWqsRY0428YsFUAa6
TKhoDc8Qt0QoR2s+0hpLxExNQn5zDaqIpJAAJj5Hef3LTO/8t7KzhBlNeekzId0WFhywdQWoBhy1
PobyWFNOR6bBv/GcF18pM87HtPcXV18fkfKElUHDBUxB+LUPflAZTWOUcUVZNqGhNynUbRDTtwMu
hh7drc/9QAczbOgNzldQLLfWr+zvXNdz53DEE+GSg+/685lWo7nrz56ujb+CuhmOkJg4JRg47ft7
IZI+nJOJpWQ00Otfiys4HjExUrDnzuSvbNL8H9hf9r5bXMeYnREGBFGhMjDoZg3S9/znRAomkNz0
SDsZsDquayTSvPXKYtpGUcUB3OspkA5CNVA5iXLbWqKNOB4rM0F95AfvsfFgUGwoH+89WVg7UCBi
m44QBup/yGDbsECBCn5/BtgzMfUNNUwhQ/D1CsbkoDRtpnL4nEuACucfPZVo1SYWbuVKNlbYMi0N
QQfLQsaopitQfS03SugPrZucg2swP/Ie/yhp7nLsZUn1LMhlB98pJsEgfHF+89j0L1mcrX8cKzkK
SHk2tMNp2wQJdDMgjMS5K8JejbGRS6kZ2YuPUioBCxB8hnqs2osfuUVwoHkRCMTfGugNRlBLdx+l
ECQ/kpDKpg4v5WFurqwVTDnsLhVlTTHzV6rAukTK6tXHwKtcyf2sHeL3PI3FGEE1JejNQnoJYagP
d6ijtzqyujolMHsW8HxiVjMFj54tSQu3zuLFv3bhLa6pApizwxWcvfDbOxGJSu2QI99czdM4fJ1o
JB0WbD2aqpX+AN9Ahn/8NDLt1glyNGBuahbvVILnqQZC7sIXLTyiPueMIEqO37vC05UvSepzqP46
LPikC7dQ+LHpH11czxagTuXJGYmLqeDKParR24CfEV1rVOsQP4uy2FVnT9f3e2o8mebbkldgenWq
bSCl8K+AmdR8vedQLl0E5Ef2KaDJQHr3+5lZdWr7dfmVmGmUUOubGHoruAeZYiRtYZw5NYjDZnm8
jRM7tqe0mV4CqH8SBe39V9NBbC9ZvnrBbcBL+2BSBIexIJV8WAKqyUhpo/OyA02BOTMtIC2HPcpU
ujfT2nXc7aK0UHWliHxmtfe0G9m2mH/qPO+HYDvcZWNTydiGMLOFmLjKpqFPNL/uB+3HC1jykmvI
fWHCCMkGtnu6kE0r6Pnq3zNWW9XH0JQ4l4SMaVX/XAFq5LXRb+t3TdzfC+Jc33/JD+T1gsosPYac
IVuKaHaGrA6ukrbgJ1PjQy1geL+zmBDx2HMF8uardWesgAnSTyQDTnvJuMpKIi2fAvybL04QGnUO
A+pVmhnBSie5F5N4xbjan5jqXFF7XInNUX0/INUqywynukDMdwLyVtAy4WOCR+egshlIQ0oete/s
h0co4UDYBMGnfA7ItfHwYIKXwhmYaMSJc5HGSgyMA+IzUDxCLx3hdipQ43wlM+jTE2QK2gMCPiyO
RDNvh+AHv1KR73yDVU90O1OxmPlzqF82YSKj4b2u+BriPvB75HphcZhjHKmUaZdsUE8NU16vLLx9
Xb2ojsYpY/vBHnw20/+SxVBNBhIRs672yvzR38paba1CeMF6S7tlgzh96/ZdXwopHpwtODCYuIif
thRlJoONFA4FZP0uX31fVpaG0FguvHpLkV2B5o2wTwaDvNVZbH2UunN/hMlK8slaSHsgfgG4MdhD
ufHURfdXGTYttcsSDW3OW3MiSXc7ih8fqoso654JCAdwggmRHoqdRtml0cfsCB3UEbHd2jS2JPPm
Qh461TFAMNCCnHAhmHCAlot6g5g5Dl4XDsy4T2uYNE4LfcJ8dA8vLFTiyW6D/HXOC8fyo+Udk9GB
7x1kLMicynt1rDSZSsS0b2FtXVh0yL8BUDaEW7rz9Jv95uFGBymE9jmHRvQhSZfvRMHVxJLgC6Mu
brV4xQdsbZgxK0w0KjAgPRVFcMTgblpPt+tZhZ8kwe0VXGOIhScvXmftG4dxwhiDeqzOQppeRalc
UfU87iibxPbwodxylfLfRGT/PNEAkGjbJyR+ocSOFgxjbTlPLKkVZC1NLhuS8fY5xRrkc2BriFp0
7ZQcObqqMm7nDVZTTtpT6jmC7bg2D1TzNRe+7VqtuZC1w7n3UzXqzy/VNTUZ6EKaf6yT4an9Oc+m
X1rs3CDwkDOvn/MzmEH8jESJZlC/K3G8qPUmkn4ij0lSIIEJAEvcYN0K2CYukTwClgsusrB7KpYW
0akKNIkvEP3v4SXp0mW2pworUeuJXRd0DbXHDJr/He3lEJqGqYr79myJvNt8cC/5w/INj1L/wxuz
ZMhQv820JZTQ2ulhc9Y26pXVAyZapEgCq4Sud1MzMyxWJ4o4cbc3u3cmaXHyYq3E6XzG+9K2BKYo
cSk6VbvoXE/jjyq8+4YAvzGueTsFG01qnaWRggCnsxUctOJQSeS+wn23hNmnb/9aZKsGToeIoIdS
C/8OBqX0IcaCzt69qEP4dO5SPOxMKvuir0KdEDeureqXhdZTzdemgnpH43428Duzrd4I2zvvLFSh
tAtRYKKekJtLb9T7FJKCtjt0aIeQ0YGL3hq4RLs1FXyQhRlmJkkKLsen7S3PHDJEfGPJitoaQwUQ
W0rIisg5LT4dDAINn/vbzVl3T24+kFZ1z/eSkJ2AOJoPnzup2eNQIfbB0Osr+WtNHg11QzV7Gjo5
abd6JMt0jqskDsZzc0RPA3LXe1bp0E6lD27w2RG5XYPKdn8jIYwaKSuaOFBeKO8PowV6I/6ZabKQ
g/LIATTzTxCpPpQtiJWucES8iefQHNWOpf5wOhR6pxed5FWMPf5NeRz2f10+zNbmCgJChdL1mrgS
SJU+otUTowBFcfdkSlNG97Rm+5isNdbXFwhioPMeiQTrlEn9bmVDz+c3pE1PmDeP0Ii/QydE39yz
UHI9DR2XSGewc4RCHAHBfDYCAqODHolqjIX62bMqTZ63/k5SVQSdBi/JYquHtSLpgVCy3IO5ZfPQ
cCpflb8cENijgAqcOv4OIlt4G9jhM5ia5Fw9eVB/BciNtRfKeFIsUKGN/3/SlmeIEjCm7fwPsPYA
ju3ynHAH8rjXWkkqU9ET3ovl8RXv9MxhExsSdq/N7oYv6fXesGxK3E8EZI4QHQATKWEHYICWwIp9
jLpvUEE90PAfDHBAWuMEL+BpEXseEqh7h6/tXHiR506oyWvidtVesy+Me2OQQmhMSmZimDH5uo2j
ZoKXLX1kGVlvi3ciXs9PKrRLzddjRF5C973bfaXxU1z/RI76GO3fJ1Jj47vSCoo85ubb1YeKX0+9
IQGY9vjNvdQ1TFkpFH1Et76FAWFeuaw47tVGc2KDOuJIjp74PXHkK0jhxNgdFDEV5hJ7NQfVUXJV
fsp98cU6z1JYInBQOFXEh7neA+Z8BocthDv6SrmZFv5muFf8gdPLJd+q8mrItJNm9ZHTSUNEmFPt
26qC0N0j1iL9P0Va26km95caVMRu4xLr7yfCZuss+fNHloxzK4yQEPf2pptwsBMH1RBzswG8cl/i
PJKrfQ0DjRUwvi8Fqjx2efdvEhjNMqJlHMFW2bLB43Go5ZruLgIaw5k1TFQYWW7HDFk6h8EHWHYN
iUhm0TtIHfvuCX0bi8DNuXr7pwXpMpQz/B1wLg2pVDzxl2LqwwcB9YRBeLtHpIIns7j9ngvDqXAN
6nQVK26z500xCk8eUMmNQVTEcttjrRcrZh6Eo0yrT3zeSMoxyE7e3UUdCHJS1I7xObUgYkKERhHp
BIuc9QvnX1n/DYGvI0UtDygTeJ9GZh2asQCalxVHBQxgbi19RLI5sg0v0/A12ex3MvJ7IJt0dfwi
e94AWZ9SMxB+ITcdHs0d1BJ340qin7yKoautkN33DnctEWINa65GgSPBzJPBGcDZoG/d6sFpDYwl
LknFtlxTV+B+1ehKD+/2ghL8VonoVN3Yq1iq2gnA3lAfeoKp9bbDI7dSWgngNJ/FQyUdwiPZk79h
nEmbAYFEl6HF9HBPTe1JkxQ/L0bbfmMr+6QoAlCcfCi5KWqmsNyfKX3jh7qb0mcYeZXnq3dHkifW
9Kj06IzrnUaNNpTUG+FS23vkB5usTnWwLnE1N9/hKfPF6TNiYSLj5q2l9x5Fl9w9vsU6HJnAEL9O
joQpyCGuaPJNKUWX99L8x1BBFtInfm4Gy+MF1ZjKUQ4PiFNfjO46Lw5UVTH+wpPro9RxFpmDHo2w
lLdb9rEo0ZpW7798EKlxx5RttXcfVmszVAKlDI1OITfk5/dp5h6mtXYfjHMjrK+UsM0AZxInlPk2
ozagoxeAMqUT7rmWXd1eOks2oo5i4dAHRLhHoxXYsNxmyJqp2zHcFtdmMhZpT3PYarwxS8xTeoD+
2MdXeKon14/oZOtfR0J7xizo2i8VGRxp8MxmP0XvUgLbRGtKH49C0+q5kj0Pts5Bx8t3SP4RtZts
XXWfNCorIOzf8c/YX2T70JadopaBQXp3PZtN4+4j5Bf9Ho9Mrq2Bj+W00xauwPy2RHEM1N2wQrB6
k1MBHgJndD6Dl6kEwMphTvopeOgpG1unAaj0EmJ2VU8WtQlF9yB0M1b7K7Y7sECdfQAnHSrERsRs
fpwOIZlNP0giAccwT984w6txnN3vBdMV8bbs3/onWqkndSP049pe2Bu5gKbVvxuyzwKq+SGOAq3H
HsWvn1Cafv8urQH+zmQw19rDz2KgEOnLhOA85IlJvu4T4ZVpgF8VShyxGML9CMjjya2Mcm2wl8KI
Z1zpwFUMjZcYT3HPkTh+j+wfypRMVT2o1yUfhwF3OPB0Q2OmXYg5KU+yFyUkaC/qWoKK2AW4MWJ2
fYosX1/EZNLQcs57onvW7OIKg7TnjlUQ1CFz44Tg+CqH+sdYT9Ud2PUnKC88S+8Xs/QdvffaT7TZ
yUDychXOIYC9ofhlCi7m0Fn1qcP/LsOZIgiV+vh/YrhfYDbZRYpDxfhXYnGkKzM7thmy9G7OeyE2
DgsuiS/E58dKZ4PBCazuY4g7EvFBseVxenlbnOq9kD3qn9ZvzzVqLmY7cjqs3odHCbyMJqcN801V
3e0Sd4IGxNWy57qux628p6F5gwNfWnv1AeRytN5mo8o1fXlOb5BGJLvn9XRFymmFKmUDaLyZC4fw
VaEwHYUfOgR7ooU8yI3tjIXVwMVhogQEhKZsbWn0awXq17IPl3nel227Bg4gwkpjS0+eoli6iUgf
en06o5uEM6JmfEKdG1p95zB5So78VAcysHSsuC9llSHDAOWUvpvmLs28Bj0HFkWgLY2mPMzH/6ju
jdOwcgMEfotCk37hHzxcfeN8BK4NVSrKzWA9dcEkhB5ECENhfxQOFVUZpzqUlFAYkILpoPTc56o5
cX7oIo5wO/JJKn+7XLfDh6Kxo5h43R0wa/3slxAduvONGXyRDSgxgFfyNFsPB7aVc1zLf8qGcH8n
TpWnnOHTJIh68gnrQIiYMi83o4TLGUQRZXdff0d792VOrWpWM2dJVxobmTiGinu8EAxXJFN45k76
fMglotFRdJsh8mzoQus8HavhpUdyn14cL/UvpglgtgYUR//YzssosAJgYzaE+j7Ij+8HKanG4L/n
y9ChkJx04T/CTsLEPSDzdrWeXDpXEzhygwKOBGvK87u+RJY32nIaJw8zZU0wjvJokRwwkwTYc4ty
0b7P3MPjNoVFg0m2q7W9JJJV2FccKccXWA0G/mcBnGCjxtiKNS80Hs0EZXazozrwqUN3GyszVYiD
/hQGcUO8IybbHgS3uSvRF9h1nUx3mYqRSSe44QWbeqk80LKbDpKZPOK/hzyL0KslzxRffcK+wV6Z
AIY8curxXtTN238xzP9mbQl0rCOrorTIuUy2CPZliAarmDPafEclL1fEsQROKaUq34qx6rnLDt2c
ADRgU8Ov3bO1pZHhhMS8yUn/YQHbU6ER96VPiG6W3MjUGVESZVuToN5kR8DMkKDQ3PUtlZJ9Yz8/
HJt900syLNua3UzpQ9qmOUGaZIf8gIkcn2GMC8XOo9rpwa1s54DbcQ5hWvIxPDGcRx26Sp7ARCge
RPWhkH3kmdZSyWDPf+9C9IvRV4qVinEpDGqiCLZr1PQezr4gvCloCuNFWwbNF1RK0zq/JM3fUao8
ebvQKg+vmFUvdcbgzsndVzpUkFCkKlTiMrSGZVJWOHW/47yB1DWeuTs5TO0q+JfgI04uDeOriu2p
J3C5E7eX1T8PpRhfKnoF5YvfLnk9+YlK6z6w4ZORZwEuLb6yWwa8/XTIdTqPeHUvdxolqHUeO+e+
cN34kOZ8YbbmkXVxcpf+KJsQrsQleig6dn+L9JDpkPcLFx3YJ9DqhfG36ePw+f82ZcRBW/OUCsom
ASfwEq3fMV1Z/RwFSi8rZXXoGxd/cphYDNhIVjjIXx+jMoTwWTBABHDf8MUcXI+C54I1Wr669l0D
p7EMxQxHUFL4u2igm1MR3SHH90meYbFXciySEziZtqeOvYY4wbd/Qg4KTS1gau6xUN/0INoGvvab
ZyRz5/3sdBTgtF6oH7jq9DN9e8WockpGUqzp55td5pfg/6RZ3ElpaYkQNIDJyQZZxlkLuszZcDll
KW87yMZdBae2ae2QNVJgdtJ8/NkZhAaYAt9GoXs1NExYW6rCWijM/KGM6MpnNcfFGPuDiCJhcHzs
bR+yIm2FpoGYeQSB6ucJcHBtHA6Yw72S/gLt6F6pqQRM+AsGfWrQSWnYWBv3UVD2tXvWfl4S+Eyg
HNjqFPY/yeVbelZzdidn/B4TdVAsY9b+7geR+65PYfLp3d9KUYdNwQbE7jf90M9/O+zVS2Ph9Sax
KSs2Gh+J98SO2IJjw1BzKhYxuxDqRLz1z+QXuXEK9vkyg8Gg4dFsxbTws0hG3OwHTmY/JRznn8Ls
ae7sNBmp5q0GVU9gyNs7J0Qy8lWqyzmaSxqfzylB2+Zaxo/9uvJa3Qkj8LnnEQRc1QgXUcElighD
/DeBVmPsRK7tynNp8LnYdcJ8gs9w89GVsOLvtChGHgkp2nkjZwt+fuEpRDKs67oQPb/RuQWPnHze
oVqdrDMjqtiGgu/2/sf78JVz75Q3NHSm2WlczrP7uaHhPprxEBwv4xuGprAHqdPUYa8Qr4z/CifJ
Sctxhoq5tmC9Sc6/zXwJBRuGqD40NmVBk87R7qdVSbI1pMKUHj8gioTXtvPX4bFoUs7SJHm0W9uQ
1YTThtm3OzkPI6dS2zJTrmWsLXbuTEbC24T94qU86ee1siphS9xGgCnaml4i+qnOqN1XEJv8asN7
zuLHRwLxCSAUO/m3rKgfdqm+KY3UkifTY2KabUySbckl7De/VNS3sLKUKBy0U+5VyMzf7/Anx/oj
U6VS3Iach8NqWMHmW44jY702IPSLcIr7XKeJEN7AJd/rnK0amvaT4m6Ys1UOh+A3BYD5hLFx2dZi
iFN7pZACiZw8Sm8wlfY43f5ChR71/ak89Jn6JqO/3/jOOhWpLpoF71sLFW5NF4K0V1lI5n4Tu6jh
9N04X9sfG7IjblrllSiFVKJ47g3B4Tt9r0FdpKy+4Y69k7Se+HVTo/5Iqq0oiE2olObFPIFDNd7L
k7FifwDFMnSs/iZihd1AyP/+tUFbb5x18K4tRdOuJ5P/NvhUs14mhCP2108I4tNY3MAfBmZvpxSp
WLfKQAMePCtJNUe3BS0AlTXjFMEB5W6v8UiWigb3564m7RlekbBH1vUONOdS4umQf2sMN4ETOAbW
oVOz5UA3yHZBO30GsXalPz5M1OZZNPfY4gY+8I1uvA5VaZx7nZLeE5LCJvpQmOpRTlWHTNcFvT9w
yFFif4jGfLPymTKUd77JFTgC8Rrt+mBFOxeb2CdWftk5UmYufaUYNic5wzAOj9A3UXYIlD7XgNW/
POxsDCCBGyYB8/KXP0WZMwjLbDYXN/FNqIr8C9mioIyQBpAoy1Ah5w2C+RI3J2Rno5zWZ3I8KH1B
e00LWR4CH2esHITdFcKgTWCFTdhThTwJTzslNmlbMW7ajgcborqVWsXhgLBaj335OX6owvMvfyjV
UuUYL/ZNf++O7PthdoULziomJsOpQX49U2oWUQYX4mVuC5M9XbB6uNEjh4+jDX43LUrB8b7vlh9J
KqjPsLXB8feBU3QbpOjzYWDuYG7Py+hZo5j0xAyyD7Sj5N/s6fBAgyTjMNTWnbvtTESjI19bAIp8
ITaWlDhlgCMrKFC842ZowQbgr6yZemKZPE2tzJIM12/xT0clxAe1oKh1w9S+DpaKI4g8qxLZ5EGf
eutqJUopScI92wlh/h5DLTbAW4N6oNwMTbtew+ENGYFyOmRxVcexh6fmpsWkzTxU8C07s6r4DtQY
arUk7r0jA7u9xsRGYVHgVCRP47rPY353zzhPWTpa48hmFgg/duOFiIyEPLC8Fskq7XZcCumI+KeT
DTF2qFYgatZGu4NxoT8nX/WjrZpPrS14ucrU4dBg2KKkiK5vqdWpnmsc6g6aJbwj7YF7z81Ub3B9
fAGZ3J95Jb2tfLDY4s/rRjhVXmTHwAphhxynCejREEENdxqOX8x3VfNoKuWSt9OwxKyUYvA3ipGB
mWQzkTMhDEG12cugUF3P99xwkzzLWyit+aTaCK4Tce1d9gOin5YWHvI8W1BAz8+mvoe1FgkQabrl
8gjASFXH3YL7hBGRYy4f/17O3RrVNs52RvvA5b7dH2p7o0yCelRG3f2GwZwrHmNkU47G6qfDnl3Z
ZqdBl07RYbouijwHu9j+3YZTAfQm4LIpqyNbuoT3q2vnUOOMZFRvf9x2MoDukl7LK+u2iVFpoWJh
fXRJszlww4MyUQ8Zi27q+KalmfzmSImqZ6C7kFpCusPZmIyT7avu4lDQq26w6TMOK8d0D3NHfSNT
CWr1kxBZ6fwhcQjKoYfUBvWNPCO++TIoIxqa2Wq8r4nV+bejhf12RdMnfMxLK7CXKj7UM5DOUzY5
FESc5h5zdM7jubjmiioJH4YDLNw4KdEO/Mj7WnNQQYZwmuvhxXHWTg02ONnd6JEydToxBFqp0z0a
VLRdEI4hXFeC2yjA26xQgPFtcBv1V5eai8yuv9t2P/q9hhYIOtjyrWhYOzHij1dRzqIUzT8miAQQ
n7uTYPyQoQVo9fNKspMSjhjO1GbWaUYfaCntWmXdV3WksjvOgEKSJw+sUipOwGkABr+mMMRi0Pm9
vD7u0BMOjHeCR4sJT6AjgfDoVCC9aonfo4gL1Vj2VeIa7KGmhnKpVKp1QsOi9o2ElNrwRJ/fgL94
GUfKXlCImOizeThFQx94P2cMd3P/5ZIG6qHTUqyHtgDksQvAyWQt2GcIQYgre0kI+tGc2VZci6D9
dFP25GfzbJ/8iRiwa0xy3noc2Mz5+ESnB2EvtXoq+ua/akBpp57H4WMDfVMvVnukQti+jismokcV
7mQb38KThHa/ZUjK2f4dLdNvyOFR9LQcXxPjDMlCF7QbjhhjIBamPZrTVt+R3NcvErx5oRO6UfYK
7vg/CBQsqQG/KahbNcvEs+GL8U+IiB4ij+DQTME9sf4VVJcWSsCR4EvhaW7Qi8CQY/XK6NJRJaIX
DkOaG9j5qBKs4CXfWyhgKakkxVUrOjerVjWVNJV4bHqGF01kOjE0tanAQBqr2r87r/73o81TfmgK
IMaRD/01sg3xNKqAmnwuxCBF7fccRco9gzu01QTsmhIvVguSkzafP/zcnjLp9XmkkGNcM0qksgYT
ZBWZ+fv0ov8m5a9yhdRqtK2W+tHDmoIz/OXCE0S361v+o02NelE3mAi9ThLbDjddddCUTD0XRRYN
2/rmXDM7aiO8rRhvCxyz5uMIsdqyKqx593ERVNLNwEg3CJOSIGL38RwJheBhWnHXTlqvLDS39hsa
yq2tsc6HQARxifsjtaWwz6/Rf/EeBbT8uweGvLOGryVph5xUJ8b6fsl6O96StiqeZJHxxNKeifcP
MEs6ZHGcoCcCrNcUKxvGmYOonvb3F6PtQP8ivKOezhEsAlCjYtEkinj1Ad/9iOxwwJntzEJkD/dO
NCfDl18sl+FJTcdhh8LVJUVnzEy1Cv7oBg1szgRQ2UT0XjJpAuO4/jZfvhk6GnAvBoGfhyuxnMVp
tjmZqDk8kRxiL2ZED4njPulYrGUtPdgyjO+uj8i6YMBo8mPDSgjzY7A4x5ZDDy+LetK6A4q2GhZn
APN3QJKdTXULWB8bKV1nq7qJMdj+3hesNG2ibsnAZUj9JtFDJdFgyddB0KdTCfm4Gk8sWlnNBy3c
vyAAJWCB9hXvcSDpk80lW4J//oLf+KCfebnEU0OMlWE5uxiRBoEtEralbD9eFa2zDVa3rBckJ1ez
dYoxW+S80Bkekgx8rrF9C4cjsClYSQv21J8EQqXynikAz1sexXHuOgl07MH8OHULXGiQXUrkpoB3
0Pi5pJ2PibTqXjjpBjy+csGJV226yIbYDlLbdxQUZT9YldGsB1D41FwjOSkjFUztZJhs5n2zpSNz
zc09YJR0SKthc2TQQzoUCyGbSPD9c1ryAYjbRQho6qRCRNAPW/N5GVAdTXmxGkp1fkHKcJ2yJuHS
wDUodTgjhUFRXdMK9Fv7UwmYFkAr20MiIuGoFzd3AK1TGD55fonrtl73EWadeGRqdYEB1X9nxd3w
h0WbdW4jfPmWpnu9iJTTvlDAzdozBIRc1wyP8DhtxLk94LXwhOzMbWEAtZp5YaZfzBo+Xchp7Y4q
NovRGd8xl8giO1ZSXwbDcVJh9mXEZpQ16hodCjYmv2uo0Jn8VvPjb7smDQXAJwEJ+v9C1IGNKTbZ
FnxlYhHfWNgdn+u7vdKNe/T9AVsBYJbiJR7XnDKt6DTArc+YMD2/7RCYtxZGmnDyuSdVe+xTwtBE
GFWFdiqEK8/FtG7wqOeVu4l1TCjfe5dbZsggpkvprQi6DJTHFjgvYbU2QOJX9Nd4mE9WD/HnjGJz
M2NtKZ9w3EOAC1mLITb1MlTmoG6uPcdKdWuIocO1PCtVIkwoLrmsagUYUDJYM3r7AwkJ9/tjtV35
A3tQzUJIYn8DtwK+WAUX/t0rX5yPol9jPASvBBRrixCDDQitD7J2lzXcrGFLTO3lvrFmSxgYTAjP
rlSHb/MC0GImOSSfT2/mp5mDYeo206wJXWP+BPNP1drlKLHqnDlzybrj098mJIUnG9pH+FDC5rvY
cGywhd3ZLw3C8ziglCY6xjyjjREzHc/kf3G6kN1cwH/+zg9PSGFFF6xTFGp5uOziEQYU3jyxr3DR
VheXxv5iaTZcSa/FcW4MHUs4QzdSFInjAYTsSE5ZXQzRdxO6XHHzZ6nkbqafvFvGFBBE053hD0lN
kGVUGsM5J/HlT1QUDDgKzfrTFmXtkq25mgPRbdjF596UCNQHbmYpRHKVWYgdAA2aK7qHPJkZnINn
WmzQon0Rhj3MMl/9ibKNIlFexuUDGfLPL/uXgJEbNOBqc1Hng00OIlkG1AjR7OTaskGPrKfLS5iX
rgKbhq2wzvjEwHQZdKsfa5cYiukz4x9Ic3wZbsKCE1CO1NLwrbNqRrGyjKNy3buB3HpCnv0oKtKw
d/TBahbaCQhA4890aRRGFe9e2EBIsiQ6psmaz20F6/zHZ0Qw9Sk3PPVSq+PbckhJz0yrQlZz0Icy
9QK3EXRW5ndYvhaXzMvfe4W6aRjaUg8mTNHMyuNKjMLRGbnBbfdqyRKR5KY3Ij0TKKnHyjUg9eJ7
KqG/O6oBLmR9jlJMl/sBDU3cfAXjOSaNSJQJovbM+9vLzBQnb2RdW5ECNUabYNbxwgdsBw6FYB9L
yitZo6B7RnqiqShadJJZ2PlNLC34s9HbPjlWljBT0a4S7cUjv2ODUZwiIYImaQyaTYnuXKx1ys8k
FSsxZLCxN9FBDrOsWug3rhx8+MaLFa96cPhbkw8Cg6nQicUxsMbGVEygQAXTS2GiPjHuz1zKfqi9
uwjRkQBwmzr7jzwItOZ3W6bDXVau1ZDAGUi1AurQJp86RrCstsDdEC1VdSkKjmQhmdZBE9cUcUzC
LXP8fDVAiNPeRenwTb1AlZkaKscO3snvuXLm0vTVKfZURoi2XSvLS55a/xFgBYNOzCneh58r16qU
1RetEu9SdQIhxlZI5oWpJ/9Nk4cY4qyizuU5/DZlP19rSLZTQuTCKr5aQ/UZptP6Ijr18/OlzOmh
TMnjRihfjKzBNpdHuUpnq1UeXjvMLJqSw8OwzOAYSUF4oqRs1vr2eJzXsYwYIJrVi7dz3ULY8sA+
RicC+Wdr76S3121Y/8mGmqZat+eJ7C5DoIeiCHY5WR+inVngUtUPt4cfPbMv9JsFwTZDzN85NaJK
cMMgCgajAk7nbCI2efy3zurJqEZDuXJypVzasJfRVQHJ6H2fmR+mHOBMGJgWiBjmC/jvf5XAlK/B
OIkIAiSR+Cm42h1oMvL2obnOrvH7XGa3fjcMWNaV6KQIoOgLj5sqdHdDpiWuG6jnyCRPm1UbbdBI
Ao7P/O/R+CxJtfhqJQfC92ApwGo37S8hMknyeO4sRbEMUZeHZyTDC1MLmRtCxnw8DjC2/XLuZKC/
Rub+9Lr9cpXroqdJ6GD1BEPJbcqnuet0kEDaVcByklW0xWKNeN91TAGFy/ZmflpGZJfZprPDQodi
d/Q/eeEcvttPeB7Hu73MusZlgI16IwIwlDcNNISUmFMSTWfUzh5RRwNS/IMC8LQAyt4pbECWdXMj
jhhbQw5dD/bWACBdToc60S3wf89vKqmOWHNZNI8e2FigJucgy2TiCv2QtTMUmbQ4u7GvzVnRHZC/
aK6/5PawpwgtErxNQE5fm7tolNQDnHkdRh4R6xw4KEypXpg5eC3/6zS267U2Bq/1a8OGbNL/yAeR
nP85B6K6KyOW0aMkmraMlcWu4QhVnS6U08sU8q5THX1PQuoo1guUmg8xzRDJ8aYWB8x5jejw/J/5
5vuAILvs4R9gy8WiXxS9QRvC6kFGMdLWgnOA9o2enPGIgYqDGS/iwhAFM2boPly/Tt0ZbADIkyiv
X0WeshtqOcJIyGLjZ7mI+WQlLGAQWnr8x7NvJv73GrDqkhYfDqlIZdQBkA+4/N736MvAr+8hHtoi
Dhg1CsuO1Q15n+WOq7o7XINrX77584jiTIWP6TiDtPm3P/BDzl3UUH4Rr+OSeIQU5TGj/g6NC6Y4
wkwRzD23GISe31qsvVWDwIbBlwIVQjfuompmSwhm6P6uycchsjbktsh+34MhvDX7eXO62kzTbiDC
YJF31fgfE8Pt/Hj2J+ipj8jfNh9hJLT7zSYwHmzJgw4z64k8WmAFdprymUhFL19WIqP0i3RMjw3R
iR0Ww8U00DpDale4dTjBRqGTmXEa9vOlnA5x88nDjajXMgt2104z9A89HG0p+7ZA6DMA1yfIAfQ1
TF2EkkmrXKVFsTWOeYK5ic6m19/u29SP12JJ/8lsC35agcSzxxDdwHPdbAGep3uazDXeBeMNk9j7
6fCLfafM+aVVfBCUwNj8i7I1p+vWBVKq3MOITpl6c863leT7gTL4ailLjO3J1Acp8OMH1bjNwE6q
h3fHEYVMdSbJt2mpWwfhLfeF2jPyamrgZzTVbH0kSLJrHLn8ySBYzl2GwVEC/CZ38iHuQaoande3
HLsEmUB6J2BVyyn6znzLvDjOFlaHRJ/vDk+GpXILDOHbrU/CHQmmFi1XTuV6oOE6qTBSLbdWUMST
zZD0X8P6KmgNjyDyPC4Z5d4wYxoNaGDmqF+cDojDYTMbg5+/be1emzNCxzflu4uduSe7xr1pBW06
OiamDr7UBt1lnBkceKrhJ9HpeOwzr78tBmiQC/TeeWZB/zFDM0QIbzVvbdOs4F1OCpnB/y8AU/3c
/eIYlo6niNhQPFd/cDg8OxozT4VvmGIOkbqEG9urK1FQno42tEtsm4OYgl27lazRSjt30tYVDx/E
M7B0sYL1H5VXkd0LloVjzqZGVBiArvHn8ymedw9diX/V+SsiL0M6uNXZTDUIQiW5jmpYvYccN2Vb
nXO5XjzWzdbjPQArOsNQ0+QSXnU9g6mqtbCVUUSiP05S1lcrHfdMm6S2Ak2LyzjUZfe8vMf7Xqsc
6d1NMUHuWfQCDFip8CIbXUbnHslYF99MiFetufIsQsUjSx6mDXCj6eN74Gfl514LzZvChf952Ukx
s0rB0xZshNnvy1gZTKRHGfZBDb5N0+CthXO4HBHn4kY+WwYhy4saqcTfqFpMbY/sH2gxJkOLKZdf
coTlOfOx/DyaXGeE84+T4kdEuuyLitekdLkKioQnkiHdwvO0tmalhg0dm9OHc5K7cPGiQPw0YP6E
tiC1nwrcCFJARWvZxj3js8WJ3qDGAqrWfDleXnlJ74XUUmFLh+4ZuugzeqQdm0jud+9DrfezxP0T
eIxAAIXv7kDvkfOTiG/bF0lqwEGN+ls/cdjCGvmewf0EgpNQcSLJSaAGs2TtQ8oAiYgcf2YzuKgJ
HJhvNdmareIwFyfMlJLUaAkVS2z07ds2XgwaK7SVUVMBlVZKMg2YDRkPY9d5yYbwK7VjkCKTmhvN
W57lpRw/MP1SjRX/j07LsUNLIDofXqw0dvWkWoRHdXzndC1DR+KGbSa1wsREdi0u6+6mD5a/Ai6m
1Rqib1zl637afdAUNZQPd39+7P3VKKsK+qaK/Qz+U8YbxMlWECakAVPcwuvy4ffJxJ07v5+AyIYO
pmyDDswMQDrBbKR/DrY/k1hDdx1a40cHn7HfJtaQjAs5jzrXkzzRjYEDodjzBpybozWGz5FFnAsd
QY9WyX4RhF9EL+XnyMTeImeYqkjXSkanM4X2owF3+DAgtZsV6cHG4Y4xkkz8s6vk/c5k074WSsND
XyQv6GqnNw8JGlqKvKVAiEvUoleM/rV6o2nk1kJqbaOL8YYclgoYeZcwVGoBjeNq6a5gGNLxvpIQ
CeLlZUciJ/A5dT/z/pWiKZz3N/a7cu8I6AXVfhokczMm6tjfQ5zIBeD37ZQuTxaNm9h0ozUJ47tt
RtfkBHLcJjJ+KWAcEuSM1WdveMaW7mLeUjbiy/C/XvGWK69QALeiqDvw1U1iURsH9WQGUcjfPQE4
N+ttNLoxVsGzEX9QgX2Fq6sOTit9aqAUQQ1kbw003H7IhQfXsxyl6LU4T4mA/gxlW2zqaRIXT2hf
VZNRPLHju2yrFInx091ndW9tjyw86rvk+/VZcQc3997RyagnPCx42lzexqxxUWmFO1SeejxcprVU
asANVzHjgk7uPv80QadxTtAu8Slnt/+AMOQiEufuYAH0hc0tZdaOZtibVT9DF7glv1x6yJL9Gnqi
GbIaReEJF/lPdoKqvKcTwAlbPHLtp6pzVcZcGyctHehyTh4XN9HPwqq6jKvAsXhoaDky4VHxozzs
U+6e/9a8ZVu2gUdCN7Tb4fF0i9lE2wVZtZ14U7OfTqDj0Vy+ZHsrbhWM0D264P4o4QEMKHD2JU4X
0Sun05o1U4mif+B/9vBeuwhciU9nPasTcgWf39bJhs1AtIi3NbcqMCP7wD5pyhUaJzJIXir+DGlV
AqIyTu5ftLWb/tcSSiZqjVVvcsSGMxTpwlPJzi9RkJE3uoYEGSBVEhTGFLZ14Ti88TR7e3p5tt35
vQOkNVYbXafXKDhLWWSXqBSrHCkBQm4pkyF3XRGdIk75HfFrrCb8XFoatXSNBGXBVzDwTUkSkTBL
tuyY1/7HH5F4XdjdAnriIFMYNwlpB9A3x8kFZpbkjuP91fd3i2lgbsNdRemoAHpa1xS1iodbJchl
Nc8BwKSb12e/m8M+T/9OHTvMjejQfu+Ya/J5ygCbNEtQqKVPDCmrjOFiIt34QWqNx5RVu5zwWAZz
/Zn4q0eCUnyTY+QFevt/u2LkvAvgZam4WGhb1mNb9QFccwf7DxHXYMTym4iHoed6AbxjisqAn5Y6
IgGSovyKiHUg7L1zxpposvCGNiE7xToOJV2ljx9q6uXr3+r1hUGkp0/2fuqgj80MomHfiFcHWvlC
vsZoFfek4N0EpzH5JpLs65M4HSZyeWABi0Zsw1yqq3eTLhBFGRmnLayjmZU39Uz6oERYUNoreZaY
lzloTObiv3Kph/3ckWS7+Z3j3ouupY+yy0w0cor7/0NHRPr7Ul6MoKCh9Sgd9rYXiBXChVJdlTSq
jTh3BNGT3AUyjXA3C+BLnVa7kAzpvhxjDlBJVCBVAvlfytCY5ST45zBXjyjrBd48jWSFeIbwlG/l
U25RiMWHNY0YpYQwvO9jA4n38CFnR0s+tG1Ymq3Pi4fPoUuO3O9krenAfZx7WxspxzH0hoOAJek6
1R028Sf4h8HAzco6rXARldhaGzL6Xu9FJ6aDqzZymNFu6C4XKzlu0IJMwH25NtrhK0scF0idIE54
i+FVbW4TxZwVaaA5r7QQjJQ6k2iAQBFeGJLDU5AoWBuek64C6+pVcJj4Kgzn60LlzZF8kBLUf0MD
dL/3VNBShs2lsqS/KdO1K8qK77G23IZMUj6KiGCUq+DPGX5mF4tZardz+LEKG/rK2BzQ+WMiFp36
kHL2LjPD3b1iLUv2PmEDgszaNhmhLsci70nqzAOgujcchLgw8NU1YAZ2AJVr9m/+HqcPPiJQE5E4
Y2qFrT4nQIkbCP6wtH8TkfOkQVdbDFX/42bbmFqpnvbJ780AfZGunzzrwQYtEIgMPNXmxHTp8yNk
lT+ir2x4ZTutJp86AD6rRILsSUDm/UgkuD0RXXB7RdPgUIBSSXM9RwN9cRxJuojVbU1AF9HXmhul
COHkBTY8eTgUoSYSGfGL9VaK6M5AeJAfhrtbC6vFrfJrXeMLzhxcwwNmQVVW3Ys3opOwnL/824wK
PbxoZD36bo5ORjnBPxThvsgobv0qr72bqOWNU29vyycUIlNWzo3WQYFQhsx6a8Nn1qKFfykT/BDs
Ti1HSikDtyQLBkY6uny0spCx3t3hhdZw/i6Gy+6b5B7jpPxk7EDOoihD2Jfpo7yF4nXMiP2lXni2
x4owjoWC8EvQrOMndi6Ang3ZNfoiemHH6hSKMRix/ADQb8ZQUSMBZVu1uGgflPtZDtQPix4AJH6z
f8Pk4fYEgoHO+00Iztw2SW87ZbZHSyu5d6R9Ykv1QNMQyGa8ux3nnQZJwq6XQCQzNXaRCYohJdV0
8gfisFvVYT87Av0qqotvt0o9vKNFS0XVZbTHsV6d41HadOCZl1YNOfcwB+kMD2hdxd2LbNW3LX7P
4vuq6hhKNRIhfMyCzZQq87RZFrK27jYH/eOrKemvZdFCVial4jC7GLhvYWrBc69J2IrjuBVYeJmI
edAFmX/UL5Bg2ncFW04ZNGzBLC8+jMkNqVKkakLTphDPk5WWGelkhNedQ31bhCutEhWYCWbNXHG2
sxzNJSJS6NsR6fML90a2oMiJBKX0oank7DN4CSTThMVeCqX9TQb0SxW+DWMakyVyNWDK7Y4++X3H
72OQaw8dDhiSyIEWbuHOqM5GBoVLYcmIK5SUG12lH8BK37F8GQuKLUYEf2HfDRF03DU8j1FY11IH
r1P/qw+xXo5UdClSZj0cgQJ4Dojz5u71jouQiJVn99CdAPcmFLrpVe34lkMZdX1oz6bRpysB0YFs
jeS6TEeoyQXHtIJ6J/tvGnFFWNQguWSmX5Yq/lciIMVEwbilFqyhlLq1/lBJ5sKayiWbDYxIhtw6
aJF2+vQ4re0I4AtQ7MNdXGS+A1rCMIbuM7l8Qrksx8cvi3aoaZL0vErAtPdXl1fTKMvv6wZbNKml
/q1A4mY9CDtx/27T7UMghI5v3GQCKU5a+KUhoTxM2wgANdC20AaP4pHbZRDToHAHWWImnWerAE62
Kg56pHYatshvv4QntXIZx3ZNFdBJhPqZ8OkfY4lYdlhyNBOMVSGH4BVok0/4LiKEnGPUzFrBR20n
Y4KQK+DD7fktX6+hrqck6DwZKqR3W0vNNg6eQ5x0qMfOC3heEDbcCTyLcRZ5wXnmVqdP2kbslYyk
GKUDoJ30iGuO2ZHBOsFtjtBm8WC8KVNjpbW0lqp4TIkhOeViV7ZyHk3gs8U8GFwBiY4wtB6p8VNX
w9oBjgUO47JY2IpRdwAJh+XEtQLQQz9RlEsqfG4xEOfIjp5KmnZkMsZk1rmuge7LuW1DlT7sYvaB
BUzVEktQQ2eIYHngpm3pUeSnWFZywvzBJLCqmX3uDB1hXjurBnJgQKoueefxeBtLjIcEg/GTiEaI
CE+xDu5fKBRpTOs6xs2m28j5I0w0uR/hC9Ucy9YO4M7j+5BplS4KlaROznt3KA/oBEDckClXDrtQ
OK/um3oyiQ7V4sGRlaPZoCtvt+3z3GmK5O1xAM/JtJh26epq4qrh2I7Vk6aNVhwuCvpiybI5N4aC
O3E7D+vKNW3zC/c8GTwYxDBDztFyoPc7trfr45HseZlS5gmRFrMR511ehWdy/VbmJBLWEOxXDTl/
WGdGkvrOwGnK9xv6pUtHSkHmXTOJxSBy7iggr+4ZJjUAOqPL/9P1k693r8c8z2g+s6R6jbTffnIK
EBdFqQv/Bgwfx30g1LDOamBBFEod1eKEeQ4684GDFI6jcge9R7WuTB3IU7GDkr6262yKZH6HJnwd
CtSJVczQpebA5ZB1XfDp1EEeMiiMhijmfGIpsAhrtUUJ1auy9zROkZk1cOsXk2LKrPd/J1kcdY2S
ZOUs57DU6jlQHVB7WHwcO0OCOmQ0wTxB4eFw8OO30dJkfsf8XoXQe8xstfUyoSY/So7hGFxFntQI
v7kvglKWrnSj5hO7xyLB0yQS8bhwYXPkFMelsErEHCj+CHANHLZPvl3tL9c3I53vD65YUOjQOve7
UKWMuybt6nfAePGnDOIGeW7ZCAIziiye4AXI+VV19FlT+hfRYo83YHxneTQIxdCNd6XiY8LcqPLT
qZcJDtYjeEh/F8m/6JjZ4e0P5KnOnd1SseZetFIJ7CAnDIiQRPkT7x27jkvYHmplIK2Uhrq8F4Eg
dP0YrxS46//fXsTpg6r96hBylGDpi0uCWFAbW2j7k8y2xgxzo7INfDQKuT0oin9lLh2SVJykBIKT
x+QDYvDQDnZbg/KIAEA5Brqkihu34IKPUpJfXCnzdv6dVM3k14q1wqYpHXYq6266lpHhPIv3N6eQ
W2zTc6NmapjkFe/tLzclaJQ9WnIkEx0TA0IP09XQ2vvl1bS/vk137PMUj8I0yBA1ebB57ssPsBfo
dYJpjC9+1GtXyTIbZPmOKHYz6ROAnN/6phCd0oVC2kLPES3GA4iA6KT5nZybnoha31sgfSdyhdfX
ISGIAfwpH8qrMJc6RYllQ4fWD+UsPFcYbs6K5uvE2WGwRP0+hE/hMfvbsuVYuD+inBqjNpKWBA25
HNjRxFbDsfLG189mXZ6L3z+uy7KbvynY0vtvOreQ4acuHVIbB9SxlrscY1dVXK7CqXcm8+JFFFBM
VDal1RzVWwNKg4rJ/hZF4hcxMTPgMDejK41T9Y+wyfpjA+cwjYINknapbYJHniNcYWXkQ4J3FynM
Y0/EK1y948lmZL04GkoAR6wkn2OXT8Py58ry0VA6byyZmPF7kSidEApL7TqRBbwsKRe3QfbBu0S7
zL/yk0rsV6EB5fqEhDimLmBP8KDZb13xgXLrnf49Teh273jpPAMNi6MvT53/3MZYLxJvQr0camYo
5IvMYa/MBYBWUKk4KryCr1w2bjZ2M+ATyTVU3Hw5zQB7AMky5XX7kTbiGRe9xlQizntD+/CyfMXq
i5rI5DLwCNbMMQlOkOdkKA72cBuqSDcPscL0d52TPnIq/Barw4kHJtpaFfUd2LE1ZlavAoH3EAsg
RXwcHw8w2T0YP/UXQodbIdTVaemSfj1ZfjEL7MXD2LE/HNmJvV0yr+LLH8UPbeCX+hhlI4EYxWKN
mJEW/vYKRlhiOZRrZzhCR7o2q1XJBt7M+OoRJ/dcNFGqIBAddxCXFd5Stdl88oK0YCgQCkXuOUBu
6zWng1umzHMT4zwXSZMvNEwk9/XTfLJuvsS4ZgKR7zdLKOcxTS8tX1U25FHhvvdcCodNrKSEXXWf
lxZ5yFl6J6Mio/gnvgug9ad4cQ3arInl3NkHJlyo9wB+y64FZObaf2xctWv5dSSowY+5rXMCm158
pTPIviFnY6vTLXm9X/8uCKWnKsULnIpi434hRqzUyCmn9DvnKICpBiWO9TpbfDcNWmis5zSeBogV
yVWsvRVlD58mzahLv8xfi6Kkpj3lnw7AiafPH9Y2WeHBFlnRluri0ruJLCuRi93P4PNekCuadGMa
2BX3tXygbt4ewmncmTbk63VykBUZG3WRX+vA3+WFyNlbEcH/XJjkrDjiizoDF/RJ7Zw4jZ60MQkM
LLcmBcmVwiRt3CNz6nBXh1Jhs7aSlEyynKFti2DQ6tfpPd5ufBRMWz0xb1Yi3VB0JlcLTdoAacfr
0LxNYGFduGSExzqIcf24tyJyeRmpThCZBIhLcLFpr34pgfD3Lzzm991cM3vBglkLhNBBGj59sg+q
9YDZWYy1N9lmsQO7IYI9ZEv8GkxAYfKSVH3burUtZd5uv2ePUcLVSOBXnUVAjuSmcRcwGBvb7fF6
LmwPVMxnt5DFvg5Os7sOwLtIGSpoB0awP2wI6Bj4hi3lfTRwOgYsDC//HloPUc2ilkST8mCbcVzG
bWt57QXuxOKT70q4nCNhrP1h7zV9Bdi6SxBjEFrW7yhe/smHrwPTE06YI/mEit0g2xMgTyHJcihg
rAzqy6lyFqrhtBV09uPUp5WQ5/W66YBubeoW1TMmmpFv/k4+qTZzssnOMhaUuD5C7P8cCVVZejIC
8/VVJPkQFAU3oITKWzUBMfam0s366Qp/JdOhu94gTCPGEEk5P1sN4tB2le5HoU3O4sRllmlgLqvw
87+Zjgf5/kX+V09prSZieK8x+GLQlJQMfE4a6iY52IS+diRhx5WKhfvct+DHtSwnJBwXx//k30WJ
l3AecGqulGEpiB4cKY03UWvmU0XbfXgZw2hNbjrEQc8034P4aplGXR5bX/99N8P9LyiEIx92CYJ6
W/fbo/ZohUm3XqLEe0crbNcHe6q8xChSDRAAeAYNuQHGCX3oelHDnePPqbWOmeJgMCNQyitkG0Jl
t9aNvdklghMfLN/axvV6clW6frSOnZAvqsYlRumXbq7ymhi/aoKcfUQd360XXaTEx3RLBcgjhL/H
E5UKEB4ltbE2p9R3zvJc0fQ74uoxnxLoYqGzZTu5h83Nf/GZ9YLqIQOpIg9Vz/ugoTeuNjFb6hca
F9Twt/HVTyDa2BPEO7QOyQe2iPoc897fl2tZHzDDpocqF/bVqyLy+nCpHLy9iJPTE7NOH/WL3s3q
2V5dcGmkgflho2CPLTO/Q3PgqmJE+ZNdwJlWqdVLMN2HsGkZrBd27k+BCPVKRe0N05VP2cUeWgXw
QC06qw5ABtnygs0xpVtDrCJD7pY6Qy2k7DnQhW1Q3g/5pz2GTNJhM6LE4ndKn0N7HJbLGg0XJ+PI
pTgCr/nHlLiBT61e8IIL65FXE//PTSTY8tXVqmCv2qpInx12SY6RLahds/enyaQCLsRimheCd+cC
X9nsT24McvNK4cNuc0ejB0AWEZ6+hEvA/902DFh46QFUbZH0XRqx/vpcy1SkEeEbyk/AsBkP5y7W
wwidj1ZdkGVSObU4zleVf5VGLBbJTtqKEiQ+vEV3vCVar9Fil2QzqbBGtBT61X7hmNbvA6mRabTD
RuXZeluUCAVweGdLwsI8jF2IlgOoQeoEOY8gZ0kA+EahCN6LCBB9a5Zoh+eWbupbn9hQ4/ANVzLG
ui6ACASIQWa7Oe8rk7f+gobWtKKuk3wUaljkm+2SjDrX51tNncyy9rTju3Ldg+WKZoWMSIEiHbKR
6Fz44/XBXbkDMSS7/s+WbRSRYFmIn79eBHP4+8BRUBbkZEAYPAQ9QNKTF8nJkyuU1a5R+zvMHZZl
NiEkFBfwEfN+ntDXBlpLHmioiXSvBUtSMUtwPW1vQ6zxs0zIzOLrMaPM2LMMi1kPqR22gn024zjY
P5rOyfmqRzsnJu5d4coehE7ZyElShh4Na/x8WnX9KC4fz9Eu39Dwn0k10XIeCxRAqyRMN3g6BVz/
EspJwR16stECsBy1vx6XtKmLMe07XkzBshT9gBc+5T/r+qyO1ldLeJgbGsHl8UABtK9DLjnI3kYA
MTmR9/yJXk97/7FqOn+AA164rc82TCRlSFkyUrQCs5pu3ZXlG7j97GJslbbmZj6nlweAB1hLNMdM
NdZt2H81KIDigjVxEiLarAvdpwcOESFlSzdJhC3GLGe3XEkThxXtPfo7uArBA9AMKvN8u+GY1Iiq
RuMeth9ipZuAX8jBIfE4tySmTKc9Wy3sdAh6G/8Xu1ACjhDKGB6YdJaPMT3yakiE2jdh+FQA1DzG
DVWKbC9xk6/MpfTpabC7eW92YHKZqXpOxnDtf7qu3eE/ozH3x8Yft68yUpI1e6hue8kR43xTCxcD
teRl/8hpZZfKmMqSB/5woC/KZ1fz2qnd45kTOj4/q8wp0bzYduPnTc+CHVj+ujHHG+t0igQMHH65
eZ1UcMB6A2o9FSqdH45ZQ0MDs30I06lOwI+Fi48XfdJnkjwUHu5BEFXNvWL4oSwgKRfvq1SrO6pa
m5aYeHTgwvEUC2XyphLcwnK4rqNlV+autFGJLKeTf8gNCkQL2OrSKAy9//LEz2iM69FWQ8wzJJdD
nxJXCITTyYfhV1uQHlCKZ1kgiMcWz2l2FrmhFE4p3KmjvZdim1G2aKDq4KaHLGomxie0874rriWo
y9FVN0sSTKXZxAHPO+XeVNGHnmMGqQC3DDx4fpB0iblycF6uvVNl3v+Cs30iKD/XNwMLgJHR/PVJ
siwn1n7AHAKc3jAo8i3ACCkNjT+vTeKZL8AhUimFYP8Bf89+Dnp1VkTeJJjTxzqRMumt3GuWFgNL
yb+WrLZiVU8ReNocUjDBgXrc2Yfj0x3RTITebBnZyWJokSoDmeaLWbHzlOlj3JYlqPSP1PAgb6G+
RavMHB2ZZCeTnAOvpUwvkYsLjkfQbGYLas0OwQMJd2JKOE5rzcVcJKOOAIR4qJm1OhKQuNZMBoCk
zNpyLu241ezEFg9p1Aj4rghuePYf6ii2buEiNfvfMzWDOCFdF/x4Wwzk7229MRbTSid8Ot+/rG78
XIlLwxY8OalFcPgbSybaIxLBZYSaQAYKRTGgFlW5U0T0aljSrljlWpLZulO2Xb2kPSdzrJbQ0YeI
X0kCsIvB+K6fctxP+WgMrwOCoUMNQej8y3vKCODSzcCGT85gtP1uwuHy8oGvRdDeaw3bRIk3BCK4
TWj+Ekgq8wHAmCY537AvYgCx5xhIwKUlZuCJC799f38JQPCQvLaBviPMR+Pkc//Cskl8HEWOAu4t
EtGAk+6yOryfxsR94G83PGo/ubRs1EK2zJ4Cx7KtuvuZdCenmHpMaos0SFExeDEaYtYhmQuqlWVr
JrwX+r7V+pRaxe9qVOBXzSvCFPj0K74IMymGT0h+YBnWuDkL9Yazbxfvp7HcDmNg+dZms/yp+lWJ
4soyPBUXDEUg/b2YyWKH/eGx6zibdJfXebW1yE+M0NHsr9KIl/hLX7CFFfHr99rFj5jqBq6QH2JC
KpDcWF68Cg5ou1yuLtMEY5JMf3pt3Nojuu2iB1Wr7QvERjUfsL6iWF2et6uKnFLjY0CLJBWIOSLg
AdYouRlBZ7AakivMisNdZZaKTkaGo/vosuFuAVyKY49rVwn5OeG1Ukrqgji3f+Gd3TG2ivXC9n4P
gHkMpMlj6oWcK23abvshDIZJXf0Hn/e9+fF0mYNg6Sjj/Zr9bIpd0hSDevLV8V//PEYqSked14t7
LoZtdOwJaMGWp1JZpBZ1GoxG6c1R1edsiWPN9xc+PBXIS5WX9YjHszBtFd/9tSSbCDose8yZMSS0
aqMw1zUTMKqVd5v3f0QCfZ6Hi+H8RQuQaCjdqP+FVW/tBKBUBW3s30f72/Ho/svb6bwpS9rQOJIj
uDQ1MurkSeamydov/9Uj03s0jB58kV7gEdrUlCFZW/N4HzvVvc+BmlawTA2PYxSTWHfb3Hr6Mwij
Zt1MbDFA71AJqb//M7EGoYthl0VIkHuwTbrNM6NDasHpOO7U3GzuAB1SpCUAF0+djYORHYAaOKUX
HdAv07OMHMuu4UUICifbMpiUDgJUGngM67ezVslXtcqwsynkm4hXyuhtFL8RRSvElbkCpSErJ5Cp
8dLYKdhs9thryhudHLNyk7K0ClAEQ0tz5arg98mmSFbmRvrXnL3QvoICRbzOc0/6ZPMP9sSSXv6q
+KyKVSKo3Au+3plzDBVP/I1c4zXv/G4K7053J0UHN9kvGn5DhLOTx2uXyPZe+y2kSakZWH07Udo4
RQ8tNG/UIo55+1t054o3mUcWctS2KPfOxEBWlqEmgn9KLJ0o3ZSq7OTpwi8n1FJc9BHajLYr0RXk
ONwtUOf+EuXJo6EioC40sDW8mJ7FJm5bHfuMu0z5xCZMA4PSXbFI+3mG77xNk/L23EAxHCYCVFZD
X23bIdxxqfKIihJ/Zm6DT3hKduaElwpaZwPKDZnT+7pDm+BSSYo7Wf3SfQ+fNStxgT27Cf0LYgg8
JUEjNzJqxy79SQfBziHYl9igZ7pu/+BSvuWrxNkIkg27Ubg/vmXnzdSRTqfeEisA1gS/eBKJ0yvr
SwAbcCNi1fagSmytNpXlzpY+uovU2PWN68sWAOE8uis6fD/oiAAAH3QM79b7nXMaWnMVtQJ1Kh4z
jA7hjbSuHlYDWIaiDX7DUSZCz7LyKpTEoSQzTCZOb0NDGpks+OJlNc6PLFm2neiCrMHgiU//yXaU
xIyzCgd93CeE2wtsQv9/2dvBbS8W6/VuPnxOIAvThMpDWXKiB96GttZQVBk6vQJRkzgODf7uOzEd
Jk+CZxjQbHgNZqRrsS5I6ObW1OdVg/5lz7tlXTRhevVtG2LqjIWf7/EDld84UgTSrETxCM3S+37z
A8JaWb94fO05HJ7SNisj8jvqIbzM3e2HcsoCW6k66Ih6vEdLIGuKx7m4+DAVzAiG/3E/xPMkL09M
UL9x7C/cYy2UYg77sKc/NGFjGz4noFFHGPEgX/VJyhCuoSrxYKThahqF6moKAQ7gnOw+ONuGSLLt
QN6XPrTNMBAeTnk97e+BNvUM7y/zi6b3YGtJNQAandMA7WUHEXfURtwQ9XHSIQiNv0r6SF2mGFUL
SJqqHNwi8Vr7m+w0e1T7Kl17YiAwcK32cnYRiW5fn2dnNLLtmsUVisibGAE2z/YfzFeCCjhoapsj
Xc4yhdGOoWmDSIIZpb96kgxjX3KvtqzyrYdH2//MzTkraOkWDhQq7x3S2JoN3Ci2cwNwhTwtzAWp
5K6XI1dc40V+InHnjA8Sk/EnDWUZHQn/not/2Ts4N5Dt3SyAgckbMLoWmoX7Qkoi9I5DcL5v/KgT
VLVFoSLLcuLVLr/sxg47xyPwD6dKvjkq/3oQ/kDjIX3DAgiaWmus9YWCLAVTVWKjp8E1Txwr4oBx
hKcYRy9m/bnME3KfhWBLdBlKI8vPF8Dd75PtNMMH1NIBsBUhL85tbd8ewhOFxVlhhyT1dcZRQY/w
/jr6hUkHn8WNh6MIY7YVcLukvvk7Z5gZQdxVHEDPDg5xHECtbP4UqZZuVt3eEjltO8KMax/Ez2jH
01Fze4Noo5kJs+m5FeWyrtUrkuVNkibUF0zrzUVc9IoNRUnm27JsiPmAN3mn8nRc1pHoZL2Y+ztd
GHsbzHOcjTSFH8WA4vpk1bmLMFwNJWJVBMshQOvZhaTL2mtf3wesSvwOp0w6m2lZDLja9DvXxLw2
7+yPlyFdlOB6e+XQYRzdvYSDsXFDzn6SsgK/xsrg+h6hPwKoYdcUGiOfYsujPuUH0PNf2nFJw0Bx
RC95KG7bMix70LpHqEi2ZeFsP6jgHZFU+Vt4ZtJ0rg+X19poKVpNeNAuP/lcFBlTfI6gUXNff4q1
aZPPo3uoBrFoB8k98smdR1Egj4VH6V/4DpGa0c7XMuY/SC6W/Mmepdok3VVqsYZmJ7EXytxxw+6e
jfjgG2sxWxgIfBL7lRyDB0ennorFJyP9vxSLMDymQ98/j64EtrOfi39jtxvJm59iV2iTYYNhSqiT
EWXcBCkZz/felxz9VJuTQ0Q22Cld/GA2w7Zal5Jq77JARYKmXSm7o+bAnPoirZfCu4Pk8W8xcb7p
R+k35m8WhyAo4XhvrB0YnZksSLBXFRF7KTjU7LeuIS+gOmNEB+YvtchzXXtg64Wpy9o+6vTMLYsn
5II25L0vzRNi6c4ZbfzUCmXf1+ariQ/y0tqrXECHV57nlVxZFuUOM8sa/zUQYXPTMA8/ACoC7hpK
7TbnZQ2mqhe8A83oad9jHHKzMTKxduZg4ImW7PufzGp5hY3sNx8rI6uB2A4+WJe8/i8tNe8Yj8RJ
7VHUY885GNSYlGjqlx7sf9xlUSThIJQGPdHWG5+23naGFoIos6YSVZGvqdDCN9y6xJqgBuTOIKxp
aaV4Yh2nmObPkbqrk+UJilAfdHwJWnpanzz/J5GmgTIE+IavXUYDZduIs6VPNhvP/clDBQXCvb4y
9PiDWfRVNlh/NMVGqwByiVwipiDAmfV2ObezWf87UzhA7Q4elomzTCE+nwAZfQc2NgTJp7/LxhL9
k6yygKCwwH3zX5AAoVp3zOlzGypVaDoyE5opp0ntcJb/2BJ5wip74rz5AFynI9rDcS8IG71orx5/
NNLkmMBHqDYjGClZX4Iqg40CwP8HLskrNFF1G0KCHDXGzRoqahlmL7TBuGDguYjCgef4gf41h1L7
9rHiJSWvPL1tfDyV3Ag/wYab9gkgfRUey4ZTx5GFEBAA2TKJQImvsV+M1mxkArn6FDApZ87mlUUy
iIbqYi7raiUzSgU9rxudmYUYWVJ+fAE82laYuHGfbn2psQcq5jp3mm4iFV+HAV4j1LqDUCrjmMTn
PjBrtVfm8mzsfoWVwSmIenI9+Ut1rsRgLtIy9pAYkBql4N+fKPRpJvGoIViht0/kEEpJ4gOHPidh
1QkaX5j4PPPYUlokdZEmhfET9UIcvjYuaTxSjRF5JoSKnqG4z0ljvFfl315zaF4u6fYLWNs2E4SJ
UgVIoo+ggOVixTIt+1ZS2qKvgWAjRpEAWOgKnpxhV+AtQ+MEKlwMbehvNaQZkoKNVFkRq2FeEgUL
l5j14XWaGeS6oCgI4Cf1i7QslJx3jOrW2rG+gpMubGCcZDdvtZ94MTxyfkxttLGs1dyZBV3BGtFD
emusBfOVfqW0meFG8P9m47k5wu3dV0CrBMUoNu9E2vkAEkBaCSghdl8tHOu2FHGMa3A+C8bxECAq
3+BjZ/SO90zvqAaWs/ok1ePkvrf5juCC7EFWlcF8+YN6EUirRRGYXtaqtiuFR1jm6VH/w7tVk7Ow
Jr2tae40LsFJErog4ZkuybuZlhfyn4GXzMFv8B40Tj9LMU3wU4hgQuuSWzwuzvOy0ZQOeCAeAq0A
11ElcY5RExuiwCsHIMkP33AIYKSpwcrtjMEitxoQ7EfNRF9e1bOr/e8guVFIYRlpUrZwUpHEhpCP
67ssf12u5Yg8eiSRpI2bLnwsFsfkxuDvyzu8At293UlG9AmNgBwvAG9qjdzxBcpPtuSTLGdt06iV
hBhYA7LyOpyi8Zo25yG7p7++UqOsEDOBmFauAeq+sdZVWyNkBV+/XmMtzZ+bWjhzTMEKGKwJsUPO
85qXeHWv9JVJf1Fx/nHKFus6qxn0vp8/qaCnGXKTdOu88FwjKKeoVFdWnPOSm7d88vMe2Y7yXQ3Y
i8pDAQin+Zy4WuUc/7T8hoqAVtQ+2T6OYNEI0Wou99HYYdm0kejEUe5+9fFskd94VzmKoPCkQZIM
en2cxqoHMLeKT7Rf3gYlrZsYp6auv4Cj93nxbetGPgM1WYOT8BJ9X9mI4dM/ymAXSSbuvk7AoPCq
UvfqvvzexhcFkb97AgY++TBuFDEBcZmwTnaSxukg/2Jqhi5uYyHeHmKgTSv6nGgWl+G5HiyQ8wFQ
ZMi0NI9lkYBDzDhzFDKCxeqTy/h1QF9qf0h6Ud6mSCA2mszre7auKh69BdTBPyz9cN9i7UNYTsoN
nj4xQb59UIw9GTvqa630/LWvWAYZGVmqOy09JO1Jhya2i82J8SOHNDBdRgpsPIAIdCnWM5Jx4odW
9NIO3bWVONUQC43M99x5yfwnRA/4gudE4l50PCtxDdtdtxOm3OdEOQo/QQV1fClYS3efTjJ3OWvH
z883DsZXmdBIRT7Mq00wQWFrWwrahumO2f/GGVCLehKcRBT/hn2K5fOH8t68UH2Ull8eqq9ehTTf
cq0GdajbXI34AlUSCfTr1s9DS7B3Lejn1ZMvzYZ14UP69Vul1pxWCJxt9FIhWu3bbMDousTqkcSF
Iert4J/srNZAfxjsOmU+1qufcxZkwsAWj8e/N7qRooU3inmbVenYnBiORv0zMFotlzYVg5BzgAEr
+/I33tvp2xlmAENquDnRTGQ29nOOmC84yfwZX96g0x5c7dTY9A2PxD3Ma2F9+zSDLJ62lByvoGHl
bSstmOgzORDhxQi16FSf9XlDp5POTo7FikFc1rfxdP0byMGp4u/P3ItgghFvHq0DKXfDIqneSja1
hWtqoW3SngDyVglEa0pSreVMg2N1Dx5T1G+/E2qqvZ1kshwucYCXP0VST78dVYYjSnnJULD30rsD
P85bBD2MAJezN9w4/uVDUJEUFr4sdrHgZDGQiZrrS57A2EgOSNz+LNRofD2VkUHL/9URHMq527x2
OazAgCQnEs2ZDii3g0pPw9yO1C0xN+DJViu6HGuV512dnU0ginLBIwVvsKsBkptlkAQZzMmQot9G
K1NCv7xXn7JLmL4BMa1xayePQQ1ksJDuEqK5AAvhmW07LApjUyeexr5OikGsNk1sybWCQSQrQMe1
bT/VBNzUU9j+b42bpeKbYZZW2vprVwIExq2Whvdnu90423iioIoYACEBDxk1Srnf8hiH3esftiiQ
VekG1aSGUjAwK2Nj4fNAXpP8j0qWCtu+QHV9eRusKUBlErLnwuKUMHhBgZLMkSRVFxILZhMnh2gx
/HeBBq/loXJAbT+8EJV+CWfbFmcM78yjXqdJuUtUIZDyv2cnYbShPBYHibfx3TuFQTapU7XFLaxn
co8TqcCvkaClS1eBZ7xrKjVoZ+F8QMP9SEPSCjIcv2RhvLOWzN0ZvNhN0hOVBUKJI3eBUCqRRvL0
o46YJfC1Dcnn5QHcbz8pAVhXdsGixi+9m4LUpVkz7frEBU9/LFQn5QZVo2LyWj5Hn9K1D4zPt9p6
MzXXqhZnfLRh2dgPPUTOjfP8TkqMI4pApPKzfMZUUNSJefmDOOqvQqGM3c/FnDBLglSGWw+deGXx
BkQLFmW7oSO8rvO9k8YviNWE9UPt+8FSSQ5gaWtLXhkXvh7ghMS2Ve9lOq9eOAkrkf0UDdMpMqct
CTcO1A7HVMypMEvmMrZ4n9SOD/VkP6jQ7opHymL+1wV2Dw8gQ1dENfILCJ9jkkTM9sX9+mnqf3aW
n9Kb0H/7uCagjR2y3IDBBkeEUb+9oLPZ1PVKl8ql64Zm46NTjQqF6UWylHm41mLqnzVSUcynGl/O
hKhPACuvyPd1t9YZrb8rNmPJ5vr7R/1l3+5H0ncoeFJIbg1P1rRUvA9l56XtcnMQTnQwpSH78UfA
R6ixfvu5VkND73c6Jhyv2I/tPD05rIQSyNKKrHWGZF8h+ncFmhMUXYRDomxTanWO+FrJLqieDZnt
BwOt2v5XNj5gm7gUq1mqWWpDB9Tn2rYqZEdl8qbH8mIT90krAtAGcj2CHdo07BbEvjzz5vCVU9+M
W3jTWqBIV9YJfwSbMmRS04R2nagYPCnAxJregIbWbm+V4RMWdqLyO1giiWzVdBOmiMR8EAulYMwe
ZKwJ9WmiS8bs2xhAavsL09l0/LXDUT2mKqZErynW6frUJazQ7WpuzekF8gOejNQEICFk0HggKS78
tTnbCKgHRmbph/jr2LJUekghqEXFV6QCUZilr5o9+5rJMds0ELUIyMsfwIv3rUxAhnLxO2mOyvUb
vqKlD/GDJ9SYQQYrBe4K9Dcff0g7gEqTahpfa6fsk9L2Gz3HAxgRXa1xkiqPnpOuLPhHJK3tRRin
mMgt8WWCD1F3xVqD/PECUUlF2oRAhTHH1kOo0KmavW+M1JnrLXYVlIn/XAvPcZ+6aoDjTdXaMSgD
5r/DRZ4auVX2ezXzF4FBLJtu8gpYF9Rm0LSNN9CDVtMwfo/flloPEg6UaiiGqiTF0Ws5aD3NTRsK
HZovnL1eySNYpYlPvVCcvnZuZ+FO6S6tcUC4eycGo/o5p9lO7JvYB2gtnYwo6b5I/u/lJJnjgtlz
7AgpgOpyu+N+PI5cy8gvXzWhRIRUnrruxrS2K33RWM2NTomuM3iWcLZWlDhf2/I+o/MBMzJb2cBg
hFtebbK4MEqFv8IJ2zplqiDDtYL0miOZx5NMg7p/8Qo4Ii4pNfDKlMNy+HwPy1rALulZ3om2m22R
KKtsa09rpeOqq+ZWKzEgWp+eyXLzcc8tRjpCM1w+1PDI+Y+iFAOnh7Grfe2eefdYqBK/U/VEPhfN
MHB5uO65EXfHzl0hJydTGnAFujR5+gJo7YWCgjRU+vchPJ6ilJ86TYBfpR+61g9NSkY8GNnVWyBa
SUDvvwi1Q42CgHC15FUFYxXAyNyGFI76Yd3nySlwsq+G7MnKhigfM+6l00naUph5Y+0h6YMOriEp
2vP5wb9qRvGpkcdjW/lf+IPYqO+ln8rQ5PfaXnMoWEofX5noQyPPHpxTQ0tjlbLtQTUBwAPuEHMQ
e28dCg6UxKS9orQZ87H9vunJs3g4w7HNP0bzwF6Rt3Md66E7SbSRNviywNUwcamywKIXwnrOxXvs
xzgN0Xu8PNe7KG2AZ2JzZSqX3xr1LsXFLEX6lrKJu9hjb4m2us6X8gxv1gN5Xlnu3r9FnxDRZgvj
dQCSOMCyljqK6iYVjEifVOH4P7em8K07y2ri+yGe4jfqoJRbjRUS0EXADeLDRdIoK1CKrnLATv3c
QwGMcCdq2slpGSGIT8d3UBX//6TouuWpgrhXOnLdWjp4MMeHBsqh+DJUD+j+OR29Xw6gzppn9QHa
uw7/6QgIVxwNBBDoRxpjoxkSBxf+Ho4YGltqn8JezVEBeByznESlIJ3fyd15nAsYc4X3BWtXIC/i
r2AjTBKsTFbr+HgszEjYwRhLbFHW9/4dmMKEHgRHWat6v7W9XBgnOpGQle5KeFIXlImweIHIRY9R
hq3B7RSteR8jUk7LINrQci3ifgqYxoqLZig7saik5sFkZpbql2ihwvmSvzmxKG57RaAMfvFaB7qL
9RxESrK8vI4ny+02xuTj9kCkLy+qE6A7t8etnRa9V1Sn7Qp4sW5Ku0CvCRlyUqlJTbh0aDfYRBai
/dAFp/7bYrfFqHlq7N4TbB7GCGChjjmmG60sz3Oesp9AlO4ByEr00DvjOs+HtLOXBM1qiMLHdEnV
FsdntOMT0ZuAJpipDl9Up/2gl6P271iTgpcIk5eqiVora6n8dxk1oRO1+V2pXCL6S38mhWgnM3yN
9u3NcyzturhKsiRrQWH1JUgSHExlI6+Ra/5jQ4rWT/dWAC0bLXJ6pSFMfs2Rnq85TnWLCUXU0TWB
YJbHnvSFxMgovAAZCu/eRfCCDdOo16VThWiPg1ceK75ZS4PGX6PAFlsAgjVcm/UHRuvOIEi3J5ql
9GiES9Yz6NpHn50+LdZObAs1xbc8gfHLRE8D7YuLfM8QTDyzwKdmXRYD+wZb8LVzRt56RcYIuY8H
RKkFpp/ek79bKsHFOeS6I83nd0uExpDrs+IbgzWbP+Rql9XN67c8M0CDsuQ4mZC5rG+SBL4+P+EA
MiiXLR/emh8byBRn2ctn932heazYmg+9IGfeVSdqYhAu/jaMXylQkEcFGxtFhG5KxFqWiu/pywAu
A/796ZOilPqbzTQAhssUcX39JQYnBw2VO3BMAS2QsNVRLPnZO5UKeidk66K2VhUX2Kv3Z9sUVcJn
BVGbYWggIJKhBlBp0lXSKQwpJs3OV6uvw7MR28vM0stvDcrB95vYGfoO8/eWd6K6QutlJIscdUYw
wVW7XNjVUYOsu728iT/fSxP6E7UaocuP/vC86SwoB3cC0XrDiARatxsfLvPRmzms7omsg7TNNc7q
8XM7XRiPW6bl0r4x98kKNftnVavZuTAcQroq8tPV33ASamrahHOivEmZ37RZg7pqB+ZbEabkXRHL
f8iUR3SpW+2zkWetaJTaS/ZFAsJdypFEs7jfbjDQGLAOaM+wrtbcGl8SYzWha28lKEwhYlGhVjXJ
PMvcZ0e9y12h4EeRbUtHawuFygv0wvzwCUWLYehhg9P14O6yD6YWXzNiotkZ5370fI85pXvmE5Lx
iHpeTgVtoV26muBKOJ4CS14RnmkRtXG1jIz1/L9P7jokPCeM4MMilsL2k+PbpefrLJofWHfe/W6W
Gb7S2q+dyR2eFfktf5oRl+q2GMSd
`protect end_protected
