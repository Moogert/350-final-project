��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h��t��
��V�r?||�o�$	�Ԥ��	&x�t�% ���kU7�/�~_�Z^f��?���i���KQW�t��c�_�]�r���إMy�Z��S�g^G���m�b!L9����4�����ƍ��L+�,�M�>+�uY��	�D�(7�}:`ku2�pt��Ϯ�m���?�N��w��;�/ch�����(����y�����=K�HH�좞+��A��|3�hΛ#�0#6�Bѕ����!y�;3[��WA���<RdL����3H:�*S�_�G���s�F�����%��Ǽ�fD?<�/$L������^/��s�źyMx#}�w���vkH�ZNs*.7v��~��X��4%UX���^7;.5��J$�� frr����I�K����"[#��#�����s��O���;O,��x�Q���ğ��� �%�����t�U�\��f4i"t�e'����Ub|��۞�$ڦ+0���<���N&�$qTʳ�_0���C^�Wg5��柎���8{ o<A��	ַ��0^AW?�n�eCNl��EĶ�Ӥl�V��V<����L�m�d�]����+�CU�8��	��3�
�_$�������|�L��x�<��t�c�l:�i�Yc� Ñ��(�~Yx!�M&��?�W� ��i���eܬm�����4B�T�5�g=��,S"rf]��G���:!V8�H;+���-HI������pU]p����o������6� �~s6��=2xI�?��`}I�������;�v�=Ə�U�5��g ��@飷sa4�������an�-��:��ф�bn�F���ѷ��J��!�ǆ�~1"z���6
أ^��tk�Lh�4�a}c+tRN��m�; ����5�m��lD�%�jf�7�@Qߔ%"�ͧ1I��3��K+�0V�'԰ң{ݮ�r���˒sؑ����I˶�?E|l��vU@��e�ai�E�9��� 8!�Pb웎�.=�]��ہF��b�yd\����T�q� ���K��KPU�:����{��m/R�X��Җ�	׍R���U����MU
������'��S/I�R#�-���	��u�괔�ِ�������(��z�,\�A��aDqZ
f�����f81E�*×�ٳ|�J`'"�^/+�/�olȅ@cx�TPhd��M�4���X��u�ű��U���;�V�	r83t�$Q)��N��W�w�����(|;���ʸ�N6e�-G`�y.��U�S�8A\"�;�qW!�="�S�Vc��Ct��
a6���/~�/����H��+����Jm��͎Yo�K<�/�b1'��
s�p��N�ȣ<��2�Zl���ƃ<T�)7[�koP4}'/��h��{걘+�y�:E��c��a����%��B�4�-���h����ۏE�V��N�e�Ж���["�
�O2�5��֜��>�|�3�ˍ���C]��`���,]�7mP@�/�� :���ݕ�Jm��g�ӷ��o6B#i�0�c�[�����Ǽ&�:�-�{$u��37��&S4�����N����e��f�mk��.���_(Ei��xP�t�/����#U��5Z��.=�t�kc�<�-��҂��5��L���7�e�-�߉��Ͳ��+�OVlA�^�~�U(�R�}�V!/���o��/��9h���W@�V�����)�㴤�<�u��f�e�[l�`��8�>���[u�#;[l%�bV��@��F癞Od���FPGELP��x�x�:a!{@^�2�L�M��f$p~�`~-�T:���9��V���n��Ҕ�����Rm�ٛ���:���۽��Fh~�{����48�:�i��g�.��?O�jz{��}y�:���|"BK�&\vn)���=mz�F�u��^$�[r%�]t������
�"	D�A�0G��Y�=�ji�p��0~v<jpΐmF[�g';�/U��OE4f�t��Z�X��-�RG��������G��ȕ�!X�=1��|e.	i�TVm��K�P�!�E�*��ŵ]#me6�4U���:�tJk�T��;�g��5=�/��uh.�I�AǢ��a8eCt�3�!��Z;q��',��-��]f��Aщ� !m�I�	�ۊ��Q?y82��mZ�m���	�/�*�b������wB5� [�ޖ3謶�Nr�r�\�y�խz���\5!;�滌.ЊCy���7h�Hp��)B2 ٤-U����A�~��o������I�ĵ�O�����5s�r��-6X���B��m�P�*�����(�ɴ6Z��g�|L�OC�$��L�^c�#���l�O��`I��ɓkvB��(�3��ïMX��ӫJ8�X����".��\�z�� ��и�p���'���##�l�b�da��ώ���2�h��O��1+��bj����%%�!�X����]�yW���5YqY�4����d�Gz��p�`�G���
,�36�h�O"�^D
,A� T�q˒b�ȡF�yP!�Nu�SP
H �.?z5�?>#]�9��'�����E����~�z���x^@�ڿ��'�w���(��fy�����d�:l�Qs�(q��a�z�x�*3��/�A%�֎h�t�-{��|K���X��F���Q�^qǩ#2~x�פ �F}����؎����u�1\Rq�h�'��S�=Ĥ2���C�0pҎ�[���V
cAs�%�J؛_�|�Z�Â$%�Y�fY7&���A����\��1����� ��6/8$-_��U"D.t"�K�>:v��fH��Wm�Ae����3VL��{��Ěm�[c�x�b�2g_����u��.=�DZ7r�U4*�����}UF�D�猗k>�����ń�E�!C�gË1�+�;�*��Dj�ϝ�R��"�4^]� ��*�_��;��&��4C#���J��oX������DMwQ�No�?jS�"��@�=Z�������J�!B�#�r��z�n������؋�8��$�ط�,�qJ��N-/� D4w���HP�5e��Z�(��B޷�9�¸E"zծ�d��<���FE;w����ړ������Ƀn���E���6�h����8�i����-#�����q��6��e�Ww������/�FA�t_\�!�[#�&�Rdq��r���폶�I��� M;xu��C��)y��ě�������mA�n���Cx�9.���%�/5�Ph��Π���Nd��<���t�N{o3L+���<�9Nh��2V�~��׳���$�Є�P���9�O�� �:�?`MlRN&�G��3:��srŁ�φD�}��G~c?�I���c*9��qP��'R2,�{��p���+`�6����A��Rg�I��{����5��H�Rb���J�jhnlU>٘G4�P�_a6:\>���ֵ¬</M�&��2CםY�N3}�D��L���b�hKXnU� 3 �b�h���m�S��G2Gݶ�8��	�<���'������7z��~���.i[w�9�+� _H_�m3�Q�����ͤ܍�cA}V�����+�vND�n�?�����P�T&�92�'���̉���%x�S��<H7�
�-=����BћKe̂�QP$ѥ�"�7�V$��_��I�y�po٫�40\pi�vj�h��ӷ
X'Mx~��n���f�����Uc� ��1%�W�T�{5[I����帥
����ZБ3x����E�$z^��i8����V(�E+�1ص��K�[_\l�?�nx��]��P�ӳ�Zh7���}���3 i}�(���X?�!���z��flZ���0�wd���5�q~V
N;ş&�K�J������J3�t��(�9趟Z��

>(ϟ���\�m7x�	G�ʤ�ze���!�(�^���Ɵ��>�k���޺>.l$	ü�0s�ݓ
�g��H1g���m��g�p������
�J�]����N���qxR�i�{�րu#GS�.���l��+._H��|�ZW�/��f�5���p��H)J�wK"Xs�N6����86 ���񳹒����-[� �~*���0�X����pB�?T`JeUe��#�_��,�Cu�D�	VB��|�?��C������+�J*O������{�<���ey�#*FVj�����	m�άsӏ�}jn[�F=˜}χ=V�����ힼr��T�d�]��&��B��M,��	�1u}�9y҄ ߀�®�%ִ�Uo�s���Ir��5�d��,�,�H��1F# q�~'kb�]xFkY���,*C7�I|�}Ag*̾�'>[=5�9"�_?��6
�����k�d'S�^����F��u�B~K�t�E7�)�M׮���Y���ȳ4�ш�ۯS-��tY�+�_�XQ��f�9�����_q�5 	��HZxE��_�-�K�)9�o4@����4�6AF:J'Khj˧RQk7�;��E������
:�ˎy_0����e�g	s=�&-kMhKfnr,�$Ɛl%�x�k��A	���1VA�@p#)�@Dx�ќ�ԩ�(%�݆�>\G�3�`WQUУ�?ߜ4�rV))�̑}k�!��"lV���*�up��5���F�c۪7�zH+~��p@"<�FH[�*b�r�?�6��=QH�'�^��v�z��� �5*jm`��["}q;�jE���ĉ�S�����jЋ�S�G7�q������`�q�^��Կ��6҄Pʼ��N�����oФ��-J���5K���C�婿�{Ȭ��l��Ux��Z3�q:k5�F�z��{k$�e�$2�!
HF�8j����P�'�b׼!G�l	Kk
�q���D�Q�b��=ƋGE9L%���D�vYXͥ�l�%	V2�Ó#����B����с����"쏈����m��Z2z�TKm��0�HX�ʚ��
=���i�j��Ǳ$ C�R���5��Y��ƍ�>�t�K�v����0;������b�����i��명���;�zR6��h?c咝ZH�胶7���v�O� ;Gb��&x���4Ǥn��af76�����wY��_�c�"�00���L�
2������XXm@$����Eie�+�?O8��繖��r�zA8w�#횂s��ϪGGgV4j��	R憨?�f=v_�E�bd}-W	���VDb�� ���/Uߊ����!V3�L�#Bay­~�=#g�tƿ���K=i�^-�&m��>��#�7ѭ���k���k��b�z6�\	c�g�v˄����"N�sW�U_z��@��]�Y���{�# g��b�Y�a��e>Sn���q|.�Z�|Y��Z9z�Ĕn�����`O�&���3��v��Cy�r����=',Vq�X�^Ș)�3b�q!��N襘����hl�5�ɤG *��x����ґ�	��N�6�g	��18mo>�%��p�Ƕ���x�	�]@L�Ԛ,+�Ut�3Vv��"��[/h�AL8_d��3�$��]�m�� ���0\�R�c19�lU��ՠTA�e�i��������@��fA�WL�o5P�S17W&4�g�1��W_�h����T��R@�.�T�*ͨYȼD�쮦���?%�K��"[��,gt%.�Iū�λ��/�MC*S�*�"!��Xs�d~r���Հ!8l�Բ����h�^�o�E=��J��)�����^<� ��]�(>+������Ixd��x�&@���x�t����:|vK��w�Z���!��|�н,仸7��/7'v.1K��������AN�����'�SEUόa!�׆7�UM,S�3-+��6�,-�h;�����ޔ��h��B���th%qpJ^�k�Fڳ��Ӱ���@�4�x ѵ�g|n�t�R�+�A7޴<��46�3à{�t��%l��'��~�c_Ql;�2��68.�2+?�[�7��