-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wVGwh6pVNdzPdCUh+oefVjpYMNMmDKfps1nSxUZt+Tnvob9SmHLVY2y73iXhlAeFKhWVMRMBFtKX
1V5fhhhn1Msq+dsMDyge7CTdAx/ePFdTb9mQlKEFHPa7q/rGNgKQ6G4T65ZmBbkteLeYU7s7Mmt0
nhTReB3FQAumjqWSONNkl6jYRqZUBOQxf/+tfsdf7GsJZqpMW+GH+L2MIsN9knH4wjrB+uDeanP6
O7KI+1DARTPmAq5bL6Dzq0uH52/mNSU9Fu1+RWajkVmkv69UIvWVIWsCaxhRX/Zih9KhhdZMCCwc
o+f5U98eUdAD09A71ZxFmyYDFudC09vo25+Rrg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
QXMXoo+8dqMp6fJlz651gvVwAcZ/o/Si81j0PxzUKxp751frb8ldqQIc7oB+4/vz6MOh1J5g20P1
9VlnU5tt6+QLsjY0IOSO6VPf/3+kpi//sNdwCSGgO+94dbUIOgyPGZRR24cuuqGSzzDAHzaIOQpi
xk17NMnFoTLd2foJNXRP8jQEWAjcY9hQPjgotLbrxVIMXRiHvC4gGbwemLpZJ6WYD2wV/68hUF32
aYA4zybTQKmytbh03n4u80pRdWEKKMgBkVR8EfhAXcJSgW/k+/x93b5SmSwhwwl6gFQEGpODtLSc
NuXFYTny3v1LbFELwkh5VLsmh4D7QtOBYKIKrUjihWAk8TNlVX/RwOS0VCM+HRMTpLRoqw+vvprF
o+i4YoEWE9NeZuJKj6OzztI1M4imLcdX1QNOygrccRKKbQPYrzJzYZycItpbRuevLem2iGrWDPAF
/98zmMnnd2ETIIOsevuVewYoSe+OV3hWD5E5Xk1klP/NCl15zv7xSWgFBXXAZZW94PN9wgCPXVuX
dc3KJl6HhZrIlVaTeIBoTmZf7skNGmRZKwCHbAZSmlQWF28YkkiZ7DM3VnOLqpDLFH1g8u7Cxa4c
ytsIGIhKroEJXfylrCQbwWpYQh9qYdAnwSLXuJHCgzbe/fxbCXDt2ZbF1N0dzKV4mnIMiw5j5QRv
by3I8Pp9A71i4OqIBE9rXdiZTMRMGoqMKaIl1wWl3hRfwdpo23/q25EvfYfY7jJ0t26eI03H2SIN
FfNN8Y+xdXrua9YXSQarIiDOBZPQq8WhCcsNZfrcoGzdpi1dTLICn+2gGvoDT/A+EjRj7wvuAfhP
Ibbm33ZOOUkAtcqknGJ2D1hWrixiwm3/a79VO5s/mhHE4vCKKgx3bVzx6bTttXt96KVLItY+XTH+
/U3F8tfVljJMnmL1K37N3SRIGNKKxnTN2c33rSEtW+0+D3UX+3JjdgGNcBqjri7tWn6z92hPEPC5
5XQgDaBwFLRV0GMeiYMThUDZXsWjAC9UWZQqvE6BpLNDniq+winHFlbXKzFw8IXWkmlmzVopRfOG
BbJujxxX7ZyhjB+KvzBTDbezE98VC1HomFVwuyVz+c/0jEDmUDSU/ys9C88+mXJLQEUqX33XcBiP
mBt1wh1hps+JQ9pg4lKvYlKdh8DbgJ8uyDRYXPydOoHlrQv+UQ7SWIb92a5CWYS0Z4z4KcoIhY2y
2zqcwD6f+FkUEwI46eCZOHi7sX8yZbL2H+w6LbZh5CpPBSHz+OYks0F6r900Z0MBP/s1x0T5TVOy
o2c5c7x/8+xN5NCncEGPYQLibumlDw8tvOnXBctoKWfMGR2RveCa7UFavoEE676epS61U2pxBeXS
fHSLYhgQRsH9BMVe/RD1hfTCYmcQw22Z/M7+9v1n7Xote+AXYhKMhIQZaMiaFwjYoYLekaropZYY
sQxvkMPrBh1YYPwGiNQir8AV3COA3NVCV9ImUQfLPLP7lZY6TdtSMDvBYhiJ+DK+A1+XeqpMaXAz
JELMl63xO09L0XOjWVEB6TMCg54yw+HAUctGDkIuJeTFk6OvBwciicLnDqI8GR6zqot2LrJl/I2f
6Ydpr+2pQbxFVfRge3C9xjjNMEaWb/cLleWMM+XP9nSEemeY9xgisAJ9x6KIQEzxYkhiNc7wDuvM
g2B5AHkpR+m8Jine61ENYs3qvNp/hEsuRRN8RS9B9uGTRhPq+uWmZU4WBG2eZNhA7MtpjNzIQaJ7
1hqqVTmKVzVJ3xhNgvgeOQcUvIMY9jsTKYuaUiBaKbudgIHNfT1KnCgeoD3mWs4zZbBXTphpqNIp
fZtygQKhq8b1YXgWAWYmwqGHGOBkSi+kYwzHtmLAp62yIh7LSKsX/zkD3vO8sASuLLUm/6vnVv0T
PW/hYU8xt7554D6OffNzgWhWv0sErPdUBUoxmZdwNw2OfNcNzplQDeaGLTicJcjeAnNLuA32NilZ
ANVmyZPxBgWuGOMvKwLRYL16wnVBJrNrfnXcUzgwGaQzJkcoliXKsFk8Y/MCOSGECw20X0U/X6/f
elGSLTArO2KqKZxRrynx1wvssZ65yVJXchp8kbD/yIYg+s1dDhKmcEm3z0ApA/ekAjC3ZfsKGZ63
dNntVRfMSua0+zg3yFi9Z5MQRtGFj/JRty9S8TXBRft4+K6r9K/WSRvv4jS3ipYCPK/sPnc6AR9a
/BzZJ7//BYliOtBoB7J60vPa9Rk8TaqM2dY+Busw9vvagpy7wCym6wrzI9Ms3Qu6qM1oQwHmxz5a
JcpeZ5ghUgvUJUFa7/eMpBgESfK0nh3FznqQrZ/RJgX2y+YHzbrxc3NttBz5rEuztlcy5zBrqjxb
woIGoOJnutXq59EQ7H+gURX9hNt+CJ6B4D0mYZQEk5jejBrR6gGXHt74vrUhg/aOxp1yIDEVTQOz
f7rdWirduDVulKPHW8/1au4Y1XOMOHyM0ZqqBsLw589dSy8PR3dIK1JQEp3mqUAB30FvjzfmgdY/
6F10vy+RZwQFROjuF/vWWKSBhlpEsoVFsYFhi7n8nIdXx1OVgAlbcGCTs3PI9KC4LkaRBPaf1n8B
ppg8VNvBCq2QFlPI4U8YniLugWseaW5olY35zQ39o15uomwkutWe1T9mIgrYYTa0mDjxm/8XFwLW
b93LGMQu0sa+mfhEdGjINUu3fApweGE5WBIVWy4nDbhi9RFjlAzMM1vGn/aaIbxWzBExNkooYvfZ
scv4cppdufS/zCrMocyoQe7s5Zjow0S/DSfme2c1mxDjOs6t/kkQCX+kNjizjqfAj5wCg7Ro7QPy
hpXZqM8l1siPS6/3UgCEBHgbuLCTDU8tlQR7rvG319MFIlWj6wPcmc99n9aJ95mHxg14Q1g1fA9v
wwDmSo//ghjz5LL3XknM9X7O+kDWt3u+3jPXA05vGj3cs9vGWnmErS8Ly/S/ZBxU7DoX1x0STyUB
6VdE5Mc0ZvZjdCxnbxKw8hXQat2CyOd5fzJLkBvChnegBQR7rwSFL+ib95YY8oxxtepl5+r9+SfM
0+/g1tlPYQJsYMupzkPXp+mf5dA93j0aHuCyiC5Z25LO8j6x1RgXvNvmEQ+eY4gNzopQWcC6+A8K
5wRkXRy+zSpiuyPPcEDQ5FmLYwF7UA6H9LDuweOu0QzFNpaZPfaFgLwgbiV3DQK+CHMwgl+PuckT
0Rp7BJq5be+QiR82TrAx94wUcQ0hj/SGFpzg8zfJ/9m8pjIYPciyV1vsrMiUd9/jCO3oDOajCKzQ
W//hCZ74Uhat3nQPGQHSk8t2uJ2JH5mizvd4TdPHLHTAzMFXJCIme1RTEzjh/7ab/T1A1lSPFNZK
9kujiYmHHXNEFArCUh8h0wAneBi1SMwftFxKdXOZS8vl1d84zF/mzkzLkYOFbg8gkP+AdLxtbFHA
MJ6TwDFhgqS/j4Aby47+hPShV5DCYotUMlEM8bodaTyFTBDO0ilIXXTCuF6zsXLcqyvGwYWt357y
T7p8K+Y89yWyweyrFUPtJ8fVgOmVakxpLhnajbXYsoRj/pGG+0XK7Vt2dVxYuQpPo3DvsFUoXGcs
tLOauTmQRvzG0+L+GDgZTBBzes6iTtVSUfnQNEqDnyDGyA6e9XqaIB3ZEVDbNlsxeHuVyNqpVJIs
oz7M8OrYbne264rJPgNlQJ9GywmhkZswW1bwan4RllC5tXtn1GMRfifxdqk/Hg7b0HXaF71eBPnE
Ya6omY5+Q4U3TsE//JVOXpwTRkUtC47j9ab846fFcJkMttrozFMMYukger2iDj4/TpFbEUTKES+O
CXxtWgeBOctKRlm0ASTRgl3apAP50siDmlO+yPSWnidybvpmfizRtdV+IpBXm4wgabOCjACffCTm
e4xCL80+ERLhHhh5bOSJjakFP9ZziQWNBSIffyVPv1OvgMwuneIFxb9MaCmoks8y4ukEyyRGnloy
WFCxzx2E6Z+AlZDO+KvuDdKnfJabjyiCLxwiMjEZfZzujA29kxi3ru5YdI5XsiWMz/gsCRZWpBDL
H1cZqCEFMWawd4aB/ZR6ZjtI/khOrWuySD8zyMcs74FmKSWOC6zbac5OKO2jPXT/bvyNwxw82ULz
P3yURPDupSJ5bo7IcryeqvQTKBRVlrKDYbxWe0Vi/CxPGbnbrfAMraU+Ypp2vHWQdp02Q3hiAJDb
hrECr7xf29b7e72VGKawwaeweD3Z+ZKGGal+O1PO9xbVeT8IT3lVxcuQ5nPWZzoUmu/wm7OleDA7
VhWdeXcFBczLOWBW4NfU75eMb2fYMAKgF0TVI8vp4FskvG1J7Ic/Z5rwVab6bcQjA7fWtFDiwkWg
Q4dowJbrZ9YJxvb6nzmhiBYDjXvG2EkEWr5eRDaaDrVaaPF98vWyj5aXzOPTwCNQ6hBINWQeTJHU
YSfLUFAa/2wilOXPmcqLZc6c2TBaNPk14IkxQxZALHu31Cv72qobciow6H1OXqH4ZDkDEzDLnE3A
meGSq2GzywQ/7Pq+N+loQNQVrlS3kItGg4I0+na12lI8pxPH1G/1UKXZ0xHhDd1nRIheQlgU0qDE
Lyw+otWb+EmI3mSmbLsPSD9JXCu/c3ppQtoLBhg5Cdw/E1MLjj3GFkQ7mfA8VzactHwpizoEaEB/
9T1Lpgx4mMNeTIFTwXLj9viNrPLDuc+rIZXgmT8t/WHbrpjYl890Apnwb32AFJbU1GBZV55c2ISD
CNPo/13z0ilW6BETal92SS1uirdcMjlkb3yPuHFW7pMaot2IB8KXIEeq8CdRqR0ylZQ5LJuocl53
VlIWp1SSCTsLnQBDSyZbGt4A+5sFT8ybMcPkbx3CNsJfw3vDuoPWGyJWPsq2fg3ONaKoWsTn72tm
5mw6mWvRKhiAN4vq/mw+R5VhMM4c1l9iEOGVjEfQKiNlMrFa3k0rHueZiL1Q4E4+jgL2PXrCFstw
idfTz3bB5+QirdlilHnneMbLXng7JwWa+lm73viTEODbcxHhqvz58Q54hbCsKtEpouwhxsovYhz2
XNNZqr1ayZfFd9RwAyrXbqUcMX9kgw0WZQwgDqam/WbjTtWovD6tYjsB4A75QDh/b6ZrDIvG6aZ8
/FcU3hl6lyLta2/IrLxujBaeWCnUv5bBE+tPM8IszV2rabHHSJDIB+30eGTJOnhSqDX1Y3RO6vmW
h2gZDLSbkvFXGxzt4Q/oW+zCRuZMl3MKBGse1M+avRRdIoG/h7c1MwGXX4+1HtmTZN4jA6ETGHR7
I02exlFbqUFpYBO1lNr5uVJEDOJyVqCw/HpNnQgO23Qdab3V14F8kzdQ+fjhfGVPwd/5dkgNmKJs
kuMhbKlNcnOONHjBUBn4LqUu4KTxNihCWBTKQc8lyj5mQaxIo2F6NdmxLCJIlRJqAGgA/asfAtz4
EHfcu+WeC4LnlIRyY44pmYjLr7jaDh+HW1TCByUexqUxdRRXuSydUWe9SJ34szaMkiapYw+epoRd
FU9/ylNTalhp7I0TJMMU4LV5cx/4uzkQ5qm9YDSbLD8H0Ytdy4+hpC6UhXuE+KOSQ51lWGA8m83w
Mw4tr3XMCc7ATDE81xTqLulJhfewe0adnaUpq73c2iUQ27KmqVTnB5Tw4Sj3eN8gwULw117tZsJw
yX4qg8Wc3JrPMfHUXEG3VRJY3L2S0IrrTxKcpjU8KgiRlCpItAyITHl2wVMSmLkFctBp+BqenruG
fCk/oU+6yla3AVpqMyXwMR/wtABJZiCerl0PqvDwYHePiaBvR/VOzfBYF8b1PTFSkSAhKpjmsJua
Gjzy0+QkwUTJP6s2zCKeweF0cbXx6z2MW/yl3t3EmcqAcwgjrKksrnr37HkQkQg0nxfEqQWlwnEo
sPNCX4yYo7BjmvJ/im06k7rNICXjJRz8Bvg8ZRHyEkJOuQR+dkrWf5uN0932BrzYl4bqLj3HAx/B
RZJeXYaJW7Choa9sb4xGtUHzvE7oHN3tP+wSWXZ18wOuY3MDwUbZxTK9+tVsbbfL5q9huSekd/mV
1sA0oQjTid7QHUeD5PlNi4LYVDqBt9c0cFS8+d2X6Y5NKg1owLc1L12AiZlHN1vnM8kbhbzqDrUf
8rH3prFxDvsU3whT48L3NEwxjLZ/iOzQy7qBGjrOwsqXMFoIc8QANbuu7ySavZvmFvSEvtWQI1/N
0zlwzhy1xWy33xtNfGky8kd3WWQ1B1mGdEs8jsmxpeaN+5hZUkxjD0K++9jkrJFwERIYJ0JGIZtk
1WkWRPeB/x1WRM+vwMzpNFTZMmWHbMZzCRdwdV6zRylGH7Kmyc0jOJUx4TDDY5wyQLvhM+pzW22z
8AXvl2moObJUkg8c50f6BrCSF8hgB1inpc8TPcLeE3/qyOHIpAjzOy38BQh1hHoiGUhNNYPJQnqj
mdAgfsNZ4D3NW72ZjpsX2Og0YQTQASgUidHIwzsuiPQFO82SK4R4/5XOTUzCWFFmZcrmRFm1ryBt
hwxUvBFYpDavHLk6q+gzsquESdAHUv/hvPyL60ySQUZ/iZsQNk5zgqH22oH1XDQ0ShuDUdhqZKIq
wUejqHN5iTa8WMmjJNotHtTR8Ji06IeYCzfp5wRgNU6Cm+4UITeO8AFhL+p5hZSsrDZSPd5usnJb
cROSdHiJPP6E8Jk3NV3wn/6PQeEn6s07CecIGp6Gt8PI2iMZ8WOyytc+NQjaZMGH4xtJwUJCwuZQ
yqL8HHCMJBg6g94WkGyjp588/m6yOzEdiNPIyJDJ4/WgUTZJEZbB2lDpuUbYtfr+5bhpL3Y5+xkN
DZJLeQ48ZkpkUr81d4L5deopWx0T9GLrAJckh/7HTJQnirPL9O2aS828D0YzwJsrIAyCTYIk/LLV
Z/dgsNotie8AH4NgpDSfuStfvCyylS3UfQXZToJbBVcCVjIL/KfiJevHeTkmZBQlbxSFZIwZCvNq
Xi2txsWdkgTzya5EN013sBb9rizEZ/75yMCk+Fl6VBgM6+FOMni5tIWmUCCnr/hGDj7HQ13dXW9k
8MTTSteJRM4i0TIKlJ8mcYFEfaKHEraUElEC54ng+3uuvdgvhVP+/1X3hmcxJOpglOwKBDc+r863
Rk8RS6Wr3aeFj1UJa0QhKDe9S9ha1cMpdUKryvcXU820lSwKWMD4sMFppOVfsZGgVRwpJvzfbuq9
u4lEDaoWDmbk082r0fRKn82N6tUg0dCWD0EzRGzcKdpIQkIFGgge9u1CZn2N8EXyczrs6kRLrqIz
t/iFOkFEcI0tf9p5euHigNm/FKPt6Aieu8jYwEdZtMluhP8wXR+sWezFMTSWoYyMY97twKLD/CtF
6O84nEu+ck3ovE5L9P0ZQjnoLDWCWfYU1vrXqpZKdlbd4gvuade8MBKRzxRAiJjfBbHFCn0BoErh
H5N1ez+rkbJMy6Mw3KWzvrA233IYwOvxZMHvvacKaYE+BjvD3F5BFFwiUH24zd97+YbwA8KMTSNf
FBx/y1mRgoSvzZCHAi9BD49/rtj2Hl7b6bPr5ITkbAgqPQpKZHTugMMBXeR7KVHap8ZOc1Jsvltq
V4uIe0EFq5jiq+qhGGR7GVT93kNRBYhwd5iobCKWx3aLOLwtTB+cGhd1G6d6jic8xNWOy6nMWy8h
3gUuT4ZyTOWEsRTFDlkn/EZ53FPEO0L32j7Mu8r7PCipIDYj4aOcLw1VU+UvHzr7R5O9WGc0sgyS
fOk8SzPm1v9andQaT8a4nrUmSfEO0FLPExAZS0p/YXesr1r09I6nve2bDpxpPa1j8Cz9qq1FoL3u
yeUkRolvo8kLrgYLlEAKo39wx7VckscayukVX4wzoZKfwOqbwLwzafaHgh25mnFuZVv295wFtTAS
s3F/V0qpKDrQtVAjFeB7AIq5tXJS+NPERSxjhmPChj8B2s7DRIeNCx5Fy3coSp0twZsHfmvrS/l0
S5VnDh/6XglR6HU/7WH4HdGcxQXvfZUxgYJAyMEgHAVEB5lp7qVdEw9NgOf0dN+UzGrn02ZzmF0A
wQalYmG/G5DHMEn16vdRrZtZOJhy9zUG7yfJzk81gWA4tNxoCFSWSfshLvV/QDYWsxgS6qJj4R6q
LnXKOhnLaWG5xulPeSAxh0pLmRN12ZfabZAVsySDI0uHQuuzH8W23jTmla8ZVb2wQTinWcGYtdI/
PpHJ3p31FGBOm3YH76owQRrnuXmTX+xbm1PqUowa98FIVC5Px6/M9Zp6JREfRYs77JlLE4oOirRQ
xX+K+b+E4pHqG6sinuOo9gJagSE+9jaMMNbbrnXLFEF9BuGMKUsCP+OzkNdkEwrSOT+fzggkDPC0
L594kRd/eLsoYHNOjyxRjKc7G6YV5zE6SQYS3S2aIoORYJFyi66e1TfKs0nVUCDcVRRNkDeIG09M
391eycHKJS2UOS+LSY0hPh0bLiptgNzf4tiVI0obOV3Dm3LkUf6sb3gZQP53pd25Qi9H9nTJwgjj
EtizwCmJuhoTI586pbc47ydEKcc3N0vjA0maDKhrvLVhXZB1/VkIlffIfphnS+cOErtV1pVNoyex
7qfP811ohkPC8W7L9YKQlX8Y01nRNJojIpzTBO4xIEFV6Mm3jUCMX8MHh9NS9H0h5Tr2CBwv9Y7l
IVw6Zj2Y4kqq0IHaGlV0BGFhXGq+tGF/PweUHX/sYGEqCnAP+VjFExEidtiloIcmI1ijG4Ixjq98
ZsRFjk1mdWLzi7GxC+9KdHYDgp2hPzCCkBXV4nZCW0G3UboDgqH/oaXGTb5YxaQGAQ4gverdSqXl
vGCidK3mQiEt4P57f30Dz8/mcV6qhPLbm3vRJDtHC1U+75yUJ/tK6HkQzoSifrz0qFjhS5e+OVQ4
elabsM1MGSMcx/eEZ3kgD0IMhux2ElLPJIvP5q8qfYXOm5NPM+MIj1WBWh8XXjJ5c79DcCNFmLL3
pSqOvGfktE74U5UuwLqiFFK7uJfeiuC8Z04cM0vkhyK5MDcvQFuemCQkdiq6dKtlZLuX1hIOgpGc
wFfD70RdNMAYpPV/Yrr4k9r1rc5RrnfH/G99BwKRnfZ3MKyMazPbq70lhM2hPi0C54Tb7KlcyCAV
Iy2tVmTNROODbwVWx0xJysBSt5HyTA90Ox57PARPQf44A1TR0QdKnP1rBBlpywCH7Tcs39bByLZv
pgY4+T19bdjL5sMYuqgm7AfKXxxbGyg1nKtDQ90UJYTdrdBefPQx0vpv00kQF9O7+9LQ0c0rCCkQ
wSPQjB8PJfdondGHWvamiw15kmsYoIA1H2Z6sb1lOq9IkYvz3Ro4kYiOn2/Q3usq9Uw+78H0Mv6/
OfmuKPcE7zjsqFnPhSFbXG+ZSTG2SOow3AradC3pvuASQdrUFiibr1akYAEaf4DQMGQF4J58BSbm
CAUigPmhyJ6AI2kQMHbqjMOk5OD1EdlVtyZ5ShRnRvd/l+AsPu9aQVAobVlLCZyATnVhstKUs7qh
lYRDlHVZnFtxhK5Wq1ooROD9HRVd9u0/VZuKXg7ygMTOoDw4pO2Epjqe+djIlkNDi3X2Q07qTpLv
AL/ccmoaYjEmVNyvC+2shx9wweZz2jgS93/Wpb3ozeZtQcBPlgqMlNMCJrs06OTGc/ZJleL8/saQ
gQksKmakyfhaHUW9DJgqxmQliAK7E+kbPpeA0HKw6oHcnMIYQLILL+CdZiy+v5f7fJ8ckLMVTvTz
m/vS2RLCAB1N+PKNBCf6makW8O2kshR9aXGLFpmxRvusXx4FVtTY7uiJRhYfIm15xJ9DPZIB8oW2
Nlm5nPtj5GTbQiFa0UO3ub3zPS1aNnoe7ZuRHiVfrW5ZTu1sh3Db023BUOAmz6lZmHWq1miBmhAS
I2AnXSk2iOw19/LuoOmxK69Ulcl0Gp2DyAfLpK5LsAO7loMQl+Jg7O5tIuQveMGeW3VLm9k53lu2
Pl/2JrKv2JY7I/aK/PKECmly6fX5gnAkql3fgvBn3DRac783GQUAcrTUawlI7nObz4Xe9pwEFRlA
Rya0aGHNvyj3wwOYgWavAav22KVlI/75v2AqoILKRHUVxxQLac+8Fs4oMmPbkfDJjgmYMXggsnF0
Pg8CO1RtFosX1dxt0qcx06PZH54NvYflfsIAo8sJCYzFNDbvQsXvV9zvNzx71456xykvJwrSQrn8
54NeAZBhzICkKXi+k1Rz9UJ41LUYK5E6MKfWkRaWBZZliDtaYsBoZ8dnFZM4Qxtghy+MRg/W+jI8
1pA4EXh60GcaJFG6/rai5l7sqj7QO5bggGLcgnd8Td/EebRksQAGuDUXF0SJIqNscLdMFWvRwope
IkWULTbR4GYmoQlUJ6owOrbYtEvVZr9PP2YNaUHCaMogifJZIJHe4Va3i8Mwtizjrvp3zx3S24SY
Q7ildxm15Kk1No8N5m3LWnQzeFd5mGFX2EJcfq5qbrdBRQ6E/TSHffz5S6MDs6D9zxzSKA91gLkI
0pTww9PNZ1aGgrvzrzqeES2lze8XMuNsTdJuWPguPQ9was82zOfmIWd7/KfPUk0l4NaadTU9rYBE
7yc5MQWvUoCfATeFu9T6Vk1qSnIY7juFXEYAozP2IxHvB3uoeasUYmfmmSN56anKMstOp5tYsDLh
uxPv5T+ihy5mYPNENA7w5UXkJLhTuVmFNSgtdnInxak+o2Q3NggU5SOpWPcofPgDE4q+P5YCM7zS
fb+GS6kGUh9vUoR5dK7qq6NLB3ewtyTI9haa9RyjTeKRGTc3uCxVxbZjAuURcYy7r955GwZIKqcn
XA9q0mBGEnh/cc+4tMHQoBfSbCgqO41/fX3E7L21mGFXYt7Gv/wDhXdhcKRsxCXI28uv8OAjKxlo
Go8+5N4t98ZCJNh2qa4F4EpALUNInNUrTGYoZ3z+MMuObI3Y/bcM/MbnMTFFaXksqCpwnDt2yCTK
jXPivY2bdHRYBFYPpcT7NGbim+0cDU1TPLSlckLBTtkekgeaLm8u7+8CFkPK/5PezIEGXCJZuoJQ
+DFWeOJ4FY2UOte1Ph7GaWAaYQboPpn9wGY4PLbL/C5Yz4NVIJxxX2yn44GiqFjzpmE5WaJaDmAD
PXR1E8MRd7BZ+7znLe2BiAdMFteKQjpap6Jk+khPFqxhFYbJk2ukMcZ4n5GKNkiSVvYtK4ZwrIPL
bXLvAGahysIQY84bfWoTFk2WDsAQKAqP3jpQFXLLeen8f2XYZPmt+O8RB6MF7peIE6PbxUachNy7
a9oOFOKuduVtQLHCqfyFkIheJMlnJ6OouidIJwW3KbXhjH4ZtHPXLup6MPBmLnwiNjoJaRyXk9Tw
jXhSzBzwP1qfHrlMBsvFmy0NH1PdlzG518iihlpV0m7wWPFjKfBUPpJuR7kJhR1bO+5u3mShUe2J
ZhI3+zUJf/gZ80Rt8dpwFKAANQkINv5YQDAO3MFywynFLkCBfqdKgV6TXCXtppQAqZ90sHiiEms7
os1lhikja3bC3eH9W92QKTzgWwMjyNb0ZHeCbBnVmknp8RF35hJMw9HODYmlHH5MMVLW8GJSo2kO
C1a+qDn8Ri2bCL6DKlWM+cld7O+4NLJ8wuT8F5MwrVPwHArnxd7kU52GFWOTJP68h2IsIDczjoSo
F9IXlNOhMEbMj3yzagsdhqbXfn/x60rpLoJQhFZyPuixM1I1YCbF29jDl5pmVGf7DHijUrDSJ9bS
6gE4xghH5cPaObZC936GkcxopSGR1YDz6GDeO6/ryxDou878v6/jfy4aZ3dkUSA0KRhr4dJJX9Ol
uqzck6Vo2IyjeX5T8N9zBJI1+1AcLizsWXSyW156rtwx20Z0NM7FmS6hLpVrIso7KqnyNU8zHWsO
I7DwcUDJSrfxH0giVDwAfkp8C5a+QOriid4wsTEXRgSWx0BiV5cTbNYG0sfYyvW1FxSPJRwZssze
5dfSG3BGxUzsYHCGV510nUhyFFJR5IJGKBZoD27/l4Tobk8Ln6HgK0AI7u519odYrqhuxmttqwgk
r3ph1IKjqOvL6qahzlR2GoS8OhFMlpTNd8/8mjkJGLTZNAdlmJd+hKuNigXFYowMPzj2cX8pTEme
TWcCLvVzzVcvchTbvC/hEY7f7fGdIVUNUxCRPsMA/pxD6YXvuvlkgr1j80wKYfgEMZaYhpPeVipR
RtZEesYbIprqYVY+iPAu/LVPg6qjXFKG9p/+bRFNC8Ov0xkxJAPrFGiZZ1mzfJKjF+JS5FgXd5dO
OzuLx7q8O8HFSja+UP4GiGkcjvR/gVMtpLppBTdFb4OWNPTsIsWPI9nyawv6a8ORKo9+D0B7BhMq
EXwDgJTBR1SZ0H5bg+I22Cx4BbQxZNVowuLxLrzuAih5JCNFO7tMrT/9cebZl2hgvSXvrDfq2bdD
7MDR8k+o6m15P+jBVjLVDQBaEP1FyBRC0zIq0d0iVLw/r0ENhs7scyo0EiGtmppbEB+VwbYI4j9G
duy+2WKPeMF7fer2L+GEMEVkppJDJFqqWk6LE2BSqbewULM6hqOeEgCSjrZaNBAEgjFLFVrWGx6M
h5HWfjr4ApjWtRNGk2bhF4bxN2XxarDEZs/9xH2Sq3OCBgKmd59kZ8au9iUjFNJdwSUwa7+fCiJr
j/f7S9l/SysDBWCg5iS9uqMjggn0OLzsDwk2B76zKvo1Sw+DzL8EfdDuL+M0PzFi/shQevRJi+6Z
YsEm7M4XwhWS2OPHqkvwN8wgRtwv/AMYA9Bq0k4X+oWfXBDmUrjF+2YhDB4o3IGSnT0aK2k5y8mp
215oSciHOYcoscSzybxAfaQZF6sCG4ddEEWx0l+4O3ZK/AhboDYddEuXbGikG6sQMV2EEQ6BTMcZ
ctSaNttUMRbLqiAOtoE8ed1THBp5nbC6WfaiIyMOzPLAOKFI87UvKKi1NRObn/LK3wwYkht5x8ae
2tJ+zcPZpIf1lg5xcM+f6yr2WDfZ28EN2MjsHpjaNIudBkldTTtNBCHHU+/7TTTyg5aCH3JQTmAC
36kGeyeB7RafU+0J/x4ZuBSIRxdUrwoMopmDjo3JPv4+G34LjlA0qLg7ZlH1AVw9B3moPX88V7Fu
va3DPFSaQ5dUN971IOZ1Zmp2iDBbgy2Vx0htLqu+PlgOMMn/8lF7Ql/ak7MGWUgSGWXAxJvL9+dp
76DliBhli7CnNjV09s0dAwvQLzZD/PqENKPSZkE1V2H+sxqgkxWJMXqTaIVSmAUq/kkqPHSBPtcJ
cFcP/jXg116Jqcu+AY1LRnMuz2og9adurjyKfXaNV1Aye5FdJEoieCiFNSS4OZq7PjdxjP0kzByg
2a0pUnW4RejZELLVVOQ+tOHmmfF9PtK8iHflB7L3tMN6Nt8FD8tHxdhO9RNalRtLut2/BcqlMpkP
3NcZ658+r3hsfCmhJVVsSOwiTqdqGIE1xeoj2fToIzg7do3RCc9tH3ErwG3U49ntZpeI7Chr/sc0
OnGfbairMZyxxiId/+y4OFndbiZryqaMNnwNfOFIqjg8aGL9vcwrVWCo7vPEve4V/6ELQtX05/dE
aaG1sOgegNQ9Payn0hGfdkyej+eJpSHCrn3KWNoLG1aWEANj8NzqLn+hy7Qb+D4t59VSK0utAmg8
Z567R4g5EX01ihRksPdZwbdEOMytU6W3dVJrj+gYefRZr85xNa5UbF6VoLwSXuxH1WToU/w5F1ZL
UPlbFhHWuqKHCeFiujujx9OQtzbR1RIzvhqpYjPO8Y3FwN/OyYZ9CWdgTIzNYY8/Rahws0vUhfUL
NAVUJjPZ913TstkC6/ur8ax800Zs34zo/DUNn/bnUY3szAE8COf38BU7X1r5r5IOGf3odoThlCh9
JYrC7LnFrdDlkO4JV7XTOGyr3bXEk1AB8cmH71DSSW1hBQAHFf/iKWf0nSBXSM8D1cP0WE5tYm7D
Zy3FzjY50qSv+zprFrsgIPRA42qyxThhElY0Dbq79uLMeroGU8Ot118Jc/jJODsKIi3+4DB1mgCs
3whysjDJBFI4xcaH7qCMsVkwlSmGqAZhsXIMB0nt8dAZ65WUH+INP8nuFFwtymlGHrkR1PIteDP9
v4vy19AkeHrMcfEpxnc1JXc6fw6lVmGvTDODAGejg/5NNjMpa2rLOGrUm7gO+6uFGElZeR8jAr6Q
+1taVyu/2+zz3+hoXwGTF3EGlbucLoIsi8JFOhy7f4DsnNah2hDwQENf5RuxXW7Z1hFI09K/kmKl
b5jOmwV1iBgacPI9rNQJcq4Q/vqx7OohOA22cv2vlJWEEeggvqGAH8hB1S4KSMUUVNu4ynjiHWxw
hEFOSWP5hnRIoGfFqSHznSoUlt238ID/XPGgSx4P0CR8cF9XxlZGe2PuHZwfs6nMBhqrQKhTn1kn
BtovcjdPvZmmXRR4b8nQP0MOgDmQRexGU1OQMem51W49bc32DOJB9phRaiuLLEpNAP2CmvNrdpQc
sol3pCJux3cLvVUy9ZeyiA4G1FTW9BKsQRma/FyceVT7Bojjbehhoi8TEmetqPPSwuUnZIC/qGaT
D+fVPXNRomRffGbtD/gzPH//V/bAdEbGd3O+2GdrA3a73BGrDUr6kHZJNnWLrCERldNQHMX5HDFt
qVfRWsYbYWqU9LXWfxkzVOgyu3TW+tlKwBuAEfWPhHpPwsbcKBXUBPtgPVuQjJYNpOJLdvhP2Qov
RbvMsi0AHXN7xckDLcPl9IIU8V5bE65/H7uDdZnoRIYJn04j6DzyuOpxejrvr2g8I7LrVlU7DzNU
JHJi6XLwzJCeHrPMQ+HtNCrc106t1i+PizKGPXSbBuZVMM9k5dgNN5GETJVizlgV49+ur0hXJnCy
aCfaB9OwK1xQaU3AlEzzKWRjc6fEP/P7ZEDWHWnMiach01hzgHtGElwflHwuLl5VWM4guVr2Blo8
txMfdU2LZHc07+9HvmtORt4b48NUAxKSTOr+7o6UadCbsvO6TNCWV7zdCZBtbVXRDdAuAif7bB/9
84G86DluNo4VVJfdoxpki88AEpJu4lMXt7a1sDTatxliFC84RUdRxCjMlUQ4N+IjPo77QLLTgUSY
k81OdM70FRQlZ2EgngkAS70lg2nhi0mC2LqalxLKLylh5obwuaUSlsdvdcr/C9arAFJjyvOZ1ve+
A2Vsn66ti4SMYEhdGQ39mgWEPyAmjqctDTflG0DqTVHSHfomU81o5Vd4D53by0OmLrumrAksV9Ql
/kNpvbV2CvhBRkOo1cmsB/S4K5Ffrq8Yo+X/SAiEHioLX9znh2S2Kn6LvC8qekfdBslZ67IBpIpv
q9U8BCi9rgv5/wtLU6lmSezWUPpMm4NJz1YRCq/6sgYLSW2xupLqiL1M35pyXU1MWMbjtjn2akPg
aP9MCm5fVmwqp9mpDZDE0FUrd0W60wDqn6Irr7GII4im+pEmwBwqRb8azblNnEGL7uDaFSCX/pM2
p5By6soo+pBRDD/KnK8SKQKm1lFyr9LCXxdKZAkrKy1asKjX2L/4lWw5kbCoxsxHOfBSRot+cVGQ
Shsg61TU6TcgSVHsfwspfDHD+YEFjLnjFGzpybfOf6QTysUD+12FhHVcQcMEJZGP1X5oIQ5GlORa
12WEds90h4D/BokGfZDbTylshSxWjTCMvYKsF2raj9zV2D7CBbf5U00lu/BDW0xR8VmIgUddgtiF
toAKnioC/NWAK0lb48ozka4y4D/mf/tXmDGQ70jt7LU5AfKxV8P4FLmRKc3L/tGhLORaEqKbGGfc
kPL8ILvy+/1quMwIFEXNBRSc8b7ORP8ALINbC0bFO3Jy+5717BGzLA4XMVM4Nj4mcxzprWfg8ZhO
u8WDtJ1flYh3486fYGZTUUN7Ao60SE77WBG+X2v11h4d83VHCwQIx0Z1p61nyjU+OsxPJPPEnQRO
U9/USS+xDdJRs0m4VWwOz+V0IIFE28sgK2kVtfAXL1lbRR2daWSYrqxAfAHWTI+j+UbNG3S7Paaf
2Z6g3fxeI4Vr+3/vCohuhQqJ2BOvsJZ2ES4hCCNQZBz5MC4lhb9dVbRoEj20T9v48YZrFl+U9nK7
YGeFo+YLdFdPDTywHbvJ1hAkH8wMpmCBGaIyHewA8FDcKeOmUWgakqErtWQ4EcdHZDR8i6uQtY9m
/FSqACRF9Tqdlfn2zNBgKNJGDMDu1Y4PgjEMZVWAA88X15ELaSMkRe0y7vdbkkzMvq/fdS84ChP9
JTaOrFvHN7H0BmkbTVuJmvilha86D8fJbIWKNlIL7oPDAkeGD4YJFvo90sy2AGNXiHPD3h+jl6PO
j4wZ4Cr+FcMDn6YfmXWOQ40VXHHT9FCQUGaNfGJL8y78Kse/DZWG+Je4dqEL7cTjxEJ+P5exFoPD
2S5hTjDewWeOM4lrKK65wlMS4/mmVvnEacKyQSBrJUAiD7hfvE75UAXjs4DQk+wOXRk7zPkqitiK
7RKJS35VKrJ08sfGjGcKGx5KovQK0+UnIl4Y5F+GqQO1nAwBlkZ8V1PBh8tJpwXK3gcNz/SIfGNI
nbXu4JaJk1ZWvPpcJooNGA+yERqBwhGupHT/M9FR1YqKOJh+EZfGNzllrjyRhkh1Cd5WPnsuXpzE
R7k778ZIztODu/MWXs3knGdOfALsryHr8tdJqzYyHDjjr3u+HDQGnaZM0Jk3ZR3vZRetx9Ec/eBq
3ttB3t1TdJo1c7GroRtwOgdl/URb4KyTUyd2YsrLZHTRul6iVm3flLhnFi7I8MmMaaM8h3XSNU8E
rsfDYsA0tHRslixNm2bqa3ZFWG5iSdSGzzmn8PMuZ4q5jZDDbU2wSxP+rGH7llVINaGhTzu9dLmi
QPStC54y1ZMooPq7gR+gwZXnNdlkKKCCTunwGbn+fyX215ASPyZL7ijg1MEtyYFzMPcBuQlyNxLk
41hHskjIX1z6AFo5fwlHc1GpspJqMHYKGjgPJAU2wxgl1/DJz7dqm2N0DuLFTSpzsyefMgHHazMt
ILFsbpm2HutAuUy9BdMlpgxpQJfyrYWCNCCMTTYU0gnMw1DBM/Biu38uhxdkIPlBGDCMoyPW/PBB
knNTFnk22Baf3YGQLr7W3Nhhy2bWxO871q4dHO9/o9sFd4qj84OuGnOYGwNLEuZxHeNFpUmwcMnu
DDZkbImg37mPQ2rWAwH+ZLMlVlaJ5SE/PUuPeQrKnhSjW9ruEWCt7SAIJwaaZn0V6U9+6skg2B4g
V9ZrhAcYATK0bG8TXiN+0n6nBA1SaqofzZ7d6m3dDSwP/YhSGh43l2TkR1SsVxh3Dzvo9u2TYdwO
N9ZXK/OcXTgx5bGA1zRYWrggp1TyDObscscS1x37NHHyrcmo50EC4UXZqEB/G/RQtY6kTo/uJhe7
IRc9XNHV1YDq0lt5QqjvX+fcpHU7psvL9K+tMK4KFIfcNp7oyFBwqOy/m89XE6Wtp5WBB7P3yNjN
Lb5ot5cW6l1ky1GD0X9weoKjN/MM+E7myMYcvZLUpVFpKhLt6+CacC5fGre+z0RoQoTF6azUjy20
SqDrHnAKwGiwkavLkbcjHl5hOluoMA2QCGN9zLoa2r24orQKTqgmt/o+hgqLCkro/8h19ykxnbe6
x7AjkZC/8qOchSpfvdYp2glvldGP0eOsnr0VXux6hyI+m9CtyYBFpy1NMGptnwdd9EMWSC57bD+A
2ZppPcLuT6p9JTb2ysB3QL5MTBRirE9dSCKEzavj2kVHmAna8Ayj7QiBKVXDyGWFFD6UcZnZd5sv
9t7Uf50fXZCQSh6vUtJpfRGFYoP2JBeAuzJU3hRdA6Ja+9n+Exbdbe40trxykRAqIiJVua0F7Qdz
FzZHzIlPMOpvw8MtGkE6AA+eCmK5BzbXrM8WueRddl2ZVMqhdup+WXs+4rjz/yYN/ewkENOXaP2D
C9k5uOJH8Zsq5JsI2o9iUUR5+n3XONH2WfYQsgi4JaT8xagXN/xvzya5FR+86T7elCIX7SPSd0ZL
opoR/PzoqnFY72pfum0ELbXakOVpbJntCw9XMhn/9ztHvpsUD2eHlsnjagkDvi2IipBlYQxcnyHx
4GTEx6Os/UekfiPHP1NRWq3jUWYyh1XfvlLsp3b9KMjX0ByANHfXQPqvRPSIZfZhaodKUDf05WeK
0GyyXhfGa2a0hjTwDWpYdNK5acOd9J+dLdeKLqI+a/IEe578ojnlFiDHMpicWglwqCjH291s4I2m
ZyvXQqHbhFSfXnU1gxRSYRE/3pAWfmPpEqaoJSzqq7lxMi8sXynjoPSYIOVhTjlyfze61UVjF34m
c5xcF8gvtQCPTAUJV5E53D1nEOeSU4miE3/KsIIUgeFs6nRXytjd+0w+9yyFbCOVWf6AoEYmBSus
8oygrDCIhUJ3ZyvGzt/Tve64uARseVhY9Vv6LZVyZ1QzH51Zx+QEmN4T6qcOKoh4gFluToR0U7S/
2LWsrDmxuTZ9vyEX+XauJLbplmKNl2g/PMjKr3IOY0CMiYbpSRgS3+NWM2gd+PEdtGzXPzg23aQz
FhsuKI8Iw3k8mITyW4yNO5UqNyWO9aE7cIQKtW+FFmeKE4GmmE2iU1NgFiW7xyaVxp8/a5VsCSsN
6xcuKZzrEbuAygh4iHxW26sgJolQtY8r6FjJoCKCFY1LfENEfkT+JJqI2xKu1hwIGsnYuTw1tFqv
ZP+6zl3QrRoyw6SEdGYT8vsu+O3ME2rum1ndh5X4+/iOpKi4LXn+mBVRyjgD33jjUKXbHTevpK6N
UwuQwtjictJVuAkhzuxgKE022+MsW4gaOBDQ3o16VvSe9XS2wwaKjwYlPl+iWVWotBuoLaPZiae/
ZTHgXgvEhmxy5cUtJ8ybf/iLtEpvaAG3P9ZILH5tCpAKDDwwObK6nDSuwGHXTGAgWvcALmA6dBTX
FDdOh2uZVntYKC+1rjRAVCBUbc+guvVIc81uFPpwSt0t+yuVWEvIUqDRBLNWkIqcHqmu2S0CoHxH
2OLsDV+x/fmuY27l5unuLnoVBAZHw4VvSVhhsh8omhhHrP/NdnNNxPimZ+YV0SJhXO/kBCM3Q0AL
sjKYtY5EV/fzg7RcYwGJneHmObQeTgJ9BDi3INJ5bwu8luGNq3FkvghVT447FWjUggqnyQxynuOE
yENJrfFsGmgrwVjPwpJkPoS6UAtQdZDtNhZNIxIXcDpd1BcMM6GW+VWJh6pE5cTZk8pRNXegpoXj
RcaunaCvPi7XXMY2MJyV3/P3CoNPsIQgHluCr5XcTKSLvsVrJKX05Eanu4or8QqnryWRjHzDC4Gx
Iv8XNqdVq/tqmoahRMMCrHNs3CZcD0xxaI5P2vGUuA1eOY+UT2JvEYROIw6NTE3EqkLQtnr7lPqZ
RWuc7gRrihk7R4R4Xe8uwvxZZbl9I3Sh12d9JFxh6rmUnrT89W/SF6JIoy/JapvioN/kVZ5JxPc0
zWgchod8NRWwcVRrlU0pISJ3MxngnlbuH1nbOgiR4zZW1bDwgbbpTfYyQmVrNgD4ISrnqQr5hGWQ
Ux+lfTXDvd7IxPRGqjs2TfwG6ain5f/FRvFWVO5oGX859V8WOygFDduK/zWBhnXrdXzoYc6CzTQk
q0jhe9CVNTrUcsiM7M7F/QrtGfXVZorXGdBi3gWHgTeWsM5XjOEjBumYFRl/UK34eFeaUYReUZv+
yaUILkIH6r4Ge9RykpOJpJV+gjlk9BkOBwLxeh+lsfA9lFntNft6ivC+kTwMTh1BdN3p57yAjXED
N282aRevchpN+Xa7BC8scZJQLsMIE006daGgbFIvLOkNqv11rcg6P+oyOQttFG1SqXhqVWBluqHC
eIEzyFg0ricdY0ZBKBvAoCSx6l40ZD9A08JYeabzi0Vd4QkWXQuyeyhev2SbKij1d1rm8WgsZMlp
xGMrqxK838199D0uMKBdwOfY5H9O34BFa5dqAI2khy0hwUOhbXrDOQVocY6fMaWGyvgH+V20il/A
YmxkwVI8sYnv6CBUGdrQysi+FkbA+B7PIfTyYVCKbc1ZxUpMrCZP0PgLqTnAYZHnIOawnouWb8+M
TURoXovXGkGLbR9yeoPHomYfBOSDy1wTJon6nBpQCjS2jdgTm3XVRv3q+zk8Eb6DDmUT4NtMAq+r
/kvFMF/2ZJAM9xVdP10he3QqxG0Bo/S29OyIJPctCm+B7KF09mz2+cloqP5xCSXosRV6VYQyr0YX
OTJ/ATbA+Sx4XJCGYq+V6LMDIkVjhoteKPemxYoRYVKOPMJZ8iOxUnM7HTtJF9cBJclcoxhZ8Stb
WL4PtOssfQ5yYLHfW8o6uuOgPVvbRjAMbx4FfQg2xpWyDgkrfVpaEyg9QEuNBtDhszj2Dr/tSPpE
w3bcI69nma3imM9zgIOw5AulG/B9mU7fruncaYQy7goVE111SA6b96jZzh3Lm7WlhgyMNv/uzuIy
koC/vSjQUlRAkWF30UQxN/8tvWrggonHSFRksS+pbSUuupnO++BPjHuUGq9nzkvmOmDssbVJIBWR
O5VPS//RSXPCSaNvhj09tDmkOSBNEkvmkbCG9u+BU5MMFzl1bzyObWEpxtXcK1THsAGJTXgopPCX
SC8UfPTRVu5Fx/zB2xuk3ee3BN6V2uUhok9j2/bnrhd7DHlwc0p3/WahRLzmnKhVVTsp/dS8kNZI
9AHUciCAH/Vfjjxd7//S7NTHcZYCFGQijkqd7QClMXw/+xWzYAHatN5OBkKavaWuwwDtIlzqqnqh
564l0fg0AwtIqw6QtD5LGcx/JOH13579bOjuhW76SyWlxIXuD/iepPjSrDzhjNKPy9J6CCkXwRpz
8g4VTiE0xhtlzyeMVnuUENPHkjsxB8C22PQA+6t4tWAx4qaMcWZ5ZNZcGQEm37dC1brSjiLBESjS
fHnf+yf8pDrughl3Ci7qJFN4jqgYoM1VxyXUNqLcDQzFJs39nzvRQqjuslIZcyzEZp0H1AdgPMHL
w4RdvHTFbzFqQBic3g5VGxAcbG8WIEzTqnaSpyXPhjcvX0iT6M17PU6jzmSicvs4rJdsuzSxsro9
gA5Dt2BWqTr2tw7CRA9sFgL6B1qxcQla4CGQigy/p1/1rHa1ZoPMVvJa2qLJKT+zDzqvWPWq9xr5
U2VfZ3y5XEMVk3xgVFENfnm/Dv9K1T0s+CPsQ+d5/6inRCknnEALYWaCRZ875ZXS1vLzovEOYN64
x6q51tcij7Xt/qgga1mTqU2ODz9YENbkvEJfOvmlwOVzuUoDVPNcOOy6LE5m5vw8hSw2YZSs0bBA
2id47alEen8EGkut1km8OaAeYByk8elC7l4iKBDDtwgzmkUWSe+Ndvj5UlONkhErakhVluIrKdqD
9YqnHsAcYlTSMNSuGhnAOeCnz5o+iaslh8pJp147g+xBXTzBZWGslaNmJFS+9Ben2SfZ7btfwmTP
Bman5o5jOPxkhwCNa4z9ew6PuE6T7Wu2Kg0d0aAUnYIASJdJHt2ahAy0ZpMD/E1be+soORdy2qmy
+YG8pkowafHzzKoqObnsfHG5mu5sbaVs3MgO/HfzNnNoi0oAWCFAX9KiB7vW89qB9VMztb6rPvFy
xgC7CCvaeI19MjKc/YVTQ7ME3+K2wOBHwgXw8LpazHZYGczwrvdXuEk4Vvvs7u/BYetSQZXmd0A3
4YIccjVlsfUgoHLen5Rjag0jUMRwetI0nGuzVHfWL8pPeLQODelBwDBw/lD3xYgVmBGlfZt1foGL
d8HL4p4Q+HC5dVOTq7iXVIJwgThNC8kn/nChHHO5/c0RoPtilmzEbfao/Evs5DG+uM/chB9iG2Ql
+8vR1Ki45Z3+oL2tlXZD5wxB+ckVNRaNw35slkNc5JY5DFSLnZwxtV2rjiyQrjMu4LBZ1eOOB8p1
aRynIms0uSQl71183eQMgC6yP0Qyp999qtaoCTlfLK7qgPIPCJc097C1gvbTA2ojomKQ+R7pzwEK
5Y3Zsc2KgSzicI6zEY8L4fV/fBOuVbWF4wyzt5vivu/knxsmrYb/SAP4veNuNGKBIWNJDwtArFR6
YPerNw5jk+KD+46d1RBArDSTWalvLkemPUmK+9KY6VogsZ7nVNRnQ08G6byUQuzgdLJhWIoxGcW+
8yiEiQ/wdiUigoa/k55TFuW3KHmjP0TfCKs/Oygs8Hu0c6cF8rGeTpFoPijmn/hYgQwDJHsbNBxH
1QIBJ7fqFMx4iXN3nPHb8xuuEDNujKW5DTRZzWaWyixEBWpNlINzJb9weB3ifC5p0FyMN+F0x7I5
fzHWXvdAW49cFxVRC3GERcAEGVKsQpIb+lailhBW/0JZrcITVtg813XYyyMTQFUuYCvVX/eQaB+V
n4CFhNR5nDVI7nEx7NZb6g8oMPFRla6rODvrjTS3RlZxGqBwPJJfGTshqIoL3hyjHBVZdnCsSRd1
5sIK8qDxEJyTpHPvlmmPW4kiNe8P0iPLBMSjBcdeWSt6uDNYRvVov6kuWMWA84qt+0KnR8/8+XR2
W724gVh++ctfeF9mY0NugrnGWDGIFCi/XO1NJJxw1Ax1BC2jvc8KLka1dMl0qHfBp0eS5b7A3qiu
mmXoVRA+taVjLvFcLYlb9qhlHZCOROr+wmIJ85o5XjedkGK3uaWXwl9RgLbDfi88MtkqDiopCAHg
He8VAAatJpNuM5cQb0bqp/4CRtn/F5rbWWP2yODv+40sHdXF1WS9no3BxcNW966XMskv5oGvkyZW
6FbBdY2JdL6xZH8FM/Gay3K0hZK8bEBeo49jZ8F751TgRTtjgcF1O9UpMEKqvlsm5gVg9W6+riQ3
yyzsGsxVPzaunJ8f6YAsmhqWbH3WcezLwmc2Z/5WbNXeYPND72c+tggS3OktUBzmxH3kVRz52F/7
F0j3INMpnv2D+Qx+1URuo1t2zR2GVhma0tVSrTQLSBQdyxKeB14Jp8nUy2IBGFoP37sntBOr8oyU
1aPCRBrV12y1rs/7nJniDAKhuXNoBfbORlgoV/VQZaeqbci9MUaSAh7BOVQC2BStu8/3M+gv+bqw
rfBP4JFp6aApZowT969+Xdzphnm5ZkBLWbMG1agl6GtgOPbW1U1xyS0e8qKQYGE3LPONTau1jhKC
GcDKtE1IficYAu1ID2UiJ6c60cw+boOuQcYa3ZNiOtfSaz+AqkbiTDijAqc+niP0U9nfIbltUtPN
LGjQtWUsSKm9P3P/cjEiToRKci3M/qscAFTrV0jxVxowDEmFf6T+1bMzpVIGkUu5LdApwlDoamkC
Wt68El71sYmXhXhxT8oL/hHmCA72j8Lho3o5wvoubgQ9lErJVk6336hDg6smMSdTA2lVay7U0TBv
9ClSzdAjrSXyt+nSLBxe9D2JvL6NpSrcdnwaC2hfZjE73NRfqcJTULSjP2eE3tEYhJsPn4D4Fh2+
SSr5zxBJ9AZbiTnNKbGKYW7oNTh4UydOGV9xSIHG7gt9nUep0bum77VG237JKwz75WV7FpU5zh5R
ZaOtyYZlX56ag/m/HHs6bZ1X2zaEkl2AU4YmzOIcq0q2Onjmu+ajt3RV7QmyJTnHWky5K+AEUF6E
/yeDfy3LQwioqIHZAvaxzclSW2zBrnFCC7Ddt3draFs//9xgclK5dNQFqSkY+NcO2KKt56ehp5lv
OntddrWk2i6QCisOdr5TppDAFKGJEhzz5IBkUbE8ITAHSiJyFo/VZ6NJklHpFfOFJ8V+T0tE8Hiu
JsNgDEFfc39zgSFEP7o0O7wl0AjzAn1ReX7iGDj9sTZSiQAVBIQ9uJI1w/c8t8VBp9jIZpt2gw9p
V6GuhqMtKVIYgB5X4HaYhtP8KcQqPwKnGHoG3pBNGnPqEWN+61xTLEBUl6pMHcErsz12XjXKYGW2
bYKRrOStV+HR6Um/cCBIXWGv0fvJL4rZ7Z1z9cCIcUMlhBVF3vDOC2C5LuBToH1ulnPtRGI6UmFd
DocHGThx2z5puNxOD5u5UrdTXtAFZuuiY98jAdcI7j1Bg48lGXH9mG/GmaDrGmy3lPNoXN3quaVf
/JJbZdNNzluUUx9uCa7Thx4YUuFlsxWwPjeMl5S35jpiqHw1Qx0lq3+Hz22SROBiDGH3VczYI9lP
HqD+h8PCyNzj0dJJyW+u+//H0MCrqjeBqEW5N9e/Xu6+/mA/BvjL97GBSAe1hdvjyAPuwHvIgPlZ
7/1VJsst98NqOPgNJ69UYd7eKzBUmYT0O7LTi0cVGhFzaFnjS1H21ahTx3talsdZYWUwVX3BZo8V
ZhT2btGHtZZZ5GKXmbvuPg4GcDV2/ayGdM7mqHXLkYgEgWHA7Xnw/yd/LyGX9+5fWJ/W7U49kqWx
uGpFYBqLDIYe1dCJNKZkIUfsKJEFk30SgjrjrI17HCUszr4aslroNaL5n0KX+ClC4xC90D5A2koI
Ni5+3nM3C7eTS1GILI29fx2sTICKNzaYNacdGYpjpsUt41tBJuk+d/4iCa0fitRzBY7qNOHviIbT
a2OcJb1oT64b7lLlR6IoSa2T7QkNx6LQZwmSlTEkhIZ+RVzZ/Q5rtiyovySBIVrnyexL3q0JPTak
O/ZsHA0IFIsjvpqvcjFuNvG1eBq6jdAxUNtOD8XD7TC2UXgUfS1Y1a/pnyy+X1M7Vv892REkSoUF
yMoUG59basDjHX2U2rXTY4Icjsu38Uza09YIslMQuwWB6QCudT71Ayt3D6YqIdY+wallioNkY4Hw
v7BsVCKu85kAq/6DVe6uYwVkVDD7TDX3HTZPVXW8h0fHzFQhG+jZWrNB8Rev57NtKYON3pmFyIKC
mpIv9LQyJVJP5NVK2wwkHI3DfEe5wwCSbJ6LslpjFAFzkXJ5z3PiQxT+Gzydd6SWp9cUaWo7HiK4
O013DAyQko64J2ad48kJfmmy/uG6lT/qBFmkNEMOGz9ofKup/53oWV26eLH2s1qAlAqNa4LkiiU+
kvsT1qNVP/TyjUEwO4dBcwDlQLyYA+JtKWY8vvhNukk7rfz0r2uKtnuKoH3GNTXwdXdeyoc8MzQZ
7VRvUZSdWuSdlSR1ALl6gbz8prw+ePXEUNBtBNK0q9Jljchdgm4MY/IOlLhTh9YQxFNgmJv2aL4/
Cdlx3Tk/SQ38NzVTgNo8+ap1BQcDzR/JHXPoFZToTwUcZM5uv3ASmWmP3DLuWekpZIw2bYu/Xfuv
7dCS08ZB/WFOusazHoX5eB1swpEB1PSfboAP7GsGpSefNRQ3oY3/iFZpdJ8wjWCmMAviD27xN7lQ
8uIr3TpZZMSkom767KxWMvkxFcmJRhp1BCRWA5Zavem9LuVngwhRCoXjY9fU6b/3QPLCWIckqN0a
MmvKnexaaiWyH0N7HZG+GlwGiXJWRMR6u6b6K7oRpR1U+V4mH/LFzmA8X8q05o9JWv5Na8Yx+nZP
EJvc5MH7H7RgMkk2iZG2vvwZgvA5H8GAABtlzMZLV/t6JbZKpJBTiyywutlzsf/xAwFXzwbWEJ0V
pe4Wiic2S0cdhKbUXMoq4ho7hD5ea7OnGeF3NkvqRQR5hG2eAbbyXdRYBknByw+D4LiM4j9ToK9C
93ZvvGJTQRWs7tLYByBj651MfE7JfO9e9UpioADwNrxQkDQ0YCDENNIy8tOriJ6XhVfCENk++RAA
prwa1+KPALA2EI0N3IKBtM0e+yNg6icjyEdeWRR+VvFVbhzHsYlyKRK0U9Ws6tqt1vijIUi3O/KW
C8SoeJ9j/69fwhYS792xrMvx37zI0uTDNDJlWFuDVUpKPpyALXOh4WjbNMbLqUDXsVm6aKOGyw9R
ABFId2vUxVHsUoUyvw/V9Pvty509GAmN+tY0Fj/lpg552Cjjim+twQU3u9gz5mWHppr8jx80SJ4h
fPBomUBvttZ/J5TrHZtUkbcLiVsqASJtK4NtCSO7hywhUv0U2FamggS6ds6vweiKFWF6/23RqZMn
GnpS2MEkfdHU0qUfcF63aaspSvr8y7xTUe6BdM0nlfulOks7cXZHaCJTv55S30pVi8eRUbZLuXtd
s6mHwhCvlmKwmG21byt+2r9fhY9GSyEIetfvP0FwLNPJJ7FkFDVQ7suAaowkso5DmFIeLY2a2T6r
KJMhwbrE/XgG05zqV/R+V1krcoyT3NuSyFd4X4Uvk2uQmf7wFWgy+F3Q5i/0tIHjj82vr3nfvDWX
ul+NlV9nDuKL1hTNojY/sUL0js8itMBECSHRh0T8UOT7nJ+43q7xNKku48+Bb+aRrwOZv5pAnKyq
UEbrEb4pRzmQ/8X/eVOhnK3GTTKQKo3hKVtGUPPz+NyfHtwxAqLLwos9P/Zyr14YcV7CBLfPjdBE
W75A5/a7Kcs7qycjVm8TrJulCGaMztLn/0n09c3bTH8tSqI6z1Qkn3Kg38jY6zQ6j7uiXMXM96nv
gA5quf/3D1xuphXSXPZBAlsfWICqRukoCYlIbWgSQvMhi399e1jls6fLGlUzLU/kbs+EPDxG0WFE
VKlZAG99bn+bvbeLQi0KbJGNNxdeb7Ux2nwM1nIh0ev2K/um+1JSebp3aoThUN0ry1MwWltFRVyc
kth+7raL1MjeJ0XBetZRtoHLcY7NmXp8u3yLKWJo8lSp1I1MFtWPG/0mC2GKUr51x0dOUYK7mj2V
cV3VfbYhyXLrLOxQ7b+DJiQd7ZHUlAe64vmRrO9CBMLwHeWokrZqDGK4hVw6utgAGTtz9D6aKgrD
Af2elbDxS75Wur92e0N8l6ZBzsAh4J2M/YDt5eYZG7gFgBlx76CRGmyVfTQr1G+Szo4zRIGlP3pz
TpxnjtY9rzVX+mgDBPr6MmbRUVs3eQV2eyoeLih4MLPtS3w2jKMP0mIBwvGM9NC4ciXZ1BbR0Xsy
zWHfVWpc9N6YQNp0DDJUDHabCgwRS/aL0bbF2KGvmqb+zrgBq6K6EIn8iTURle/yPO2XX9QK+uea
UsURtvNDAe6RTwtZHpWfE9fmmYIFWxtcazGT9tXcMcy9HriawPFL3KLfx7VzKmKWYN6M8b4rZVfm
Wx2GcBMlfP3NxYvHbuQm5p1ydFvttCiG/70ux4jsRlW/r7Jp3RrieuDMzo0qJiAAQMID0OMPCVK7
TVJJfnkobzF/0pUCXqAnxsEVNC3qYj/LkSNEIzIOGHYRw6jMZHak9pAVY5Qvkjyqr9BYqJgHGcDl
ZPxYPj0hLNZSEv47siHlZGl3oxHepf+/FtdIkNrFzSzolVlF2yHuC3iIZPePfQOfB6LZmWSrRV2F
oxMVgVfuZha759Ynwe9BaZh/ispFfJ//PQvcDS9BhJR6Y28SK5wszaHaURyBAz/d43R2QSKB0KF6
FrwsyJbS+IMLFCIA2v5YYrX782gxomNkpG9VAp5ffFP+nPNWXitl9fTHr9D0sMlpolvGhPddEfvB
1VaVHQqX38LEwkyA1Vif7O5/kgNrGXpxbs4y3MoGjRXD6g4bGf4GghwjReBDpd0ZDtTzeUpiS+Yx
vWjpyn6qr2xresOpe4DjbtpepLpmuPQ1NPfxdQHD7s3w/dm3WXqdCP/e3Bzy4K8Dv7yvJ3AiNZYe
y9R46uz8NQd8MnO5MbOQ7CQy02vOZpQupElu2TVCrNtOOUqw53xX/YoGawFr+/IASg386dx2bqg9
qsQ/15+m+X8LWrMVvp4os+fPZyvlosNtW2FAJXy80o87knV1k8fXop3y7hXjUp+M/HaB05ib2JGz
YHlL9fyNhKMDAmURXJS6UAedUDcLqWycveFt+LX+6VpMcfaBhf+lCbUgXxbUw/jZxyTKvhCVBU4+
bjB6QBYfuDNbGSblWQ5EdfUb5rqSVe69m4GwCzBHsONauMwLHSp/RhIrCm/yrMunO9lFTx8RpUpk
QTFOH44sH1mJt7kNHiYKPJvcYRSlLcyab96FAOE0uNbnO9JPwJPWdriG/2j+xqV6UAjZs/HRHHg6
8zfG4DFnnef/J7NLmeaVxNGucXBsal/UV8OMIEOpYrCf99fG12ei43GCvlRDG+S7/3GJ8AT6g+Z0
wOxsVGIJJ5QDNr69fTZEoHndcITh7wtJ2yu/Ga72M5la2jUUfMcv0g3+NsiX2Cr/vVAPb0vieieJ
58XLURaXfPon78dhc5hpIpgsL0woreqaRm2cK2zPJ1e6ECEbYV7lpISge0mF0BfB/5TVReF0MdGa
VEcGNyFSW2FZp0zuYurepeX+vv2Yi7vfC66DCGS04hSbjRjLgBQHH+/QutoXNN8/bC8yiCmDeI06
kE2strvQ4jfOyR9fV0GmBQHqvRZ+AknO42SHFpM5cetMmZjb6JCW7sZOZxLhMgga1cK89NYzyUTf
svVOhH+YoNH9kEmUqFKPzYcnjSmUqamWg/5obGsM/WItIbOLjbFEnfDpCTG2NH2/4mpuMEstu/2F
Zlqd0BSbnCHLg3M/ywN3odVduASsQqBTv86bXCX6uRexJn/R2w58IJr/vbKzCyFC53YZCHBtGpDg
ssoW1AEB3R64vgmsGP378UQIgo44iss328u+oYm9q9pjO/UHmz0pjQoce8lpfJBts7tMxIrl7pMD
sapT3eFuriKJ3ETVGvzyRiBHs+qGH9oCHlqTaLl+tYe/00vFpJspIrZFPeGVEvmjC6S3E1w8i60i
DNY3Yw5ich8sjIMKqQ4bnB07Bnvih/6LCJgmjSdiGOTlRyN53B46jBi2qYwRHAuaPHwIB46xsWHi
NmSdq4TaHrSQY+lt8fMS5HO81XqYngg5zl27VDHQV8bvq5Vj/rCdB4SVeoHr/xn0uBya+GDoe/zT
OS9DVQ/aaG82psV7U1BZbUWtx5AUXGDQF5l/UrqRrvIqEAigCjKEW7Ch1OHe32h81ggTTAwyAWOi
beq4LTecEaKPK+Woa88qHcdXn3/RGw6utlY3Pui8U4zwln5gAkOaS0taeTITYxQG3JaJD4RaNcCX
c3l9WmUvyCZsg/VVGGV6AmrQnCQwh64gWQ9obbIj3gqdE5OKGnVKSM4ZZQZaH5Z0VfPcDkszXHap
zOUD3Rnl8qyhtI3FUI0vLHv5ge0gE1rVV1r2Oi4DKTV15a7CQhriRdfy6MAy66MesI2ykyjaZIIX
9qDLP8Z5kOhjDkSluL1SFh7zhMbAgVyMwbaC1N68708HKB2QijB65rPgactw1IbqjWCAFFr/gzY6
5YgZc+Z93+HeLNrwP+2UaWQ13xVkN0nWN52JNFU7ICWP1X7PfjS0+8m48lD5Kot73ks8UzX4mEkR
mD6hgKo5HXnLCp8e9EPgURnW7REc+voOCZxCDhHqngszkJ4jQOnFXeRZpmq+Nv5xa+mk6A0F4iEd
yhGCr1eWTKAHFrRWngyDYi0prWSsFg/tNv1kX8wp4QX8VMFG91gH8kV09GxKFbBLuj6bSmTVm9Q1
u7qnUZJUQICvqEYWdjDLwNhea5hRAZqHgLXUnQAGMzQghKZEt73pb0B+0Pg/xj5eBGHsKJnG6JjA
BsO1J8K6l1rQqnYyxLx8jat+sfyfAMJnxUG03cyQlEXZAuL2zAyeRhdPI1kDoJEzEFPKUXLc8G2F
Hoeaayy+GMPCiRoeTK7NEHTYBOvwhJziV+LBIafy3SjEPPkcpAmd3b9ptNib8rVW3rtajPlqTpm2
gEJUCf14yyYqu1F2rWAZdzstocruqVzEe9klFdSJzeqhiyDtw8Xa51Wn9K6cBvwFF69v54rYemZV
Wwc6tbJq+vZx5iIR/ekaKWIKwEL5FvViChbjctOzCo5AL+em3dW1rKp0SI4/6GzPsyRZpuvbi4//
9ED96DtvqAsRvx29LJzShbwcyz+jKepMREVqpY/oGHQPDeNNvG6WxSx0Bs+FfHMWeiJ7dKHgWoMk
pLPqnye6BAvZdjyUAZrUhGspX00LV7s063aw953Xtr9e5qGG7sjjOdI8HZA4IE4bC7ZlB7kALsfq
GylwV2p3Gi2/oFFAM4UfYFnE0z7IZZn0QqYYFIvsQ6uUEdykU6T22YmJnZqbFhUPbT43TV9hk34n
1yDwBKW6c5eZDwi0dd/MVqQviEwBS1CLNh01vo6Vh6GLdJbyd8MiBfIfMUB3D8xcKiW65LBQCIk4
TsTAPc3ilONSAx8yiKhAB0NJKB9HL5q3zXzlqXkKDzVlhB03kDS2/51LROt0Lwl8PJaioTHUW6kL
HD2/tyiCE7o+/Mvxd+ltKkDSyUZb+5EnkTB3F8j/JoW2cSIRWzkYXLyoB7BY4Vn3WZKFhXCzzm8u
sHry1z4PPcVA0Ah/MUcXh3XLNX8Yrxedm+OUkiwmByQHQP6ppuLUiCfQLEesRO0GnBnEttbxm2l+
dqnQCIjYhSnCg46sW41R1ycREO8WJdefU+F/SnKCwCespfZ80yXHeX/7K/Bv6KQazzenKDQ9Bkdo
v+vfhM45PpjAjRWa2iwLyi+SwSRSbLwmrJxHg35/M4l2mfONBUmPRFsAknkwnk6XV9aPhIU+RWeQ
N7vED+F0vfx8PaBRJXYxuxY5qqA9mTUw1hwue+IaKQUebwPa4gL+IFR1elMCXgM0YV5revng8vx/
gZIAmi4pfpSpH6/R5ZYL1FlU54gdjMp/d9h+wrPTWHh6dL6d8TZhurSMTZdpJqoqSKgNYWgp8CDY
1G+dP4v1KwjeZCwYQZiOHjIJIPoLcuxy7GX7Yj+tcXc9jyudLNHkO65KclU7VZkUypjhS1R1b4ZL
YAr5q3vZroA3lNA1QosdLDiM3u9sNYKIO4jQ99puLlR66luNo62zBpQ2ODynHYsxV1ovhnabKXno
NIlPNzUc/C+9YuWoZOSmD+rXH4GEI3Olws7Z39eYg+I21n6MKyXRartDlEhit3gCeVvZB8UK+CY6
eek6TGBhaFDaq0VE44FmRn/SeyvvFOMY8Aawon5j3bj4M0Q0hGrLiUSq5X3OuoO3e9EuTu7R9lc2
JthmPLFjm/IGA6UnGIPwXBnVPAcE3J4a4ozCQhoKBoB4vqGs7lMvfyNYDjd8u3zmXjBsdao6oc+p
qoDNbzMS61OLmdOy76Wdo9Pmr/87CGhiGmHlvcDBoOWnwOe445c86ncLtxcMmqpQturJQhs3Mh9P
cbb/gvS3dy1Q7AooZVGc74a8htv/fkpAcq7kw4qDGWc9GeW45wJuxsb57Bh1QiWf5y9Q9xus5M0M
dwDdGTHxVdGn1wESqYlZFaGKeGYseQcMAG5C9iOudjKHEd3vUul8VcA3I+eglOVSfHLZqimilNQx
nVQ3Ljgm0VJ3+8MxkhgLqxH9yxMqt0nAXj6EPEx6n3jjKif18PzImMHvXjKkfdp6Kxi/xKk+Z8Nh
R3YmVTzE4s1utZ0S0M1gXIHlGiDlTsiN9qdtXFlRJTPrnEHlnrdzvseR6g8SprSfJ/9M6imIe2qr
z7+L9gYgtB7rXVwlVxPpT5WFN8UI7WtBl0M45T2FoFlTALPyIi5vm8e+8pXX/mI3OdKT62MLsNLm
QdYbFen9SDwvb8KLl/um1bXGKLS0VGMbQQvJMIX8P1I3swmmUmRNq749g8UC6kCrEREBULw8FCzA
lzp/u+XXKTRi250dnPyFciNEeOtRlrWXpocGBWpJDtSfPSa+231q1yRrwzMpA73AA2hluVu0z1Q5
dFbkGmXyR58txriww06ay/c8qNSfqDJ4DjcGAK68BTqi4291r14o6iAMLS9G1cIURnsQDyxKAv/Y
6XUc2z9dG0/Ag2XuppPuydeiW+NhH1g7PmcMcDEMdQjQ7xAof0xmEdNUiGxNQwUj7+qwJOVqY08K
beDedU+LrWQJfvBZKtEl9JyWq7KTvusjnWgNuyfxlx1WeM/ZWaeKmxE4PluPF3FNNSudvPBVfrS4
2XUNkE0GrJ496Id4DRobSiMY1v5y2bRCrLWGEgxwram7GhcCV6AKZ3N9XiLxcBLjM/Lortyf7gGs
bUO4ExX9DfuNKwIcXrz8HLI+pko/St+F3YcBz1/rxfHWsxI6JkTQSQmXRr31ytholoIMAaSYDypz
i1Nf9I18lNPDioGiitY+5T85w7Y9oCVDgS+9MiCh0ZYjXy8I7G/rG4YBss964sOZNvZVTMUHw55q
yWNfIAdWzBajMZKa3Ae4GpA8dh0mgMc4Vxsnt5AV5eQjgSmzrSIk/2QJFkOS/1lcMLNrVOAcgOK4
pUNhb7nriWUAPlqpI2vRsh7W5Y39iEzZ3WU8E9V2jIqNbKAvgLWY6+10QEZJ61x9upV0EsdBfiyl
H7JM51noqBAKk+hd7FJfJFHtiYT8bMty4tniOW3zWXgzIKjKiwNyb50FM27ptExzKx5qQL/FzeqI
I+m6B7xHBE9GMiZCOHCqV/CiDHDGiGEUepzLqsi+C7UiotTZJsnkP6epaeIDFlC4ZOnu1rMUVQTa
nOOLFepieDgVD8Zv6rpbOFTw1FtRQ/8mEaP53lF1ZlprNVvHyqEtde3lmdzF07b5JMvCuYkAJVvE
CoaRMULU+aBQFhYc7rCLpTrd8myVFrfsxej6A2cgNEcvEalAUT44ZIhbPvTsPa9Lq/K/LUr4wIUq
zs/LqXiU680nrAWHp0x4AEkNwOH6uEG4J5FjaCc39v44JCGBmbnApE4/qnWYwjzWY3hlsJL9LsuQ
lmdRMLoQ1jD7PzyOl6dAYAnpQaSY/K0xHIvNL6q14rFr0yD+jF4o4GYFECYQr8dxXmcYPBSesXUr
054Vho1DL10HLoxsCpo79ZNMHtuAepZlLR/Mho35gK/YGTpCCgeUsuwuWq0y9aSwMP2YRuntiR/n
AXOm1TRImFIcdT/uyJofIUw7r+u49xB+mxSQXKRfKlBV/iECP79IR0n3Akj9RQ0V6td7cRqYC3Wj
VCoIZ0OI0Gs2NPj+Cm5gay6XJ5k3n1lLvbQ99sUz6kiTbH3wQANr6hn+Uzr2BtWWaSBLUo+H1g7b
W28n/3l4lqUENdMONLWRFouvKTcx9c6+85fxsdP0gKFErg1RFqLfa7oV62wHGxisaxlfdZNNaL5k
ktCbwUyAcH+ECteklTSJcJx8PiFxmzjr5r2QH/y7gjSEFoO5TUg4vj5y9cK/7hUocqRusmegEwOF
7irx5s5VKq04baPas26WMJpZpoXtR/QVVKEwTzVjdi0R+IFFAun0a3FddOO0B14HM6Ipi8QOyXXc
U775s8xqMBZVGAaEeui9NTf8Od4fgM1KcZGxwA9D2no1eWjyi3STPprzx5spwVQz7g+XcGz3fapO
VIhpDAtAwwzOBmpzJhoTGJMUHJ1D8hfd/tfTQ2WV4FPHe9C9TraJcIXkV/huKhazXx8bKqQC6xz/
z36OuIEmcer3m6po2iGO0QcNxv3tDUugZrZZa0e7l3BjKqWfrOxJE27RIhKR7zWyV/6xGTWQwDAN
F991wzwFrdpv4ceES8xlBGposm6JtmQTnO0Z77O5xFyuYzjX9VpzdAeq/udG3QWBE7kSJGuJCSRh
NFULOzHfw7j+6yd8vqV/LfzwB9UXy7nr3wGuSvtF8vcCBmurw5blTkbSTeiB2qV/ujhQwIe6HBzL
rZsqsp2QqY7LlZv8ERpKQgWFM2Ov+YEqZPfDdNwWr4wBjK+Dn8CkTSjXnwESSNN8Yb7zZuIypKtd
3akVB5QVxH6yNBozy2z7RJtHMf7PSRA7yp9oGeKmfz50uEYtUDPmjAqYUG89lW/Icggce2E2Cxy1
x6DqY7GHEhrEDeJRJriZa57eqb1whMgBCAyXvzCV/sT2nI3gqZ9CSCH2kguw86H8zuNRvdjXbIej
TG0B00h8Md6W3EwmPpWbAtBUJHEaARhKZqRgam6oZkHHKLJi/vO0ULYn+cxcOUuj5SRd7t3VYYba
pkF/erXRa1JS2q1WQNwT1WjoFhvV5JX6bi8hNL45eUAM4pZjl2J+BrTPlRc1+SG3g1MK+jHAlBMb
QtW9Jfr9YUpYhgSNdivoT8+6PNXUpeWhjrh7/hmS36XNr5TWKm4BamipfFc9vlcFhVHGNX/h+zhV
7fC+1itEch5/Zmly93unu1253wEUl9Urin9EmwWIyi9fAHTU7+FTnyu4i1qSz8KBwFlyaSgBUlZN
pjjZejBCQXlHtaLfM3/sAWM6L6PGW85S5bsE2U1jcDv4RDzwyLX2a50BVjgArMYqJ7PwxiBowEcG
Za7LrKdlQ95rE12d4JjCC+MV4qpAJ/ag1fsfaa+aNJAOPjBtBW1Txv1RgzraiQIAlYYNWjJ/hdxD
bJ/1aGzBbsEx+OT9LQTePAkcjImX0KjZvY4GspA9JQ/M4IAjGwmhO1I9IJJ0s4g7ZBHAU1u/bOnn
zU+L0lajk1xsRQkTnolkM1BRDMkefCtpdzuq3AWfc0CoXWyKZ/waqn7zmDmqvmFc5w+lIARlijKe
ivOupLKwTzjQAVQlppk+XCAcLL+MEjSJhr4pdtO/KHoBEc/B9n7AzgThQx6qI36Up1qK1BAM2kC8
AeXeGhA267dzWO1F9gZ3R8mbJm0Uy0ORRb4hKFxzaq7qFXjPtBj3/KNhnANpAoYKZ2yi9UlBAhHM
OcsSik1MEjnjSUi/qmdi/O4fG/iXfRVTKNweqsNBX4P7O3+ZeFNHzlFj64yaDwHo5fpV9+quSaVz
HErMZCYd/DD69sEx7f+hUWPiQp1Siru6TlXm5rEWk31pl142aPnQ7Bt3UFlHEivCjDckD7Zfkv1X
+hmBUCZrBURl+Rs2M8zpiqrZemrBkp6mTl9QxLjQRbcU8OjNUwUW42w6qfhVYVtCDMu4RpTrLeyq
jGlowO+VWN7nzueTDNMtZMTZpBWBD1OYHrOXMZrlgQ7gYyBnQPDDFeDwprvBJf18k0/b9H6bZLOT
OxV7Vqt+n4PyTgxFRUiRdS9VemV/Jy+peIXL19Ij7N7V7InOK20QNO8YpjU2WIyJLDSMxVEE5uhB
64Dy5TrXWHNwbQ7gyjS0hrahCW6K7O/pTwe7/Kf8AVCZNxPBYZxyzahvGv8G8ULkh29tfNl4EuoV
lT7yvWnylZ3I8fncsCtEe33jVMSmmwX9T0ODzcyZKalKcR36qwTcQn8yTtnI3L2oTfO7i838nwoD
coDxYOwp/b4tDKtqfAVNi6v0BBRt5gYuM1VaKU87WyJ3CHal9ZaWjHCxuvpNobZQVWVxmtu3YCN0
0YNZIUB1Y0jw7puW7CdipGTkiWjEBhLh0VniD7OnJHMI78SkgBTYtoU1BIN6JO+2iVi9P/7uF+5d
dIF4M0JW39VY/42iq4JjESkbBSjI3YIk8e3DU6IhW3LrEZ/QwNf/biOOlYa4BCsw8Eoe5FdInoPp
vcwmsVdVxllXPE3ul5Npr7XCimrf/P+DfimNKyCzDI/blq+A9otMJl7hcFM5hz15/e6StQdLuL2K
WltGhKzaYEwMMVpZWeJFa1hgflrAzuK7AABjEP4U12NGfeXfqVTOX4SexRrkppjnA2TpU8f6GxVE
mU6VJNzczEF/SxeEOsAy4t6MvTXfMn553f4ok/GhW37AWrwcRB134ZMant5u+Yy2qQe7K9ianN06
Kznec/Uxk6yIhYy1GoAvc6KtyE7Sx/ct44Qt45D1yEgY4IzkkLIybXd5XVDunAWG6JiGUU2TcMAv
w4K9bjzuCNJjOTJApnvBavlhoQ2sATWsrn1FBtPChnBYDAyb+LrT60ZHOSxHzokm+kuzX7npH0J9
pYKXRR1/8+AC8VZNwQOUcbDv598T6HbsG/L37Vne2pf0Z4hdPJ8D+ofPTiGrBuC3C6tpAY3scqLS
AsNJ7UuL90CMHYGj5sDI6wWnViHtUDNiELf9YW+5dfizaRDTnvv8lMnmaR3MPgqJqrYBint+TLS/
q/Ux4K263p8TntbWB0fQcWFvPjW0BhS2Mvnva7UIUG9H6Ttnqu8mfmDnMOY9OROnyeG+acC5GFRy
fKNWX5XFykU+h1ZwPO7lDMUi0yNddsiMwLPGHSOW5OVM0DNO0sLnvBjk8kSP2kiKMW++PbeaI/G0
81eWUtX2ucfO3jWZVQ+5LBIGk60iSz9Jf2Hstr4f3Z3m7ui2J6/31mAXvENdU5lIcj0eN6CBg+cN
aErCLIBZ6RLu1jiOGdh8cM+ICWTZhP2DhIyneYKX6vICsZOk9lul4yTi0w8K0CgDAfEKA4FQkkgK
MyFSMphVvolo3L0hcgbbVX+ZxBHviEo9wPcbuKwl6JTaEeoRr+dBJfldejQ/ia0EEq8K+Hb71Ud3
LdiNPPKKmKB4gNu9h2iZgT9xn8EZEyOVMYUSRDJMtXS71emiJLNV1EdgTy9T02nQPVMDYPJEF1XT
JJT3+veBzvMD0lY3wM09AKJe4sKw6yMKYXx7+9oT/cz5QqGaRt0/FzQLtgd0DGyckyUu7P6CHXTc
/h9SGORaMaYcQhu1cNBUgKVXF4aQpmTkWItUKXsnOT0j/WC0LfbJ3mCgzA0bTk/sNUmvC2tHMHTB
5eSmSl6CNyead6D8FbhcdJ4zYL6bBWxb+t8VqyrZA4nYrVEa09bP0PYpqHOlWPtZzjp6OVdK4R5W
9Vf81y+jhVe1teA3fg4zW/2LkezoN016nuyLNPKQN8f+79+PdPMm4YjabsbOavnkPUJbthmUjmpX
96eAkDvMp21mBfZ3z7k/E8PToVSCht8aPb5QErLiai37WpRNMUxhsFhlI34ei+/azaqWHFniusy8
MRnzG1taIwN52dpGx24kphUO3AjR38h+1ilAjM6z36CGwam3Ms7d0oMEtzmDByWC5dZQR/sHRgl/
V9r3mJswLVV1Z/MKWUupzhX1BFjmFv8xdAgSXKgpI5mC9E0Saz31UlSbZwNwNM2ldxUQhCIq9uxB
QSL0ZmAuwWhwtf8o4135UeK0rHcCze1CO1fNbBKcbFOJDJRahtslc6sthH2Fb3cmI8QDcLXpcXWe
nwM8sfGwfPlpN4Owcnatn73H3f1dLTiqTX2sd0meOb795uOsHoA37E8A95gKqQz9TOvo7fTnRz+g
Hl4Syu/x13UloVA0sTdpOBScnEp1/HOjZnSsaAtp1PPrmriy2q9drhICq4J9TvrbvtX+loFme/WR
7NW7JvkWTdfw+C4csAAryw2pI+h779hPwh0k26McDGGGeda+QeNe5gMrcEZT05PTN8vbAJ0KCrI2
msqbNxyncDYNg3soodKy3tCsKf88DB17T14I6DXY1LWVefatbgq8WgFBtlM9SBrVvO6INSx9k3JP
Ndsgkqpt/Y2r1bdqT0ro9m4cEnTcm647yRXibZRB+BpTRTfIk9BglvWToHJ4/5SyZTPM4CtDowTT
afIPiAGB9pGgrXZVf4IBffW8VH2ipr3QUoJN7uMIUJRbx6/F71XEflGtdgdkZ87PNdpsqLC3XZVC
CTzFnXG/mhYgi/1elL0MP3WvxYkyvB9TNR6dAVLrmCd1pmFCO1PRfNgV8Kw2/uDMK8CbEE3KhIfh
lNmkTME1X0FBZ+183AmmwIQT22QoUFjBY3aUse+JnQMmE9ptWyNQnnSrYy8M917tYK3uYZigUzi1
u4zcY3A92Cebqd+8khaShtzHGNpPrZNN8avTwBMlHqbY4KpOx1OqX+mMg7mhBksiBrEZnvmbHPYX
QlDFbWiuP9ldB2YZ1D8QM2ffYkMOS3OO1qZBRrwpcu8e1wjmB6SA50Q+Jr8Kz65+C+zOV29au8Ly
j8Nd8WjpWgzP0sUWvvej+eS/yRX/X1IOdHhL8FPcEjO7E+z1JSHe2cQsB5RnS//+TrbPxDYNzeSG
RH3WkLc1OqOg2Aw0JOuNfzi8f9PznOiEvzXY3sgA1glR5GTAleY1NrNcI6XJo3hp7hkc3zS12FCq
yKNZEOdKyoYmcuGPaxM/Rh+8GMzr79Hp9uMtL8l55MsIVWL4xdBvhECwBlZcvbiSUokK2WTqdb0v
dgdcTzCdlcIRuFQZIywL/UQsT8hUqihyuA5fQEhu/wNMbJW8UTt5LgmC4wOsQkd7RjUxllfn+qwr
nhdW6OZESTfnbEC6o7MV3VI8bqEI3ZcyiC+VKwZ5TuDi4gTqu4XuvY8w19T+EYqQZN8pgz1YuQKL
vBsG9D8db1UwJH7830W0KCGGSboSyOxPR0yH4SXGqRdT5mL1+4Pe6YsQbgWPd3DdIh4lw389XPsa
GZpn4us2cSi+I68QOTTEahN7IkOPlyru+E3gFhqN06f0AK+NJZGHfaICgl9zOOKmgpVoS/7Eyo9u
c3v3EznKHTX2fInpguaQfAFtytpSCX9xY9nfZpiyDwTTL+i09r50ZTDmFpyDTzy4Tko8+78a+5V0
LDIIkq7WhnkvdPCQiutuUPuDykCu6jEUrCdtCozuVSslIxDs1JeKh3JC9RUqTIZ8ZmxL/1nDv4Xw
vpXTSR1qufIyY5y7zKzj9kuH0dEogTqoRnZwmgSzhwVu+E7t50pdYIeLHZnfwnyRPdD8ZPrEitEU
DmpSRtjq17LSMfbwVLroPXUs5XU3uutkeLqytnMNBq5Vk/7bxiFxgaAlFhVAh+uRxDhdJClD/rc2
FD1VPUS6Wc5mHL1lswKIVsPDnQ0l3V+2GzZWdIkJhRlzoXhKdoW//cEVSwBWyt9p9m05Dvm524Rj
148sJ+3Xr9QawlXzQShACtDVGEwN9INaYBuqlMg+J3HhykVHfXNDsyhLG9YFwdYua6+gHv4r0b9e
6g23gBaWl5/gCrPdF2urBE1ihKCI4hhaNX14SmDai2ixxqGRYHtXuDJSVsPgEptBAPqokaXQxHq4
tD5R7P8JyR2w3bLUA5C7W/199xY5xXatZ5VYNnTCvacGTsYoxPgbGXZN5rR0VgAFcfqVutcBqfs5
z8qnm8RzoNzIwZ5KxIslaiEiKmslu6DXT6shvyPc1aw3Dnd9+gLByBIaJfXc6y2FAinvjGcvH02b
ZLxr/GK/uwTwIxIASZ8Ncnlfgv7V69bod3PExyHXNjO/k0c51A93Obb8cjLCX6DaXEhl/aflUKgd
hDsm3cpBYby4a7Bk5NH2FCf5vGY6HE6CtblqAiZbvVTqYVTO7WviA/n9+eD7n0enwS1uGoFC9rPu
rI/1C58vhC0IDu/22iDO7fUCaRdLyrKb5Zw3rVS+9BAcLg9PkoWzoRSjnrTD64MfhBROALbOku4q
s6OeRfnyVrUm7ssz5EG/RorODzC8FNfUr/0npjwUUan7QPdJjzkIMJLag4TaKsJCu97SHNa5cIq6
th+0xcxOETBfcxaMDlGqgONFOQ2kx4/ZNjZdpxGPvdkgJ4mvtKkCpkRZ9fY7+YKZvzkAErL/zYUJ
88iGxWtn7MtTh/k/N5FZHHd6/k5gVGSIGgSX6wu5qyOadgWsCrQ1X/08SY9yR1UZY8q3u3zcVsEQ
VxtuN6H1cwoQVxHp6KwcC77xGq0wVPLthUxgIyS+3yJrM7RTXzco1NOsjKlpTYQt4AZOvGfhDGW9
VAsO0Ve6D4Hsc7H9jefT6ZZVOuOZssjs9gEmfXpzGNVOb3iHB1efUZUHobnYd9TKj2026SZT4DEL
lvOxvXoY9wJY0qkaGUM8N8qTBicioSRVluyVqBTxxMYUyma5y03y21J+GL3bqtdX2RdrOd+dTTBU
17hnbPavssPX8q7yrYAkyvOWEkSHEAZVTEspOdCI1wiJXzS1StgtZ3aZWbQ53tm/V1Vg4FMciQ0i
R6x6JArCtTLPI2/bgMO+HATLX6ttI5ICk2JlI8aY7vABl+VnkBL8PLR7z6/NdeC4zCu9eZV9qc4V
YiGKj/dQWM017ZaTL0lbLl1hlWYBBlOUM2VCD8Kmz4EdnDMbI9a8o54y4NMeNCUv2JYAL/EA9NpU
akxF1lEcaZSqh0xqGZ8OlBLA7b43pdnHjxd3fWr9uOjXfBpKNEbZLazju27UBOVosCqz/6NFRvkk
Zb3YwkfTWQXGSmLQ2MJRbNPmHo8KspmCCZfOf3UVwOrzrZ/YmoGPTOhsq/S1qmekvSAlqwnCv3hS
L6dcyM9OdgWZRxk0iVRJobhxGzsEdRAIgmEY0ZvNN24fH6IjOqNKumA+hQ2EJ2tSno2V9MO/kPji
wMZN+hE2G5pK18tYIbJYgTH5UAZQYsYbg/cyIydJky19WIlrUBwmXUSRZQX0u1ATXeszB30MMPwk
4wNxQnQH/V7XMLgyalYQ1VQwYxwDJVCN7LO5ypnU9xPLppdlgnxl/5d/gm+OtnkZPSf497OCbsaG
JXaDa4q87uvBS/6XYvDDJJgGRBncoluxVu2vqD0b5hilj0ScYG0AtNObDsbgAd9Zl2eR7euFYKJy
KlWyEkaoi2Rc70ByFZPxGWmA3f0YHQhcsS7vBDKaihLdTYvgrjn81pL4OQHaQEAsgZNb68rB0NFX
+7hQl4DcJLo53mB+Htl7dB50iqPu7dgwZaa+vJjnW71kxb0lXgrwFstclApGiQfN4AM0CCJweDr5
BNG8abKoK2l5h8el295zNFPFhXWVQmb9YLhooZRXWW7J7YRo0X+raUBlxbA9S+cpSY3lG+gbRZ7R
mz65o9YM4UgNY5/QGjAogd0vKSF09G1pWcjzKUFQLnCiiGzRLXk3WBQ+8VBp2ptBgq6XSAItB+9D
hpUNHrF7GNMFC9pdiE3lRu6hk9Lc+COdNgLu65ufnvzZM9vvBWFp/FfXrdXKXEA5z1q/qIGf33r7
l50o7QAVM5HJGhAX52kEzH9McnrpsrrTDgwIxtvUqSyrGaW7/TYdifuIdTAV2/LkUT6gKOuv6Yjs
XzAImQBROYLoWog57TRTkcv/tzfJiG82hD6ve8/ywLabqi2S7dCK1ujYRaaZSE3A9c9ge6fA/C60
LY9s3E6ki/QLCcLISuboP871sOc6UlrqMcS1WSHzq8SPRmZYkAlhOF1eFXhNd+li6eYvlN+FVREL
/owtg1l0hN7S1hxUcc/bwqZHqsxU8XnA8S7vR7PgicKkCG0UAMfN3emNzvyu6IUbQVSVnANTvHgO
2ugGABag1uS6W7cYtKdHcIyCVmSMD8dBVjGNOStM7zUd6FT59MqfPMGmI6xNSGJ3doIpNEjGfK8F
crh3UdDaNOw8wp6f3lA5WD2Qq0dx3ejkVtlHgyvaf+O+9YWH3vUsLLfcNavUOb0weTA7Fw831xbX
4bRPDK6+cRQQBgsOs/WqzvQCN+/d6/MT9RoX33nOJaJ4M44bUvZc1232jUG+cz2w136giFzoFAnW
suGeb9oEHsLIjDivDbryJKvgoF5Jy6RzY1O0NKh7WYCc+huAGG1OWFq+hvBGRxurkTfo1b4ObEWW
FKEQS9kyPWgrQQukUJTyodlOpDYT1TrAP+5bBc6JFBrwbNolX/d8+Y5K0RyonW2FH5fM0UrEb76W
968ooHXiOGRndD5rmO61GAkMG0cEaQ4XDU7jtfigguTaQ/C1lpyKF0EIp1tU08f1V+6wvEf5z1wQ
oYQMQ8PkARp1RFXJO1jkluAQ0o1cUhdeB8gqy1XK9QPTHFVYC71DcdD1clF4uf0++ILjkL494zJa
/rpytxZYSdXPaGPfuMXihsiso4WvC/zGxflJ7eYbHKeuv9ksqz6SdLAOzO3sRM8WDYm/6q0aAHKB
3T0lPvfbrwijWBBLRY8iDn2tu2OgDceUCL091AdkBpNL4lDvu0TaN3T+Ps/b1nLqC/q/EQueMfV6
atiC7/SyTgBQIl2W1pKXn+OnnjJXQSC2wi63i+XpkToxiAhAKbm/e+Kj07//X02bSJd7I6iT3wVr
OWKAYwqgAH0f9rMqzZukluchgvUwepTz4fjxekoiALTbzNdtAZiq9G55wawthD4XBA12zSyQBltw
ROj9nOlCNLLnw9VRzjJ8t+IYzACy4TpnDkSwXw67ztE1HcZW/pLc7PY0d2Sc23JjR3fucuTlxoCO
wTtmqAFuW+YQBcoRkxmBUBPUlCBuw8Wgt+sfbmGOvVsmcXke+cpctpSPWxQ+ZGaVIfprwHnRWpDs
airfBEK+ft3+I6bME0jqGkHd7SaFkNO8CKLSDB6I8Q6NIt59pfYaQweIt2Sm022RVz+vuxNiIHjV
PGU02a2PIeqBTZTqnBRqi5SgoBS8C+9qWwLuXWjRTWrmrGgF4JYCN0c88kU/zOscBlgv1SEwH9g6
d3E63TuGBqFs8mzuKTVAfnoiV6SAVPk6tkKKy58V3fRQ3nGPwzdj63vmijM6QwLMVjvw9QTZar12
RV0HzhrjzwJsOAube+Ot3yBs5kTQeKguz3Xl4ZX2FJk/H0y96k33rfOe1gpVRFy+KNqhxqEVkrdc
uNMjidB28sS3kTePVIgirKfDN3nWoGeu35WZyJsGfSAfZl5RYC4zKb3nFrTRiglO7swcCt4tzi3w
w/ma8nuBkD5GXJrD8RxPp6v0YGxIhwhLuWqlCE7Nr2rbP7ne9A5igklHZz2NkS3YN5NSpZVSepdP
EvcYYCTrwMHaXj3IW+KJOmbXcELXc7FNM5Gt+Yjtk79Q+pwGxB63105igAmh6aXwLFTHZKtIc23J
9i6brsDS1CU/dXhmDnIQ9AishtSb6IuSwXkzPWQWoX7j5KNtOMQXKZABImlBrJaRWUDvihaaxJJb
18953LjKxFm68WwSfR+CDsN4Eeq8V894GSr5sPaei0WG7mZL66zvXJtq4vWCuEOOPF64rJbPagIh
VQ8j5ddyldoYcNIukQ2ALsx5+gTe2tTkiVLebiL9nF4dAYuUNmHlau1LuAaouEhWCUlWQ04CdztD
5hM8/RBZA7d0+s6RWe6rXGt30iiAtsvfIjl2ltZi3Pt1a9tG5PxQIHt5xywnwEiPdvm4nCcnS1SW
66c8G1F/O+dGQP6Vo/vlfruni69rgI3qN0+7xtNRebBVRF+Dzx9Sh/x7d+/4A4hIQPt+w0Ftgle+
vWjvZLZCNil0gPVw8LmK2Rm7yHREG7ExGrIRwumBSSYAo/Z5r5VzDFStM4bke3KXdxKVqLM4Hznr
zj4NqlXl3WP129zUwiZ95VQ7ge1vavmjyZ5Qj/toU0S3FFkSjlmEBoEBbCnTbe2tO7O4aV2//LqQ
pTpBeoPapcVBvqsdJdcAIrZQwjBepMvPNOqtnsRzsB2rsNEdgqv3VZeH4GglOtUFfbl4n5uyT7YF
7BjOzH8hG7D+dH78ddMrvcyVF0U+HJalEvksNg5/RtzTMRAESnuj+BsEVpzxBVop2t/xvTj0IOFk
JCaq2y4uE5w39vJnaYOMjKk4BUTxJRkEvc6dFOCYexD2pbzIEcWsKBaki5jx1r1Y1tTgNL1Crfc9
L79XysTblMToGDMtHLX7z+M+ffkP6dsBfbu8GBA+gnmJ05EMiUlf5CRW+PrSIHekAr0RbE+IgsXc
A+kuJV0L274JSoW5NM9sxsC+tqOJww4UkOYje+1ZadJkLVGLx1I4Lfzx8zcYjjufMlONBjSIYY2B
ICHKNeS28s/hFCph4m2Eb+svwSQq5yGkM1LIhxhmpLscLJToUIL0PWmVPLSjWe8I7xv0s612TlDi
3KeHFFiqHpdzRGwoP6ZCN6DOBP3tA4HO9Lhnr6lXr88lRBpeaiwrUx09UFynocsVqvXhMZywtheI
vcYpYyTgfuSdPBtOJVl5mw/WF6UVxyyl8/Q54ZlWq6Ctwvfst8Wuq6QuSRcPz6TCSZYqzPtKulMb
N7Su77H9gPAzhU+pbnsglEnBwhRRHB9ddRj1Y74Jagz+3mF7RdK90MYuEeO1WjYlEHx4F+ms741d
HR2Co1XAoB6NhXLdSZEXg/s6C0H03BSje+0BOxONhamFY14mn8yIFU98JDuoCZ0BN+9NAze0xIbn
SYfW5kcTAQ6ceYzGueKSiJym0zmKiMZZ4+zYe8GRcgok3g9DI0DIh0G+ufZ6gnzLHH2/tjpwVrep
3IJTjj/cLj9HU/6mGY1t935b5+OM9PYUPHIJ2gpmLtaw5roW3Lq7JrqUXsqzR/2zjU96QyYiGFXf
S2scx/mlPU8slYrVz5EvdSpYgIPSRjagZWif7M4oR7L3m3JLOY8RofNrmFkBCKr97z2wLJ3pRehd
dVDcQTXUEefOYSm6nnI9eyZjSGNuXofUfknpl2ozGugIoO4GRdMuBn4gvxwOizjkbat5lU5PQ7IC
gf2p3FzBUQlxV46uaxnWhOZ4QnyhlcC3k8CV0XcxURY8OH6WxkJXrbRyq9CaxrLdRW0/4aKag5oY
JL+WXgOnUEXoEpGRHAw5hSQuLhFY00Dica5o5dbQj3rvP5aI1BLADTbWFwTumDFLcGR6c+eBZM6e
2qi1AlQD73/b7DefPg68f99qYuKBvlPimUcOPG00GShT58ZD701IBdi+o3oAIj9Xu1YQcJW0aPG+
MHKcG+KSBDVlN+qLtkpLK+tXG5TEldlXrhlIhG7cCdBMcETjSeWHiyUIw+064m0d13rVI809xQKw
AkQE2cY3U2V28WODhXKqZUCkzMMVDquOpixHlp8ui704GycnNRE/U5LxyZeBWCK9hGPEqUwzNHyS
0vqkr1FmRn0FTnba69kt6vd2El+sRvzZAuOb0czzm+Vkz5r3Ka6yFunrRXoDXf8yporLfU3VkmxX
rlPBHA6Ejp+jjMWHPMZnicmXUQZFp8Sf5FLWvRh4DMd+2ogEIhpkf9gHPecG4r479U/iZ3YLsdAS
QExk6JzJOMnzIzrJAZHSz9a2r0sq8hs63mdUgOQ73wIocYHUblwJf0OroxWJYI9aTOPp9OjEbaCA
2T0d1E/51ILXs8s7i1Jj/otfN4hszOJCoRhkB3tazJH4P9NH3Bws9jxQd5M4NE1yV1ffzjbmZtXp
YjH5TO/+wgbzU5OB2EkzGHvvP0xYasMS41P1ow6fAVlpvLTbjhoPDO5dBSgwcsibT/rBYbwHhcqO
3e9KEOkMFBFO2dJDAy3kahNM3g1CKuK+QY/edsc/TPZyE0NpTbWPuBQy39ceu93HJjR7aXrTlPQ4
DW1t0ZWHWPKrnAclLyWirPT+Syl5GjgNOAGaqLve8AK5351S5vADScE+A0CYyPwhPcD5LZI9v3Sm
OP/cWQMt5/wxiqQfHJS2qIcSzNMStyCCy9n5VnI0IRfhq/mi5jaljNdMZx3Qjix6w1S8CPKUBdMF
4AmhwzPSjhA1SbZvcU0wyF8n1PTfCBx9KfxJJceTCbuwGui9DXLNFgAE8G/W1T+8UEuvB9w8rzFb
uHL5HRHXtFuSUaDypMiQ/Y/noVSZQ0uJuWLXsrXXipps+tz3GQ76q6tO8CJ9zh+aaHT46wsP2Q3K
vg3bjSwTdMKxL4fN5eiwdTBb2V2F9hnWQaAWglckrM8Tq9gylJWE3uy3jtJ08RbB+Gk+MSOPjjqK
yxDDW0FL3xgps4pyrChIGuH6CyGg0wjUGKt6/KJtAjeUJwix1ljMIj2d/3yf04+jVagGr4vhehgc
mZ3jAe3TQsq/TmRmJFyN3LFzo1ytdsI8hxx2nRyQZV/tQrXLM6SKbuui9z+aln/pdUFJWqNv1OTj
VWbhP+pDgxcGDvOu1TdBtZscpFQ0udee2aRIe6U/6V30GOMpPn8Z4tiFWCE8US/oMeRlfkPoAb09
YuP2FXk4eCEVars4b9zkrdRnM1oRKwX0NtayuCfvnV3/ukKqeVdPyKEc7609tirXK6zageqiHyX/
iT25yP75sfTWveqoVMlNm59OGBcInoZ12wPkV5ovyXwQgJ5CSh523YzsSWOE739qWaWkcyqYKwtZ
VA6SyI3Omh1vlsogDntEl6p97KjeVdEFjhVilCA92Kf4KxBxOYgBQDy1+7VAyXhgV7AOLu49tFWl
lDdDzs8ImQx3PTXDNeYzGVSz4a6fafS0uRjzLOB0nkC/pLy6Whh+exjNfbhsJZQoLm+IC0lRctb4
Txc9bZjDQbcl29beiVfsUBWXtJJHIx8Nk0GEpRmjqTglmIBey8m2oZIFimSeLKAGFnPD8I7g/ex+
GttOAPdYbAO1UPeKvfskWhoY9ijWjxC5av17caoA0GnhzrId6lADPlJpSpnjuT+wDv8PcbZ8Td/+
w0iG69mtcxu+US3I4ZcjXGZLc0kA8Pm0Cvh74XhdwzcFsgGwz+FqJSSzDiHwbyZcM5KAWiKMCdkV
MYaOxAIL92CiVjxvdjQunDe358AE9kOVw4mJISoqW7GjJ0BlqpQ3lB4ew8BhtsObXUrqGUlvbPbk
EG/FPaLJhkBXfiGED2H8df+kiJfm8Wsk4faRAD92rAEHasIxk/LSrwybid9adEhowI0XA2A1csqG
jM87kIWQFzgEB8OgjKddZUCkI3QpXQLIx3TGk6LCkkNcFoXTzBoo/Tw5tnHNkDCoRjhN8wEsqcTZ
LcjHQ5vTZySkTGFJtlJL/hogQMOGOfp9Rb6nFyQWbQnRlvYezolPYAxOS8UFuhWpE1AYxeoXpBjc
NqYVy0aZB1UTLy5i5dqc6Qie9j67pOYeuoWpgnAQpp4GMvxWipKRXcS08+ejhlDLrIag3ag+Rk6m
7QvS2GsPAEoDPVc9iLtoyhAZsEoLf+J6cXeW1txNd5ESEPOebVJkNlwpeCI45nkHaNkpJAo8rLn/
Pe1Vw9kORHcxeTZ+9qedhVhra4sqy+mA+9tFY1b5RY4YONMTXae2XxiCfGbyQHWnPHcLDojFwGum
UNr7DPNf9yts3BIq4KQl/CJ1aT/f99bqVwYkWQqelbdpc+SPbMX2fCHEHaRjw6QUPqIhRPl/Jxju
VBqUtsyubEvPTp4+ZoM9UW9FYTRKG8mnGWSqcPFAKZYLh47iq+8GYbB8taQDqDqdzmM8HawpS5x5
8Vs4N+tdvcufla54DDGKzFgpFvUOtF5tsy5/HfaaI4PCP3kJ8DpTsRuvxQkTbZYRBkypdogN3U+K
/HR8qnjcnXXWf5rLVJtCyeKgKSbdf2SHCLIDfBTLR6JDwOKNTZ3DANd5VLmqmrDGaGICn3n/JoAA
SEhAn1gJxlQVLQ75KUKzJBxlcvJdk52BApo3/AdSY35OvOnkY+7kuQsYjsFjTXTm5x2K/nIKEomM
5dZxLIPnG7xbaR/CuL7egd42HlC3vOtDY3gsfooXo3PbJIW2MsL062eX6faKaKWWznmM092Uhck2
LrntPMdY2emxKTZMu56ZArFYWBf0bRkDKR9f9e7G6fkv5DQII22FdvRgUNqfwIEV/wbf6OS1y903
lPN1/DQ1XvfYbdrjtKHt0XF4ZYZZPb++9q/6crAuuUgEykLul6fQV/bkOH+MuRSwEKyjsbz4mk8a
qHOaKtNaPOVTU4u1DeaBlBTByhea+juEa3wELh/neeZxEU+gTyRnUHpR+BYspASms4DJDwULCc6U
0OHSg/dPaw0UQowPq6WBPz3T+YdBnd4a9zzY4/XMK6cUNLKHb5LjYp8l7f7VVmgnbigddjJioVGU
Ykov+otjJjMNb8OL/DLLc5MfnyxHTaJ3lH8Nf2BYOWYYzM6MEnf/A3s6dUYwZoWaZw8ywaFzAGLB
cKGR5EyETnxvSg2c1R/QxFYNGUSUoldRHYoJLPRKJWMtQGc84ucIaOFvTxvTkQISQqbZyx9c653F
e2CD/F7/6oLhkP5NjcjuMXgG6CcdO6DsA94vv0JmBpxG88w1GamGP1wWU38LzD6ATKXqVQLRZhnr
cP5DppkuPVTIgcq81Bq+5FbmyVfzX0aMGlH5QRjNdd7UvGHAmfcjlCxF3euwDwNez3pFO2Np7R58
DpclewjAdaCOm1n/FojrEua5p8eN3zP3TX/vE2GN1/UYKWILccUqn5HEGWtuhnl96/EfzPEsp55M
Ki9XVUrDUEuE3wHfHt9kR5dm80416qR22Y1U2JZkquh7l+PgY72m/Z8tqK9tFzxBsKTxnKDiyWNL
/dXZleToMDKUe0QMMs8LzocA9+JI5wim2+V+xSB5NUgZ2M6EbJdkvpSNG6INaOmBqmR8rDuUMzTM
q9oibMRiT7qNfZBSr8d741dKYFHcg3TrjoMRrETfeKkD0kjxRWQfBUYK2pqum2tIxRi5e7JquVjU
fBcuKgrtbeCFHLoSQqRdTxuIonojDQu499YnT+qNTflERtIl4f+g7Upcd83LfpQ/+hs070cXuh1q
Prn/qk9GW//fl20SA6p9YHTxcL7YL0kbQhqP85+bmzYtB1H5Num/d/vTSUwM5eifZjXBXrYb+tuL
AJ8A5/YsseZ3i+LyNSOJROmwy6F71IznbwzUjzuzP00KWSjwdj9JCtaeF99Xomy2LGqn1BrZFNfZ
kep24HlAxKkJFtUZDG9lJEqVjlLp3417O+o3ScW39zCg5iFPtPMnCFoqsbg8cdYd4xvSZDqmbQJ2
FsGFb1nh+Jfp/i/5vFGi6mrADosQeM1ZSpD5AwDe4E9Tm0WRgOVNetYo0vLb/uP4kcWyH46j47M3
s0e9xoTbmwVXXskxFf340EmK+Nd+8fnxR5znlF/H+PVY5d3Pqb1hDlf9ZNhpVKiWM8KxNWmHBRVA
R7q6Sci6tLw2U53QHHNHcvd5pBJuAxqekZK4461XiR2y3L2GKLudUZwe70fIDHMNgBe7Gi/V57HQ
GCzSwEieiZ6ljk2XUzsxffQwX/0GPVzITtAWBSsFnY3w6sXKNulanzggiO53937GUMNWQwNGHeTH
L1QW6JA8GIhKVpLKoAhQ8AF5kvZ0EK+kuXDrEB8zeIkdnlqz6ZiphPnfJce9oM/baKj6fOBsyHCv
wxSL83DcIDbm2F2EAv5+0ZlCtJTM+Jvk4mojCufnehm2jmg9TS6+5W1veUDf0eFaWl+ULn6nRU0B
e+yFw5wxR13v4BgV2lWJIFRGDDGyQzWg4oJy5s3cpxtLdDn1UAgSJcLlIq2QCwZxmiHAtm8SQyHj
K+E4ONrYlu5OjRsoFOAaWgSOt+UiycdofhIDW5M+xgJkGypE5JDWfUIzYwy/H0ENi+X804eSUWCI
wRpBl815YKSzwCHf4abxuJNkYi22qRJBh/7+Wv3EYQqQ59yNzAbJ4KHJh552TET5+2jyLm/snOsD
KB4/8JX4Q40Ayb/qckXmt8AZDAFOWgwAZEkBR60W0oYlgA2zRPotdRf4lHShCYuTMMlaHPKEaYHU
kCN+SPVTkKQ8fknKuc2Y86FjiuMIgZXSzcuDdwI6b3DEAJDQmnC+eC2cd2/YUWUwcPZuD2Sgn/GQ
UIhzqk6yqzFTDrL6P0wV5T+KJRsLNZXP2D9iCACXnb1x8SmB0KDN9URo8lREfzuh57QNm4GeFGpN
jNX0yFlzI7XEWDJW/NlQgShrFwfb95Z2FVwdnHdCbDZ0PEui8jLD7L6Tz1XYTUyvUbH251KhdVcn
4FtqyoWB0l2DlHpiBHJj2DoczCFVHmZhgANmQJ0y3VmA2SyM9qRQz6IjC0PIPZAU7MysOd5eMrKy
/hIbL/G71FTuMuhJyNsESrVtx4Jc/TUfj6pTVvReG/BDmvM8JsBCRjE+I5sFTQQyKLGMDwd43ZeC
5raR6nvu/t3iZXgAZaRzluE9rEMZu/PyoTr2tlGDc9qKkIKFQfemgFl25HArfpKbV8Y6qsFWl3QE
PQqHzsM01IbOc6XJBD1xVDxlYpi3exrMia8ZxHoZTKWAxKB5vjyRQBGkb+vUluVhOHPZ6DrY1Dtw
/9fmUQx2WQY8E9kBARzyI+rhP6O8/1+ckTSEv0BrT80GLz68VoT/KhqTz6nKc1a0V6y2p/JIcxEC
gm6ngVz3DNDI61LU5mDiLUS1Olx/sfd7tuEHrF389iKesggkYcZDPA3ry291hE2v09zYIzUlL6xA
C9T+nsv6Ja0MXO7sMzKBsUuC9wrkp/CMDyBa32OWc/QBvNGm4TEs+AD5T3uUwRHkRzW39+m+uIj0
D4bwKtg26CwP8nAl7FtqlA0ftzU5ncqznZCFS5bHqyy+zB/fdyFp72ypqv299gpPE9a9mX92IOxB
pK3uYzgPYrI+Jv9lr7hU0GpuKHsF1F0orOKngOAasBDaY+nPzoegZVWO/dhI1XlrKbAjosqTa9+n
Fdc8fQ/QiDerYQWzocxUZjYuMAlFwXQBVIJ22MOFa+iyBPwfxWjTVAnp1VcbzTWR/P3JsnsqrBVR
vu0+stjgK0/P6acKC32hzUUFUw/OgSkpvO1OL4WtKf7TPY9FVa3kLGKLWVlYhU1tv/2X8yYLsy5k
aP4UhK5GAAIGTam315SSYpw7ioHIyVFZddju3mJcZ8FS+ztlWRIClv6qUHJROla/TWFv/Nj+RppY
K9wKn/Y6GO8m/xefjZcVt4aAFKT8vQjYy4jkf4C+078eMwUeQhv+dQG8Uum5kdUey5EYZi/s09Mc
b/PUEU1ZnLSXSd+bKZc1ffOkDeEcJL9YWw9pEt/9A0a3xFTKXv5eU3eAf3P8p6uGsP9YyRDgWFQ3
Jgv1OtHLxic0ZybZGGRl6QZ7qwdBB3aAF1XX4BACwiZhXeqYE58HVHkVyg8p18VpXnZpPVsiBsiQ
zYmtCcCwAb87G7M5sSLlQQMxjS3rOIrynhV6cNilcAdTrOo3JiqOS/LxbnfYxt3+9co3fQ6CHU0J
YFmtBjx+pkm8fWs/i3DDC0OoGNQ/VbgPu8HysEFQj6mv+FFCmPm5qvCiv9I1VKrFiV0viw3AURgz
i9hsbtY40gu2xOdf7o3x96zHn/0RTz1WnJ2jaXqDVWXceamy+w5xUtwsWcvnvcZW79vTgea9CD/u
IYPhV4QCjDp4AURE7Kpm1bmhrJ4OnGdAnuBuXvKQHpjXUcsFci3WV2PSO+GGOy0ruy8zvo7Y07F4
uBf8g8D8M7wOz2MOt/jWfAPgkqLe/Mke+c4mDUKtLARfeHOuiVWlidQ460XGk1UwVvaxHuSD1ihq
F+eLnVncIdYjaMEQWDZPSikitgJ6ESzyIK5ZkemRbnG4WpfMDXkKdTo0pnKOwLPklZZDa1B/E5Ak
0akWp5ijgU9VR35EB3Z0rA0Uwgw3YNIAYucGKICOXncXq96f0MihqLnuIKtFvHDqkQRjQzJlryYQ
fIyFZdY+f9ta+B03Qf6OF3u31ViMnqwIJRd2ftCG5B1VqjtKGvcYnVmkI/TIZrc/CPKYufUza/V6
sSafXLERNnxwowlAurkdU/5/RXT2ehZ33R7oSXNGidg3pQg9Qc/u3Fze52KSk0gE045DEN94m1YE
Qp/ic+7QN64eelmenpYIBKZrPcyd5SB7lOZ06osblbSaUX+5A+e86vs18gECv0cgEq4b1bRg2Mhe
2veoFadH0V+St8R6PBQCpIZQUaC6QbM8nrOOHEa/20N+U4dTz81TnGhfe1899Nmbf2fK+8X916eF
oVw23fg/jyg4fuEjYUc00Vrtv8Imwusd1AQCcZkJlED/0qOuAsczxpzLg6ZETx2DEhD5TnMoiuor
u4yuAQM+Px+LP8AvWfKdFOKUzWJCE4MC2KLs1tjXrvXUOkJiHrLmXa4PfUanP2G0CXibIQY/BFWP
9OS3wkTTDWmzxzjtbPuFJwZER6H0oT1YIG5krt7xe6q5urGKm5Y23VIDEs1njyce3OLXMUY4/iYi
uMaXAN1gvIuuPIdMtTP8dLVYMYWI47y5MQ0u1CNM6MdXxgN0SwTwGFxQ2jiIY1oS5+govQqsSYbI
EPGR11QsMgKlUOyVDlX9a8lZqNpFEpIlGx1pUXEDBCDTIq8pxsroF9dB3fA8ajFVtJlBV4AzB7db
JtgEvSKeG1CNOcHdddKV83AtoTBL+RYhS/XoaTisp8r5aON68WC5to9pzOWvegRKVEtNISUbeYr5
vLke7lpYMmxBkMc8SfdtJ/Lt8C3P6f0MZTY+6yBYtuFBJVxAaGWYFTmSfJd+NMMFNg2Ec4WwLRi3
wSL7ugb0Uau5AvTKcWYi+3QDaHi43Z00qK0qwuHEZUlBQ7meAk5dKUk9CrPCF+LTuPUxxAv0Z+pp
ZHOzIBxOziasAGdx1ZyeYnNo25K7xxaCnPnjaGWY4jA9HajDWYjOztVX8tHL0uGWnvPGZ587Wv8I
3K5ow9ezsjhCu1xNYg9iM3Y1CywJQUTLXmddJ/S4EV1dvqmT00vUt9QLjsFM8GwJKy1C16BOY7sp
yFWWBf93o0ks+sfmbw3cgS1CnXPwRXmmL7PMu4KhbnQDGPeqfAq138oS3zUHJpUBg8YzFPQGTgbQ
EPBkqxIlSR2g4prn9nazgQXs5UPW04mJN0E28P4oJ0URj0+ZJwAM13dmylHmJLTPEF0t9fPZvxAs
QNjjCSrQu9k6iOPsLypv9Rl9hBrAwQMWTMcn/+5pJ5S+5f6gMX/QHOk1/ygxHsaGuqiKJb/tZFCj
WqNEL6w8/FaC6tmHECq4gqyrNHdLda82soBqZFgCdLYsD69EDWViMElo3a0UH/3p0D4BmkSt3E17
Pwh7rk7yPUznuU6LgJKdS+4FbccukzHEdmBxVTlss/+UcMZpN80CfZ3Vm2mViNI5Cp4wxbhWfCXM
PFsR5pwnDt0Pbn3Y6aqHf05K3BrSXqCWz4i/m1MV8zYc9WJSxNpgoXpbP4xlruaoMGpATXpx9LGA
jP45k68iapzoVCpchryVc21zH/UJRGyOa6hsiQnKhJElALa32ZkihrSRk5dxb03sB8TONeUVsmw+
aveagtjJZ1TfuUamxUX/ij2dtkVUdzSZ2g9kv9vBYxeLaZj8MhzQ5QOpBDj4krvf/dFf0kyUCLOi
f2+gsluHqD20Jw/czrSgl9PLuFQN6eeaLUCIuRFGT7AhFePNamVI9WD7gj/ZXlRinLrDm+IHFTEi
94N5HGJdyGbVrmTeS+av4+LCDdazdE5cHe72DZ9J45/iO1ssCgGXEraYA8m5AB1EPIbGqi6ko29Z
wktzV87Ar9bTGVjniT1yOmY1haX9jrJPO+v9DT1QgbVx9EMF6B4Uqf/bsyfnxRXmh1WpVudinDyz
3huTB8i7flL0qRdNGhJu3CPwWrKFyG2NKyXwFi7x+DsPKRRPqnaoBjTAWdwdkAmkctatBHMWnc7m
7hiLFeFFR8+TOEUwK/MiPOsu3Tvq/6Rgfj3/X6TaEkMfbyBBHqIpx3GKspZWFoGwI+aDXzRaxNhl
OZ0FcRuQ1PhCVd2QtslqNkuRGt9xdJACOaw12bbIY3UPq5f4LhqCzO3PvN6OykGS9AkAe/jQphfS
nwPNzTbycughf0sFBheQNOm6d/dkDzZmfWf2MIBLfBPIQc+ZaOgtvg3VCpAMzB5C6lnBzDWPdZgX
gOP1g8QHEP9AQlcPkrfu3UBXy2mXNBQMoEQZtCAVHJqR/90cDwmGPsVUH6VAQhELo1+xC6L9cEhe
YxADQmKD1ExyRh5MdQYjSPTlUkoPPWXDuD6VPvnaErLJW8obBf14anRFyzPH8ZUnKK7VdMPTtDap
1p3d9R+5px70LIbWdz73LLKSoprY2ZVwJvRTdoslVRFTldprzNcqqwXa16ENADaUwgDPVmCf04n3
cr44c9t1U1nDWJCEcxps5LE3etou9/9nRT2tZ9IIp3ErSM8TN16s9TugDDYegOD6c+dhSiCOE5Af
khb2r4Fj+5zHdiWZgdF1fgQch6kr02QpxszD/14D4JMW/kPEzh0Jo8tqQzdf2eCx+Se2f2HRZYz0
ft+B8T7K2FYo5R3sIbKqE8l1lX37DfIvlxPo6C/7KizJSzYwxurdhbKVN3MHjXflFGc5zDJVl83I
PXje2fQEjZpzktDb5ujOdb+y/7Y3DV1sDLJj1i2IBhFBxGKKmWQmA8Fb6to7zWE80m11/aqK9bRW
4RomXtNSIvgs4+3w0Ur3P5GkDGthVvIsCIcaoQDO++slEthxLbyVyDKDlWel4l078aJ068UgBz7o
6Kr5H05/PsY1TIFWNcK2MUfNhF3vH/wojZoUt2fMBiAjNkVs52QyheY9pLCR2rW4UmpWSN0ab49H
M3R4ZJR1u1D1YVNt8FxGqFt7nCECHWA9w/9U7VYtiVq38wF6hKDxBjV79ABrynhuSfJq65a0Z8an
hRJ2Tw7HHmPMLiWtJ+1xZ2CGmAuh7r7BF9w2Hd+DsAYj5FEdufZbKTKXzP6FU7KX2Ax6sJiiVVcG
mGzEGtdX/JNx8Xp/RT1tVsCcm3Fe1JxxDKz4BQ1CcEDZLiuc7PsbophY+gUNNcOBywht9Iutf8Gp
bwKKZG6KYDAiKxaALLzcwmzcb24lITvmx62uR2wAALg4UiW2xoKcTXBYWiigjVos13BdFy7wS0m+
X0NY2lY+ydVzyrKkg2RDq5GZUxwVdLtC3ac8PVeQ9/wqT0vvIVQp1U6HbTBhoHZ2h6tkGtLonACe
KS9WFFvTigImDXWSD6S+HY2HQKQzIYimyjhMk3R67roFHKPwG7jiMrMrJk+baaSg/OG26Rgq+xx0
zrZYmF3F8zq2mo/E84gMksO1hLX4zjLmy1FDDh3Qv+p18g/Zdx6Ud2Bd15mYOsRHi9RRkS94WNYR
aou0w2v3QzQe+0kPnfvseq9XorgVn+EMx2ciuLkuX5/DYixyW391dIhkK1qI/Yw+naLY9WlgEMWg
WsUVbTss4kuklBobot2+HtGeQhy4NKigXY2H6iyvD2nw+cpWYc7J8vyyKQ1pGu3sgrNv/6HMn1DV
Ydutm0PD6YFGaQJtx5TFguZhkKCokO0Hql7XUeChVRIK5O92r0KJxqZ/Hr/OhQimayUBbf+CVp6X
yIywNxJP3XHKojFuNfyEhbEPfJkjRx3UKo7QWFcUYGs+X3+eq+jr+Cqnk/IqKPyoZ+Zz7MuS0W2J
nE0GhP5ezQMEI1ak+kzfKVAelUWhWsiB12lxopL87A57ZY7qm+pzSK0fHwHkHG4Gw4FJ37IufkyQ
5BkJ5NHphCH+KGPfcGv6+fnp2qcWP+5jsVvmjLE8iOctglts4r359tn/Mwz+4HkUBtxxcHpK7Go9
VY45tqBE0YvvPU8tW7/Z/5y/pOVnG3qo2JUY/52ul/RXZbw6+mAB3LfEgD/cv4kZvvryXu85B1iM
fFpgboYCjHWNzsC+u1jwkuMtf+4VKbHqia5lqNjwc3buV8WJsZaS8uI3+bjf6yxSeWYy4AOqlRvz
nYqUzatuq/x0IPjBEuvQcUEZsFzKq4Gyg4Wh0ldxh9cke3jRji7eBldEjuQ9sjv1L1MztBvDtOvR
8U4W0jRr7zuCLSWtY3unX4GiDLvw8A3O6uCC9xG9JzDqpCTCoxw91K0DUpn2y/SwtHM26jNyx4Cl
jQ+XZZTl2pCPj+jZgdq+4YdJzx/53xqr8gw0/+puEglQ/iZofKfgci7nuYhsFOuMq+si85yhRe/s
TkpeMr/SmbYv8/6uwdc6TDXDYtaA5wGMDHsk+lgxuZBbLnPw1E/SIWHUD29kThFdReaTz8awgDil
SiQgEdNVBJGA/iAe80Jyhtb/BOCREasIVpXiglHgOWd1szeO8wD5SsO+3xUSQNnL5uDagLrv2OJs
ZmRtYKF0cpCCdZAlez4/qpcOsgS7XNukVgbDgKwnbyvWv5hLMTHy1L8WM14mwErVAym2G4YCyYp1
0cpGYSP9ChCb1g7eomfNtL9bTD095asfqtayOX7kvfXC7rWcepC6h3u3tMRRMIfkH0oD9gwUKdAu
ayxK7n2UNms7HOrhjU9iwziEqmN1M2qKVtJdthK8PukPlwR3Uml1zMPqG7qJDMvoG97Lu4mRP1fi
lqUVk+D/3IaH8Zu0Cff03FmzcQhROvvz0otYUhpwT0ohpNcSa8PB8Rt4wTPN8P9Yhti6bbyw/rhL
wo6eQSQXXS/dGWhU6kvn4N7E/5qwAmoOdkl0xWxAEjsJ92BRpIIUVMTl7EWinORAsf0CvYfLv6qP
YIdqSVbABiBtvtqVgBzu0dQpQVG2zeX7aUb3PKi8pQCXIFnSLywXx0frTZhTNJS+4sHK956875XT
m4k1HYW0Xb9meYBSmaEKLeC8rXFSu7U9dwSVcqqiLsd/wHtlnUQ+fLQLYR6l3r8y+VUXPjO4IxRY
1z/BiH+bxB2Rz+UWB3dQwShc3HUgg+UfZIjjea4IXpx4ScFXZzNbnQ13qwb6AfUXXevCH5OFDkCC
3F5BIFl75l1rJvfH6W9It7ihd23GiEe4iucr1tiNVT/7B0DB1oJikOsFhAk6vLSlEJKgB79RKaak
NG/uMHM8uog/+mI+3qtq8KiuVL0NUnou6NuuSNkX+tQj/7x0yDnpYFd+n6DsBL3wTaayyf88qc72
5Lbl771fVeGL5T23aI5G/yECzUVW0eZGwle7lAbDAV6ohCE3G+VD37sIWRHXk9VY3iAQOy+cXpH0
q+6ZoAJA0WM0E4sfEZ8qff18zYWOkbvS5JX8HED0X1kRVKS7wqHSLIzS0kgwzFSBFWks9e2GNiVx
IE7/MumWrcZaxSeSjBqHP6hKCMoRc0KFFAzVd7vsYD1vMGizc4pytl44T8FLyakcczA+0rQj+YgM
RAoFSqvBcEvF3Q/uGlqZ+CMXJmBPirgox3v4SGlbgP+L8YS+6TGy6576Lyv/BwUc4HheuwwcWRpJ
utfcNRW0k+nwKUgxjEFAdoRFbZtWBKJieWVfIuODnO3biVgzWrBJsFcYhahFFHOKhYIj2IGhuCjA
4/a4NCOXIrViVbAsUMpvNi1HBVOEiN/RySiRfNDoiVAkN8KyDkqT4UuLgJAujqxOEHmW9rtFW+/2
eLq/QXLSBVZUdOqBgeKHySnv8nIZw3C5NsNegBq0EgPSGmF9fK9h8BgT+7+CMLagl7vomPHJUuv/
qXSGRLShty5BgoRObzfrT9jT65vgRxYhabNC24zQgSI39LwcsZz765NKxdj8F+Nbzm+qv1ZQE5+A
l9wTNNbXYjBk+0twuxOscnbWZMS7EaTdvKMvn542l6ZVQc59uz5wPxsdtRhTnvIkL8fIgIgOJ/ed
eu72n0ove26v7l1jYpXUH6ZoIyA3tvnLsNIh4l8erQwb1a7+wjQgGpnIgMekKbZe/KxTcPFcaIPw
KyeVcsxUKYgFIJlKS0y9dAPGkTQH/18zsqeNj7JeOTIAjDgm7zzKP34+MpcHA6ePDADV5xLZoJtt
+rtDHMmUhrjxqTU9nebdgyFs1P5UmCaeybrozqfeohww44SSqwtKGAJkh4qLX7WGy7pvNOTCT/V5
0n0g/0VXjztKxS05JLatidUVPlm4LdeXTSFGJCxDcaTO69BWVoBnwWpxWNkHo46St+37lCSsWHbu
sbJgzzQ3h+JMr4jroF+uDOr1ymOJZmpcZyzr22bXxoVZHw1NxQE6uTPyj8fu6nvNoY7iX9BPrgsG
FRbaRr4Bzng4w8/pWvHrEyML91N17d0W2YNTSNXv1rOjcZTEj9FdJbBs55Hv4gx1sCuCLhNhRXjh
btSq1wCr7Y4FnyOiKsQ8xeF8vpEZRRRYj3qhE45tynSVfZizHxYDp0BdqwSebnrTZVxg3xdr+kOo
buJ0QL6Ndgt3mojhdcYWoazhfo9jCr4jDBuuhW+LDHNjZYkrXYYrrhh3gBIstgt6vV240cd0s6WD
pJyWF3RHR/tRen9nuTiBMzBPwHFcK51mP1bvvpsGK9hrEojdhDBjqxmyAooW+lW8lzvtzgXaPdKn
uiAOx/QdWcXSMzIwDKp7cqVt9K6lchU0btMB2GcLWQ/38IEXugz7uBkku4bOjlE3SbLY07Tq1OjO
c+6Kau5M6LSRAvTOXpr674LV78OIwo/82vw72Thxzn5LIk8PAwpIqlGJheplEmvagJufyNIVYu70
RBoJdciOLsv+WHlyA4vtUb2fQ5vBPHjEGydz46BbeP1ImSe6Clu5lL1D1VWHEKNHvu+ncl9aTSe5
ZiOZtlrJuh6rpOGe+KfDPDwUP9oBfJNXHJhOdGo7/jkG3xDYtfGDy059Pm9LF8a/r+J3oq2hAjSe
tChM7Q/rf6gFIi7Q50c+e98Mft7x3TLH36MTebbC3hwf52eoqpgmjjRMyDnndDZlGX7XKDaCxljB
K61FnxYumB5/ug5+g0lF4rc+geKwtd4BrQkUnhDvPgXnP5z4zCMl8Gu/YPkggA37Ir9fBVkDTaR/
5QZHdN8KTu9eZc9IN36ScXjem9B/iLCS4x0aiycEQ6I4YZJ68f+1tgmh3m6RHiLo3e3xBvvPpSzI
VZ/Hlb1N165fBVrNjWcHt5hH0ps0rQGmAG9nl+Bzi7bqHq9AMdG5HDb8xmc4KKvdn4C/uZOKaaEp
13DKAtXxD/TR/WYuhDocv2fwXqabFIqSdfuxN7QFS5wrTf6VVdelxNijl+7Tt1CldQ8RV3IGkrIq
NToe+cCYnE0fQ71YlNpuKPCh3Eh76DeIEzLKXxt2dcOqbty7chNjE7CxV74fc0NmkEqZUnBMlDp1
pUVVGQuGvJrdhSGK9mmgPMMdHJFz/RdOV0wYJrC7z8EDg7Ysrl5EMnqHpJRpercXr808bjqTvYhS
VeBkBzP/2xmXuqc7vDBlngGxiECL41h7yrWJd0jcSu5Gr8WBhUHOt7jc+66MqwpxM0viVMxJdM7Z
6nsnqrUOK6msZnnm4y96gZuKua20gRlvuTMNS8k28uHW/d50LpPc17dTTv8uoXL4LMfj8XmTgW/o
ufyr6Q0GMkgAaZeVOwggtT2lC5ZmTHOcnUx5gJNgSX0lhXQaAWFK0heu+qrR8Wxpd8FMObHB6cM2
dRpgvZ4M2B4zVPJ20XEU7yhI9eQ1XTXujC/rt3eC1CRe2demMD6d1fyyqsSL8tRAl6vkynIdKJHq
atc8mZ7QS42uPRntD/ZpQLQiWFO7h6dqYotNWXTJc5er674efG708IHhXwHEGz6nzdwTA+tuTt4I
SZ/kz33/8NnHqsPbItlguc/Z/Bh0u54wqZCQI+EMZDS1fFRGCxvj4T/KibCpin+iUCj8EQKe+zFZ
4mn4iX27t4BDzltJVAf7nswZtUXC7wGILCwFhaThQv6t6UEaQpxXzwAzX7PTFo7W2uWKMCpvTPjC
DE1nsQQzp4HAwji/wcIf0lpnFLraHEs2FZoTlSIjk4VGetpNdMp+KnTxsGCiXWh1irgQcHIvNGD5
9k4/bCAHu+ZW/cPnnqL+Wryeh49kpgiwPXb+s+sx3YREpFSw0OUmpWYPA5upHw8Ph9o46/BWVBs3
w9uFHoXozhg4QbygpeqBGaX0WnG8L2cV/JcwVYr2bRjYflJSCTlTzuGphiNW5F49dz5xkzLdjH6W
ySLQ/nxyHeDDbCcSDsZf40OfszRI8SmJUoDagZi8k3cTtjEl2j41ef/WkAdU/DUyLCdh4ftZG91n
6GGobPU1YySB7TAawow+o5O8m06cn0g/tDCB+3vJGRezHdW2hC0TnxEFs6WyCDmP3U0rjRrAW76I
W2M/wZiffXtYB0FARmwQBgU3e+VfDWViwPCRPmDoLSZ6DN29rE+tKeE+6JNtYQjlVMQHnnUxeYnO
9PDB3ncR7b2CcFRhEfCSEcbcTCvnV2T03vpM8bN19ZQl++DMtcfXlOZoEdkr5E6qxsbqDR2dn9c5
cDrWjiW5oillXPJCwzY/yTmheTGQ3aFexsJyq8HP4qbX1IM0C/7IzvoyNXvLhEtfg2TBPcQ9cGNJ
c8u4ZqutQJPaF9tBLCcVcsPuIjq7iZNBH3iB9P8r+V8I5hWlsnE9OLx839IYbfQPGUAV5OB49GmD
1nt8caRFdQTeWA+wGmZYBoBnldwdZE6V+JBS1sBkmafkHduitmO6GU5U/sNUizW5TrSt6QA1tpkE
zi70S8iQTwneSYpZj8BVXsof7Mg1ErtEayW9sBEfDOhyNgOu6eZPuofltSqEvyRe2wq0vYYI+mpZ
IbEOg9eYpy4THNY78FIfkFJ+M+zggY3Mb0u8DKop0lscLnA7MjDgjfcLgOIvksAimoIg0WkkD9Ev
aZHibKDKNHJaVJY2tjDlimdFvzK6uJpx8BOxm9YMOmW3zvceHPMov5Hj5kY83qA5MIkOyORnH7sa
Gx89pEoVtMeAKQZxwlQL342Z2NXWUoRXQA2eiIOzGwmHpBW3puPCUvBhuwdM0Uimz/hmzVOHQGMZ
HtivIWoAh8HSjZKlLz6MAb756HNVNBQF/uBfTyTOnabeDufdKHMWrmm7nm9T9Y8YDAX4KnnTcKCM
O5gASGJP0Pm3G64jyCJewMu5UvKKTdtGDWfx2YPHGNw0AxX5ci52ipsOMKukNCiSK0yHUDwx9zIe
opsvKeYPnOzkkoI16wJOj9N6AWVYHg2KkbwhTqGGlIJqgX0csJtJXKJIKt5B5RDej/QEIJXCroHs
SKpnxgJWRj7nszewSq1ZqowQ+8J7SIxJx4rpB6LW7drkkClsrCxn3FCH+Kq/RdC2sp9tk31NygRq
fOWqedxT49PFKVmh8PZxmHc4N5fCqLR8HJojkDbz45Z6OJfz9QeXHNX1OFxmEjtvuMOlhzK5lyOR
NZcTzPAq/nqQQyP4DRjtvdCytr+ulY/RRlBkczqrDyVGQN70zCXZiBfA1Z4kioOHWipcQroLy/Fv
IGdCBbiIAul/GYK/7rHfMK8O5JvqrO9+tfRT2w39vMP1f5FDIlUKF4Nxd/QKUakhFsfL8k5vo+s7
rqiXJngRqZyQWHILQe1FsbEQLXjFjJXJSo/6xe8zO6bzX4x85dRwyjKEYTYVt4kMZwTd7jpe+qNO
7DU6GeDxgar2R5tWLSsUCx/7KoH0vhPYBfLZlnd8I7hAqDsVPQlOzjxCtuM08k/nL0nDO+tuWk8W
Yyja6QlYEHvmHKrAdjSZmjvLFxwQRSldObu/eniPuRpmYoQrh5rpjEscwo2QbLJaDWo2qxZcX/gH
EP+wMltpObX/CvGkYRCCYy21TnQAYxviCN/xNLv3q3VmnWk0eGgl5aZwM2toxD+IpQYTFTduo9vj
osGkNMKGu+/F8HdNr87ZCOBBuLr49GDuDB4Ln9krXDhEJZ7HvL13VCqvDQfCqCMzWPNSqdTe6xZp
F/OnTBLm8xTlFo8PtPnMRtpD9y0xeGey1ekeRhbjlOb0CaOiGXF5dZZkF8YHa33lOGiv48C9svCU
Kxv8NRMiGdC1+yW3z+Cu8rd3gUwy0NgfO08jTSzg//IdCxjj/xC9YUaS0XN05upoPpEQfW8AdTE7
OM1TPOVid/H+pEBIJmR/hphfM8u8MPb2TY0vQ4p18pL7CYdCUf/FcD4LaE8dyYdg12wzDvgkmXD7
ZLOHxP8lQVJCHFqDTwTjCbh9OgDEnbSOySxKhPsscTIqxOOZcX4ysF8WgDZTBY/V3VS7dppAQ5MX
fWth+9bvfFjB9Yg6eTpwSjVl4wHoTVp51KoueFv25aeos95YBPuih63XpkyPHDeCoa6TxoW9r6VF
DU5QGlQGmfhPz/DHNOVSuOeNqoHjJXbjdVsXJ2ii4dQr8xZ8KDPo89yEPP3TTdatooup6Pm7SeQf
jopsLUDGasobwUNHB0WRAGVRPfkePLWNUgbUFzI12cQU52/CCLCZyJOC6KJZea1dIPghBoZjtWAq
uvAxfFagTzDDrJkVLnAN4qRnfvKEeGdlo5jFf1iF3GLWjoKUlGWIFAKvo8tBwXuXo2fdYtCC+2Dv
YFH6rfCuSl+nFKwo8zSV6qdzzOeLnNNP4cKm3JSH2APsJOdC0lIa5t1GT55SygWNERKCplPrBlwe
Lu5y/PYdxmji0NJjN2MtiHEp9T7qLtpKP4d/Ungfz7FTLfYmwpa0dcjVM0fFdTWQBnBaylZogBbU
n1EsTeZokvSJI4BUahlb00cTks/XjcmrJeFbNZXto4Tg99nxvAuS7FZ4wz+/MTfx16C4PivJvOnq
T8fhdj4aTjquSyWlSYCgHfFLI63vK3oUuS97SFZMXBtvY9v0cH1OSUWFgF8PUEzksrM6gqXpvG9P
FnLCooIKW+8XfXESXT1gWWmdvdiW7WJ9htC5ZKxttKqtF1Q9fHrje1TruBM8IbvzFxhU5Gyt2yn5
WsxImEG/mP78rOw3nW6ua5c1Qy4dYjPLUzTcbIMXLfxM/fUOTjDapikXOfV+0Hj4v11688b9ZcmM
l9YO6W3l6EbObJea8T+TFDahW2g5i4cwUM1/QALnr+xGTS36/yvo0F8hU1RLD+rnVisgGtibi9QI
KlMPj5gVa2jClQQUbtNQ2AArNTYjGTNcD4Vp+fgINIT40miAoyxoO/RaaQ78er631dRtEGr9X1Ij
pZFb1AcGkaBxNVZJVVrg1obMHiTOxvnZZ4a5/kaQG29+aNtsTpiRIG5+LrNLGe3jmdVX/WO1/DrD
27eIuclKTMOpJRQkavLDI777smhD0qEaqJZ7A2Ly3MyD0sLZ2pNEWNvhMq96LXQblLUSzFTADXBE
3LgMS6cuhjb4LkNLlD9hlxp2BbvMek51FP4fbWyzgjJcg+CCByDm6vyznsBGwAa475r6PCGW3jYx
7T7LE7fGD5jQAyKI9xQPWSnKFYBiOk9DO55LDEZ5yhUq94/tnsFJ+VdevCO8hKN+wMg/GgBcRQE6
RMQPfocisOomAk/hmyAlCcbMHOHczXfgKr3pFxtvhxtWJykHjsnBJTzfd1GXWZHEQe7kZvwOAgYB
cTDj1wbWaqKmjuLrWU044DmDC3+lS51qqca54f38AzZUI0foMMgVuZP1WEYCpFBG75yy9YO4FHxr
9np0kaCdevg5BLWVHP/ekazwasb8KcXu6ebkLCuFoVdxd2RJ9kFBjUpdBlswBJ64KX5iB2RLJ1bh
EIHM11uvjez5jdFNnPQj62rc6HpYQZYaGj3iQ7kylncpTGJ951Cfy8LYAhRrckxydaI7x6IP9MFB
d7oC3VXlgDnIcZ7Cau/ZlzqzM5r4KaptoybetF/BqGKoPGDfgmaPG74HsBNPEqvMp/9oGgSMnwTB
mvVU28QYvsNCD6CveMuj3MVee7zCKbCt7/Plkzz952l1ajOr21TgloG9qwYUnsVesgwbiv/2Nszs
XhTjHvrFcueawcsI1AF+Vbu9yW+YrpjEgYdot5cINtBIDppzEfeIRqG3OkyrsATsrZJjEpftUls8
41+veEe9UJR0SU/7bIW/4hVdXIqp+qi5adtUhODhh8M/DIf7ccpKMNyFkJ9F7/9Dgt8dj8cNY8hS
trHYxSo1kfqdRVjRNVkGnK8ELhqeLnrSrxBZSGAkMM2mrhq0appl/c5PEzBqKoU2DJYSmiomvsVE
FV3wQbyu14LBymnhZeT0sDTBKIUcdkcBoZA3fpoQh70WuuKFyQeOFWHiUmtwizITI+RYVclvGevA
6sIT5QX0wa1vX3bJ3Z6UBhqy4GS7exqfiqla4HbHFm/Pas91+dnvOQ2t40K1sVLV/87TwT2o5ct9
8LL9z5gDY5p2z5ccI/SEhgkBl+XrUpatG6lLOkb4Chf/8kTYSmUJUQTrmQtutlLI7l7lc0BAu5gz
YAOm1KifjQ+54AaN8h9ewZAi/cWTaf19YMK6Fb/lk6VFRWEBWI6HRI7lw5i8bYoPJxzkuwl/zqsX
0RABes5ooQbhE3+Urt4YJoBBORmdVidz378OaZ6P9tOzfd0AKpvC0qBkAsQ4dh6/SnmPUbovoYbt
RLzYjYLxddwPWRsmt/A+8PFoYYUUkOjHOzouPtoOMHxoCAT1wVZ2HZlxl9CUe5RoVWGYTL51DaIG
ZMDqS5rj0o3r/lO7jpwV0TAWdLFF82OKIfjlhR4qPg+ABKx4QSF2H4x5icjKhs8qCf6YA1n5dEe9
/VHaxnRGLJbxjONo7lASeuFcqdC3Nx8TlWNvoEYoiF/4v/juNrCMpBslyByGBaSczTYqot4OFF1M
U5f0u5t58a3OEKYdJ+kZwJyiC8Z8eYmggntC0aC83NnwOtZxYyIkQGaA2QLywf1jTvcbuopPzaEk
vcyFMX43+ByGDpEEhnhUFJ89MUrjYVSCW4VmEYLe7uGdi5zG27lMH+WwAjEOELAuCT/nbNQf7OQ3
qn9fjq5SQVcPLiUhhutZWczHe5mwopZEhZHDCPO/8FeCIrvdE9yphzo89DikegM1Uo8IofZqQW0+
bKfmZr5iYeEJXEzK7tMeuRz6dhikHLPDptT0+mP/R/lq903HwAcFcf5QIlz4g0MEGU01gJ4nOnet
GxFXzLqrERxd21OdSa2VCHbvTZe3fNa7yY6IkNGfWT6/wISbUvuSCv/9clXPLdrDJszylATbIavV
B0dBaw5jh2gKpMlDPwlYw7EEhBpjzn7267gap5Kz3tHZY+WfCVScx3q0MW4mx1uI+pT2Ox0BIej1
jfZtrybAbGmV6wpl2B+S7Nz/LZ4X9YIpCpN063NtH7WFpXP56qhaR8cWsgX5KUh76rGZfYOfbJmM
NpER0kxKoVl4DDJPu49dWh+/nE9B66QyV5Zhr7DUCmpumnOXRPXo4zdg8QcIJeLjKyptEQ4M1Ohs
WhyF//sDj2lta4bjc8xauedOPQleWuuoWgrjmgloy/NUM2ReB2/E90Dg0aM+wycqtBnRWA0ekifW
0/DNz3Upt5iR13jA3GR2FTrU70p7dI0rg6Uujji/+1c7JavbkYEawa1LQbv/utSi+krb4INj9VHP
14/6AMglID+qJu803AKJNxuLgqIBtdBOYrLprwKVkDG/hCshCPtrpjtI+t5BfoFicvCkGwanM8Up
adeZJQsuLXLvLa5ewO6aExFHr6blp6ObEoB1I9dauNWiVmhrQ5UISkAk3r+hKkKmhtxblmoswd4+
E5HcaChaF54eR7xo1pKEW16j2Aa9H/+iOgEYwWzHx1Trq+VQv1SeOyHYG6KzLmW1w2MGSIdA9IJa
u2oEnGRjhlih6k/XmmM2XYXQwSus4P2LrNl7WLHyT6DQP3Jy3yeo+O/453I3E09kYoBfMgrx2EbM
6oXKNFvHLuaAHnK1OcnqbWGr/B1f+Z9QT+F6L/ojZEDND+H5qJ+fRX8S2MGk0di62cjDauRdiFiw
yJd0L4xbaT3P7TdZc1aG1PKqZmjACCqaOP53orgdaSvzGNZX9TlrEV8oatwWHWN113bhlCtWmr8k
xUqJcLedpXInYN4miafJI6bKq/vo8kmHzW0gDwdzoaC5iau4NyVQKecuffNX+Lrp7RMGdPHqMosk
1PDXZ/M/mDcm96mvsUKu1RrJ83zfflmb13e6fGg8l0UjOVWRWCQ/1t+Z9qbnh2kSB2tqtYN9Q/QO
wlxozNRu2ObR8h7D3mu1qY2CAMXIwZiuyEZu04aR3AqvnTDIykOij4cmIzcXyxI9cK7sjFBH+IiY
Ashl5dO2Kk3do0o3ylODsWWfzl3tzVsAgtVcdOFpYe/nLoqqtwecoQsT8mZ3wZJcuHdTJMFHC5hZ
C4xi9DO/e7wcnBe2EhCSanPE4J6xrnEJmiUFSHY6pGpuCWwowMdSkqE39zkY8OWdWiPt8RbzFY7B
wlgeIILnp3yEFaWHpi8jlJ4dUV/gVfrmZuZf66Hv58hzKFCKo0YyP5K4aG6fD5tmlPnQjwSBT2Wd
I5lPWuOsnrhq11XcM8lDLFNvm9g4gYdLCHnhmhgdeM8k88bJXl3ER3Ygkz1O2tigIfdi2DliTJ5V
6irOTcQB5kRderV31lydhlDN6vi/XQeIHwSsIN11cAALcmPJ5JoUsP1jCI7PoJ55wZXOHTIonnBy
02rG/4sQwlh5+TLsJOSsQ3nhAddbUr9NHBqcb/Af0KB+wV5OBkO56cyK17t2+fMp7DppXm0N3chT
PHOpqHNLbfY2fDJD4VLHSf+NW+HLZqK0MWOutChQrxzQzp6i85CWzXHOOuZcX6qSct4EiAAucuVB
haC+B3l1wuRM1Cq1Hub4Vgt4HVrxOoWJL+Twlhs0XcbojZikhbTPyFZgug6+8qn1wkAR8KtVoMkk
VYhDfZ+TJdJvRffW4Cmkl6nRtKM5uObuMeOYTYu1I/JmSeYJQTK1wsVTL52/h9t2A5feI6V2Efuz
j7yNC2baxAAI3UyLSnprDcTsK/g4lYzV+mBeJ9NJC6BIkTdwm6cB+KF4RjbRjdSuzI1wjgxMJHxx
22kDLyF3QQXzvgPKnKGWNd47k8LRdRumqDeAHurkqZK6C9mM9c0J9ruDvIi0ZZFF+YfJ56GcSsM+
FX+rkSFun6fqhpSJ0iEuljOtQRNbMsgk52y4wFqNUbxrQP26uy3WLq/MFo01A676A4eac7qaBCIQ
Uy9y8mWj0tvZyI8nBMLwuJB+3Sa4aO32uFV09Sd1WdMROE4qMPbOekxW7bM/hVshua2F/4pUMJ2K
NVbst3CUFI1FP2M8NI268rFSJR+OUJ6cx1D0OzqQ55PUynufdV7WFAnGKVjlhH9kUEkV6benENX+
omWp/syciCWz/UFkKHcBVwYf3HhPAFBoBa/zweaUGIcn5c5+VzjfsSNaNpGbWs3gScGAt1QBx4xe
Nv0og5TiTJqGREsh5Ydj5uUJTbwNuDrVPHgfvJx5RznmmhF98xrv6z9WGF47/EbD22cG9BXs0Ru7
AlhKGRSg46kpWkewFztrowunHV3GVGza8XDO/lM9HfyqNot4RJhHSayBSiWrMrpiGrmBwGbeireB
z27j8NIBVS7uT7oyUE5O8FO39Ww4KsD1JWskQrRQ3vHzZZCcwvbhwkobpacWE2qdFnTY+8G+7XeL
fpa3hiRrMTz4zA0PDBMZMjjYerdVFUpONZEkOAfXsYiKMFcuIgLg4ZDLrdYUAtuU2AAjDmp4NGpN
edJSLNxOUAheXo/p8Nv5Cxn8ILn5G7Lnj+F/46d2cHL7axiDJu73QdMGalB20TMOUyRbk8ys+0R2
uclXyywtHpU8sKIajKrKRgVwWYOgwTw2xFufhgdHXsW3N/jNDw7S31UXrxSHY6vL2+xI4HjjIJNX
vu5ZeiTf/4TPaHcv2GxePn85VN+s0q7/DFWvgMMImYUb2RYcx/XZg0eU7rxQnkTnwOjN3TrHnN1m
I2ZhvIu/0c02X+DC5R77EzCMNAzRimfMfdAEG7t6ikBwlcok57/mkykCyFAU36eattCWVrIUgJIQ
7xZD2tutDXBbjKFovTgxNOxAS3KGCFitfyTD0HNTADz25bZjRbP/0lnCxlci0d3Eo+CfhC5Mk0p6
RBPLwqtxZZ5zqGubPaui7foR3gwCR4Iq0l6Vuazm3bMKssRwy63OA+yQ8UyaRIldiV8bEmzuUMwb
/KBFUaRfjseMI5kBAsAWIz31BQ3MFglhTvApc47i1A64wUO8mvuV2ktETOfCb5Km6TUnTKfrsPoo
4c53p3Q3bIcNNAcBnNDL8mrkLblLUgyynDsgCd+cq5h26+skX3+OZaFtKEED44VTdwjQKh3mBm8w
eT0EjsAPkbJ391TW9gZqjY5gfoBrj5Fr5+2PS2mniGU6jou31P1z3g+M+A+iUaDcp26M9O/IUAiF
2/M9A4nLGbXnTb/ZtVn1OS6XkZCvA0jA1fVf93eEOaZhAS6+9vOseqJ230vxyfnquv22SKom0n/N
YIYO+kvBam7Mi3FuOaVhBbW3gb43js5QK1lXcXkCQdpfUoflM1pXVnFN1dXDlPLzG2E0/IcriNAK
PfZiixTkSlSH+CXwFjhrWParOHL48ApjIaLZXqCBXD6Imt7mloF6mcOzEOKNUWa/IgvoU2duNd+8
fuMOtuquVnn3rlsy9G/T/KjT7AfMmzqbdYVStvpAyYar2ycrfWA4YJVcL4DMjhIjJA/MITOHGxAN
DINHSrsmUDtMrsQsSOR70oKzUdOdBLbxLQMlu4YSNxyW7Hgpmf2L3p9Xrx9UlIwFCSZ332I12der
iBqUPaYa6zpOI2FqWvCFUMdoY6rIvSUpL8lfiAJoFqsYrNh5uj6iNO3O/8vM8CSxnEKH00T7jWMM
3hR5GiNir3ys8CGG8tInmMf3KIoXwRfU57Kdtrs/QYmH8HPOxZ+DFtaLrAjyeacEfj1RoaY894Y9
LfE191cxQlCEs4YfMX+43wzgnT7xJH0RL3pMrQWj8oImSJoDFQ34YRA5zHpA6+OUyXOjN7vHmtaC
Sg+64TWM3gdXsgxf7ug9VBi7VRhGzJwpAQ6Wi98nhM6cYXjWznKrQTajzn09UTyzzD8EIuNsutgB
5UorC7cWFtEeHoZzAXIHuw23LmH55NpempIaTYhG1rVRBLcWWFRTFodn14VBq0AV1wpkWVQHNCah
S7F5g5vvOoUBRqvVblt9GqZX/9O9WljtoBiUeo9bE0pqPnsrspN515Z7I48xDOB88iT3V3x/5fD8
IecSXQWcG+nuPRDseJlQ/yAVHV+4Bh4uhF0HJbX8uOZk6rSfCXObtGB3VpP7wlyizhOGsvMlld1v
rIxDsOyyWxm2cC/RI3KvpZzWNTQR9RYQQ95+/ycGmhdxb9jBfU7qXk6HNUL7vqPYOpAVg2oQvFLa
/2rx0fdkO7dQuFYWw+1qgzHLUxtF9fBtSmv5kp6TRcCpnUriOkLDrTc4cS8iYI101cYREn2lIdPZ
kpXXKvkfEONIzV8QGihuodolLzqHIolrv7hS53/9w+Vfg29dftQXpse5F8icUIg3kyR1E7GhPpn3
kdvCGkP0xF978hFmJEzHsNPFV2bPIbbkxpKiCOJPQurBeKjxVNxseSGxn/d8MwZ7JMLh1VLvpIaz
2Q5i5ur+0tCqPgq23QRtLE46TggMxhnZLtIvgaUeVZg7D9wPWne7K5RtYChI8fy38fZHQKX281/c
4AmBMOxXdR3V7b7+crtDysq8iJYlwzjpp3icvjtghNB7BxHCEUtRWxutjxWxOB+1qMByUi1vW3wr
11KJp9vdeqVENwI5LPp5pnv59thCh96tpDKht3T12abfqk5uBv///JEnplShflVDHeeOSG8airGR
Hp74rpXDMqm5/rn5/i2bOdaLa3Udaz0OLkLAar25rX6/Ck8LrTL74vo/bZeyOlLcDnvBa47Gix7n
7GHayqBxVeGo3Hz61ortugANtiFOPnSxV9PDt8NVaKDIm6j1LZhGRuAUZoSETtRmczjKEaRgY6Kh
GXVufJCFMs9CuV88RibCgfyUQhO2EQX0kffI7K7oPUNHS8p10nTYVWXMLqMg4UDz6Myqi0gdLSau
3dGsWSvtZRGKkibFBUcvW9+fi1DeCPQyw/pBO+1bXhyQEMklExeKwfavmHIvbkbA5uESh3qpo2N0
VjludJRzyNUQv7zhIA4AkridOqOXhsZVyIir/B6Bgm1NrrQDTvQObeifBni+vTcFNuzEGPLbn9ob
aII2LfWMeOAUXw8+5EpdwQFvyZx6KElrTTLpDyOpgdfxmysTd3zyzcVOLNDl5mJkyjgXaC0PvLfH
iFL27Z+2cthGtd6TzKPRQ2MQZRKgr2z248mI/2IqR2g07/J2rX56jrfokIrLZ2rn2uARULS1WLFV
JZSbnVJCkEwWEpTg1xM/66hSY7L62VJCib8xtslB2CLG+D0xsLJAwJAY54v1Sv0mVt8APa/3LeyM
Cp7MU9/UMkGuFpBfRtWMi+kqwfSk6b94sCs8GzVYPTM+6s7w8c/+ppox0d8y8clipResIOJVf8fn
9xQnn7J3UJv6itqK1PctR16MAjiruKyZ7EziJLnJN74n/TwfM237DGwuM1usRhq9K+rV5OVDq+MB
p7KqBpPVy6R8LcNSNVmWuMe4+o5koBxwi/q+RyEbpmluu9t+KmveccHRbMARfTPt/ELNK46KhfzV
ZVYEhNlBoorHhJ5Vw9RZ0lJR0/CMCLx+OH++vDBmJshXUjOE9O2cpKElX9av+BreNqMQ6MhsmCiS
lvcu4BlX8I5zjK+YG2afVA5LMEOjeDEnLWMzTVS33CjBTS1753ltouSnggwPZ2pxQ3ztKS1ifH2a
HEqKIRFA2e0yslhAr6rT0pLd0SIo0jnl9vM9Mkkj3pw6Fws1lN3Y2mgdeOFxeAJ2JJFS4yaXgqGg
TsWaqfwP4pxkcfTUssbGK0YCkOhwIMQkyuaplWsU4QOyj+bQcxvGyQlJsofdKitElRamYttBTck5
nIry3rUbeNuQQlWXKUFnK5NnEfVaOuyE9lfKt4Tr3+2nUIWMbXKWD5J6Uij8U2EpnEDUtRPlQc/6
9k2xOdNMD5MLBnR3fE2JmJtSMXEbA4vOWBtl99u/Pd9fbmaI1MDMMmN/tc2yq3VVIzQqHhKRWnlQ
uPMrh34ge+q1sL4YhatDr61k0Q0MRmlZBdMXMb8pIqU9V1joISFqgTXW9GjKHjosf5RC11NmFQqg
QOXVkKsbMOf+4oX/LB7g16pq7VfsMMSSox7pzcIM+Oe4hsXftl5z8N3IEG9WMGtbCmhjXRWCwZhn
EAg9+Wpvt9yoZnucFLXKwiIBTHHYbCv7g+Rx6y6ewaShd6uaQpajI/c5n9j6SbfArhI4NJu7lGFm
LpN1EohexuTKMg6vyQu97sbMT1/wawuQkacTNp4MaOMusb7zzfWMJ3WtBBkwvALPYckR8D3O3Q84
pNLLamiw4OybS2ekNDuu/xFm2qEb3BT1lo652uxbwDQGJUimffNN6g1iOPD+uthpdlUuEcEzz+nw
i0OuMvftFTSTXYARPZEFZcoHr7zHUA6dCiJZMjGFNlAmR5OdXE+w/5uIvlzwnumtgZ/uhPXflMZQ
kt9Jg8B6V83q/3M3UAcvO5ydi6OhfDn2WLcKB/uknrwPcbkOGEs4FG6KWiRmsEyNtGcjr0ytAsGh
NZ3BB7uhbV06Q0Ifb2q3bZYOxqUyMXA87x173uUJ+gqEIwrUQZyDDw8u9fQEphNbr8VHFzFIMnJd
c7vJMl8LApDGRQlLrjvL/Our9Sx7eQ38VsT8W83f9j2Cwip4jzpelBGYroPKbudOl2CsQogN7BF3
OFJqgAY1nUUrb+6SVqXE0n495iYND/jMvPBLUH3WJZOnTOtuMyMOgoCorb+9FsDpc5eLMShkN/Bg
lLIwXL/hpt9YfDKQYP4XMYHDqrAIX27vbk6r+6b/EGfoDfwbKErQc0ZDRY0OIFDY34eybYRk3KNC
WIwW8DeVr7h9QAsCtKYxhohUiqDf9qou1I0Hlc8Td3bA0JpFMNDW09qGB9JGiXkXICMEHv1YXZwQ
3F+6qs/06wDe332exXu7PCsFLdRnaZBV016aDw3ggB5qJGsWFFskWX/HS/nH3CfcrxFgqxoMihJ3
/CNjRGyMHvEg1en5NeIGpBuPN6HUrOO3D93bnhKqyKSU4SY1fjLzxQ8YHTjXvGqMx21dZ89Jdb73
vmTAaiaPyPWSztdGU1vRkbhWrRUyly7lzH83y0bFnjmZq82rNfDo+uDrM+921btQgQWxwoGYs0oa
eeoi1cTK/J57X6XH1OnTFcB5sXBLOSrX3e0ZJ0TMHPOtFGfVrPJ4nxhOdAzdPSTmwvhB4/zRRVRN
dAG6JFU7g/BFwuhBM9frY96lRU6Ol8VZsQTpWX4vAfDwoGPHRVsExHKtlenuS4xxQN9S4MLhjPwX
UiKwOJR17MhFTvqrNfdjvLjHlWXo0YbMN1P7uBJkRGvhFcilZih45+TXF6Mo+1naVeGI3cgSH/bT
RduLjYTA/de5BjBVrCKRRAPQx2znd6wwW27w+YYKiUpI1sKca+SKi6teRp/By28Lt20NL/8zcbBW
vXvbvqF4BvbfIkDL/+fHIlNOV6YvkRd3vjuX6pu4vcCUQw7etwduSHIm8xOc+z6PUqnp6K2F5PLs
MJg6FZhwTA08yf/PeFr4CTqJhDcWVu1vp9A8Dgfl+rMW5/T+sXOxj0OZpol1c3txrQnLJfW9hdhx
Nhsf7JMwNeyc5rr1jYHApMCch2USZbJcONwFGtk27mPq91HNjul62Yqe2KIZ6OZ5vi3VtV9Vkcn2
qygZkqO3c6XngYG4u/RTKjcpafRr62GCRkHAM+m8Y5dbSKGt3dNQgj4bnofpqlxfPUJiCOIS0jAW
xxRLktwGtfYJCOM0f25iZInAAoxT/MxnPHDP9H30BpHnL/yJNHZ/TXp0rIKwxz1tZo1CPrwKS1rN
o8wIRvziLqtNvhINC2UjlP1CC3U+v9vjCksr16/moiryQpGr8ZYYeckItkUzrQ7RxdEEKUuaDXh1
ykeZBLSfFfiaYBHA3WgeHltuGNWWJdA77OjoA9cn9VWB6shH3HJIVvk+RXLqNT3S+vHx4xwnDYEb
IuxDBzt1TqpoWoI2rDnSvPUoDDi6Ux17yMNuIki76CcKtJ2qI9hOoc00yBlcoJHTYucm85oH6HGp
3hbmetJfrMV21WmCuOGgXVQa4UHtwiLQgrpEcw6KQMJRHmBbs//MFI+WhWK5b0ESQGdn3LcIJAJK
G1Vbwe8LR1RHqlliPS+oPMHj0Bmxw+AXFx6YQoBKPVHzVecgR+0cQoe/hvLxxON3LIDW6ZMOrVhx
2N7BmJKKHcjpC4wSlMuujEpYX1s4+U1aVukPt6nMW+uUN33mBOK0Bsz8RquEr+nZFYRebX157OFr
dETo74PAQqS5Iqs86WZFICk6vZa6eqqocgcbDRLlyt2EE/vpJdFn0ANEkXbwjs2CrlVajIEhEr9a
IHrPDjmsCNzFoQP9Ntzy5nyLvPYK+onXKXB0/eHJrsZngh0UoTl85a9NPUDNv4JClp282wiR70eN
rED0eVtRocrophFDqtOqbAplKbk42N8zvZqVo6ZRNNs2PhE9nAQahNb0snJ6MkHNcohZtDLAXQ6M
qU2KiZCbteXRXlK+e4qL/9T84ztTCmvkDvajgL7kjTHE3Dw/GKo7B06n0M6t+6mRMcxiAY6v2gkS
9khk3bQXHASjxfGlONAAmPHNFsS0cm0APw/iAXPCzlgpU8T+s9FAGAViwDxUUkK+0c3O5CC4wCh1
CcHecMAInxY2NHahseAyVOtc0VQ07wTgSD2OKcNk5wiawR6pCDjn0ADpZBVn3k7DDGGF2O7cLmaf
CGSBhH7AVHO2eJl/5PmaGW5zAyg2nJXsmORS7907nb/O89CPrLkFbY/fSUSezuq8Ktdt3GwXe5re
QIaTnwbyHVE6897mkNvxfIxD3AKudHCs9uXRjE509OOnmzRxcKSPMqpA/dfQDR3xDTXmUeYdfAUh
cVIxVtM/X5NrZ+SCsAh0PXJ4BEB2xc2Y+l71xUrwEXAEhVtA2YZDpXn4A7Ec8GQHa7bERSKT/FGx
ZjO9yeBmdQO0YrRHiFiydxh945VVSx1ubw0e3+nlVj2XI1oozN0pSrQu6iT16V3/yYxdfL/diOyr
SJcIFxE+33lVrZw7es7lswtidk+p7TfmMS/mvv/8131OhjvbyJZAo1LrVnMzvidsqygk2sU0Wpav
RP0APtVdmttYVqvM+ccabBo7UX/B3MQdcGd0llzeqej7Mu+OgQvmyfCSLjCjpKgU6GfeCn7NkQCb
Ygei3h0bR3UneBOl8+wi3eOwAduB4rutKKKOY4gAiC2Z+qirtWAlpD4FqCYKlSxY3UvyNcNqr/hh
ZwAfPcs/Gy64z4/rpdkpvX5p1sWavHDh46i6jReojpQELaf728N+reOcSl8IZKMvWqWbdiqaEqfV
eIjmhAxnOMydURgextNYpbbXf3oX0Kd+E2SC+V6KNcYqqhB1EydMuGezjm/dQ/mwVidFQqn/cC+x
adN/f1eGXs7S6FdWnpwPxGxjqZUAdjyTk3/eCXBv/DbIk/o8y/nY6YYv2kH+OUL1DptKVkajyg+c
VUcWYc5/t3HNoodTiy2wVZUMOqmiweYLKj3apTRMrpjnVAccAQPVxYIWObng2kNx3Bc2iIxwPNWr
iNaBsYJ91OPG/5/G2O/4eIt4piGVFAjHqt0J8SHWSrDS4kFiUftWhWiNFzYj5k0t6qDOIcwmzAfN
H1dTewlTtaGgiNsaoQMX/lj1JEOm1sUlzHwMAR4OPKUm5GSDPxZGUxpg619Z759UBb0k2mITfHLm
lvVEKapupy+PMrTk1rlzoNuAtWJAH6XhyTfPvKo4IRVXvATCXhNH6LmqxyLf/DVfhUqPhILhPxIb
N8fniaUYFMPSxNddDy3Q0o1rby8+oLGiABFpdH3hxzoZ5HQgsoNe5rh6BwBeNdDPNMj7sYZFpVTK
z8ig2X3XuZw7eI6LU4K4mbgLMaw8ABjaUNhogUILNe/dxNRJukZGPfIFsxe62ZAJUittXawYhOd+
9ef55n39iKWcTU2pglDKdDI2vPeaId6buDeljh/YQPLmDt2boczk9b54LtpwPb5WrT1L9kW8oJ3M
VJVGS207fJMIgRngDh1liRK38n4AGuf8o2uQ/yeXrbjNu2ujauitjRDHyDs41hieIF1GHug3Y2Wp
MWUesaKB3f+J5k23MwbrsFXtPiHPQziiJuhIc/C/tO3nKjHxksjnLRNRYTH1HTqBmjsoczAfeW30
IQLbgjvogpbEGe+WrrM2HpR12BBdrkZXmT4M1ep2A9IIliplaMhmiORKOwYhSnJ20W2+s7VQ2KPW
VZmTYcg5qIHJ4jpC8OMoHvnwBP+lU5bxWPrp5xTbOr1ROcX6jNwcHFUsxIvlO/YjZOTLAkW6+MKf
je3oDSSesI5Rpj/XcsOF/aKiQOoSiDbsnqyh3QapPxaexoKtIgSKasfARb/D1kbprzl36G0Mx+Og
c5i9QGEgRaJHQpoijf/JE+amm5y8+hMO/Ga96h9donMzncFAKT+0/O0j2Aa8fqWYF4g2mu6MNedK
4wCPgwz48wVY3+/vIRxeyU8f3rhVkoebwiiSCdiDjqNRsLVa5lcvNiMtGx6JA7asw+kOfT6Ol0iv
A7UttsYIXbuRQ66ZXm3l20Qc7BR2m6aLAI7PHMU5i+hdbKihixj0q9ft4S4qROj94YnntRnLq2Pe
qZv3gD/HigCSnn26okwY7oqanZejI6VcsrM79ls4DU4aKvsGhcWJGpf0B5lxpRPBN67+f+oChDVW
AKperRK2I7YB/d8JOzKTyP+00CyvawlV37Vdtd95jt7jmLzfzb2M7qjxiaFEvIo0Y+akaqipDHNo
0R5yM4C8Kn2GNuR+H+rNDV2j2mDUqxnZ2XAGhzj5OopqjJqCscme2BdBNVbgJTUJi0wJNFU4B9RQ
bydwPVunmcjvqAVykgNahJNX6HT7pK0EDaywrFhn3HKPuN62F++SZK3rUaRpqoXIUK6LDOpZmfoM
4NyXxcIJi+51s6pSz3sr6aaACwEC97lujX3cWFkxgXOD9RgA8+2wiHv/1PWbkr7zQQlH7zEwD5mI
c1Bzra7F2rusQ7F6MaZ9z9D6lzydBugy6f9PQIbPlNfdf987pg09eal1J6KkMwd2eqdYkV04f1AB
b64uCqujFlyIJdyF5i/2ASPgM8rLy5uXIWyN7OYowV/0slFhuGfKKQiz/ZREQxd/377JA2gx2koM
+5sUWY3hMIUzD2mNQEdPW6OoCq5H0KjAG4D8DN/DjpvbmsfcHj9a6+y5B26uxt/6PKhiETaUPtk5
MyOU5BSOWFRN9DVHew0gqeDJ9y9PXJe+lKI5TvSUuA5BxzAh2Vp6IegrFDglIJY4lSyrVBfJG47q
fox+GvLw+zyZQ2Yxt4cbRAIuMM/47F4GLkGO6CQwBtInwju5eWz2cgD5Kmh2uZWAwM1dVNsi+5s6
h+YIfHpV3+m0BqKZancltWtpInSFxpif/81de3YgIJDSLis7ipWHKeTng+/r9YGaDyjSQtpmgJrA
cxMQr6kspXtfCRNaZpLBuwpVL2Wqr+/wTKuLtiqhSzmOfhzKVPTfrzrL45SF0ja7mO9exmieBtdK
UiPlfUItJnZzXjnQSZu/hifT//jj2ZNk8OHY43n2Q4bGIxGNiQSjbmaeqJb0OgRPC1scjLCGuCrc
12QMZrUD5i6sjDddUKKUpGlteY8ypfNvwx8+XJ2PSayW9OpO0ss3TiDDwDWAxwKtgXcSXhewh1j2
WNpJvfbBPtCa4mFswUius19KMYJ1YP7ksvdB9ef4XfG29/QXNcvgzIv3LVr09GhR9dZew6nQPshf
fUpGcXzmeCKabmnx76DA/VkBl90ySUtyJzZEy/drLR9oS5UNeFMsQSkWHj+klCmd0pWP2SMbVj7I
bAj/uN+bHH0hA4giMfn4gyjaaKK+AOFeZXz1myTKSCe5raoEABG4Mnm4v2uIN3+3bhIA/liWKt0G
CAAFQ+f39Z3IVUof409mka7bdIFYqtCt5skd2NtXACZ8LKLhygQXShnadJUN+XxomQfVGm3Ooibf
gKBWXt7awpFHoAxZzc2YJ+T4IfZeekRTewGV5LrCDLRWMswQVtu3xUOd+oF/Qnb4ssNAGEkN3TC1
+o1Q/eXRIClPULxRHyPWBg1sXbx4DIpczhhM3996DqmxYoodATvlbWQE6lIr+UhvrOAuKHPO+OqV
0t2jjraDODY/RxCEPjUQXfsWSdpHDCvvGWwMuhISqe3fLTmNV/YhbmWCbOQjegX0Ku4TmOEM4mbs
DXdbCG7dsZUMURtFl03ILlJDAE/wjuGvo57lVvvLHB6nFdBuVUW79SEdnk1CuhQu6nJp2Ji4xPah
ihWLkO8JZRcJmmfWgJ2VuMJZW2S8hbLXif9zPp6fLmFfJsMp2OBANvZQMPjhXbhdByLUFTjq0dkl
Sp5sEzUm2o/ScBCA1xQSelPY8sXV4px9ajMHzcNbyKPVq54zcAXUZPfRA4rAoeA5oBOuBfzwY1w8
8AM/WzyJmpIjZQu9aWOeeXkUnqoEu+B+sQTST7a/8DQTvLQk2l5a7oblJV1NYslCM9iSb1Lk4Ntc
jteGlC2vYxeqhu/Hw7SAwo1LiukfYBgXQHoXkF6re6rhRQudpOW5zQGx9yb9pl9KInenfGuqgCKI
e9snH2invF2z0390WfY1sA2ABy/juLsmtTB2T4yGRN95QLL7j5Cy03BYh5PxyBxnPrxRklyMqnU5
y9mXu527PFJ1iZTjlplMgLCL7WXUCKVXankBu3AjqLvToL64TijEhLuLrSY7ZWX82EA4uFY4Hz2X
kBOkSZIw2V6vNHgFByo7xuUzlX+2bn2v7UkmjlwdzVoV6pWP86ik8jNpc1dlf/Jb/kz9ZpuV6Wlw
wvS7BW+s+PpxcVWZjPKXIKXx4kfsLiFU/RsWOrkH9T1lr0daFL5r4X/ke68uXDZc7jvT0QkC+vyK
vXKQbKC3j8P2KvHetFMwW4nosJkzRJpNXldQ2NRhf63z7e44RAZk2bePKu25m2ChQpNLMkfRTZ1h
WV9+QqThHeKNMpa1NjGc7smlV/onMmMupIQbDmVEaI4/GpPuRW4nRtiY75lVsGwZ5GFo8D+qslLt
DRxiFrsVa1V44JxLiGgegwI7jc0EzPFVrk9FlBJhNj4myZGtr376r0j6lZLxNe48CLB/qoSmKqU6
CgelVGxmSNLo1yQCUpKNpXsYxJZv2BQE++y3b0VL+xT/8BAJ6hnnm0WV9qcJBMqZwSiZlVVJiTtV
7Kbtlk6Iriz2o6x+jxhTp6VR/WzFmQnBx8V3vN85/nlS5knetUnQZtWpBEPw9Gq2LgT1qgvQwjw+
F90yPSdlPlGmOfZHMuhktkUeoV57x9OmAqVdE+rQv5rIhYDlyA7hvw6Kx5KtaVTpHaYgrdz73hsr
Gyv5k3/niQFPwu5w4TVDacC3rLWiUqb086W4Jl72t0SpZ3TX92vR8stswq9LWrOeXvp+UfBo59tt
CwNJ4HYKk90E0dHxhHeQzIkXDh/C+K3cbOMz6cBoAYVimtQukQ9+0Y1TK/WmsgZKbFadBrWmIbGX
qPFL0x9qY+1E+7rf1vVf797IK7mQ3FdzmvuXD5elP6bRIz/L4yOTiYaS8k+5h8e+s0RGm45CFDOE
7gpbTkrYv7Bm/KDoNyECFBlZq4U4Fom8aEjGfNRBzmUGDp9t2Faz8mYBZgIt7Xj2qBNwzCRQwx+2
orn05gcFT0HkIZsCg5bg7PUMLnmTu81XPgMKXkaq4LpsHVo+TxkWUzxutGtSGTZfG3Cg2ZAISNXH
5zlDuJVDBCvfd5a2w1UV4zbTyn+3qaG/LM8S0c7H1LPH5pzEpRjKdzIQ+xKY/rciU0Aqxe9dv13t
MFO3dMSe+uomU36AovAZ7rm/QFPitcL4wWy59IdLb6wvuzfwWLdbUgJuzzFMR5ldBcT8fo3zHfAL
qNy+CGDSbCTxaI5zBYQ7MKCa7MSqbzY5Cvh8UlvtbFY4jSL+/lLprRRBo29CJlB9IoY5vM9YK3nN
LyzwpoQ4++eAN5Xga6eIMyll8e+E12PsMw3+8GpCVDtW3CM66v35Hm5cT3ZFpLa9yLdkZCXEHeM4
svwpdMf3a8mkfDzgfFPOTt420jyz6FZvlJGA9kTba3CsB+bccPjXsIsbgAqGZdZFbaQhT+VjDF6Y
BVfe+KWhYDTbqdGop+WLgNDdBn9zWG6jmp+ZyWkfRL0O7g2Q+f4PyUyeqP7B/DR1mgxR8TuL/oTZ
Ic7Ek6VDsQskIo4YdZtZrs2IIrC/rBdKW4eIy/4tvu1BLy2gsXpaev3m4gkcEd3QkbfLKIwRI6uO
qjlxexF0Xiikq5DItkXo4Iptn2dwjiQ8G3tAix1dyoObHPW7NMAfn3gd1SBssBHIpBfMVWA9TGwQ
Wo38qqhubAWdrMLFZN2d5vNwpLqVSnAEWwy/F5YtSH3msH8H2xJvklUiIYG5prJwa78cwdWsb3X9
JlZEWU5R1Ndckwu3PpYRMGb63ubiBu0SC2g1VUuma/WRCiIN8T0UojdyoUnUfDlKe1W+osFIsPET
XTz8/eC4r2kQ2C0JPOZ9mxSWTYQKZxyreKrUs15XbxdmJ6L7UUxiswVtuiDXNrCGIF1DRWn9FOLF
WyZ5S75o9+Q+miyb6b9vhnCHcH3YNzS5WFeKUaUlwL2QBpVoQqmT4rSQROiyMbPYchP3iRQpq3Bb
5lKCIKcxbuEevXAh0846Cg55v4fwbMnFrVhyag/7CiBAsT+NabQGk6pDTkwpZZ4yuuSDVWmwFMTk
X++tWkIRN6c0x8diBSafh13l1R0u7YtpLNLLsEvcxO2ZDsOHPxGgveghoXg8H62mviPPZrkEHCT3
yKbruKhu6BfOEwDwqSygB1hULfe8CwCV4gACWcpCavbBguWC+aFjLeCvxHbjFVdRK9V71uHolgAb
caFG9hk0x6AXUg9gAIH+FQdW/P1W/vHZHo4gNwJEg2lVZ4IurqeDVFDKJ/pA3TN/7+FDjbSgjjIx
hhqG08fjPPBujlikxYOnZ5cRI6zGlLiQnG705Fo5Cj06c7vERuNrGm8lNUiwrrME8/ob6FFhFBE1
uhlXNcJgjH9HWE/VLaCF7jWO8XesdZKRlX2IgtRT5vMKkxYOs9AVQVbuZQptelf6bzXP2PEskrx5
HRhgz+G1fi4PCVlekCx8k8aGE279wZgQXGiIa1TWQzg7GHH+3v0XFcTLxqP5b9I4+vURIgEs8hww
646u7FMpILhD1rbGu0jNzpdoZkUEi6j9yRMlWSw6c2p5Kaoe+ukG6UZmKckZuy4JkglqLWpT205S
SxuGe1z4UAJrW6rmSXk61LkKmkKFNM+jVIE6vlsp1FpPh1WISxHbPqmA+X+tvOBiyB5WMkh6iSA5
vtmxpLwgkoitM25QU4kXG5W6qonrkgQBZetdtmeZ6g9lVWDYO0g3UuolsczwulD37j6Ikav8rUNV
lMgmuD6y5bv0c205FGxrC8b8x+BDjtlJbJkw+gpzKJtgiZZi8gi1IodHHru7Ckpro0D8kJZCm04o
nkmIPbz9aMOIgOUzill//I5+mElBYDCm10Gdo8pACJreV1GLDoKfxlZlx02TYis03C8i5RkQfMRl
wXKB0XhXNnH1U9IabSz6GTe28fBOlHfNHWODpz44oSDcFmfcrLAnghkWvlQ7/LVpnzrdXFB7eK2U
D/X4PYZcwqJ/9YwzeozDVxaQtCQo75I2UeUCqu+jLmhFJrxEbr09lkeq644w95Fo6d/hIChzVW9b
yNP0Wravoblwsm1FZvihKH68waH8oUADa+R0OVvyEZPwm7Az8Ks6WB9rZAV/8d7dCX5fg4TGj35B
ZMY/EDFlwpvNzXJf5bnU9hSpDMvclpusKBiMo00J6j9pDyvck8trntq95yFrwAUvIWRKy+jaIgtq
6HGqRDgW55aUA8DOzIOPIdfQ7qnZlGSXnM4Wg7dYQk8rRYMLfkpREaePZyxCkAriWCOu+MLhRmP2
Sc/u1cNOn5ypKgCz0/erAYpCjlsct9lx+MJ6UrTexM6h5QLX0ofi2W7OQsQRNWh/S/aN/pH89uu0
gFZpy52MMrN0fdqlSwTFJlczARsD7QoXV6cfqiKNad7Z4Wka5tAOQKkolB+qVlGKtlhWH4Qq1ORx
OF+g4j/dhQHdPH+Z6iYG7T6O56twCpuefKySauvEXrX1G+/UfZjf8D4vSdlU7qehLksKaUUQjfeu
q6pRyPBtDMWYVze2Sx3xsiiikMzGUu53gqP8l5gnUcaZJvJWEwaIRtHhqe4BhcMYZu/IZZKIwpHs
SLO4mTuE54p8H3sCfDxynN4khcR047xZowpewlTXpfzFfum3R7E5G3LNyhg9w6VZDDtzxMODkX60
GfvRWzBuOozS1+KLZK995xyh9TOA+AFelNgAS+WnGsbbicLquxhilie82tARr1UWlrimwJ4JK7Sc
a6Sho2+qrDFKDj/JlmjwoKHTSl3vu6twvCIccIzu7gVASCoSEPeOrjbqOIxRG0CvSx/DXs4eK98m
CBf8iikMmDi8+REJWdIBxGT/rOsmvdPglVKdAKKvLdOfDWwfRGwAqWeEoP7tEHoYQz439weWJI9E
On2M0+yVUjPSRGoUHg+bvFB8dmYFvj+qsD7/jvMwhxHM4HYwiQnjPJvUp2giY3IFRZryYQhb6GOv
k2GVuUOJx8T3Z5dcCATve4TH7LRFgtBbg//mouzCGi/+gyGHGI/c8qtgdcEhBYCqXsuXocrGU5j5
kjRt9TQBAsFTBXt77Cme90z3SHrdENjbrQ6vFlX5Pv0z+Ncd0lDs6QTJc/mAxdR58wum5VO6f1gg
9QH+P6JJ52iGWQ7TFVe5pN7M7jmOduDR7G2YHPdSO1bZgpo+ekcqR2kgRf/wRqzKuDwQFpIU3t3f
NHWWYFgFwQrVxr6F6cby7R6KvoGLZwlY/iPQMYXYrSVCG8fqRzerj+JVX9/CugmgTG6TlSGUzwKi
g8zq2NwvIvsZhWZBjbE4B+FqCqEFm2BoMeK9spodlPeg7dnXJQdARVuY33FIgV8uONzs/DptTMWo
hfoGIyz9wxgfuQWQU84B+0uv0QsSiatbK/4tRqE55cNV1qPFVCyTLC3JTDkgevmYMsoPgeC3IbE2
lXPAnJDjPnsblqNTwVtVJHFbVWquWp1V8zpru1BS4sgItIdf7lg7FJjXUWx1XOlSpmHpGcOMTxwF
aOB1eZ2a1cMGRRjaeC7uXp/Ty/LYE6ReyzN9bt1VQdSUkL3Q9WFgQeg+wzaWQbpgqAKOe8lmUY+p
hZC8GxN9TtScwBiGqaQD5++zR66/kSu+LCG+wBLaa2j98uRCuA9VR3srRYbGAcVNGKPJkHqd9eu/
d20c+CiapNtN9wI9A1LQe7mYS1ZRGim6fIxw5oGbkPwCK5Cg0OJAQenKqJHy/Js1bKcCXPp3Pw7T
9EiQ5NEh0DIAoQf6heB02tx0H5g2PE0sVOZ7oNflz8xYRNnm8sPfXuntUfchu+KuggEiiMoKQOIJ
LKpbZj9hQJ06OzA0c65834Cmz0ZsudB3oObjgQUMtuNKraHx0F3/hnwp+YpBuxpgk/OvWoifOnRF
/2j5xxQsefvnGpvFySIJ5v04YWA2/EdUwvRsfn/S4Wm/lhus2v2FIqrC+D3M8862NWXmnhrv7LsK
kD7+VJD3uXINy8hQKOYk6MhvR+FdeOAbg7th6TB5MqgGJJormxDHFbfwxsaq7ucSlmZiEYI6Su3P
AirPUxPp9gfCnZkoLo8uKx+SqdDzCx1/nu7oBSiZZ4xpzy3EHgKwiaib9Oe0rjY+BUFR+yGGhS1N
eYJHS0VoeceNUelHB01gVR9w7c9lWtM2oY5jRP8+MSmLzeQmmrdQlZ5cpWutZYc7k6kTzc5ky3sX
cndklB9k3XR/XT0lxclqMxbXF7saNMrgD+eXX3QMUxHvSbEIzoc0Qe+vexox/c9g2WAzyuyEPeTI
8BFSZZCHAnumzYJpa1LfgJHr0mY0/9pIcYX8/HdLcXnAtyJ8kY7YQ0+ujJ+Ylm/5CrJihu/SauYl
q2/Y6IE0iKz1Ro5mYxE+Kb9nYnFT2yMw7GxD50t19JKRl2O8WPgGy6xHPv5BwL+hHn5RupwjX9X5
tjV6LMs+/FpCbDe8dDPiwwaDWebj+PNjTpU7Z+RZa46VSBXd/uoV6pcGOfBNs9+ud/Nj6WBEcIwq
E1Cpqiou6J6ev1LAKw2DsPjdKNLV2wM+nMpijZLW4rKUua6mgpPMcJJPqzujW+KhHuzBlUyh5PQJ
W1FzTmcu1KZXyEvuo/Px1bI/SWzOeCyte6vmDOvH6pghs0HzJ1tWYbP+Pm/XiNhILwfUzCrk3MV9
9PSKTDTWllaccaFoGqb7uzrl2K3VbXthW/AuDO5lackjrqopE1rFmcMsuX2eTS26qvm+j8x0emHk
1GpxJK33YFzme6PRx+GjwaGuvh1KM/zs6ctgPQbLTg0TBJE2Iu8Wj+pfgXGB9mqoHJ2Mdy6HjA7w
/g7Bl5IsvQrVldbbH4jFIUucVINOpnN651JPaMj6jUvK9VShoPti/JOiG/RTATy1AEqB0h/YyUV0
lcIfqoO24/zdCOVvsvrs/EXhofT2PsqNJLaSE4GglEg4CiM+iNqOywaqMxa7grS2d7qN4IDktSQ0
8KBgSOJWOerjj5aiUJAmYi8055ocRPcCIVZUrbjXQ3ttd3BJRwLo6jFgpLa77EcfuFXv/uVLGPSA
eb1bWv7yvvfxni3jHR9W4e0RAuXrjEcd2sqbh/U7/4acgdMvVBYrb2QxAqdnzdHHgH2DRRoMV7v1
EZEoFBjAJEGHDro5wo/tqw9jkvi/zDS+ihT4UNTTjmF/fRYRIz1bn2ufKZqGqOyrvGfxkUkmdONB
Cu7GA99gw6HWcCBzP3ZuU93OlLYpI9evJG4FDpHzQ0JDQ6iOVTS4ZQNWjfXofN0wYctTPMgi7nMI
1AgyL9ppQmdqdjWAidxU0SYpI9x9GW98OPwhP+9qXwfxwTlRiitV3KUzH5h3IPBRXAiGIYtaJJFY
rDbpXLL4Wy5vpFkNQePouldFdRcnXSp1o3jw+bNltLIXQ0gOAwcSt5XkYIQJQjcxwW3ZlViNERxz
ytdm7CmssH/wuG3oTtpY92nIa/0+FOs+BKLEEuiE1JATqlrxRKSQBb+N14j7L41nklGc+mkOiniI
HtZ9fJvADXlDFFh3eytip8Du2PlUCFHhbd5HzFtVFLH6Tklba90p6H8gHTSewNhd/gaPx9fJHzJt
OBaKHypu1rNAWqH8Yrqx2no3YWPDYj37QVAocbejGBBhdVgNfdaBsNDUKHPw6KywQbOKZ5Wm+BEY
Pav34dKPZSD9hWFlw7EAgwDHUOik819PNM+YyE3Y4dtaRp+IDZbudcBDlZ/iO1bS9ioI1XH6w2wF
hkgf/+PQ0GoRdwaBm4oUXYxH+RzMWsR7dlIbxu5ZV7nq4VfU8vMXRSqV5f2T87ElH46zwiKMdxO2
z4LK3fj+Dv2zynFUmq789K9DjPi7yQSGs1zoPCZGpIj/VaiEYx3Mk93m5wcgEAMPqL6BrM0asUHR
iRw5ygDyihHDwU3dj9n1U3nXdRrqQSgAr6ap0ar2NRwIFwhUiAmjzVvrqS4HV8k9NcwqPpfPUkpl
9caFffsgNBUrCfKWtToUTBdbvqUje9ncduYVcVBltLdivpfCpkTq/4maw4Zf6T+XmucyfrweLv6J
+ldbuCVSzNdWt+6rZRGAjfgCoZF+JrWaq43mbsM9JIPh2PYhUmw9D4x++JtaOj8FTQithWo6+5kh
HUHIvNPsT99SHJkd8Cdn1obvCrc+8sFb1Smmdyq8xCQ+QQXjdGDGshR5DbTuLxBUqDZXKntzRmLR
41uSj6/wXUcGsb2MW0moFMBaZMJmqnpxyrMuVIUHt0HYVmhsOxw8dOj+xijBq9Thd9aRIR90LVwZ
Rd9qZkPF67cpsk+U0QeihvTnrJ6MGk+eBGOPawsvyFm9mQf5Q3v+Ivi6EDEigty/jnC14Jz0mx3z
diB96ntEH6u8miDcL3RdKVOGfBRgveKaQTaAcTmXsDXQ6Ejw1iQIxdC2sAIuc/d1vczELPnBT9y3
8/qd1C+UvkqhFzNn8P8IO8ZmbIPpjFo4k7TFiXDPi3cjC7OmD9v1PI9FIWVmoQmQpTzl5DBjDvrG
WJg3mOihW5VgrhjO2sAsPxnQTULTQDu/7E+eZTN/Pi2EPwEAph0ZOlGL0c4mz0io/icsBl5Bekab
iGVTM/iwZbUPRqd3ck5CAVq/7/U3NoRSfyhmueihBi3N7alrgCqCU/IoJfycKeMkUkRqjjPZHXwO
16YJ/7PTfh1P82e0x/j1EG61jnqRrZZYGEzS/DH3jfOTwpjb6SiaNIIKTkVj1nejl6/E2y96ubK+
4eAmHCVWaI/ddI1EyzIVEzYSLjsOeSOYpvrjb4Zmiazuf6DoBOkPmTw95eVnD7gZbjinYlC7rKHf
n35Bkhl3CEhSEv2fUjTcPVPmN6vA9kEA8LTlH5CRw3e3HLOMP9hREkXJdHXO50fJ2hdHPknrurgf
9abhbtUXkLN8HpNMxgzxupP1FlSwF0pjwAubF9EsmyvnElojLqb0WzVR1S+XtmPCwcun72SMqrBo
R4bPFwIYcffnAV/rVl6SqZKiX/f2KmpnnRlmwrAlnz8DqBPCou4AcDwPhhzTerkAWo41L+jI0P7h
9PprDc7pjBNSo9TcJfJdaFnfa2X7Ui/FzU7Nt+gwPy8OsmUYX0OyFk1K+gAQ6zdozaoYd5p0npEP
SVUKSMOUU939L/dsPRjkocG9yGxcAC2IHXzPOAyQMus/HEumzhCzQKdFMkIG0u0Jsr9ZzQj950Ph
OTjSaH3QSZuzeCSRHSRWTEEG3zP9rgLK8/MBxsMW0lmjmRcj5lMED2G84+tbGCuPqv23rP3oNolU
AdY5bCDcxY3+FwvzckdFrqWcEghZdWcAfnwrk6tHi9a5+Ov4/iZ1HCAd4OvKqAfm/yWWZ6uvNE6Y
GeJ0zBD5i1aG8sBOwIzMQiKpp063buSffyo+Uy/TT5rEcM6Hn1MTNVPooIAxi4YQKzTNDd7Uy9SA
+N9FTwBy3CJggu9DPxe/EQ+98m4lePXOVEY3Q4OSROcI3p9CniW68Ad7W8kVLJzdAxXXr4uuaxte
IOC4fzRjfnje/MfkYrOVfFoYR3kjNhVxOe9wy/JgkAqYcJck7BHktK34VuSAwBnl0Xw8dfBGB3G9
fYTjXwcPL2dMeBzE9kH3pxCegu4fTm4XblFnPPYvgShSm17ULUGsefbqo8fFQJEICfmPKDcPalAu
PKzdLSifYFkRyaDfTn6wNieWXjLw7xyXT4F3QF6691jN5CmKucvfRP5R9sZKceH0gmJG5pTs7AH1
lvHrprpiQJQGE4+dnSbL43MTiBjZNVl27LcmNAPTM/W0LVQuCumB09GiyAoZWYKdv10c7l/JRcx2
6IlqegxYJh/f1GNLVLy7DAmWOSk0Yu46HGko5x5hUEBkHwoN18ViSOpuJfxxXxWHvE/JPMCxEk8x
sBp4oIHmBMX1Fy9eHwwl+72Q9uFVjm7nqr9OW6hbZ+bldXlUijCQo+utxKqxu3S7wedCA5oxgb0c
QQiyIsph9ewPlXi0HKRwlmyohLMAjUVsHtMmltDNdzMTswCBmiiDXi8xQc2uGiAB859Sr+QJvIzE
zsuB0iMjJm4PNDaMsrMZbwXr1Ilaek7ThELqZ1WGEBjY9bYkThZJVOh3sHU/IyTq2kcj+ePgYwG5
9Yl6uf7Dv3f99/oDc/39LUMARzxAYf0qDJL7yMq1vqmgHKIfQ0eS0W1gm9p0afSikw6lycsAEJKt
ziMDJ+a41Ax6NWoIbtA0MUwGi2I9s3HNeJv3aBOZaU8FCxR9dmHllgxykEwM2M8rDQ6U9gnRRHol
I9TAO/WOcRYdA4iaHbN3VTfn0By8gl3LwPtaVawAEK08ZUdwPuT3K/8VA+nH56BMJHCocuYUoRTU
8E6isfTFnuUgfs+UvMId4vw199K9q5nZRqvMMasQI7vsWjWXvN8oQHPGpRuxXwPAFux5ku3hr47A
Am9CzMemC+vIAx1J5m6OaHr2Pc38mZ6i47G40lSObRop1LpJ+ciha4OniFaRY9vX79R+4DvzBfmW
pnt6pZjKP1My/723r/1+IemwrWhk1huc7AD97si4athSzqX3oWaXHOIrnkgvGJ6YKP1LM7ewyb/g
G2/EG8frCusQ/PjInnfsb1OhBCcUkRb2xpOYmGHQL1fysC/6Iv8YIqEP5oTPp9vBA/OQGbDsJldE
C14hPgxZhssT+tDQy52jAW7hvoWpCTSLBtT7jwNih2drqCYp0yKZEvZqLXKPTwmpaOjavj5KNkTe
MW/o9mbmZiW8m+G80T1ubvs6J/WBAieBMdxguu8JozEafAb17Wk0i6Qkj2i1E8dMAy6YQsr2h3x0
RiTBlbaE2++4LsDMYM0c9ljKdfzZgxunOzkwHFxi5LMtgEBtmgVfXk2aM5mKaGQ0ZAHetd/9MYqF
2vRW/XOrOcNnT61FBPIFfx/alSsU/uJSh3Xws6zNuGtobM8fjzXblFsq+XEGfYfYWoAMC6aQbtwz
j2vm2O3mqbagfkdVaTqpH5h4D7RIOzUkSMzdNBaiBAyeQNsBYIbekF+rrPnCv0FoXf8Dwoxb3cYu
bQ07VuJy4d6MHxwwmjjMP0uR1o1IvIkEkHCKR+7U1KBAw1FoiVArea0phoPsRpP8LuPu8LyndzI0
+6+YMDgN15Z7jLBAOxXN0ZT9CG8r51zi5uXYSk48Z6yfyhOYQINYmq+TOosbJE3I4aXF+sdxwO3y
/fJekqr0CVOxRStgGAYe85dLqUrM6afBcx3n6i/kLxsIuKnaIpkJpOkVVPzKr6aXPwEfBOQFRq6x
BdLn7tDYHHBetVQbI86vn4OCaSBtZEQAuJopcNebaxXlfiEW8evd5Z8UhUWTWsud3RraIF41F360
hbPenpTCi78STQXmAmOTbM53H2qQ7hOzOMyx3By/R/NZOGLaL6i2PwEWyVVILkq/pzeJ2IGQz/wp
jrwgVK1/ubc/6Fy3UYfOEReAmyj/iImLktWtaGhpEssJbN8Jr2zuzmGPY0x0xNpGgSImDDtfaSXD
6b2ls5mQS9FUuB+TYqAKm8Lyql+2CXBSQa5hoB2NiEK0gbyXYZpzIaSYY9GyP4fPPpMH+npHpUSo
je2eveqaRbp33mxZbTpjZV+4fiX4Rohi8podU1jy58Bv/4DprXg8JMlqsb4mBhx4MLluhC8SIqn+
108Mdj7A17UFbwtyl8yZRZb5ttJLD8WnkhuRnqbzJ6B41jahlXxZBuM0I2Y1a30kTGerG0xpRzNP
FgJD9ZJNmsWEPy79ln7hJd3T2tVBzVwPA5fMfdXAXsL06BMQ/jiAOXLI6QUg9HgXzR8ab20PzWNK
LSvlqT941Ghmmqs2v2rCVP/9M8IdWwdIr+DGWw/oWVM6pBxq4HuEYOSB4rWyXxr3yPjLPhs9jorp
mTLewuLbAU+qVFkW/vMHeGJyC+ir7czfV8lwVC3AD9XwCODQJNMqhu6N8CYlEkTg6wU6A38gUbVt
Rl//8zjpIQJFcyivgAnkPz/mC/trT6YCO+OCWz+EyU8RRxknM/EQoBPEx/YoGYVShZanUD5MPL9H
xYurpJ4ysa+5vKjakrJRDP5Nvv+iBK/Czj2rWLm57M/JGXG+s5nRpNS2YEFbWiaGJIY1R2RYga7d
j1KUnKyEAMtHBlAYpXiVOShx37oUIdKyHgOS1D/nRgr3HiE1zdoO0XuPOhBxP7IkWjtnnG4s3YEI
5QgAfmty5RUfJki0dyIlrrcnRwsGRBGsaUmLMTqyaMm97j4gQDP/6WQDlOfwevsL6MT4yJaHPqEX
MXiqp9K+VUsMqV7zoFqS3/jFvtsF+BfxtZhVV1f2YOoT+62umwODZsuGme/Zqdw4NRdvSTdq2888
1BuV4F91I9Y8Q/UR5vvASO6En0fghLxTjCCvAGIAITxR2AsJhU8i1IKrISBknrSVpHi2ytxbvu7h
OvvfcN8dtXH//0eGJXB/9O50UEIOLjaSyt+d6ZCgOMUItmUfzX7A/0BD4/aMgZ3iMuqlufjf2eeZ
x8iXy/WaKGRfcpKhBVtlJ7tRnMPiwFx1psO/WBVBM2igedKBl7SWX82/mgszcJyuZpoIPOOhF5ZE
vsVbZPCfDPasUhagMcxzneo6ERACyyE/WWwco2imiOFHah8laemTKgpBsQf1JTM/68gINRnd702J
7Qw6wFDipNMkS/DHlThFVjvGIsPMRsZBa8FrQ6Q2w1lfMqahq/E/T4CN2hdSJ+U59sNucj2U8dUj
ozHSUmhCx/KZoID9dpraRWhtXZEXxIDr64QWHf+sI06j7o3gV+rVXEXdgMBZwWrBFlNR1S9dQSmS
7bhL8LAgMPod8CF5z6x0DVQG98nH2xtFSj0L6Cb4Bxls+eViMDHBHC6WR0tsFRXlr1IafDkunanO
MStsyNqbAyZa8vBgOfwAX32FK0pgZKJTt8mylwFLOLtIKG88BiLXQMoWc95jGnY6LO8EiebO9N8z
nCiqrlEbaCowC4LJ/ciibzsogQk5iKzqAmWZ8IPlb7XqL8qpgFgvt+TYytgXVElXNyBoMVxIF2Sk
CMAezsgrQHlX5OY0JqHO/SLh7RT9p87fIiF2KeF/ldPjBfyUzhQulYfSJXPDbXf3mnnYtQnDw7OB
f2Fhvg+c7Sn05GFBt+M6sB66IZjI3KITQFFO0juPPAAvi9mGVab9B1tM7g0df7G9jVr7t7sUS2FP
47nAOPbBowkkGUlaRWL0r1q+8IX/KlBV7MzLfz8JrJyWJLXxPAQtTSSgRZdwiwNZS3MLn09PZx5F
wQ4cw7XEa66k/buVkNkutp+0Fa89iMI7udcRc19xWXxn0Ezf8rDwineOM7D5QU8YoHifwGTGcQbT
TS94RyuuOT7Nxbiwtv12jwDtjRG2FZaOUmcmUSzpfoVAIJrhyZUUpyUJrYWx+f3Inna3Hjn1Bmc7
X3gmdvwTJBvEYWuebwLKNyzOpIRcpkI9WuHAw2jK4LbsyZ2i1ggwx/q6hxNKNJxEcIb9teX9KoBH
Nx04uiBVR1eLFSSU+p6BwRXQnypWlHbm1sFjrnf1mW3/nU8eHGkA1uqbted1lJUH1ddayadb1BVy
2PfPNDC8wXo4fZeeaIkwnv1I7ePIzrQ+qjhWBZczuDhUTdWVltFG6yRGj6mr5Zy5InKY8Skn9Hxo
9EwR0Ah0oiD97FtsSyFEvd8qoXpaSUYRmy3S8J+fQ0VktnUX4VH1xPBFDhfaBiZVB6L4hapNaOBX
PQuMoqC6gVaUZ3DCMHci6eAXxAzczOp1jQzYFnuO8mTOCrji31Kn/ySYNJz/5b5z1LeUWQMqQ12M
80N25yU0y6RoG7Tq0BXq7LljquKSLgp1JY0iz3QdE4XHbVI2e/b5X6HL7b3wFF8e6HwdkMRlzvAR
W3rloz9TVD6Cu1EQEpJcAt7wDwatS0zseIXTDadJFktEfUsv25phtax1i0g36Ar+Dp9nIpB/oXpY
/vda8JfD5nTCrBt00ZWPXuGpTQ9ViRgNPHY7uAJDg7aQ2ZT3L56h0xnHdlHjuKVMjO+4qfPP9G+S
a5HKd6MNp91oc1UhDlYVnjdqLNialVuEohH6Y7LhEizajgbZ851LuCzRjHSuB2p9cc4rGsH2qKB1
TplQm/h5Uk6Oqyh6mvBUH20rs00jzLI/aYjCn0I0hbDPhhn0d0alFgC/P0PTtG7Gkjp5qArTeXC+
sPoHTXZPEAB28dUgYcmVFKk2Rw5kmyUwzbbH2OXuXnkZ7LcmbX426wwAg/LKVxMkHaBvg7a/yr64
0pV9mJw4cVvK6tp/sHBkHJCIKpG3vkn7QeazBAp9VIwjFDaFDbpk54Fn5DXGkO57j/Zuz7E9d2zP
up1776780eQjMIdfsxojI3131/ZuSqgUrGmHbeSHXLeC5RbB0Jz/T0d+B/G/MhrnZ5ALFrC7wDAh
gILyjDFpOF0/YJ7DpYTSfm8kteHDlJkdNcKAPTrPmEqUmxKpyEMZ02wldI1rgkbs+8LdZz8QYspy
o3MVruzEu9Nz9so8kNqPPRTCan+dHY3+4EjdX1K4ruJSct30Vll9EvuJ8b7gasvShNK2Tf04AXsR
Qiml01QDTFXEqPrc/mdRWfXDz7FFylvx0TyFoKZmB0+Pmuln/7Y6QSwPGIKKQtOJWpDhflLyrHky
AuLAjqNUsVTCQMnN0waAHZjnAGXccPx7cRWnjb/E0PuYw5dUuVFrmtNxM4QDVnrV2BWdFqws5lub
TstL7DGDI+25NWqAH/OG9JjkBsGJiBLq3qYDT+5+0OIobW4veddaz4gYL1rZUjjI1IU4gIM71d+V
N/6wLroen/AyXreYonQdzay7SenJoS3njXb+33PL9ZAAf39NEc4qtHR0jsxc6dg2x+9XUYA4pEJ8
01WTDcUvhoLSrYqc/LflMW4Kg4Ml7BRt1qSpnsP04KBkBVkXSonwqr1Q+tX3rRQr0iL3LCKEm2ue
i9s8RHEIuBXEaZNUVpS3XWI6S9kQri5vqGKKvij/CocVFiBqfshc3+Pw0JXtHv+ZQqZKUid1yg4X
0PwXSXqfdkzmgjHm3L6LNqiPqv24l5rYnTlWeBcRtfwkxRZwk7s6XfGUhaWghXryNHeTsqJ50uIu
HYKvC+ZJZi1o+9C+l5N4lUX3M0wjOT2SccwQpkgb6I7awFkcxHoRFcDuIUDeeC1SGR3alrl4ij0m
hYW7fymiR/ZlYBn9r0966zqc7oCNcHBvyqnWrvff+N1aMYh+NqkFQ6iQQarCmNU7gZDGlLIcHzX7
aYgaaY1mZr52+raJM4Jho2rV1l7yzdI/nG/jd0bSSNzgbTud8kv8R08/xSmrJav6pJpAxO/KB7L2
ubMBRb8PfZYSc6p2iG6FT4/B8UAb1gkxKSTLL+cyGoS8yalqmkjc8CXj+F5XsalmjbByjNoRAxe6
QwqNWf7hpKf4QNnmt+XU8mzZzNqjOLAe8En9hqNqFA4ozz0CR5n13tkvFPAhCuYG72rC7SGPi8/k
LO08Rk6yK/TDmjjwUfcpEGl0kzXuNEGFNmN4UWHtZIZyidR8pihM+xHHy+Rwu8miauvE1lwJF8Tv
c7mowSsV2QIAm84LHECZPWkC3eSdZq+NFim+rfAXcWUMJNlbJ7LJ2TW9MLQCvN62qW2cxYRsEGzV
e7OcpUVhybD45aB5qhFJIHEKJC4j8K7rASflcVy/zG5KLzWaqnjfRzGXYcL7x5ywAskJLQDhBRZm
pYCpQMx33W7pYP1pHA/1mY51kWR+QZ/hAPa9r/ZKd8/OC9YNhrGZcRhtnzfu8OVBpEPoiU9DRfMa
adNnYgzl/JOEDzADfR8KnnzQejjnGTf/MoxEnaOuyfGbEdPLBDH+tpdsOC0Nx7yGpIahZP0wSHCv
21n8GMq+B0bVe5UAAYMdmVBCcvS1qYVViY8sfZCAWvYIU/DUMUrVovdGdL/lm8iC4KTR8S88u7v7
xkJCKm2CpqLGcTJfWMqtaDbCygWj/ypz4WCdvXvxSargKDNQGqwSx65JXt7DlwVxx86JuDtpAG5k
pzn22Hf98pyo0aj0l5u2jzHnoSAyVJpv8MScSlxb6dgX8GPthaCm5DS4wXEpTXNzmDJN/geMWA4D
4OpFjFE338BjiTkMCkz4j9AAr+X/zeegtDlJWaan1mopi2MtksPOMnv/omak4uVYvuoiwldTPCUQ
OjAZe4HeK/W8e0kky//8XntWzQccwNTf+nolXXVqZVQfM4sTdMHcvGhzqInosMzrgAo5RDCQtHhe
hgxb/NSQAmQ0yhCI0/tx9AuYWLcz6jQfFOa6FDvCNK/3bMAsFSCplXgLBaCJtF7u3bv0ZqBTogmj
LFMkUWWUiPQS5ALbMJ6bigzcBuT3cJ0nL59KvkA/lnZSLzloAhwD6s7St+Om2tkdF3nIJlSmFE//
E29bmbecxfR3wvor4KOQoP0OSABLjkVzF5mBhTCCFNaAMNMWGy6kfLteKxo5221DOb93Gely3dcz
1JD5ymP51X81/XwLrSV4KfKc5AboNI3OqjFJEkKHo8e7Ts4+4gR8xOUnHDf17RQDoSBmmFh+I0BV
GHRFshlS6wVn0Ny/ov78U5BDwjl7SvhRMep8tXl26DZ9T135dVc66GKOcFyoHuAbYxxRMwKdqsTP
ehYC+DsVXXlTsy67LpBknYBmBRJYfThGbW9abH65A+gLHhbV7UcNqNhZUf1PuLjS1JHZpzi4lNB7
it5BtGIzauNLFb0B0cJO3yHYvD1Vw/JKADzFSdr8OherV9mWoo6eyHD0giExhfJqPVzgjZQN8ErC
qMSWGYFWzEotz/b1zMcRaVxw6K74usZoM/jq2xc1C/yVfCZvFaDPPnBXiDFT0mDI+RZ1SN1DOBrk
susqoYhJRCGaHJj2ZpeIhIgmwUr35HKxXQGdYkdGJ/jmEVQnIZ1YGQvYHuseuAEdJuseBVpNt9FO
8hk2vREGIO+liFaLasKBpj5lRH/sNwJKaGf7n91DYuNVsgFbgQRglkr5h41KSwOQ+dh1cDOpZLpO
cN8EApFGTmbluLI1pvvvGhwH0sUL20L/JiS40n9P7O9dbCvkMlKL5fAVJCB7jBOQ6FaPHlVU/5CH
fz2hkWI/uhiOx7qbt3lZHj/L1unKhZt0WEtj5SjjtonBBW3PdCShgCS0Kut0HCJ5z8KWBPwpRSWE
m69vgJ2/LkHyVv2PA4jV0nQNvOsJoTo6UE4f1BQM0sTzj04oFx9MjwOKnQQW8Em471Z3lJchheGd
RSiN/wxmWZj35uMdg3ifjkGOGJTuKhD6Z6HuD2/M/Vp2iHQVU7tT+Zd8l5Owb6/ULSBfAVINxp/l
8BIDlqhlDRG0zYaeVwBxo4sHE4/7LiIsSp7yiLarBY/jkCbyBHmWz+w5mRfBiI+q3LnpmvQ6eShX
3XsiH2C5xogdOB9vCAUHMttx5y0xs1VLlBTIYNGDx8CrpWqy2Q9/IiI2N7LXoUcA7Jw2oKZKxfYS
cFZwjrOwAqiNvyyWOJSYqLSsN+qisASYFfSaLVzCFL+RnaOui3P5OMwoQdRFx3XUt24jdMlAuM8Z
XX4/lV5zDJzFHIsZK0urhZv+UOOe8EchkTAruUi3QTYq+ziAnyuHpg3FoJlm2M2YNfzDVdbyRCNf
Lymo6khlTzFe/tMYM5CXZCU9j+G7SPR7izYy1pSW53Ra83OoJYXyAyaP0Cr3/oPI3ee4In6UuPYb
jETP9Hz0yG5RKFrZD9BIa/+n1viFp9/ABf6hm50ce2Xs89U4quPqv7LC8/jrGEF+COboo0Dpivcy
jpp3aq4rHegsXSq7t5di4aRSMna+80jXoZWfWlIHdYFtAqSUr2ocV31VKZhj1GlkTuWHJF9pZ1iv
zfwJySuuoZlJmCjZOB5WXdcPmR3yb8OSKrUmLMiv6dMMLXslPF72aup2pUTKQunIxBsuuGR02qbl
eDmZE8YiNAO7U9eBdd+gwswDfHXuJaEc9XaZ6MSuK7Uok1xpewab3FpPEXDuE6p/Zp1D7ojyW9LN
pRH0dMaxxBMKWOIc8KR2CtnTLexx+ibRFvnMETfWGw3GiChvTfkFHPGlJjZzxAWOYbRrIfxwzNSv
9nDfiFz0KFtWLiW579cidfSE87z69+DWD1hjYsn4yiIdwwUt0QNsAp/hu+jS+do+H6sESk8ATicb
YyWeh0HUDm/k+odzMaxUBVrfSoLKo6+VrOhutQAP3pFA3RJrnWLEOGuhzkpgUWmly8I4n5QI2r0T
9iYTgDIgpaFrmYzAkWWjRaJmx6Y/FxuCtqQ0kcmlorQQaCj10NxyIqUIgmIhRER+mAZTCCp2FSe+
SnKIgnAvjvzHDE5S0NyyA+9kuix0fWdGmo+puNYFm6SgApMWLKYBbA5Ek7ZtngbtmxA4PzkOIhxu
SC+ILfRTF0rh/29vBdK6J74gstCJTYiiM6G95oHcBjE9WYJv5r/N1S5hd+k9tDTDXr3lWIIyWDdT
3QLpJLpbAjAVFGho97mD6F0IRZVuzDnytuu1gKW7jtWTe1li5SjDhptjcsYh1tY6qBXslUYnwg5j
YIVGje4twggTr5Pa/13NwN2OGOwOEN3JN3YjQ3Sq46rz0OZFSfo28utRapza3JmT06uM50TsHuGg
RGT+kBS0RN8ROPdT5TToScUDdXuqLtHPY+3DM0wunJUlzdNf6JFFBksYQER9kmmuUEFSZT1mSfO0
QlwEUEcCl0c8YWgdlQEXQQdg/IrTCXy5iCURz5ep1aZDFpx6noiBmNt41029XfDSb8IY7T1wAn06
cSVKesMUF18b2z/1OWq/ndsQLp0WSBccZb8C+wSaGbnph5ft51/EPjeRrN/BUk88lZ1JT7iVaVLG
IqErIqoiXQz7oFgtpWmqUPZ6pCW+ZBXLov8Cf2ZnL2Ui6VxXG0P/VNNjIwooQDKXNP6rF1zCjbAP
/J4WgRRgG1T7QHM7d647BMmyGgknIG+TcFsdjmjtZCtgVpmD+eDVCEDMPSkIAjV9PFbExazkDXu6
BXSjWak62qTxIU7+xnlmw+zOr8fTkc2cydQRplz6wFBK67aTMDht/PFUCBKlVUBAYvFJJgaMalvM
fEL8ZaHU2jzmz+KACAOY0Q48JWujLR/Zg/vg2UCOhkncCQX1XpTpuJPjLA+NTQ0Eb2qtItGAh7co
Qox7kXB7mtiR4Uy5QQwJFwp1XCpdCzIGUFgQgGtaPQgu4MshQU5tRTFh0GJf9DSj7z3Nrxc37H2W
HPRK7n0bnkT252t1hnqfNXqD8kn1LaM4hwixZGBAYCOObVAjegFBA8dHAicC01/H292QyL7cVf0M
KNb9XXRW4zIutzeiiShLnIJmZ+4OuwQtd4bcjYizOBFYdHt30+FDd67c9xNge7J5M+n9N3yu5Xb1
fKNdjGBeEJPZrC7HX52NDPii6xyge0QTmZutNqRx4t7hRgKCLe1q84f3TOzDIkbbuGuFBni4PiDH
BhfwnKmURzX16XdL1O55jGzny6zEiWmhH74LZboeBj1CHs5aFWL/G80eRQDRgdTEHS6hmOeqOyIk
/pI7hpH/BF1TQZHuh2dU7FlFKWuML5AYmmtQdH8tfAm1X0QflzhsKYCKesgdDWLiCye0CfHiVNOd
LpHxA/GVY7nya93ncuHYHPjcQRwHteCB0cETGwp9lVsU9c3WdxAVCYPv7hsUtzpF6qIhI4Wuqllu
bow48nxrsMJ7mHe953XAnHOjKA0aEDS40gwtVz6iTGrGOPZmRm6wPEJVq5w5+Y3YCmAyxxlMxZPg
45XBkJ7pxApGxAzQyMkJlSPW7/zd1AmozMZ299hHx0Q0mKdh7Lamdb+pHTiEFd2uaqFtvCoT1j49
nwv3jDNv/wx8nB5lE+74T1HF7+DXR6tvzk/Sg9SCcWi6Wis6LjQwDLIMJ6PkXGGBPx8r9VGJLTBR
MDbU5JJI9zhrl6UdaaV+Xane53uoKwmbHUX/gDBzQPI3x0S8hIG21faeMQj96ZTBGEjAIvAJSEdf
wHw2MPhpefff/aO/8+I47YbaqLjkeHwzEybvfOpX6xg6NXR9kRuczllLKqriTZ5SOYOcPJ81F561
WRjBoJQJLh8dQ682avBIDShWAoOL4/eTMxFB3KwI5fT/1qbd9+8YJTj5JYNq535FbEBY/947ru/l
QX5my8+gS04EzCOodmwOjR2aF/Krv21hFYlwuZYCvr0wltumwdwBFn5KmsLrru7xJPMWj8LBM4/s
+wU6tpS6/NW/+hEaTYLur7VwqggUW8pziFMX7E7UH0RKyWy+6hEIYlsnYTFKu+11hPcKokDUcAUM
RfbFUoYa93+L0Ney03OB/w0aea6FcmhJEDLL9z7Z1ugLjYqna4N2WUo+9SmDsjiUV7Fmad4+YmOZ
C5lIRGssrRGxCbHz/v2gqjnW8P6qRa3pAWk/PSKnyNuL+siArN1PqxhAd+XvyghDkLEw8rCqRm3Y
lfoUc7F8BcE8g+EZD5NIizv/lwkiD9wwa3tezqHHMewfrtYDxHOQPZ3nKvQquKESMU974gz7XHGL
IQtHDVPcK0c5ReCMLGNF+wclmVWHQ4JEYO5cIz0Z6dTbttUgXDJoYrayJ+DspOwH847W2qbgYvAb
by0Z1DTNTC+CxEMM+MJd8R6QeGO2hQywyXvjFY0xmfJWovQBTLVJ8Gw5DgzH4EtTjBEGOBB0GpAR
d9fYGb/kKKOtDFhlMhrH7waI5wvjI0rKSd/74yGTsS1P0L3Txqms4ablYWIfDd1IVVmbCzrw8h1y
g0Qzo/NMBJ76xQt/WaoS9Rul8WezvoHTaFKLZMYsfShQk47PJtVBFJQnViyyL7X//eq4L2AIE0qW
y7PQ5KNxQXUg/2UotOH+XO9iPe42/zhO6fxdNd5lH0OdoEJ7qy44Kq9LLuV2H5FLaHzNz2rhrziM
vAKoU8m2w/WqTBruuIkLjuSX8jofxq3njKxUTIXW30P9/LrIx2CFZCnTX0z/0MZZgPeJi2tJjeT6
6IfxZCtcCAGDdnnP/IgN101IftSs99gkoYN1ZnRZNfe25PjB0zlSXriopdrL3iQGzLXSESp8ZZQD
6Xie1rGQjAglDuZsIk4xhnHTpVkHWHEDH/T+UYC7V7WFgEdmE2xGbz+2iYZ7eNwYcW98+8DVdJoH
dk2PXA/6RmxLg1h3e5IyYUSd6BInilpYR0p8W5qLJp2JZrm8ECzuQQV5BvH5p3NIkJxEvboxdp03
ELsSYElJg1sWAxjfj367VTtD89sRRuGqk53La/aGwRP6LOZfhVeFMvNp1eiPl02ZQ/ihSQMXjyTS
bG/FZqH5LJfaVD3Qbum1tDuk9CWK1aqMLZVDE/b3Z89YcJ3d0Z4X8lInlEUCzgHIoEPIeMcfTqCZ
AKyVQUCWdMQt42UcNM1myucHqY7KGBIXWX9mPtBP8vGjVp7Z4GHeRfzKARUoTA1GeydIYLBc64bQ
VKLT4pv+704UPccBzZroYXBRNIBzXMu7HJT3221z7CDfJQNyreIOLf9cBHz7UHdLRZl75N5GUBy3
kjVegeoTa/fg7oZ4fOmHBm6Dqn+yf7U6W63b/7ewVR63RgSzPNbE3i65W2Mo0h9v0qYQCjOt9OND
kzTQ+CmARsvrpMaEoVdzB14lckFvkXxViv00uM/yWqPFzGPYgdeBTYp54erCz4c8ppVVDTuduEn1
DddeMbEN8oq0rtuT+tDuWyXP4ayHFjrHzbmLFrtjqZKeu1oPmGBa0TECE2xPReKU8jDJvF37iAXP
pj90jLc9U5+DdtCJAOb59aRqmFDWDvx/BL2qZtEMfAgor0vlE9Y2r1XmW01XyE3uuQQM5H7OvF2m
rdiLrXfpV6d+bkdOqE3F5E9g35HoRI6n+Rk3abT5F4kfKKR6Viu0KfYNE0GO4yILUGBqFyjaNXfN
3u7s8IROHFmKcSmfaTIzDRXPXnyNLDYT8uAg+kmQ16bVH8u4AiRqdDHSZidbe2iEHOBkdgTIg3xd
NIoV4gCKFXQao1E+BwWDAdsimFkc7Q7SDYtW2WTIxyvzalAPqk9pgmFku5Mw3QHAanBD8MrrXRYT
ISELO5L/60UjGsWZSuJeI4wTjpBcWRWNJmTjGHlLGmxyHhcjiUn4MhetYy9VQEb5OXP9YZefImPR
ZDhrV3bjB9K4lQUrgPtT77rPtJqNp+r0m+EQcs2l9kHPFNoIn/rGxaHYgN8oJBIW9YvSs6cRjmmo
lVdGlD0VOLZtZi1jK1VYzSq2f1cFRtzsST8raXmkQTxTjlkTJWOQG6Rq0O/+AYc/e5b4HUWDQe0w
it+/glj+jxj98pc7xnOv0Q4aJcGsXOuF6fb7qu09MoLdm43/shv8rsvN/Bz5D3spSWpqVOwKycaA
bvB3EAwvHSjFzSN01zya2yGQaAs7OBDcACVmji9JkykeNinbxI3cy5UwXVJlWV9KaSpPh35GETBX
6MVNktaseoK4SmWrdX8JdIQmvnVQ4hT4rg91C0UYVcYVW5K6ON8boqXIVuzmOGuLQYvOpYXbPOek
1J7ggP2U3nHbyQdmSUac3c0VTkv2jT+xad0y2dhiTqc6/70kTdPkS/a3Bn2fhrZ+4GHo2QUPPZz+
w/KpZRlgDYmu8eF6oOwNfoWvMlmM6NgvHyDQ4FQh3rIneRgx091n6F0HwKADW0ymhLny1rbXSlGO
L/TbVwZU0XS4ZWvM519dZoyzKe4UKlQuGr14mgrEk34DEH0iEto47myRzveydHbaC7EAIgUHwxUR
0XBgFeRropsvbowZuJ9E8oOifKGMs22iKxMFu9zU6bf2ujtoUtLoFzNm7ve1WvW7SiXf+0mwUWu9
aAbGP15k8RPtI6PFOWAHFFImLnOxFQgS2VInXJ+jYJ7xUVNqSkj9kYdSAuI0YECfnChgTxOg0mok
f4AtvMQ9bJh/7bXL4LDnsU//YJRaK5RoCyIK5IUK2eHikItREfSI1yV3hwEbfjtr/Cx1kLQbzk2Z
WDWp+3CACrWEL4ynDiyD8M2s32/lMkC1CuyZCMs8EvkI/veXt+XlWNCPsOW65rOfzBsgSGfhAGRa
8xtZXhxyd+azgZCgOkvrotamyLP8DCVmQE+Oe0zqQmQvoE+zBgKSu4WlDx6JResjMUWcYxlqh5u2
uGjMjyTzXVFt+qZwshvHdZcPd0fVNdUEvkbB5ksncJ6mc7pXqURft2IwchHavUSHqtN63svv+PJq
D0p7YskwRm2uLBY/PyLhnbavHSFVbB2Hk299kUwJgrbIuWzSw7YoQP++1QlNZvpdxbWf1wdF4CNF
3TJ9pyc/Jr96/9xnXJT15gvNhfqybBBQx+32ZiZlhPSI1zdkraJI3Pip82Y9B4nrgRAzsefFnOXP
TnfAGJJpaJFOuti1kYXxoBub71uYAoTj09tonrsAf2EPChoMl3dn6wiv9sTemOZeJScYW+4IYXrU
qcDX3azmV2piBv/UfuVPSoPU443UX+FF0w9JqKK/ybFMao48D0s19S6j9dG0vHTKdAnDOizNNFQb
0WtFdG24slCNbjV8AjmfJMxD+GnPB6B5tFJ5oRxa4xRIZVz5Gd5NKWweUiyrNv3Fi230dh/3f94R
sJ3pXi3XRrk2DN5vsOOEXijCL7Nqve+/23B+vCnzRrT92DbRWRAlqsppTKlSvNcbwmhIO6/LznmW
xMGSW6AphfrPcX1z8awxOFnEJ5mlIR6ONLKNd9KQyEDB4ezw7rZVsnOSEl6R/dBeA/MpZcH3/tY9
39QCcXjr7vncVV5csFmXRx/GPsg6w2LRRcfUCrI2GCH+bTav7KtG+gj1rC/R0u7k/vc9qiHHOG/W
T2f1WPcX5o2A76BbO49IkI8Zp0EEXvlvVfTHKieBRb8tUQVv280EGeDBhuKWN9b4UA4S/Wj8LU9n
Q1MSl2Zq+BrE5nnFcm4ZkANrLU7sgJVj357QOzf+LdOa6OI6ZG3X8rVhKQCk/xlANbDmortuxVMs
p7sO1+ftPP8KimCydWh+pd8P/XYVGFeGYOI1ed3sXBKmMNeEWGBGPnCBBwtNAK++1kgQhRnScjyu
shz9rmIf4D9IR1eu+vdkYX3ZVyuh2w1bU4/ELtTfmyrnFVqwz8YXTqsUVrUAWEIDThPixjgVqLwz
S67acg8Qb8dqJrDvYd4/YkL9Bx0RoyXORm6LoObtdGghl805TH9QbKhvTm18H+ivLR+dm/Z2UznJ
zVK1ZeB7A6Vabl/B9qKBzIHraTV+4DdQNAzAK4TOkGWXfKUTAwCKTRE/MM70H0YE3d8JdkHckIwQ
FRJQD72e0UNsUmP0dCFRHrLS3aecSuMM3oGaq/lphzXI1m8ixjgit6u6FSqZ4C7u17YbQpU9cxxC
KruYGnvJYu/DCot7rO+qOlfJoocRDZbY/6XD8S1+ZeDxhgXuKBuYhSNVb7vZ5PoDxYmiepgzUuRt
E+0IZgHvMMSsMFNKnrt0UUykvtTPsG4nntgW8ZMDmZ2ed0e1HcpCJ+AbQmEsW3VbaemK26cDh2v+
mzV7TBNXU2i8v9hIIKY7qn1dqphBQV7UycGts49Yg55N5OtxLG/zHh9psv+3kstErfkslk6e6zeG
oiEq7jdPY7XeGutgTmczH9llRInWkKg0nIoUb2N5F6/XUtvKoG8hn1FVSc6oazwd649qFwXZX0vZ
W2zeE6N0D/OOiSy+FL7c+V4I2BEosgHKNxcqYNIHhF8IM0d2rhU3dHhPpNI0TfKJ1cruguZtomz6
qxS4o86BP+gqCULpSZiup5IKRVn6tKaHNwl64ZwzzGN8y65kSjGXOmGyUYvgTsgdt18DOZEFnfS7
nUW9abLOAPWGfcFqiiV8eDIsAh3xMIdvpftPHLYTV/vO0byuiLJxVobjpkUKnVJkZnkKmgBycjBp
UguE908wb9UAVmNVMsUN1TnjLaTDf3ihk3fJr42x89jklXKo5xaqlrUdzOcNk0xrsc+CoTWbLiD3
25sizfqSX3y9qm0XbvNx35qwzVINHHosHo3+f6asMZwJrX1p/5nV1+mYist0jugeDFgg1Hw6QC4L
k+uY67Ba1rZIDmF7h8i0KDgiPQJq4jfbauGxtk2lYeCNPMBNQJLhBZOmymthiM4k2dBPI77wyf7S
SVjh/sdCRJm9s52QL0gyyzytA82/MJt/CfPDdOy8gcHCaqXpEx94kF3rALpTVK31t+k4YdOHhWaj
ukBsKqlIjAM0CnU5lvcRDXzgELV3UWD54nf/6rEbwhKTHEXcjkw/GR+QGyHMqnvNhcMxwUevb4fH
mJQnDMVk+x8gsElYgOVsyTRJGua53SDkykJUiLmKZALA3pM4rUL+QBp4sli1Ql7kaHyLY25I16Xp
YITUvSrkT5jT3U0+vzmAXAUPcobMGTs6tIJvDDZzkhCjWn9ScFujia1eyw4MXVX4qzW3wBFvyBo2
Fxv6JRhzDSxbsaAc1BXWhHjYqZVfqBocBykxGNBEfVGPTqUP72TGwjUWgJDVU9lzNxtgAFJt3YVl
6H464ygVEXKmQT9aFW2oMQN0n74omSHBwHe7l7Sgpa4v8dbFXt1q8RTZyasyyTQrB4P46ESIap5+
TfRHil6+QdbtpuwROzR1kbxOHAwCe/+OcHX2xQLNqceB3tVodRxKFxJZciih2Xv0l0S2j1sHpj6+
06W1iv3n9rj8ZAL0M8J+EpQtEIsJ4y4+0XCBksgBncXyYqZrvcjUGqy3Vy6un3E7tjUpNEc6Gy4w
p6BiIh6Vr1izl1VoV9X9QFJ7v77KRG62e+0hRoQABvXjcUF1SlvyTpniQr086Msdrbh/hRxVPxJt
pSu1qvu6ua0Nfd226pPfuRujhn1R8thliEv+obMvxCbt8TtZ8QvInY1dgk0x4cKG0ZhkDiZPr+Hx
uRsXimvvMrfYdv6X0a51/FkW6CgTqGIYLJYF77h0rQNuOVb2/S9HbEPI9nezoWaMkS9EH9K/RG+7
QqCACe+kBELZ2p7y2iYfkKpCdpKeRlZwnrVm695Rc9djq28t8nSY/RFjqK+BT1qoU65vRLg7LsWO
txAxt+QqaLtk/OzTZraup48s1EfUPbfWt0nYFc89WjxeUXvhIF5SDZSBHSA24YZjDCWN9o7HThDi
PGThsdWbKA50yK+ElDKtmu0Fvpbolds+cudMIMdcKB2Wuq8BVFZVYEbMV51Rsqcy45w8d5AR2ZY3
Y4r9YJBUk4NXunt5zbux1jdtJw5dgzg1DpIClT22WqGaw0VHKwvedH2CMQc0tpgj8GaoMRVFAi6p
4QWxLB/bk/uvH9+C/su0lYBR/dFBwrSOj+RE82kxzAkXgR+YhrniWAYa0dKvM0sf9jhOZzKX6txs
sd2Q63jCoY6DEva2MILxXq7oGH7fvamnCVkOSexv/8lORl94pcLgem/sRjoHjGduNtSM/s46YzQR
XB/t7IyQhRuzSOfgnt9VP5KPeLsKvYe2DT1UBEBeARNV3K1iSU9xuHY0Bi55lS7jR2nyzhAIaBrD
SRfDWOPV4HgD+M6J1xbWU6ffvGC0l7Ozgd+BdSHfiY+tIFRBBAkf8dmRZY9iNEvHnpexAmlkwtWk
7WyJ0qsdvlHt8tRtxsYmw+VMHLC1KaBLL9dJJFchJcFrOwiUDHln3ddJAYV966C3TouTSrubpEGr
ZrS+Ebsjkk/cha8IbdKKVZMP+y0hVQQoReSusWoQSjdJ/bZWf/ogCPy/Zrmtv1rYrNj2R6kEO4vt
syb6lLh93VGxWAcOOfqgKu0m1Hhb4mivnjuLMyZq9oFbAMkcpvmRfCqHeIdOWHhaVzNkc/2HZA43
HLEVwdPH9jZ3fvKJEADg3SXFoSHoMVLGAdnAwrmXQHEE8fb++A8JCsaAQhSlV3bOapYfG6aiDK4q
X314PugthbeKRildbs2qs+J8oySzInbI1iE2pZEJe6mNWJe1WkiDCFyJXseBbCr8YHv42djYeJL5
LJAID6fKEyc2uEtgr4MPvPbt4/JUOw7BuTgD3BmNcVcFfGrHKfoptSUd/2h+ZEpmjv1kAIlNxBEK
LBe25lZZVdfXfgHL2onMGfkwMu1HwtK8aEJvlBqPWddvvTklJjnOFM3wUxBhhjQ/TUxHgusySAUG
qBSWsUJXcSYZiQ8Mz+uFlryeHGhUFHGgF22wm9Xnc2cMnEORTrqJ6CgpHH56HKBOZgxBlNpSyJdW
2zrKvqGb3sbYahCAc9l8FsprB5UuEVrUb1dQAPjF7YLdZZ4kl6pvPIwQu1JrbY4Ik8rDGQaBkfFv
FgrH0OP+dM6oGRcZOqYbcCLZQ7jCiJMdN8VhA2+2VtSIz+rLq+gWWW8g1LN8dXkqy/+SA3+pC3Lq
WfaV/H8u3/RhTjBnMWntuGDbbB0+6zrHWfFETzk1hR1rad3dByiePGci+gRi+af4L2Yk8yecRD3w
kH//xZbGXEM8aRtnR4wAF1tiCZRcqNg8TG2Vjtu2TCHEucewXvhAb6bo2HKgPVqTHMC6GEM3ckmt
NAsTp7xyQCVE0zGIflb/d7URztc4utrGtHXKnsoUrc15k3Rg4jowQ78A/v7z1PygQV1JSwbCqVUP
MaDQPs1q9Zh8GChrrBcRd1n5je1vlKqNxfdx6iAJHctZG/Rvl23K67jhNWookrMCqcXeuBn6lRU5
TYSXluOyQcbs9vT/LcG7pzuLHJSKaeYU3v7peBrhsa+/8uXTHNBnuMCgAL6FxQoWEDsqorhNx9Iu
Goo56kYgpUKmFjHdAKoRbJ4kzlZNYGkWGGhkHwWjhOxPP+JfJeOLPq/h+Z//f6zM3lRuIKHiknC8
EaysFoFHP0wHmEUiGqx9IIFl5F+iJJu17NVaN2OFIYp1WQM6GPSHj+C3RkzNNyMypDCKjoFVREvP
TL7fDslGh2e8S2FXNDTK3Ym5x26bEHPL68W6jN787aO3wQTls132+H2n31IMhDziy+6YCWxle8Kl
RO4zlP1BcNxmmbZvPR/cvHUlYkA4u4QABI0lqldl/vPw/BZ24gdz/cllo/vBRlPTp5m9IiRt6SEa
YV0S68InzvvhWJBBCddPnrCMAv62woc2tzwFTe4ffUPvXTUy55fG5h0H9AyU6lamImyOF4kESVs7
LgS5wwqP3XeJoSfMuzb9G/NX0n/gq0h2xV+3rRRlJ5TTMMNIC/Q/tFi3kzOKElnN4qhfb0yrS+Hj
1NC9XtxMyEP1ttuuuefvzEsmy6k8A9cKpVCh1/xlGlbbweDNpOar2sjXw+U3oPK2/pnB/kKofiQ+
e+AzM7akNM3WKhuiP/tb1nlhx/lOmfU8r/d3ISBGeqdmcmPVNgYfva4WheDBxt1ptDNdCHYpMH7i
pWx7U97LO8+vJht/OoIqMFgO8TQX4i+++0JM9LkWZsbaDEGyQFyRPBOLZgoHudxFk2DJM6R96eNm
0EoM+JUiDXH70m97ADKljUZMIMTK6JEbxFtp5bymzE/2fGMvvLeZ5lmxqqPTIkuHhC3gQ8LmT6AX
fbgIjyGvmJpd9m6FNFrTlNa3z8S8/ySKBlVVDulkicuEQqaODVe8mUkeHa1c0NtW62BojLEMMr3h
V9gBhbnca7RNLSNx6LWjedvrXqGNGdIK2tV817yKFGPjzWYxlUhdcBERFblvIBfHj+sBkbdOYq9Z
7DeyPQTOLlfocPR54jyz2eF9h9HMqv6mkizjnToMXTmellG4DtPEZysO03uaqGWHYl/y7B57Sopb
mqS8p7glWLmc3oDjlmQ9x8hAY59A1ggGnQOew3Bpi5Zo10y1o6k85wvOhhoN0DYCQHjt13ms+oDU
k7PgQSLmCt2bb9D/8CQVZhMlnmqBh71qBCEZWNPSeM69YJGe3Jppn8Hf6wSLOxHzcbbHkHXVcNtx
NG6+uxgPUu1110mEsYNTU9oaIAFyTzasTqWhaXlVygLjyhVEjXuqbd0PAbsqSFwHvKEybxMoA8aH
HkC+X6uPsd+YFwFlqcwXXfraHmK8PJVfVLvKpubIEM+AG3QIk90Jcf8XZdpm7qVvnJdPMz+i+tfu
1cpFVJFCHKve5EG4VJMJNLD3w+CiUgGpl4NSyjLJyDymv41OcCRMuIr0dDMz5XVoph7TV0YSxZrI
4YlBQf2nkTjHGIp28MFicwYahY49RZTo0e8jcL+L4QAlSqPux2ALY1iqASjhlCqm5xE/SFl2EGAw
abx1rTrEfrfwTJEQ9MQTKX2StA6t95ohJo3QoJi05P3DJOS80cMpByoXBL6RmfYYSCxvLQiniePm
zkfQgk4VK+/z/YqUS92v39myWYIpCEZWF9D1WMStcM0UMd/K3+lN9YWiMqQdmpjaeyiFEF/8XwJ6
kS9RtC3HIdigzDwPt6v1wSqAuyPHpYFC5EwqfYG2QOLgLQZ4dwZf3XabmhlumZpUytK+LM/hzB0V
NNP2JIeCTj7hQR8fKEWsxpG14kXIepO95OFm6wfXIm15Dulh5gOyRkQNA4/e7p5BkdgyYWf4TJuD
kyxsFVzcbTdd7SPg3lzqUZGNXr7jALh4Ih18+SRUYVFy/BruVgDYu4JrDJiHCFCYJOEKqZA99bZF
9wFbuAa2b8L1spAw70UkwKQddm21Y54k/pfBYHJ+v/FPUub7EXRQgtX8oAsAj4mQY7uzy7SFwHCh
qVRWjWVXZoRWtJKZU9CNKRgdu9w6WRd9DJq2beWQOu6ugjUWcjFnLF0TikEjpE+/QLrp4mCS6FKp
BjVh5F9i0UyGxo1nyIuGenMwH6ZjaKR1YeRULB8qPxl6o3DLctLoUQUQIhM14U5w/Sik49NgJr/+
mpkVe2mdTjK4iT0pV1C4v2JnIi+xQ2mAYQG3Wm7zfj4dcGBd9hmydVhANcQT7BfBUwkicOjFbuon
69N1NGtg3sPSVjZ5UnjzoEzg5OZBV1irx0jDQQylyEWAA8w0etwVELHr4PTdw/ekge0B5zcxPYw/
Gyqi24ro5YOacPXMaphvz1uxxz/SgyoUFqT79R7IDFrA/cTQz5kUJnHu70MuS8v7n7BksNhqoMrD
vEf/11iGf/1D4oRV5PXBn6pxvtLdHSBnMkKChE8zY3Gc2QR9/5QoruDZsQwGECGORMT/n5Vk+Vo4
Thw+Jhmhn6R42TXJAIwvfYgShCtUafP2ngEsa8aqhdZgcA/UUVl+ogcXh6avOSbYeKJZzzgX0N9s
cbKdbQXjP93sz0MdnypJNlcVMQXMl71f1G3YscYcGx3RjUTEA9odWMqegE9hPBdCriAXUtXCEAW6
5SHgNoff8wXhg7SSzDw+i0q5m5f1nCbuL7aaxhj4hQe8rHZwsf6XxWtEhyFoaZroSVc98j8PcbIO
bSr3u8n6j1Wbhj7zzaOYEFI9LOptEoft+DHcTDNO8rrqg9uDtMml59Q64655tXxsXI7jAm5QdVyX
lzFdN1Vr5MnWi2uLo6SyxnsZhfVudFzyQlCWoWlwBg3NxxRARmyzz9sSUVM8mZwflI+nZQ+J9/wJ
RFsG19XtaWHZmOePpsE8ybUOSRhXXT1bVt2wN5dCbfy7b1nV+JQ5pjDi679EQKVIosrnKe4csL75
walDqJ9GLUkjtYfL5VqHU1ORT1oDjWDqHc1hVBQEYPFZ/d7xa/Z62r4JihdbAytqkWhgfs2yc/nA
w0rtaxmh1mQd6jZ5fc25F4+iHuPEs/3E2yS+CmzKB13yWvl/S8uvQE2erRl7M7NoXjAKbLuvxrmI
S7R5nT6O1qhMu/PVIWH8VftGxvHs8oIxRyKPtcBJw1kVn84NMS5A13yWjezSzDC2myAXB81v7Z3/
yXV7CBZJMY2308OiE67DoWzlXzUSQHTQ6a6RWkVtWYtRzS760EuW7LSO06UjlsKO/glb5CYC463t
MoFOBq+Yn8VQHD5/M3zG7C9tpeoouSfv7nHunwCUckEP+yYehoABS3Zrw3xVC9vBdV3G6yaUn+ku
3HoCShF+VsRzAZ3sCypLI9YRz7KktBUD038Kg6X1xN7+6vdQPBFSL0Ok5Pq+cXBWDck15MoebENk
9RhiSNToz0Ctlj3Nfp4ZhRez3SmZopgtp1sxa7UKFbdDwpyoIUpDgnqUfpFg1Gsui8r4+ax1PTaF
oILgP1/vlAfnEElQiLTMGqUJ1coZKZ86x0jEWaGYWAIFKPMsatuAT0/iZsfdxXN0dBztPpDesKcu
70BGyzXJmf+QNGwYOlGFiGrPvtRPjoeVvw1u0BG3HRYz0E5ywm915u+GwdPSW+q7lo527bKW/6yE
ckyd8E7pjr968tWHzKf3NJX2u0OJi2+TMxB5QN4EE4PTfofbJqVBW3PFXcBwAOntsIQ0q1AYVGgq
w5RGFY+RSbpH5QkM9czvDFzX4W41jJsAavC1YY0+CQnAANdBeNdWYD6gX9RBFbtK+cZSvkObJheB
Cd63e911mki5D9ZURXdZHdrdGVqu0J/3Ygx7EIeQYXfGXYbFIkAnfWeWuQXbA0vyHrKPb+77/9Qu
jfHZHQS3aOZ3RilBwKjGykvfDlDEs/XqTD7N1fy4KX2fjHFgw4dCasyARyTuj+xBVmoqYwj+LagZ
sBWQEhwCqmJ5lUrGOn8aZbxOUzDP0iN6N66SrCx0155BEsk48PaqB/dIK0OUfO9w10ZAjjCC6yMk
8deq6dF21e1Af0CD1o+yPz0XaIeviTSNQHmFG0QfHdSbJP/ygiHxkQFPBZ32ur0d5P0QWudX/Zts
qKLxEnpATuz79bMS0s9W2IP5dkIwsklL7LuAIy/zFYzDm5CQlyP/DfOlKtmZrYAy17Jx945bh7n0
VeHkj0/EZ389fdJNDB/B14dhzifs0YfP8EdvxiF4wyn09n2qIfclh5gUyfhW/LQvyZZxTMrB6xLr
Nef52kIKM5sX6Cf5n4p151Arp+BsYdCe+qPCQuauK2ini7MKDGGT8WLSXgQM+9SsYyekc6MkzSP7
UL7teS9huQWWLrWP6oY7NxNdOCh0EefYBvE161PqEvN0wrLNFXZ4yAcMnJGhpDA+kmAY0/nY3WSw
Yfoo7szxRLSLPwcVOaJBWC0jFNyBuk3mFcs+Bidl2B9FZpIkDyCgGa2MYUOlR7e895QTudlppt2w
iAhNSCSSx1lciVLDyuJqtDrpb6zVnFDg5H+wzUuJECA8/Mnuyqh7SElMz2Pp4Z8jdYgDN9W+5EOV
AKjL7li7ng5XyOi9STer4g+jhcATEIcLUOiGJOj1RJJweZ4DbF1ZMSpgAmpHl8X469IIpTy4wFEx
fc92ihi+JuTePpWvpw4yeo3IIqdibIqQqE42p5e5qnXibWSzhXMmtRqI8Uo/h1IRcKxM1NUWm1A7
1p/+56OCm6D267oY5hWK0GXih/249mdeSHrdO4EGutXewIYUd7Vk1hSBFs7tsXPgGhrNuf860NNQ
BxhzP9wFDZ0j2segw+XJmHE7Jy3lrbsQDL+yQsMRTyfSIqsFamUBrUN0cWts+07ksmefiGeRV+oL
7kzh0MF/75yefrpx35mtLdRKJrpMjnlrhLx71rcDMm8o4P0F1yJVHbOlC9LE1tZNZjDBFKWz1w5o
+cEICkkrrmxd13MPCsyObHTMw+rqMqoeS4JYwk86VqkSOaYSkoSQrKCTmcRXX35nfdV5sSXCa5RS
nbI1SAmkxLHxTWyjDufLGQTWOgezVTL/wQkcm9hThqB7soAmBH3zXZysZQIJvQ2A1I/BqVcAtuYM
x8LtgS14HOdhhtnNx41vigQHDuPsjOE3yCnC1DbkMZRM5lUjavjt/jeEjfMwGfXOoY13SiB0tk71
Xxsr5YE/agZ+kr6sU9TzPwS2fXqFWvpMFwgbc3MBexu1lR3bQdRWo0uzuoBW8WClZSJwyCaJKqP2
snVj8DZl8VdDXr839l9RrAFFpfTqlx+uNpxBDO6zvmlTJhrvPG5Pg79exG1quKcRpoNGSl6Inw+Z
TWj8GkmNXX4K3JE9YiNv94s8wmOvurxWFRDTCzhVvVB4DABwyN7lrAbS+Ch7hGK+fR8vqJNfFWha
Cerstjhorrz0ab73RwxDqDhpAYUK0Pc4EDd+b7uZha5LVd/F1nl1B5ozSZwO9C4wJEflh8aparJ+
Tnc2D/CLMhApE9cHf1r03vygYdVRFBs7LuwGBnZEmgHeoNCSqltWtULpWHie9dU9syakcBo5K3Bb
ieiLaYgRsBCmySlqIfEcBMZtyXTgeIEelYc/9AUly/trOcsIeTj28gw1RTzrMhBQ9QgeLUrK5eIT
S2aor3LFddh4JPXHyIM45kYCAp79lyODerZ6xokIf+i2hZ8akOHToUOXUsc9qkIVHCtnwaqM2qBk
L/GpXNNH15LYlkwvZ3dDZlXu7YZVUNrI9OfY8jWZ/Y19MnBEEeIggnkc9jhqChGH/Igj7IsDbCiq
9p8jLheVBuWdGN3V3qHopAvQu0bZ2QVmERtjWSjdr2f49MgmNv7eCd5ze8C0KaMQlSLq15CfVhpA
hfhcy4ZQRrk4+ts7hAsaZ05aN9l5+A92IcQB6Pn+Q4QT3hB89pAN+CMwuJnDP3oepwLmBxYZxn1D
FcuNyUB6ktciIU26IKk1bws3PeS1zf3B54ydT+vaTUg79HUQtH/qKyh2CphpVITMQp0W9w5mZnMJ
VkWW4VXMiTuXXEJ4bYjhi/PBTqtT7o+UPnC+/z2hwNrea4iThfpdetTvMSSsDaq73PD3eaKOJit4
mZArZ9ch3Le7toKy/RnOTtFixQvBJTEMfj4+xWLGDFjGR7oZGLod1xZH66YKNXn+4Z02nXqXlKyF
HFvsfeA3/e5uKPyWh2Vtk7yzIm6NZEdzkQMCxjUJ+7xhPRh1Ay7e1aFnTnV6AkY9yZxvRNwx3IwN
ky98Th7uzLDiwpwwTMV6Dmo01yXZxklvbYkV84xmgczrIbHLnjAjzywUFHkUM8Gj2HKLHKVX+Pt4
ahTniRRd1pgV/AOmZME97WMVuILhX09YyA5dCp7/0xseDQVm/YegkPg6hMa8rWSLkR42Gp2pexs2
FXceKMNU5ylElsz91lB98agjg9RIKxGIGkgBla25k2uLUE3516tAHlplWR8Z8RFkj7c6gx+cJlRS
/OvHP74GAH6RtwRPgKG3A9RNUv2AW69N3KVmcopAEiZDudFUQeQFFIJ2VIJKcDg6X5i3jv0Eut1i
CGJI9v7Q1RuxSiwDJbp7wx8Vv8MBCP8ZkcJOcKGXZPJ5wrV4flr3hoduXvGRqur93D7PejUNdqLc
EPZLBKO7j2dqH44kPQs5bEeTMq1PckUMxKA1mFxuok2uoIVLtkihi7+3fM/iMQs+AQK/W2tDIngr
2c6YJx40M0wugD8faDLKd0b1TH7fMuKyRPVv49ZwZ5/Xt9HCpJqraFZ4INda3RWxM46k7jndVvg9
qZH8iXNho4bKbMndbrJXXGG2sXoXnhHmZCZxP1hPrrNSKS6+q/0pM+yF39CNCe0fNiXSljy666ri
VFZ/8ZWilsdHQ2yv/z72Y6e+gcMQOgnVb9zE9HOFCxeXC/6z31DMiN0GJCYDHmqn+V6e02RLsQnO
6bBplxoFP79pqCoHPrkv64VtRNglbaGFdq09oumayNpEj00ULwcjf98iQQqx2YrDUX1Of30GDvkY
kENm8aR4zHoEkk6HjMmOGcv6JnO7YpqxSZdqaA/NWM9HaLMVeViAIZRNg8PSIDK7Qzd5ksTv2ho1
w1/x/migZkFV5p+scVbatlNwJT9AqpRLZLfwvxvj/AMQxovIpff+xNABHVG9RWBBYKpdaZAjOMtE
HXCuyAKcAcQpM+y6mBdyDRuNQJJr/sGVxLajGOVWmnfm2bsRRKJYTR1bcGFbSSwrO8xUFXqBhKtv
VM5G2vp34p6O7+HJJbH4QPagtn8mtkKi9zbrD4yqd6qBiM9Ka+dZo1Jc250t6Mpx1DVvK3Te4TOk
ne8iBmxQRhZ4PbgHwg0HzTXSZ6ykS8W/LHhk0kpnGCIcsCYAtJxrS+MzC9DvUddZd5hNzPUZ+x5r
SdUYONneefBNiciPqaMafX6ZkrMlmnd7IS7F2uurR2AotT5W9EunLkjsH0XuHG6ZzbcNJtZ/FPiz
zUG6WSjkhIMi5b9yVdoh84FQ1DYTlwXOJSoYbuzbMEhC+OWnAXg/8gMShz4Zgp0GB77Jxclj8VIR
Z77aL38fnzQ8+KMAJO3wzwASW7llwyFjOKtRzEV5RcZPAynDQ19awMbZ35aY9ye9i8kJlHfROgyr
MP7vmfwxSbrhbv55+cvtgINzeSL379ElADg2fCabV9FEmcqgdbHiR/WyQ1ipncI7BRFgbtpXmOrP
1/OyGKVkASQo5wxUvcvdn++pypxP3Qz9aIrEedO7bc/OFvgB3UDz2w5OJqzoPqvoGPwRlZGccs3g
pnig+0/Oa3SlYf9HM+5cVvgGsS3brPbQV9H8GObUoHvHexlqQyGC281JTd+/s3fYPdls5+bPs6Pa
Np5yzB1DobQVoNC+XNhBzdFCvf0961/u22ju/qH0ZgrCdtUs9ATqs55iiVIvIzTmJnrUJd8J7K/p
EeG6J3p+hOY/YNeMH8TU2RI0ndT1rbdEF5eabEe+XfGQ8tplfS/3XqJguW4NxRYaQHjBHy4gIR/c
PsK9eF004zSv8fOKYLNrJ5Hw4DgQ2okxwcKBCU835Ccrd/5y/fWlUWCPdzSEHtQGS41UL/69dxda
FRVfmFECZmAugEg+GWT9G8fkSt4aTFMdnvNg4wpMGSEbMDi+1a0DnNVjECaxhi+M5ghXsrn/nmjY
qQZARJUF7PyyOiGOt59LOGLAImYkzE/NWPL5IKDzHuTSpDzy5wC4lhoCR5i4VgkE0f/xDHiBjECr
MCkUS1duwacra3qqyBwW48MVK1R/TJeOdOyC9eIi5Q3y7FSQf8UuFXwHR14g/XoGUAt5JpzS7AR2
LgqzKzUpr0XM9XKZ/8HsN7t3idylh2E5jfh23PXWUCQeNLRJ9UqE/oK6amaJE6MDEZrM/MpwZMYZ
hlg84PJpG1WRuKzEoX/Azs17Ou9fc8x+Nu3OgyPbq1qrkOIr9X1auEpHzku07IjmDBjNZv5bbVoN
dfZWdfe8zLh7kHW542Pziy5WIXG+BzMTwc2wc3PWFsf8ZYJ8Bg4KikFZ4F18zANMOQFc7Y9yWZGU
nKoL9gALC90XILZCmbjKOKeq3bA2+AK1TyLT1Ygmr6PRro4u/DCb194GuNwNR4HYvRTEFOlyX/0D
wvVNPGC6zUltZD/jzGBW+cIhjaf6/zXSiYB+FKPn2UnR/topsbOhpfeZ79gfwrIs6kCe+gc/+X8E
Ev1+sUkYjmbRds4+6DrSq9z/8hduik5bkrG38EskU15qY37GjmLjSxy9lUhXnouo+gFXaq85IZzJ
ntDmRd0SRVH8NONv2Ng7qQNaNtGnOIgX3jpIVBRGMDx7dqV6bFSifoYNnBsH2YK+kS+2tkN45byU
fqhEICZOA/rMROFlgEzTNZeDSK9jya2FGgIKuBE3UuLRHZOtwROuc/ud4PTPcib6bGzT/+WEtOdh
y3uZs+DexBYjMPBLhUndhUnvbl5u7exZ5FvvSdVz7G9zdhrZG1RgknBM92TdE8FHPY4LMjlLhuG+
dSX3wjKqwfiMaEFBhQuDHZfg0q1ikg+QMwnPvI2do1gStDzh4AoY7UM60is88Y7G7OmUhcTh/xM3
VVkaF2CWCvn2FmH3LrIAWYmxB47yqC8FIV/Pxm466/0sAhYcuCPoNBk8WYv408Gtom9B+otVz0A3
v/bDe4QEjRTpuvLaf16C+XDWnLBW5ucQy8dY5YcaAlnv7Ltf6b0+mX6amNxjwg3OIgK26qYQxy+V
V503+WjTJFPccAAcz5ShPABNYTvUKXZ2BFgddsAqETNbbN68Yi75QFZoFNiAgy4LABnSCzMRF8p3
p6aeADLp5FFMm0a3cYU/zcFRpf4J5colILKgZNWTDeQsZHb96/VVYahgWkvP9ECz7x9VTLu9sl1/
FjMbN9V8xRv8wJX+2mwgKQ/Xkc/GrDjtiHtQ4CmVof9oLCBPsQ/47n0tDauad8+Y4rmKzpGDEHs/
cdn7kiQhWnk6IKs2skYLMFSy6/8ELqWJqM7NbNleHdfMDdAxmkicpY92BNjM9n8TAPaFI6xdx6ms
HxAA+JeiAJSDjFN5Ex8PocIOTsruVH6tAH8Nc12Wuh60WnymQU9bflpkXVrEzSoR4SKQxGN7E21X
+T7p04kumc2+XcmuPQc7S22yx6Vg58dvuJSRqKFQEQ5em10kj3j2z7dz9plC3Y+zZdRoumzKEeiI
SHBzsZ6Mclau+7ZqMHdaYxanDTtb87J2AdwBzo/iIcfq6stYHAgbd6YUSjV8dpOkKefV6YrDRbDW
moFcuU8S+e0cd2UNV9mSnC9BRwwuSgjnWBylx8qsK2Y9LuHg+KDqys4HvN6TXpJ/0KRPw+EE8QPO
F9qKfwzq3fjIYztAmZQfBVXd25VVjX3kytKGgwSgkcVKuJBJ4II3vWNXTcvutURpgYDEhl8B3fj5
9JXjm0pmppaw89dOAH76sd1HruGhfQ8LSi67ZPCWbjYSJEmCzwce8v/8DFX7v5M4eW4u/IDuP2Ig
XkKfPwk7fLNOeqBkcdPaIr9cAoDZLgoDf1E49lV1RloPNxud59lBIRpn787KnasI5i9x6gOZfR+1
hujkxsBctwgKzVl+smichxergJFy4KlNh5pIy0vD4MG0ECie9sqJKy98ehPi7O8vuDIRoL+lAOKq
1Q8IE5XIDxOVPSu9EKFsYz5shl8grN4OJcLvwN09QOPaJZcze1Y/0AOhEpAzwDtGMsLIW0hiPPpT
gu46R08ffHCJUJmlqtEuBuBa0vRNpyVUp8cH+VPbk6CzTlwK2Y3xr54lg76RXKjxBj0DTSFqjTg3
riVSF6ipkZmzuMCP058LxxoUa83urF4f6x7ncAFSPqDTY0eLNKzEjRwya8C2+1N+4MNfdrWNGy5j
oeh2U0tdgflpry/a3AcSs8/OljIPWllCIJfSGlPj3OG08dw6U/bOuSWNE/iym4zOXcOV3QO2BjgG
ckzdH2DBWnae4bae2erHPob3hZaDlEKJKXX1D1LzV7SgmvE9gLpJZQfhOu+Fh4OVBNy6rGwQQtVI
nXW/N0yfxKKjxmmI4g6WHA6lvWOZjurpeL2YPuMHxAJJ4d+4tPsNh0KvtCe/vmwZJpprbY1bWMcR
/oEswWEgLAj8Nq9Jlg21/gIt2RSDrmJ7ptlGRMFxxnxrOJ9mFvYHu3NPBqJZcWugOJhDEL/7Nts5
22SHSJGCpHRUc2Ttyl9bUp6xITLLhVmemopG4skT5aw62FhY5iR8KcVs8wKEsle7TbwgTHNoqjNJ
RICsw4VXKXXQ4jezj0l9szYFEqiGoQHrpKgs8Yy3/E6sd+iIRQUU/A6B3BYoOP+9Bg/xM4sf4ckn
F3UvKgecYufLheMaUG//jsBhFEzTrVTqL7QDuLY3vPxoEmJX96RIOcAaAHM9td+VT+lFHtPZ6WNO
vgzGZJl+4nrj0TfbpJUiUyVlWlA0hjYyJbS+dZrcT/MPmBPfeo3/UJT+xwSFs4B92OE5MbZwKbLD
aqo7UPzQP2aT/Dfu7qOIvkH6FuANFZX4Le2nb57JeSi//HX5WLhKMWcQU74FqGhbFYAnCYanXfNx
6G74PC8nuzLyWz/l5qKLaVIifLIjZ6180mj3CZhNb8wN45I9nWCa6NqMGxp9Zg6+SL3s22UfO7xJ
Mx2ci+mQzZH9KXF3dtWi4x1IRs8hLcggD0AAZggowJXTlXSRHyGwsRtaVfJGEf5G3QYDAxXyfLI6
00xcw+SwEWyL0mvajUrzpbdCvBc00qXNiKuqXv46Nqp779bo5xGtYItwlgtbsUzNSAW54adgtzmO
ApjPjoEsclbXm8lKgncVhO3/WKkbTRA5YorkUZEebiOtURUcL8wA4etFok73nID1GBRKBihLPqmH
1u+aL2dGlDLPzWtWk8FYqimfmWEdoqWZTZvEnW3ECpxlZKHxT0P/TT/iBm5clxpJ/RseKodKuc7u
tMo2FQO/T06ANmNtNgDzzc/YcLDikphPm08U7zFhFQ6B5jYFzKWPjcBe+JpBOC+4dSfw1b1LQNFn
tWwh1+P9m9+C574se8cex9fwKozDErjTShpUqWDid18dUbKHgec6Nn8eTzhg+AYsSNkxMuwTk2WT
NOFmGw95tgIm9jbJlWt3n0vwVo+BEWiM3mJx70a+MlL/TZbvyUtjU9E6PDtDIJWMFI9ya1o/mqf5
F+CucH6HtfHkTGckdRIdblrYK/6dW3JqUHVhz3BVhUxoGWfre4wjtyKWYRy5EJWseeijeecdG3P/
jO9X2E8IQT5U/4vRo1E7uMTbYN6D8o5BniPqnUAJU9zbJMaHvdRColkF0VFjHiRXW2/RmCrGSdah
R36koyL0jOBycoD+vq6vt7lnoo5uIFP6lKH8AYenh5SjoijT8S2pq7bKEz4V8x8lqLGNvpHr8we5
b0SyJps9XB+LPVbyzl7MdjRLVYXG98LRZ5HAHuqv8zvrcP+4qdmxEYKWMoQMrUFZF7rHazS1VmOR
sy7NQU9fETfdmGPfqnlZaZ/y7xvu5tklvNYYA0BJxzOkLhz5ZwQVwOyNfL0otxAZqWePNwjGY4zj
p+yQVeDsdE//Rjt9iSF51jsfvCo9WpAh3pOfVi0/OuTMW+64xw0BguUcikZ0y9adx8QPBXSOWjBH
aBSrlPXkXqQG6jrxchZ1yBMWFUtSGUqLAHtnC/7Bykker/SRXv2bv+cu1TUD2Kl9cwksjhuLwj25
gaMyQMI32jxZtRbpdmu+tBIO7gGwgn4n5JNXEQ0ODmvJe1jIleGCshPMRsCbqwc+bqGl4jW3G6ig
Ju7D0Hsix1+1XdAYxuHeqLfjgiPxxvCvHS6H9aIlJUi9AJO95w1/wqfzQahVe5Vrb5Bk+VvQa4m6
doxuLyBDMy9AGKtdFc5o8pDFH5ocf2i1B8Yfbk8q4Su/JLe0pkxV1M7BhDPHaAGyDJubXtFDPOcf
EhUh+jFrISS+dsDgUiEmWjYo4USVVEzGgju5ygLxOJsJoltMiFsKD6pcpRnFLG/Xm8Y3KjG0tuBL
uxCC//ppMf0TUmjlMjgaHUNcXwGWwZ6xW3Nq9gnyE1w8xQPSETm2u7FNgSoZfkHBXoqCIhkVaeJm
gzev5ktS22USRV5Rx+Y17TUkFCd30vFGoK5m//En0oNGW+9N1zVQpKrMTxRuNE0GU06XE4A/KTbq
fscn5ASzeQ+HxudG9IQUNDAaaVLXrC90mPkAJ6i2GccVFVbSKOX/LrMFyBp5/2cT4t8oKUmUYVax
T9UjueCiPBi8p/8Wyjnocl+ObWu1X+Hq50TR6fT6Xhq9QYaXzyj/EHt2Dmat2L3Q8/b4p7aw7sRy
PrK/GX/I9l0NginYZX/CrnDKsOFFL0VW6fsEqIzfW82CEsv59L6OQM5WdDI1AXJ+lNwXKaImIdSM
rhfhL94GyVKpBuiHPTWlOYVQD5YbnVb7jpIccX5YyRSa5w3tvZuk8noSsGnThraEMejKdMnms4k/
xVFZdnGYrXxqRlB/SrMZySmHzGln4WSKzxdXaGcQ0t9nKsFgYa0qmf3NKT076DOV3J023BXtaoNr
4f+UvOhavN0j+KJIOVfrgdrjflkmnw7vpcoObHfGB1yzZDjNkYbJpfR4vSJbXMm42C4MRf87Zm9T
tOV/2QM/aoTmNvZyB6PS2oj5NmcA6m99DhQ6YllGj4a1ZjSvUqOdyHq9SC20ldpASg/il2NErWP9
Z8VC70kCynynqDMEj11Nb9j1FVkpxY+DwK0tCgRuyQBjWmylbECsd2KZo0Xrc5jgJoqvUnyHzpmj
gp2sAldlaJtZb/NQ2CGZqDebS2ss0g87TR9spvGAQOT4NpxM9jLvoS6gsxolKPVqEZH0DmGRzVvf
lJl+fNVHyW+FkklJnzyGhVjt8zO7SBWUXgxbxKqe9YZYHNy/IMkd2yWHnrNQoBPEXd1PrUWHyiCI
P7BhhuqnNqj1G+z+DgAZ+X3OJDy8WDuefUxLurerTWmto+cK3sXoGNna/e4PS01DqiiOhTbVNB/V
V0syE9G8Q1debVex4kFDA54FHe88qYVLi7P6d/DTUeqhE5P77F7JnMFDpYppf+ZsJ3ZeMAdz5A31
lvE2TZMXCuff6XSeAi8sImYJG0Ny4ZPBE/BAR9PpJokf3cck9Fz0qg8Enb8dGfv8HxKCh6w1XBQU
tGunFqpUJW0qth26Y58/rJSJM4Bfpn3WQAZzCKSCcsf7Uk+uAKcqLf4QprW0SrilaIBeOxGSJyfT
R7/5y7Qh+kOr6GO8ZsK/fnCQTUo/ftUO3KUdjTwxKlz5+tW9L3sgH8R4x118Kp1Eu/gBju5JIKuw
jW9ArkDJyoWmfbn2lw2h0z23ngo+IpnPVdIPiDkZzMfVcnHA71iOrt5kXMMzdAKf7R7iGuU07VJg
gudZ7v/pMp+Cbud5giOeAw3SNMgQ6pygJR8d6i6P7RDQ3OUcREW5ZJQJWakn2XORzeNZPTQj9eye
a4CAQWKderMTnfvldNboj8zfhkaC8nQ1QF2xJaLTbQnv30s8JKsUE6P2s0DtM9Fai0GYwlR55wmG
rVz45xRRD7wufzbh01trL2UnphJRFqybIoBKZ1NklKJwopr+5wq5zOb/g8AHY2WzKuev0yTdEYFI
Dp6txq+kwyAZ746gh7Upt3UiHbe1AmhoPQ76SlV41w4uuMyLGrmEAOGJ9vxK9/3xmP//a+W1xAGj
JNYWwmksBoxkcB5ZxXzCIsiYH6bd++e7OuyH/mLKXqdcFN/jNVTsfdLHMXBNGBa7/b8QYgVqXVJg
cDAIYX9BgrI7416nfeTZEVC/CvO3X/k0ymy010SZWK6x7vC1ZffwzOl6KCYV+WTuBU7O8OXApBET
R9bqWzM7H8LctrJZpTFtADBckQmn0w6AWwqpRWYOw1/SuYkCkAFyJc+vThzTSlCnvuG89x716F/W
qQbZPwCDXdhZZONYnv6jJgeC30TrnXwyz3FUwF691AHfj00+HlWQy/xNDHAWzBjSeXT0r1+u/1AK
OvYMZhy6srfhv3Ek6XbRNprmAfTKxzk0RwXoJuDY19hvZsR3Qk8wGNeaWuOqPrhlaLulSqGaN6ri
4me/V6acmXp4fIxGFh1PqtJgBtkAqQzxBbS37za8Zjf4gcVFUcM8H4Ddg+SRtafOHKcubTq1ZiFp
r0g8caGESeHpWJE21q4iLBtYY0N3ujj/Nnld48TV9Bf6nywiSsUi1+MWzCcRPPFhyW/wNUi3VCua
uYwy9Hkg1zWJaLrEYepT72hrqzo/kC8fBpSH3n0tzSIKBDNx4A8SbH0brG70BN6zFf19mtaHwAgW
g823WgzIv8IZFh/RxXWwI5tjqD3K4P1YxssQQ+s+Xmj1PDLSgYRxjE2Pups+x/s3usd73cb60o0k
QOOCi9UTVUzjBZ1PaMKF7c2m9KtaCYmEn3uTkZvYjvnY2vhJCG6Vj9J7Gf958iv8d+fs0XIvQtFT
8BRzt8mBHDNWXKm3d+Zl8EtIwI8RD38s4WSJ+7K7nwZFzF9NPsf19lYUyf6Gs8ivB7MAzRjeRO7A
hIJBY54pKdr8GapGAL47brbTsCHwam8fuFJSCJ1ZInzOoIOdSeoMwombpfHuwChjwR1L0ZuVi329
90kTN7OBgFaJwbIITe0lzLoDR9PnA6ejJFwVfxnXNe2TNujG38xXhawJdwME2jwZYzpsoE6gHL1n
mXDKjgSuEsQsiTnsUWiYGrOOF09P2glHcmf268oI129yO93+O6IOwqowjW89GDL72GQ/4x3ZXxZF
mJBffbGw/7ZsuIDdpXPCvJkUysyb1MU+Kf0PM4DaRV0eLbBg6toRYazZwBIj3KJc/E7P2ylwQSB1
LZKqyFE91oSN8OpvZxd9MxVk/dxGRSZqYXiMfaErVghIdi/XMjL279w3uVc9nLPIHBiHoXSJOkJF
4hGlkXvHxks76JUn7U58uuTj0mOp/2o4eDRohEerrlZIJL0mzIl5bK3BlwJSUAWWpcgXRAKovq4m
U6Qmc13JsJJRf85rXHmBDtL7Y624tQI9m1rSbUc39EmfpC00IQXqatx1pspM3h7BhJikolUz7m6E
ABQWL6MI5Oui+ZrEJA5bAEXTJvWYVsVwzbi1JWwlitdBLXP3f+LUc28gMKV6bICMLibQtY+DJDjV
mxkUvkbuiNk52+wweAxKJvJabs/A89+vVnv9p3ktJsLXm19IF7q6rVU6UCFvO17Yorl+6sd6TaI4
2X00WhBI85fNyvJQaw5EHVL4nQFbUgn4VRqxk/n2UeevANdKHseSa3gfjCCQVf3KkFw60IjNtX83
svSu5/JcoXhsXQ6qDp4s6s9tsvTY8X0yRZb6Kl5OzNENhCClDHgyFsDiCRODSFTthsTvWATbo2Rz
RzDRYvsU0AV2XwwhH0x3QowJcX+4z9GW3kKT7RyysNUDHlUuF9UT9mmlo8Cvox9gEUcb4tSuyPJR
jkA3iiLr7hfwXQDnjPDUhbBd8f/RWVbLXxwNjrtftOXfmxYq6MvhDpF/4XQWIrov58nGh8T0NAHQ
+rtkN2LnjtZUUlPG9At/wIiQAJxCuBeDB9wxvvtTzrvyNSdoKynH2coUPBKHhE0Mm+3mq4Iz4rCl
LiOeaI96zCz1GRM6tHojTTTQWj/TePeUYzvq0Dlu8dWbW8KLduNKFiprdjGVH2okZGSHQuANwKGD
0k6l3twsxsVhvjCebbc/ql6FhBRjfF1Av4U/CnW9WfHp+Hs262X+KaDGaVSg2TsrWdR0rF9/VP6d
cgR49TFsKpVpwcEIM8XKQPPkX66jNlVlZbSMwWSXOLlqt9i3Sj8FmT2F1bH/B6b9tlcc3vDYx2hg
zEGHBrMxW9INkUchTiGaE98HOUvDcJFn34jl01JJDgY0KTjr4aLwQ1oK2GOPRlRB3CTOpAuRZsIk
hhpNg1l4BcO6ZzNGjtWlh5e0D+khl4GEI7WUuI3Qj9aV3ToT7OFVQSUxLAB9lxpt5bxi0qY2fs6D
SBRfGTnYYWxY5Q+b/yVY0XP1PtN5YWfD7e9/+xmXALlIOx2KAFUs3gRDc+FPPsdfnMVTVPErmfy2
DMV4LabvwOx2ncRjlhBe3Fgcu7XghjtNEk6VHrgs2yFTXe194YJ6PT8jtrwRflmkTlV8MFQk5wtS
A4/VOcCsmoFWtRB2Otsc4mc5Ym4wnPuI6hQqTURBPfivCbRv+Ut0+cz1HnRv3fdmaQF/iyrlFOvb
5rrOAu4vQ5caWj64dRVQNi23JJF2jWM/ApE5XVit1KqaiwoPQq2bh18QeQAi6hzntf6L4P8O1cus
FMMpCPm92VgPJG30irpqHvKkWVX8vOP/MOM3p+m/NDY3Ty+8jUb5HUneUsYWDq73w0+9KxbQYDxY
dIAnxHINp9kmx9tNdc9SQq9uw77QLNV2jDiDBPiWPoF+tj81Bd596efj57hBO/ZSKZmYP6+R2MWQ
VmIBEsmDWd3g0gDMGsI03FYtDkdbcXxycbDuURpOpV6iIV6yjcTtLVBR9y1/IRAfOtiea1/ojmmj
7H9SeKLrrEu8H3DXOef5ppojpBYuI35xpUgke5CV0wg3cPy7d2jh9ehOW7Q7kFQYNMtRuQKSdpNo
bGpRiIDOtvY5OrEqEubbHePrHDC9m0SPOIN4TNDrT3JglTB6SxGniEmXFwQnHjf6aLV59JSnf/Ee
JdazlQ8BdLUJA5Q0TLfS8ygIMxN0dDz32iyGBzxgDUlg+7onJIrSroUmUygmND04/pr6NXDzc0+Y
E6X1pIYn2+AkIDq4GtGA6hq99ZYBJ9/q2fxhkAIVmCiyUtaBJJd92OVe0d8qpy4R7xDmYahTRKAM
OP59ITm9tjs6c6I5/CCyBa6iQJW35eobdwPCo85jDhIGKgdCg/ZCLks2aWZnn8UnKM6ZX0oGShp4
L0/zYgSFd20d+l53gyFIiLlVbTtLw+73Ifc2otQZCBygQIiyCV/tv2GulgeiEe2yaiUob50TVYAL
Pr/offYVAO08XyYpb99wt6i00fm/8+YFqwzQGZ+BnIz9KJocERd+dZa92MmWR8imgQP9rkO1Dd7l
eUY8trkepUWeCENn6i6jAyxgO78jVz4q5ZOr5M7A8ADk3CxR2fo00cXNFMQDUy3qTFS8CTIvPDCq
uFhHvBbVGm+P0u1cWORFwfnyiTZ5bgGeNW0CxAOoU/UzruV/EsYxO8IQI0/hFx8hnOt/n5jdwYZG
N18CVQHpowvojs0+FIvLjR9+GKzXmjQQl6nuuSaBqcJC7++pFTMRWEWoXWR+o3Wugq4cl80Vma7G
tlVc3J61MuLXLCren48Q/QBD5arr2DafuVnrOVlYtoK3GQwWY4uUyLt++R3yMHD574GwvlMUYdS3
xHl2ediqwF11gjo3fWfGxFLqckllDgQKBb+KuZ4ZLe1eUp1etzLA1EB/vbLGfvLV+vpYizaOtEEb
uXsZC6mqsXbmngrpzkhv3oyeSB0SD8jAXPH7Bo1oQwhAOYRhryL+DdgBwIACWLC9rCzOj5hfmswI
u1rYMrObFuPoIwna8G1T6HsSBntcYEQDs8xMrDtGQJ+4Fsq1cmgwjxtDUsjlllhrnuhd5NhLWHVw
UqIcJjWABx9CA9Sz9165PBj6rHO/1vEjjqisYvj+BeabsrKJwRB0O9oaif0Vmx/Wn2Nt5euyGayX
ah+i1qYa8BX9G3fwjInAEkzmFVRwvAXqZwgfE1Z5WbZqOn/7sjPfSskR8apnW/0DWphyybTCXNPA
DWzhSdCrM951yCxHBK1pieB92CRJaXnPDK4WlR7bpZVsXBRl/ZQgfQLTpfSHqVG4OnGkO4Q5mOlr
D7xicqUFJ/abVxFJDTq6MYAY+K+h6H5z/F/zERDIwJbToXRxSDZEKBNFApSs7Ha4IEiq/zy7VNfv
kl31fF9sc8ZDKSvpcA2jpoouqH4TvhfKMgmOQPR6CNQl/06QMbeHg8pu93QJ3lVAUyRsceIwPmQA
3RgQa4aM7Xh8rto/2H2X4oYRMncRv7FHl9aKq9J3T5qjyUO9l/vcZ6SgDvRFVeY3nooUFBQAMsLP
pA0RtJwPsYQ9n2vGrcQQf5l/ojPuJZ+3hM2eAVUx5p9Y3c1IqUalD+wnqjwv0Q8jZVPQuva1xbGS
D9DRiPpqKyKfnrlDgP5mnm55nMHb/QgHRHLwd6fwQPBtEZU4TPF+1SLoxFgUa67iAKKpqqy5trJY
hQivTQwMmCrq2Cb2lHA59YtuuaDoMkHI2KKNwIW865EgohMTGbXWfRZkSvL/5dahSPobNSqITqsw
Uz3q31z6MUt6i4ieV6lT9n5E7lA2aq3o54lGxb75CqxJMBd/4QBBwCV5ONr3ELQ2a+7FnLdw4XlI
JLvv6/+fHbARp+U+oscAaA5duIn/X63VcT+Md/WtGmgINfs9Nh1kf5ewsG4bsiZ76tniUpqMjY1v
IxDCurR7+gExcGjKsrBhOtnCDG2f+MiUthLjXIrGNb1nrev61+dLqE//h7gkfTcsD/WKECGYq+ik
gg0O/kcEsA6Wrv4fXW2Ec2De942bGkuf1WXEAA5GK6BK1xudWzpRJMZW5xASme/KiRoC2WnCMgUo
0oYCk1P6xa0ivIY64S67r1KoR1hOO63/MPhi5qW5fRCV+F0k0XtT65ypfPtcacysXFNJUhVDO1QA
ENagqxAZp/Viipfm0jDo/1hn2zOrIWo+KYBx2tXBtllnWMq9Te1VzIEAMVfLaRf6hyvEeBfoBStv
plupN+mTqq4gF2HfIMOf0G6bpbj1LODMdS3X9QWO4ZC4mqNp8X5trqC5OIeDBoYVzwIn1pBO7zJD
c2AqWxePprFD2MtkzMrXmW43kxx3JMBHQQ8WvAPGtxUbR8j/tu4C9HRXWBISN5KCkiUMobQChPs4
VbC81SxHDbOx9uBe/nB/nuNzhOQ7tW9njFMzZJVOggCST9J3sABGlHlGD1dTrMc/ieXs1JH3wJxG
PuWT/fktH13T8ijRmSZwwCbaSEYduXsiCZnAjFpCkYKgbYkPgpphlc5ixXXu2csICfPrWurK+zKk
vzJczS8L9nBEQtgnQP/j45M4hE3Jr69k7SJJXg8gGJAZUdkpISaIXi16C1UMTV4BPHCGMrklMyoO
bHkbUbOlRobc0J3fykskS7jVm5xubruJBCn+n2Kc1P++imnglIC6o7AghOp9MFqu5tJhnN8LAzRD
GxEj9NgG1bzSlGanzWdCqJW2ohplMcLgbptsexSa95VD+ovufaOrZb6NOYwYKiCBSNIZWrr5KJUY
kewgcGz8J34gHJkank1XE4jRCsSaOstpbKFeADmNI4MgYMwMMSjp9D2azYkttPv8r3Vd3oFF4Y9j
Dg3ITfI3qAkBPMFSQHzzsc9ZK6foxupIvffa5/qOWHKMHkX3QEtvch9Ye7R02IHD5S3nvN+kvhu1
Z375gpqD0rwOWePzZ/wkESEw2X+3UJ8sZSp4of61MA3AF2GIBsUZ6v9tLeWqw9KvG76za0qC0dBJ
ENGYibZ3G28w9Hs/3asDrY5GNLzX3wPiJOd/dEVhK4fq/EkjJkONCuscT+HSFTW/+Yev44xDjC0Y
z0WW7I193qePFuSclG5POX6Dqedv40o8qsmyCs5Yau4HcbqMWGEvv3H5QxBXpjOBhb+X2+7J5SXm
I1LfZva/wcPx8OO7Hy6ml6GJmqNp3Rt1oDZgFVG6qsZTHLR1p+6+z3fJAgch4HJ5c+lnUeCJJMMb
d70VciNEKz8xmHzSpk08l/AbNM/9RkM2kvPItIbhKohPqzpirR37rU2Eis544kKakyQEGDbDrKGJ
5L+WsBFXwjH40R3sPivw5XA+63ElitGu2n8vkiu/4rKC5GqXm6PNjeveCN6KlagTAfvNJC/CyfFn
h8+o9Dz2IKifls3RCHcoAoxNSpv9sKbs/UfmwnXsX7YX/fs+hYL++rgUK5A2FrY7mFmucDguN0u1
QK6mPDA3nb5x0Lq67P5EtIGgVaiLJ6Ab+JeGhG09URdSBbOySZIpmpmClX8t0GhuQlkUbnhD6mtq
tGqDIzmhqObGyGTWfgut0fSvF9AupQEAEW92UceQu7quf32fgVX35R3iho4BBbnkDE46PDbHhOfV
dfVMcMy4qithC6q7OVDaF5ASaNoE8YK2MnpeDOErhz90jeiwSA9Uwd+Neg4ZOhosP3Q6Rk8JJ/l5
XOK1YpZ2tkSZq6SzxQsUuXlPqwk9BezZiQGNnN/FZsTAA5zwPF1H+JvVSdMD3kCG6/KB4BDb5x7x
ICWdvs+qN6Sc9PH3efQTGrn0+P3MnULmMns4cc21bX342/w4eWMtTgm34n8Mg1Vz7X5LyCyTiDHf
DRG2jS3RZFJ5X/iRbUTqXnEu0acNKvqrmX6/p1aOKhZOd91zjHw3OAPLXl/W23UgxnCcrjMR5H8c
VfCBySah/c3ZpTQpL7l6U2BHgENOZRp9wYiJMv2BWry1yLoUtfWffEf5JfZ7obsO6TZaGbFSDKzj
quCxb1l9/iOY4WKsr4XCgfvgQQKAFhaxpV2ADRg8cdfVvkU7ZgkgErkh+BuZSz9fGkUnr6u2ZPYs
VDXveragR5yPVvq6A0B4WHb1e98NsuMS82SbasNRynD3MyDjN9g7b7HkIPg68D4KQwARLdNKfJmh
T8eYlp021K7uWOST8jOnaOooGI8GOcQp3Sj5ti7iKSldYw229X1G7sBLStxM29NoqXOkn+gH5rn0
rnU94W1QcsEcExSf8gNZOE/++Lw3kPGNW3Kv0wN0cU6PXNDDIzBMs/s/LRYkzCQIOZBz0zAM4Lhw
2YRupcyaj534LqZAMk1m1k+IUg69zoAEmYO4sXBCkDaiU64SMGvZIPpVJLq8pkIhQcno1nc2qYX9
blefbVFvyPXBAd7lLcPY76GSco6AWgDIOtGWdObyJRSGPWzk6DZn+3DKE4rdaT72e16KklxL9r+6
zLFPsQMBnxVn1qePaezRnFWwJ1ryM9dzEpBkRZVJ3UY1fZlp0tc8E2Q4MDeMj9VpDbPiVgDqrGK6
H83L2AQosyPp7umDu4EmQUDNNTar/zeZCXCJNep6/Y1r6S16GEnuD7UzToTwVBN4gRBhLSr8bVpS
D98C9n9Je1Xz0Te8vfysf/CnkpS5wXNijNbKOe2tj1hK6ZTt7dH0OmL+BNDF1RUQzStKmxf1ohK+
nQd3FEGjv+X1EbHIqlcfmJc702Bj1fh3K26ON0nUj5PyPCfUKlc02cv+kvXFWmJN7MIvhrehCvbw
NNAec4gQfEc+cCeAMVEotE2PSxnBneoGyv1w85vABSFwqdlgaU644T9NudSXN+kv7fT9kTiEcmOJ
e+KG3KtIyml8zLyUIPgDv2ZViLDW4QcybI0zjmqueyHLoMDbVLqLmZpbIjdIbPMrtv8Fpqk5hAGT
syxNlRE29lXnD6Q6ZtIYbZoJe5Ylj5IAB8CIsxcaRINbViokScZnDEY7Ttsg9RewZ6e7rKcPIoIu
Z9lU8/3K7/SvmVlvqePuv+TfMsO+9Yd5BZZHutKxwC1kKr+ud7Syfq3fwxLM0hqLQwIf4KnCww8Q
cJ3lZqtfY5A93/cev9dUBwl36/H3Ix9AURXxn4kGPPcQWtERjhHRZU6QCKqF7Xlt52JNwMDcYkqE
fII4wtjwVNSRXRldGedIlMLiOfPh4c3IAZaxHdkFbKqKAlTdToW/DxjvBvorxmB5B0c0UcRi/kli
7suDgWh+i/Kc8wuu0ixXvG/E+u/OV/sZ9p41BIZFhuavHIoZOeQ7sgcWCxfaOGUBvELXOFV1lcwc
fLQV7Xw7j27ywoDVx92tTBx9vWcpPn1EMjmD1QQRKj9DaUi0yyD1O5XkVDdtfM3Wx6MnjSOpx5VL
Y6Jm6GJyPqEvmpecbgz0zywtxaHp2bEMi5PB7Piwa194GlHelWCL+l9Ctavof879yd1YrHmMSd6j
DovTb75TFPTMmTpfim1fu+x5TFsYHYFvatvG4QHXg7RYFlBOa2zpfVN7DtoRnUEYk7MOLv+T0OS6
Kle2MJ8CAjJZkjJ3LvrDGVqTbiNK60/qyKOk32ABa44cdnWJfK2qVd564zsBtWHBWQ4hGs8Bfv9c
SbZ7rgYugRRf8u7Pn9n3duNJEQlCMEhFWVH0PuUrwfF4eVpQcFdJtE6f5eUt8F77ucAly4uLA5+D
uAFh54kUXTyViVVo/ACDDKLn9DrS+fRD+NikJI1rq+D0140j6QgPRDlXxmEPNpVxth6SCvoGw/X+
czunSKQ1xHb572fXSO6Qprnxnna3B2lJ4WtHepqUNlPV9G2sD9ljDeifovi9kLB7h+0Y/sYWjuXJ
w/PvJi8h3UIb5ixaQzD7+9L411JPM94Jhdu/LR7ZITapvR0qQcj65Nju6vucs06GcmoUuiE+gEcf
eNBMkgQkgKHng+/KdvMBm0aOncTfPxzBPZN3qKjDfGlzqTsq7kuDTImGChs0SshvHnhWMiVLUkK4
JqhUjdMRhQLDKG5T3A2PTO97KB7Hs6/fItmxQs3wFOzpAOW3YJeOh9s3JeNLuiqVYpsPgXtGn1iN
15/DlVmYv47D5EqpgQpnX+loib8zRXErWoC2DrF63ldbQhAQedKfMxzNhGmajI6m62HeWezSHIM0
6DxbqcfBBO6RXymKL56vfefpLEjFjzB8wzYEgCZNTMv2m4LDbCGBLpsaGVLbsvlGWSUoSrwVDFL/
z/yoUN7x0pDmuyTef12FVOK4z0lvY3tm0cJOXicwmyDtBNoITsnc5dpbHP39qPVTJ9fBWLixlFUe
jjkf+JZOLkxgzrqjNiJX/rvsTpGDH7ecVII87TPbh4O4l/ay41oOXQoHLOsf017VwfOckHdBimte
E25Fd+gWillrzlH8xRcVzNxMdBErMlottsMdj6wcVR8z86CAbwRfwVQh0LvBCJNRUyUzTYGeHApk
jDxRQag2CSPpVnamUMos4ec2g0LqCaXF//tui8awerblsHxVrEp2Yk6yJd86w3sHNZy39T6wgba9
uMH+mZ0Mzlhd4CYHY8BoQRwFik3/OMzeKJlJuAB22PN8UygLlUuSJ/IR44JNfPg0G8f/ppBVb1P4
vKJOdPUI3RtFdPvmgMDEFlwizXH/92iTGwdFY7aODpSpV7+oF2TmuyB2Z5wwb93w9E+h+RpHfDGb
g6cyRL4VIn6FTARYnaQnooPUN5NvgRS5svDtxfvA9d9cwTHARGtkOpgWO+c2JzMpYqmkGLjg5wfp
Va8YG11VVEAIO1/+CNhKGZ2RfVw6DZAutCF9uxhwlGNYcFumsZLU5aIeOcjxMiDIUFvrVVtmpLSt
xBU2YcMM5BaElTL20vtzZWIfgc2kPfNjRpidqRY3/lpPQBGY6zI8v2k2ABeKdvYvoR9bHHN9S8v7
dshzAM4fPwBPJHw3HBbdrr01Oodqk6LlWK0Inurzap0IIokLhFM1fiHcPLQknt6lAh8XEwcgYuBH
FSV9Ba+JLYnjr2pE+YlQlvqYEsBdflGSTm6ysHfqRVrFMpMmCGsojbdZLQwWewvwbr8kTwHnkEOA
CEjAjIfevc2Ektjasv4950CN2Hn1bQbk8E6Vtjyr4ZAsT7Kzxsnf5PzPUdsw1RZAq7wt+V0k+mKW
gBwHzGLUI6pkR0/QPPmADBRQJPfhIGCiwYZRuUIj6Ojle+blRhmX99DXOM2PxiZWP2MPdqy0TbWo
npt4I2GA/+sVeXYCYS3i1Kc4wTutQy0ZEGiiZiK6oeFWtUDwhltxWgLVu4QK0FFSnID5oDtzMjoy
c8RLYKCHL57ESl1K0DaQVt7pMZYCpNdBWe9/eqQCMVIg4t3VxD3WMD3wYcwIreu5IdV2EMRxBvIG
kByXea4mY3SpskI1R1yAjvwmX/pa91pOQuPOds5L1ht87ZFRD60OIDpTatis6XqepJ7i6XWprs3o
VUWuvIi3BYhMNWUdDN3TqogPjl7xBDXgAkzUgLpsW4SksXt8sy9YMKqsNoUtUbbEmJwT75QrERh1
Bsbk0c3w+INU+Pn17ccYM2XX32gZU7AeUaZl7nl1DIF9PV9hXSoIppAlAcV6jf+CxUAEjGbaCz0V
w5UBkUERwWe4/OmIfOyFge5zTBj/+LjgZ02mCUTgbj7W3CY11oqvFuS68glRn/7YUSEKPGfv8NKw
cpxU6lG9Owv+IIxAIpBB/lqFYeh4vrcZz8QoJtfGDvHK65WJKPBNoH2v99D7LnP7jxpWHu65foYk
nyYS05wYdscp/WqIy3+PHs5xJTB4qqIzsxhj8mVUPf8U4A1zIsWZWKVUiJH7nA482qICNr4HgVG+
TseD0HWSFXvDIFkFPftLL4OX2dNhwQson46EeCDb7YBhTqqd6GgE62722FKj0XkA5yO2nXo3wjSn
Q4cQVViQSmd9Oqj7fdppl9xySIC8lR1f1d/aVOuUZ04G/dQ6G0JmwBpAe3jPyirjUjbvGlzDoSsu
oT923kVHR0O4oReq3zkR9A5/XPrAWqQFf+NAHJePpH2XYKKvr11tu9AZmRMS1MA7VGFtHktu1YmZ
3Z2gNTHxMe7/fLko3ASt+7W3O/zT6BpGh8TqKrIE7/8BBdbgKuYV4o+X4ekc86lMj9pKMeN0C7lQ
NPiR+VjtYrueAGg7uDdYqDWwhwGfup4y519sPhunYMlb1g/kWwqW2pxFVrY8rPCh6zGM4igauMGN
w0EpQ6QiAPuRWLiJSzj8tUgwvIwuCRXE+3dyA/qF8LMNhP3LvqJQZ8BFUqXnHoHsqTmMTBjO6Kkt
83/weRnca/yQqLw2f0LZgzrIS6mzfv3gxBT/PczH3YCurr6Hc94wBstthENHqvi0GeehX6pHUVTD
/VqIPxr0dFAWFKSxxlB9EJT/23ALvhOe6LzaDLm3cHI7tXW2RYRr+genBqriQdGPBLH7LT2BIeOM
65lxIm3+ViaznG77RgMst+uoghk87IMpfSrQKRZOauNfslDqm/dv+kyLoTZ+PmhMEqoLS8/KjPGr
7y4P6u60ruGdjqjB0c6x65G7Uo9KFKjziNqjEbpaBJTliURoJf4r9p20CgDC638Dke7MjhEB1+wK
5zI4hiOA+n+nvwSrTXl64oCkDPDRDNZ/yfuGIUAD7PUT4DHJ83NIYA3FY0WIaAPqXkTTHGFyFH8N
k5Mry9Sj59Gdee4CbL1dAORL6elCOm4qmdqcKr0aVlbVbNCmr1P3P5qRcgjDDelmtZqIwH4hNPuO
9KJ0vlLem0muggdkIqOZevvYTNMY+GcsXeqhPrCLQ2tQyKf5M6AcGR7WIlOug7sLc+Op2y7RMqGJ
SZtDz9RSojn/v0Hf0ZlC9fF97fy9/TolCtB/EYOceAaZugW/7+8+T/X63p/aA5HVkwzBY5yFpz/l
HkVjaL2pZZn4P2BARuLJF/0FTRgxguBa+OBt+yFsWPJfNFcfGUzK58PR/Ozt0K/CVLGrv8PgvHAu
T1l6IkvDosS/U+PvOLRoUgID6PTww+rt7MoYZlm62mXVYM9zNW7xji9eDlkv5taYcDyRjCOgN5jF
rdcUpwJnYs/+ItTEzX0BgsBGMK7gC+3zWO+yVowG6HbvV1P890M6IQqidZsfgPm+h6lmQY5sLHNZ
CNOw/6DaT8j5SDxu75kLW5MkEGEPCMLH+IZiuFDDfarykWWj0MiB+ggioQMA5FR6I//H9ncpiBOd
J0/+pUJnJRdiAu1S45OsTJr5F7LNR42qrd3XwGZszaTncUg6sexhQiSaOPJoUQRW7H1q8gXzpgVY
lTHY488pRC/yOgC0N270GnQ9XWcCU+YnLreQyRcp0HWxSxB9lNMlSrzamgkAYUNYJM7O4y1BJfcy
MgooH+MuEHBcfTU10XWXdOyDxWwb0p3HqlHctGrDKZeTnTEFse+j06amk55b9FeIbFCnjQW8kRUe
4MFRXTN2b6w+ewiscTKqypncRH/Ca0Hied49K9t1XzVMpm74vmgTfejCIslJWb8iqSK9JLQuZDGX
h6qf72phd4a86ez6hDxuYUtW/Rvo3ixGYygOdXo2FjKu9NLdxU2vOvTpTZBMypOiUL32bchEfNQF
nxWrfLIjlyV3XMMYzjNv/sf3X6TlmHaBRy4U2RVMTjeOHV1fXOFA1MrxuP580idS7RyxayAoI9iR
7BeUisIuXCqENL1Aq/D+6YQSCK/3zZJc/u1yh4PLacAF4W3+koFwXGeVlw1V3+YfFbFp4gc/dKUR
0cH0dsFT+HFuGF74cd9RtlZf6CBt9QM9crYejMhY/4Veq4Qb8xBS2NSrhBxR4Yzd6/yT2HUvX+D/
tZgr/kzFT8qLHE9UqUcwnIAYNRoIJrAj54IK5PcrAv33Xcu9YFjkg4+R3uvAz6e8TwP7H7wtYOnr
ZOLUDg7a1U7QZ5KCZqyqK7kYbUQj7qRg6NOfjYFtO64fI2BhLtIpxg07CwbbIQMYxpc2Gelv0/9j
SN8oryuiTfVgkThhORF0U+PIxU2Fv2mJdCmCUD2Y9p1xs4rISHcEQbiLT4vCN12+zDf4YWaK6+3I
aTqIK7l9I77N07hMV+nDFGt8Ci5j93GIUEaJLq8uycs9/Ly1OJ/COtrXdBZqr2shfQuuJPsCvbPs
z1LRXCf8qDCtamTXhRb5pll2ig3tNo0Yj3agunXuj51pB0DiTKtERAdD9Riuo8XYQLCvycO+Pkwx
Oq/QG+OwsGwfVRvUJmCsHps9jmT5eqjZ+APOAbIFltMVfF+o2lF04kR67D+WpEktW9+V418wnBP4
Gob3wQM/ghM/fdeq+ngiyTBSUxapEa3JGgL+BFhH+bFgxatFYULmfUKCTvVLCjR0qtRjVZFVWsK5
8eI3JmceYFuQe+3bbwIgIN4Xv4jBz41PsRAtgkAJbqjWKsFbyLCb5dtbyztmLSwa3bVy/H8AMqu5
ekoCJ7c5318JsI90/jzOIUNYMQS9n94y1UdHMbcEFzBpph1aIYmb85vo6a+4VLxLTxKAhGsJbhiG
J0y6YC4RHF7j1B0zgyJ5/dv9STJLP7HE0aZyVJvgeoMSIZrkoWNLols/3T/hR0yFGUyIKe67W9j+
dsOhz7sgUSKy4+W8tBXTVUZ5LDuITyQp99oK2arDZGyurtq4XVcx3w1UTjSPGSC36dMrlBTApk3g
LfajShebhUtXzp919uSoL8WAi3iw++YrI6L2fqWmTxmcx1tk3jqrdNjlTsJayBVNaCzZe8detQF3
edQgt+BS5h5IEdkXUDhaC3/i5r+P8Jns21vRZz6k7dEgNwu5hALCePAYg1vcexTZKYW0Z17wxpe1
TTW55xg3shV93xcdBCGTK7PG+SWab/QHL+KKkE3Q7AKU9zi3O9eoHIGnn6JO4QD9NjukqjUK76Pz
Zp6c0Ey9aqJI4N1ldy9MouYstkmM3Jv39LcIVvMJiBoGbT256ASs+8y05Cu39z559HozP6c2EiKg
yXpo5lgpkJaedgOJSg08a/BsRPkW0FCSbQVMABZFeEzPM4/wQ+4LFuKlIpLklQ1GcktTBB+Xw+xq
sPHoDi49SEL/H/4o6p0AMx2UjIHYNkNNmPv+QjFkbld7g7GZ0RqKBhG+xM3w6QiUnECvP6gVjVTd
M/Z2CfP3/BL8dT82FaR1UNbAc4MZZ0PGkNAuo7uhJEgCc1Wcer8jMWTBZzV5JBa0dMpCS9b9DxBi
d30ULp6v8Hxf3GSILfszwrKdEtMJZIOQ4TPLHJHgjkej9VmboUHrlqA+3852uwv03iMZlQxnJsRY
lf/zyky8ibco30xDSEfAluK/kSYuAufhNX0CU1uZ48ZvZYcYydQwoWq4+93VZsazq+Y7ZL0OYTZK
8YDODWioD0/oJQ5zkkMKUni/g0GuM/n4pVpJxbFyKIWMfAxHSSdFPdZjTqBab39gku1nDATpPsQQ
7KhjKK6ymaZcng1IAUFNMRaABHaRQcbFiEj4F2TJod3Gvzp+MZtjMJtbgE6t8sKN+97davG0Pn5d
hceIaoqqEIe0CHh4FrHiOhR3gEzSqnoyM2a1g5+ZB3BYOWvQobAKwz/N/6cdQXIYXoQr90s+LNo0
vd2Gjyv1ZakpmeU4nrfOvJJr7E1Tipr/g2dpAJJnG9MgaV9vKf0vK2UfNnImOkNt25R9Ll07mh0G
hKe375yzFl3pZMjK/C2PboCSk8xb2hYzhVEpyH52FI4D69J8XOxULs21xgrn1yHxIs4B9MWBqftN
c6/PpiBvPmdCswWG1Qf0l8GpXio2ULCivrFi8eKcKKRmARKCtDfU56tkjKyI2mzji1llL18ZdRCj
VmB2oAQhENiPMJFUoOheNZ8yoheufOxZfbAURiLTbLbuLpfWSz9a/qYwMvyl6WzZaZFikOaxU3hH
jRX2vlyRk2NRI1frovX2ThUg4EJtCDcp6QTwXQstCifyBzGmmrPflaL8WmRouvr2DG6AGDeVFEqc
doh7RC1udzHs11jVd7axoLMXNU8WDUO3sh5TnAI6vxr0EiSO4/yTTWla0uoO1hOgr6ebzUs8k+FU
pbvaysuFWeYaxWrqv9LiPNPBzwaRnhJf2w4aodCYXTgdRvScwRsvZrx04wJCmlZIwzuQiana9qjm
i6S5MI1MWQGufsZX26PoA1vR3+gx8y5Ulb/GBEYH2xrq+SAfa0ZvKGn9l15QToP6k2WIrteB/Q4L
pI9iv4Qj6KgnmwXz3QwNgeT+edYQhnUQGPCBzYHgqHlcG+bOWeHZ2Lr0pTNUgaJ+emthhH2q7OYK
xCGIhsPE7bCVUa3DKh1ITcQH0Bep93NWelTZB+rmCiV5091QTaPY1M9YKHR1iPQIRVUTHTeHyn9s
zn6/+GAnj9tQTyZ/FXn3vSubJtiXOINvj8lSaBBvJnkjLTGhpD8xm4I7Cm8YP5ZonMx3l0FXW7L7
q7omDZlziUg10SDV5EqHSNt1bIfOaA3dBTVGxPfZDwOed6yJUci5hu0x6TSBCQY7faqejFrG7/NT
CkLP380i6e3HoNgQaEY8lry6phLMbjsKHl/zDxJgwGPL819vKd/775C8xfreUAwidVVTkMYADlt5
sqKj0R/exiH36IG52EeqYtkC/2z4hSCDqilJX+Sxt7791U26YghK494qjCK6MVgyKzzI91CgV4bc
6HFnBgqd/tScxj5RcvzAtkUwx+NXzZYbgyuj0zPprbqjH+/Z/hXdzbfQZTXYHAMzBlNTkgRxUEDB
QSlV02cLly3IxITT9wHZSdk1hsJJuo+XtP2WxXd7QMA+ArSHRkc98gX5A0+5AnuK9RgSogzaAZ1c
CpwyfClkG0I7lD8pZdX6eNzyJEShSZvyTSdgkG9YWOczQHIiei+3iiTaA0rL7iHKk0OTyQS3JUdK
f2LCfz0iggcZcFj34zQi8VIIZqzV3Du1rdp14grYWc+3Fhs3KiojOh/mVvnFv9HgGFnKEKl2XkJQ
EbMz2XH8AuGjxyriH8BG2SysQHZBJbK3/pvGDxQRZokbMWNDfhMAvSoN6NWekmPpb9hj5sb6JzuP
XfTLiBmm6ybbyjJ0kNtjlrlxGiWjPZ4irU4SaWXxnwxly568V6iWDDKjwffuBuIVpShvG8wArQem
fbpukdsE7tAT8RYH9s5otAJo6rIg5K1yvNt5SmYTJAYud39lMBdi1iX7QGIwmOLQD8p+eg69pnSr
pIRzWWWhirJqwDQWM9Nzn6ZF6h+nm31ZfeECB00/WN7eM9q9Lp/FQ2HcWLSGsOU+uQaUO4/hM2SD
pr3bgGCXanx0qto+rK3XnUR6xhN0sNV2jy/aZKddq5auzhCbTqg/U0GbHddHBLTGycO3mDZt1fdo
rh0M1BA6xiERDm+aGV75zu0dkJgTCPH15iM99yUse6f+9hDpFcD1H2PcFitGQ3f2yiiZ6c9XLbkE
OV3zcK7ZlZEAwdJSCihM5lWZ1VHmiyLznX2fmUK/Tss9nGg9wBaGIcHYKPpioIvJty+tW0y/9r23
vCTAbtzQ3IifokpxgUdkIl5oAXzXI6nB6x6HB/2kuOTw8uEFerjre9pY5vlNOGLQATZrULSx3gUk
AIN6WDPcGGSH1VkQzRM13KIRac7EhVAko0b6EZeEsdKoIzjhpaQ57oJvFB98C8d2WYW3d3c7Cwo+
FxACk6FcKG/FPd9N9JGO28Z47AnoOHomyjmYc6gYtX7OVBnrpx4nFk/YnPTbzKQooBOs975Q2nrn
voXxgmwLpVaCnnMvWR6FHmmn3nLkOK8EgZypikrVl4id/XfjXZ+RfDS+FLJG7GEMiqJG2uyf3Wee
Yf6MN8XUtPgIdwuCInDJ2JDbrHuzfocPToX7bw9Txmnk6VYsEH8SFpl5W+rsiQE+Df3gyfo/hk/t
GawvjOM2Z5CX3033OHMLeQ10/7uE9OH4X8z78jKLrhbkemR3SjE9ZnVRhR4M2L5YUAvpS/A9lrSx
Ea1RG9P4CipOsdsAp8cTKUrl3P7kqzJV6Q75woWrN4dLos5cWfbjBxFw05dzInoYwMmqeCXJC8a4
wXKTv6QUTgIKBjm318qR3VaHdMsmNxrIoZeX1wa7XfIwDtdGNzS5JdnUY5vWouxsuhbPCbrXhuMT
EmiypaEA7DxHo4lj/GyE+2wdwH/TCvBAhBnqjm0hJLTP+vz/ANMCgM7SXbnCURT5Tb0nhp2qbWgy
nWvrv+TfoR8olAP1Zqz0wZqRZSY4Yt0ci7rtDp9ed9aCKZs8iNAcSSOtap1G6wgTK1QuUmhf7nIb
Z66/zQ5MXkSdKZLSTQNAOrv9G6yUtSJelgpx79V13N4w06KCiiAaLSayz5NwPpAxX8CRneTaQvgq
RRRqsYIQcMCt46i3IZoi/qGwWaCaKVPyaeirfiX7/jK+97JT2ojN0wnqMX0XEK/Yeu4lKAfZj0Wb
3vAJmvYQZ2fV2YnBX0egBBBOaaziA6rCgGY4bkFbA4hR394kZ8XYFGWkpscq+unyAoZFO7d88vUp
Z9ERmQctCw6Uvxn2DSlwxWGIODuOPvFHouoFnkBHbfb8jbl9xZWmdh5vSTM4L8jpP5xuRWDf954+
p42UF+TQpXSYWTwP5JiU/jCcHwrpIif61f1fisnYRPXnTuSa8sX4LwfiveUbT3ddxhUSXF60wrRc
1/i4WtqUqqFYnwggcgJF9/O9KgtjlGvhXFz2U4OWCVJiJ9Kx3j/Va8MquOoA7zJ5jXz59JbAmdLb
fsrEoTBPcGB/qFepUB30UEdm9EGhUvu6zgguSniFBcR6rQLMTkNXeqTzaALavOu/LUzLSS684UKx
6QkCKYOFZqAlia5SVZitUPHn16h7EBXRIcKJ7j53ys1ZTQAr0tExwDfrfp7uVKChGWBjgSXMzOU2
LFggtoKKvSUcDmD7goGm9QgEzObExtVdnpxo3EIeXs12dmwWjFfHcGMfrteznOcNj/MKeXjBj18g
uyO0mwWsLO+1S6XCP/Cn9FJkxWfxJ7FrrzmY/QXxTei6am1v5mg3+BUBg9ezNueC1Zmui01t5D2V
OVJ8+kOgItdgKKk6gmH4kLxDTqDlBCMxUvWJaOt4B1caNBj+AhGMszRm8tV+boIMN9aAXDn06kry
OWud5QV5nepjEYPORW8nHeJyma46M4rwPhFw1YrcZXj1oyjNqIoR5Dc2TOOPvffDlsbhgQSCyj+v
1Zqo0bklQVHEJCQ25aDQUJtdtHWUKE18VPyhhzXel8Rx/MG1cGWsFquhIkoZJaMsCNahvPs7g8wB
6+mnra0vb4C2LYlCAQV0M2+wg5KJYKMCJHfHQHx5hssPrcysVO1lBttTriJxwiz7RgPJ3OaWbKNp
AdTpAaKUfuLQhvs5UqhMOABDFFaKk+zQ61pVPl9AXXIaH5qrpRJa3Q0KKCM+i7u6eUmY6hO5Trvi
ys0Wv31nDHtYy9weEHyUYu3RxSmxfb+Yh0hqOE0AvLHORunH55sYzdagbomoAw5DdMwPga1+r8nN
hc3HwQwVJ6ddqMIG7dMb4jTexQvyq9WugC8K/GSHM2XnHuJjtTyVXjPpTVMc+8h73JZBfNdtzeXg
I7sSPqxJgzYMUk1dqUyQ8mMYlvnS+R65DwThFMcD4hQcbSICI7hU/Z91ml3LPzgiByDp6Ria643z
Q2MmMMgeg+Vgm8fbiPce2cbN780T+bgTTl7xPKu0pfFw6XB/pJoImpdpFExxv9B9R0BtRlJbESGg
A7Eq+h6q9i9m9q8sY79m6SMRn1lJg/hNRJSi3hIgZ13Yb8v/Gcb7ZXQVb3VKg6+6cgYojVf1x+xa
QK4PyUgw6UQcNctshq56qA3rbc+by7vvUanKLJ5/HopJ8oE5TdIvUBXl92vDyVxD2bYgSgsZEjYx
3x2oHIc/viImYtBDdsH6CANWhSKIiLc+A2T+Z76Ty2VUqG+gcYHv7z2jUpk6k1IMf4pmNiA29j+7
lrQ380Fh7PJUFyETmJFQmk+p1V4ikCXedP1LLIn1/kSg+bCIhs2y07Cb9K7MbBHLtNMw0XupvoEl
fnJHlRDIh1S5ogmBHEH+K0DQ91KAlM/teX36J1MlKyf/uRwEslsK8vop5olKIzt3NygS5Mi5PTKK
Zo6+MNtwzIp/lIf7KKnbcv9ViuBxB414EAGN11pDRSpR73mHr/+s42B9a3Dsd9t+HZ9VL52E4VBS
bmD+IwHqCZ0KBEDpx3S0wkg8mC5A3ns4pWUbbxlQSB83CaBkTrnnxbO47Q2e3AsRvNjg673HFUYW
Om+wfxDRXoWcTOl9SP/iyDW2+p5rqPAaiRo9bRgp1d6Vwbs8ha8dUMp+979pPyPFj2EteHatn3jH
Z9IiQW8pYW0iAf4MGtDgp9o6L3Am0IXUZLp7V74Ar+cPkA2x5fFubw4rtbNteUJ6DUkMEaxMQxVd
RTeDrDmRzlalE07dyHeuojkz/HsHnu3hG+TtTGZ2L8Y9qeqjjKwko0g5RCIqqie2XLOWXJezUUP0
Hhp1OdFTmNH0Pk811e0XoFhX9Phku17eoIJKxTq9XkZs7EumzIwGHBKXz61cOac4FHwki+cV2fU8
J83Tc5nCsvb7kEsMfwkwmlzwTEZqhDNuSfQit65lfG05rm4nOI4cpjQGlYr7J2n5Fk57Gm5fyWCK
04i1WdoZ5ew6XTJigMcoM4G1ANFJg2MuRfcT7leQle76/EUhHC+Kj6sRdlKNThcGaa1MRjC497/W
+kvgmH+i4kMDk2ZUsPIeS6nvPMow3JggAL7BQ7mfKXIuaXse3CXtPhXPeCwhLjdN9NCkTKqwsEOp
XGStiGtEp7Rud79v5AOFd5F0Uyk/lU408YtI/6VUAnT76glFdmsasfiFv+JsUKPso1u/01C31Fj0
R+rE3nTcUGx7IQrVP+1o3JmlWLCBkpTMbhBNjimHm9TEoIKuJl3KmoaA6PutQ4fllY4s8UM9sURu
B8JQkWFdFGorUCvKlbtA0qEGQwO0U/+2JcVmo78hHau1xZokEcbeQIetQbfr+Kua6pdcLP5N0XoQ
RuJXGxYAgginPEPaydjC7z2BT/RtB6beWhotLOHCZnsiysTO3Dyl3yI3mcVE2MQOkMTwIqdFtaGM
sKoF75fgh0US5zztMpXC07xcPdJJf6rxuNWd3JfLCy+2HQ2oc1CcyNLDnuOEeW4II5MW1dF8UwYR
vP7i2aLqa2X12+m3RuWEFx9WZ15Uudl18ZJ77RIS96XfkFXSCwgYGY4wF8fSnC9uT5OTOsKMVSkF
ARF9rydVZnnGT8DS1AibvL0bseOJPo5Agml/F0NvfSMqauUqQLYeNS8eA6FwmRtval+9GUVb1VRg
vpzW5fLDJIXAIObSmkD2spWuErUoiPbQk5dzy53DpTjwuWKDuGi2bdynn5rOveDth4MCSh2DLEuB
CFlsCrjHXi6nEOxexN2BGyn+4AqVM2nMkzfAmWfTSGGTgARYCTM/BDq/M8rpsUPfGqdP6Ml+AZUa
97wVYOeB0kqDUZaE+GpdPrsbDvXHKjIy4LntRVzl1zcBqEYKc7g52jmBbs5ncbxJaYcdJJ7wPK/D
nRo9MXc88/2EmROJc05vkxi3oS+fmUllQ3EwSrQpXknFAunqYoawfEsWi7oeQwfIkjLTFLfw2vq/
YPqveHKEQqB15QBO1arrEgYPbZz278sOeZhyzEmxMVi5Wbv+2UqxPw+CE09+tQNbP0YEW+vGAwqP
4OyVsg0CLKklxzZknM/KzvqXIjprggu7AXfjVkvtvxl2p3qzWBeJWUxiOPg4MUfVNdciXQ5pI5l7
MlzR3ZOrUvgRZiSJwPcdQO4Z4wTFAh728xtDJlnE4si5/4uz+IsyrqS8kd6bijq+vdjSWbMixmoT
SD3i5h0yUb2gXo+FR4QNsgF+m35jrglXKTZAiav0vM7dC9wbelBsbjCsAW/qNR9H6mFx671Uymnm
w95WlcK6ZdmrCEkKaA2J+ZHlbhgPr6GWgRpCyq1zx9Ecyfyri0ARkJpYtiOlv8W2u7xsC7Nwqo4Y
xV5YmKqInHkafapkUFLeZNqZzgZLD1KGBO1JZgRFhk6WBGy2iLGpuFtvPyEVlXI4/00Jgmk7aLqM
ciPlDQiNZisTbnM566uYIos3pGWk64Ir721ea8noSwlHVxh4TwKUBxx3aJ8Ethxfr5hXn9HlimSV
DesP+SKs2FvXg9yNilRDaKHR97NxqDd8yPdjk3hcseOgmoJ62XEq9SoaiGKdfznT7KIbD0rtIdLg
T1ETiAvvXlcw02CM3fB366OVxQ9okd/jWEk34TznhlR9oUTvJNyRTXJ0yfn4k1PJw4ZkREAm+GPf
/mCyeOpjpCSF3EtViisHRsqYUUuo8AR3Lmc9kC1RbKzKDiAhctq8Gl85G8V8Y4v9J32rTl5eA1Z2
Tsk6l0MyNeIe3XyT68XO2eQ/uUh2BIQN1sRQYEDkIN+TG4OV4omHEhprdVbpFmizOZbXq/XADF7n
YX36cuNepi9HE93CkUvbUY0Kgg/i0Qe35A1T0y+V4tSOnzffky/gDRygBERr17Jkl980oUDHLK3P
0lepRaUwDQLmEGWwRH8GNJsG4auatWvVx38BmuXWGxuLPCVlDafs/59wUX4fD7N07cbGbjODhhBl
IIiZ9J4EDva/6hWAOr/5tZSeKTfwjyCnGiau9VB5v79t7Sn1CLRRTsgTeU0dU1rKGCeLTFaobkVA
ma7JxDJi2Hqiqi+hStiyGuumZvtcIBSWDHVBn8ZgCm5x8mF8/3ovNXpX7bq4tU5xg5bysgt6KSET
PHZaNHy3I7YUqqu/F2VCHkC2KZxzZ+Pe1lJ8/aUgdAHs7gCdTVs5nheIZkfCm0mfSy/dGSRKGYfd
rVrWTcnorwQK5W13MhXesJOhG6QKvGfjoclIr3gxqDeBo0BmR4gFR5UA/BE4RlnC4kOda25m5Yi8
ulTgZBTISvtzAoh6abtYpRq48JVsUtTGk1+YSzOmhZLJkG4QT+UL6+JVgSQX/IDJ511sTQa4tjD3
G0+4bd7K8aK7dhHKKLwHDkjjVef9nlzawqULWtXJz9X4UsRjZqVQ7baOInBhDO94zkxLzmaYAdDg
co6wMP/Zvs6wyJ9xPi8IBqWNrF1H2PKb96yrMktcAE1QjmXWbKc2Rf+DeLYVBHgxNRnruYVmYG37
eY3Rdd/pZ1iYBVxZ3et/MYmKExHcUWcgN8Q53vlsTfoTVJOokMJ4YPmmWgT9eJuT1btQ7l/7tLVf
3DelZ25VQ/htD4vcAAa8cJLpZl5czVHiswio7wcx0GyGHGp5jS4t6eNRUsaBYsUjf1z7xYAirWlO
1T954a/4tWxbD7aZRQl6lxpWeJ6ugQX06tT1AeAv4buX3acHGPnvfSY25vPX13ZvLfFRvs2BUbTy
+iLmTRTgVgFYvhem1EYucCvlchCTPVbGAiWMfoi/TipNS5WsxupAHHG1b6u9OpRDnPb5/mhjUMQI
kgCcjRx2556AA7Fbgb8MZe92II17iU0BwPUCn0tJ9xiPp6t6ZdlFuxEeJ7KHOlreiv6qCVaUBgtf
CHcQnFJhwi6V7JEzJsJLYr6KonfBJd3R3ErXq8kBVQnI/CHfeoD+qFAZYds1/cBRqOVG2WurQ4g7
21dh62kda414fPuZFeTXkFhhEmY+d71gyNld4VmpxsMmgd8tQoPP1QwebDnWHlbl40p+Bsi+8NP/
FKdD3Xm8jvwgEg5Ldjspr6cn6+WtUcoQtoT13jquV17Ciiqv9Lu/WoeF5A6gK2Lp51E+9L3/fhAF
qFWTejA4sE6u/sRNnxkCtErLktjDBBncNXNS8BSnwQRYDwr0sn9p/UlyqNOH9bhV2fsIHr8af+Qs
O5Dp80l5rP91PQAmcLk+XmtpzGuuiSE9c3TFIGaaI7JCnrAh0RSHpIK5EmxpnfSKlJ/iOR7hAcn5
tHYuTUDZNriRHneSF2UCVmr3byOUg6k81tieoQqBNN6LLAgwwTf+MHxpMJDG8P1huJGrTD/T8+Qm
zKRS2RnbJERzgJDvkkPhIlN0//MOmr8NOIcbPSgw20GFLe+vDMCBPj42cfwXTy4f2Wc77+8VHGHL
G4GdaOUzBk4+X9cWouHjjiSNDNVX0dGJBX8VDChsSOD8rCWyo8OgWGEh04SPhq1er+6nvBctFvhF
EoBkFyGbcA77jWbOLdfiw/KUgqExgyI5vlXYzzl5lgdjL4gLMJiFAXJfaPEB20ctfumBTpOamigm
xCiVtnRwta17hUFiOw2UeaXLo9JH/DKxqLsMHZY5RbRG2oTFJIK/halWOIuRVeL/dCAvopwmDt+D
+Ja56gSlJuucksXxedVi2Fimx39uq9Suq1HkobI0CeT8E9JrTN1nO1ntEsLWA7SrAVSyZv1fHsJH
au4VkqYVvimn1h29sI1L6x3PpHsTTbogKE6ak7a72Xx/CupkBADaa7EzAXD4QA6NJKtKsTdpkFo5
AD0AxGFgRrjPAjufsr9zVLmhhxWfde8wFZVc0PCMbSdFXJXzBpXtKbuoWC/itC6XKlniAyHQNVJz
MrdYFc1Y2SCPrjA7Ql7W5MmuT2oaKWhft5+yMcQeFLeOXCJpk9lIOf/3r20X6SmeH9o/puEe5TZa
Tgz19ogJ5F6p4bBAbs2Kiy+S71HBRvR9PdsKEdThzNmsOS5yQ9ed6bguSk0QEudlcrXksZ2aXR+r
ynzJ58OLOlabGYIkXJQu/6Vxie8a9Mm5BcTl6yEI7qtJKqciHBj+YYYD+W89sxq5ibNoakjdqyOC
6nBgbKNt13e9XMQ+qEGqX37Zf3XobAZWrQI+n/ECCs1yubHwQJbvWkPJb5sMFwx0h3fNinATpMKk
OeG3OO6sft617KRSXWqDbgR9mU/rbDvrTfBM0V9jBe8lxxR0iwLxkOoTqB+Y4KSalwapX/i27wau
nGVCogwLSIZklcCmSZuOzziHDLUfap/CU4xd0yeEWnLgyXsNEkz+rxIYarv8VZ0k1ZpjGxfyD3JH
0PCyu1uwZItzDf4HAMsZEF8jR0nrl+WHAwqPDqjl/nQ30ruFeIjk68TgrcDeGTd7i9qZ8YLZEeCL
RBgVrY5nYDOs7cqmyFTPGJh89mQLWPYVOfb5vMtbllj/maDd4LGFS3z46LwlB38hJIoodtgd7Eqh
morWH1buvL9wxr8fQrVeaTdClU70roI3aW0CK3+Z1uAdP6ISokhB1U2SVKIxYTQf9zjjCvdOgC5M
FAAX1ap3EgzHhOjns7GlDBPSW1Ps9xR0hG9yfJzrRTiZ1ChYkVwvrpGT7oEOgU+uHdux73slgf2A
l10O//sJwum6H8VZEz4y5EAp7lTCD6uebGFLp7/4uU3j+ngKuC5TSUVkJ+jkjuyR1Mqlb8t3Rj40
Y5H/Q0g2NouBdomjVZ3qtgbX6VlZ8gk6cEgrL5xspn8/iXuzcpXQG3x9rqm3CWSCzpQeghoPiBSr
7VLqshqh3CnLpuZQeoCASyRgUNg84Ivpzbt+TsEchZbTZwQInthSZrdzvjyclN0wPIbd5GpMfreO
NEcr/BH/tOUfmzO9pLJfSIQIv/cjJcBfY3oZWBiOiPQR5nRBxKQHzjlvX3AwcWwuDUN+zKlPzVyP
2fNRMNgQJPFbQDDxron7Cyn30Pn8tcJtebRip74G8VUjimQQdP1YaxWv8n1v1A5WMb80Cn7jbznC
I0yilghNnZbUwjS+EUoqn76tr9wWGOedUcr1vVBkSfagCfh8yVTAcAqn6O0xqFylN662DO4itEbB
qXPZ6hqMMnYHO5hl+TAY8YYaOWGLau80eyysYH+PcQfhXAB3pJmutDt8crRDR0I0p/o35/AwyIJ1
9TM3Ys21xLzGc10S0splujmK1ErGOIvbVqUlNcaUCBsptz3TL0PvC+sKCkLkGfuYWiJUsINTbIqY
7t/aNxzW5kHei/uJTFzmYlVmwltNwqFEnfUoDWuKHDeAUt3RFl52qJq4YVHgvSv+0Is7YVwBouI9
XU3RR5ZMzVAf3cdCBQUwIp875wfXRjUywV1Ffp89CwwxbQFWQnCf0NN2CCxOfTlRzzAZqhKVme6H
BbSLbK6qoN+3SaahU2al4p9FSYKXrBB00mdtEZX3S4p3YOzDm5FlmZdzRUzUCoogkZX42thw8tM1
E+OemdRuCxtVRrmYsmze/9hTGZfU2sbzM7wAOHSwKeVWExnPJox6Zyu2UDRpMc2Kve5KnjuMg2VC
jm2Eb5cHCyYNnxw2dTRHqzyZ6+OOriXr6joQA/G4i0V9CxKlIInJWdhOEixXwGD2mob3Yv8fRI3Y
bMjrwdAGo8BAm9IkX6j6PC9pVuMkMjbslvGShzgDebduPXkirSwuIYuYW8WwZQI8aoN4wTSSW3m6
8eownol7p2AsXM+Fo69YSkA0exWL4NO4A74z/rFYMP9mOAtmp1AcGG7hQsUyWVrr42/9EmCKtnWh
G/jdgDbJXmChtHP2w1zbToxZXFexsSuz6uPI8ESXScR6UYRsADE7w149HtWNlhIatglpdE20Q5kH
lK/5h6e/+aSz94F/ASr2LBmsr1XbxJGJLJ6QG5csFJrlUney3VuFjDanP0qzOGl5V5ypGBYoQYpI
EuFnrYJuTR+fG3iC0FAO1Bx974utHv8hzozi3iGZPhBHYGzOOdIOyPPT6tgUscbSoA9iulYfvCfr
ePvqT1Hjen9TljWllf1UwOuyITvpTS5rLWqFoPisveXn6Quq5aaeFsFawdcdjm2JHNe0pWTBPEOQ
wMKrDLVmVZGpoEACZ65ot9AWs1E8z+64FadsEsD8Un9FINqXWlPNek6Tf3KtG3pll0eRSRv6aagK
WBCEwmCyjzNdHmD2+wvIb1mo0yPCOfuboPjeGlHa4xlVu1izfQu3wq1xrkZVfAztZF5jGhd4E0yA
HSM3CeWONZQD+c1JePHklqDVAu6Y0bmdX/y2qgafBD/Rgpc27hZ6bjZgLrlZp9z0+7js8q/7m9OZ
5RZ4jYhzZXxXI9rPRy1PWJ0U3emh2Qhz753aOygiq3l0KrXGwNKCsIM7UtHUIvvp2c8463Lz/2f5
LqVYzJp6PQxOaVVjSvF5ixsxJgFcBy/eDOCY7vNT9MMiLBJ/sUJ+tXTyjMfghR8QFPgozTjZrU8/
ZpQ8yIxUPyNtuzDI4ldDfm0j/yQAt2S1aDXZrLPdggBlOz927rcjuWLupeZ3W429KQFMYGAoW1eb
Beei5C95Vp7wQm89hWUxRoSqNfv/62jZVSdtpr594rHLfgDEkKnO9BhF4PsT/rHXuP+iVDQSMwRY
e7PEy9ropSUD0DDsr3MaKo0A3WpXCTb9aVMo+NcRzW1RzWNWxJtKKWdrO5vm/VisD5N1HNCDdeS/
Ki+paeyHJV8bgZuylBh9B+Fz166Z2MHilse+is2fAG9FHfXnCHsARBqgUyyHqfP2LKEZdmTauwCB
vFRIU5y2ttdMugDjjAqcq4GEgHHQIHCE4kQ61CrqCzB5T9yvNpHsG8zuamR4tEHDBOLg1rmniGdM
mS/u4xNB+XWV5b6u5Mh/kfGwcpWf/jS8PjasBYVRGamim4td6zBTVRSDeblk78/fXgUm9omV5YmQ
C70fjMcnc3heDOTg3eUVFXCouCyo3FuYExV/wKsKq1Pk/XOC4pKr3qQfU1GXYBYo42QklwfcXZWI
m/dvRZykopA+6wN4XV9N/Jx8maCFifrrVWpciZX60rT0urukEwbHCFJlN2qPoLMr01mELljl+Tqd
7tMf9JZlGjC6UvSx4E0Lni8ovjRVMVJXK61N/tGVmc/C6mmS8zuqA5euJdcFFjrLLCa4FQaITFya
e3GhtA8WVXHLBd17Mrc6AXDv1+SwEnatBc76NivWRFBoOxPtYVZzBwIJ565xxcW0KxJrPsf/n7vm
evLDtoViEGpbUYkUqBuEMPYkTG5ZhdCxC2fo8bHuG3qzAejxg3A3LGYlBrvWWltD7ZHGPz0gIk84
lbR8JX46DFi44Xzx+WcFgf43Lhx7KGnWVPlrxsfnqNqajpsTlFh/suu5TbRSsIB047RbmDf8MYrK
lgDClGj1LhdN0mheIMMjcuzg4jDiXsvNAK89yiRXZJrRIYOR8l2lPJQzYdnICDgVFm2ZmnfRNNzb
S2Ubb9nbsHCeZ9JUvnrei4v4TdgWjjEVV4HHNeAfZ3KBRNumUYregWNFj2HKoTmfnMRiXHhs7a1d
yKIP8ytUSYXUJcv9iJxgFMbsipu56M9y4MTbIdXoasMfcIhQl5dIIyh2Y1dYVrK/+LNgycLDspzR
PeEkvcCBt6ptRtv3w9A8JXxOD9DCImjDs2q6DJ3ZwMfBEJ7CeRM9mXxdxSyr0tUS4c4VrvNdSk32
6jnAJjiMcpT6H+Kpu+wj0KLt9t0DLA6neT0SQO+ycWVWAYxZyFY7jmPsi4aGGiaLBvOL2Fc5nKvm
um46cbW6wmYV70jPBYTXkkOUeCRKg4qVaB/Wm8lWLvjJyHTEPtitwTDOToOJKAlBE6ZhFCuet5Xq
FsFCy6POoDb6tQxJy6iXVLm1oOOIlDkKyVfuN11cdFZ1eqZgVLdh+JJQO5nd4GH4J1EKFK+iekAl
rei2ZUw/uiUbFiOF4vFJ48bbCt1x6FZ/LD9RO7b/AFtue0nR1pboBrIZKBZKL7xe7PTgwmXR5pA2
IggNhPWU4f656FV/J2Q/PHkpgbY5Nx0CKcizcfU5TdMWsMLQiI65FO11iGSz98ilj1WtnO0E3n6d
664swBJaH8exzEDiNa88fcqd5F41RVttLUQgqaYRYOZMhiEunkocngOXNG40/yo4E+KKyx2bjjdw
Z5m97HMWCZCuenCUeNsR+AuHWHiHXLlxqUUNaT/qIoZUIVkjTJ7MfhliWzJIY2umhA0PZV9eysvC
B+rrHxMk63TqqYbqU8q3Z8JTo8B7gfKJUY/zvmovPmtESwngy8ni4nVNNBAGvwA3OZsP20kJPyiW
rX/q8DLalCPLOUPT7v8giUKInOKrMkZw0m9dZaF0uHYXM70A8LP/EY1QCY4v8IhwKLvkTOoquNSa
hq5YUzRMjwoJpYu7GumlOL++7sIqPjb7m6QiygF3gfvQHfXk1mUeAMX6OsStDzoXCN3MYcmNM9oc
6j25XCzhnce0MuWU7ygkDKYDjQ7eGtOvVdXmiKO5Z0R/irCdklwqV/mCnFXDAm1d200kZXDnPv6J
vnWbVkSdS9zy6uGSh1D5ytCw1NtbqDMlqTJh7Y66HhCxvYzfkG8sIh4OYF+uThCvo2ZiL+m15hdQ
sCjSTA11l+noXrcxixbxyx3kkQS4JOopAcnSxfIzzIan349oQqjPuc970qHePT2Qb23usgWpOjGd
zQbBPhIHqKTqbRePCXQhzBJ+2lbRrHZumGiyGcI1P1MCXldV3RJyFLGfQfaYedorMsyihre4eFjW
iZqhBlBJBsnmkFJ6WSmbbVKGQ+6O20/cXjYUP9yDuHRj5KfocVI2mEkAeE4r8Z5cHWUq1Z9JdCRe
x/HWgmE68Nw/DXwF6tbvHCPqlQ40E9A1UwgGVcoS01A07ctMoREIILL2fBCXxUcctRnm34B5cuv6
0v5jSfszPG4N4wpV46C5w8toozIOq313OtzSgj3Puk+HmAeeU5iaTUk75x53cRKSGKjqZ5xGEmd+
NiiTZ+Va+0C+qPNF4ppwREcJrcTU0A7FHYvacx9v7etbkEnO7/CZnpXGKEZd+ySh0Tbz78lwzm9L
dXEeYxmZ3cSXw3rxyJngpWaUf6udAw8rf6syKaKqYpD6z0XuExni3NZgmfNkpn73Xz+fU6j499JN
baPJ30rJrql5SZahrcBh9LyGny5iTUqDtwHoig5Ub7r5IFcnjmju6jL5D1wS/tJWaViNzLYoHqS8
Nv94yPV8cYYx7x+sjA597A6XjkyHmTYLBoN/AGWBNNN9GH/H6x86xz0q00B+ujH7v3AQoibyFrDs
qORRiNyYSOVAwkLZqVOnh9mKP84xmhQ211Ahmjgfk+GmZMA6NY27+OTGqBwhJT4BtgnM7wKbsLeb
Qr9G51ffCiwM4BHNZgOlf2iPN6nKMpcc5S0cJlANWnJLjq0543vheJhE45/iFMiVKsr+IXfpHcwn
aH4TK/FTvCswiCPPPZ5G7/qqzWjmrMQF9xU1eyrsqLNSSBSLUX73LgONbAThgi+DQGIh2xWgqKA1
LNRlri/j2mwe3JXOpJIzPH1gJx1HJuWs6zyBy3pNqyceR1a/mp7DMHtX1kPXjaMyosgBAm7cNFpu
xlkLzoHcLdvX34fZMOGiQIP6kt5VP9bEYFIhtw1dQwcAAFiBCmw8HNV1NTLvUAb7tIfjXYFN4mgD
0B1P2UVec93j1PhwPtWGbaImcO2aTxUfdr9yXrNUPBmBoLtFwrb9MAvKqaTxh8A49JDfy8xU4oVS
AyGdZOHjWy9+1bwirpvtv1RR/XxAWH/IuSnJJBacvmiyL/eR65dCK3GBVRDojo99gHp2D/VtATDz
dTzjraEllKkBCZ8feTxidIorSB7SeS0mWaRFFH6bo6ZpIa0gppoT0q89UfnqIdSQfH5G/zzXeYlq
2Ql860WahxW1axPI6By0ZubfzKjB3VfRA0h50q+lYxuZkizNDK2zhfeEOSk6bK0XhaSXvr/O7qS6
J9102QeKw5DQWXHK4Ux2x/KwpNLsXy/1oVv5OEY4RIy42eqostYQXP1DlFJXpFFU9Y8q51K/ieyL
US3OTXOHB32Tdb4Z+I2KKCcetoe3f0v0qGBvP3TvsRXvF2NNwxnC7bFNOBVwtfIG2dbaF+MH/BIA
tGZngxRYKV4JDuBmW02L5+utWfS8dbx04TSWb266LwVZ25qVHf9/edDw13qCf/YsFnPHSM1tuPzr
wnOGI6B9U1IackDfiONrbwL4RFpCqlypo+LHTV8sAhnxUqLX/ANcFwKyUmbPlp5XdkYx5p3BTVox
49zCSGT6zfZVzV3nYwMt7vhRmpexg/u2F0QLDSLm8nYmE+OX1rU1GChwl+EV0acIdwSC6I4DSEgI
MlQkr/7lw+13V17+P1bIy/6n1fKqfzwNkiJly+0MVIx/4HhUEyr5g9T7fd87rfc0J27xsIv5llEe
tCPUmTybq/GsDqb/v1QramQ2cxPaZhsAHPe2VjPnrg7Vpf8VT2mjAj7HpqyjmnDk19tvp8THugc6
d3y/qnj+W2BZ2NL7PPnhW6JgJpPyOQe/6O9qe6bXHVtkCdjs64uRyo69vCtosoJniRgMo+ecnjeB
E4xQHrBnlm4E90njaLBpHqjzhHOYtaXjnCGmrm4SDtPb6TYgT7R5MxkSZo4eHpca+hbyaaTfVVfS
9818DnBMa6tVqOL6yLNEpqYb3WgSZVSogBAnUun+xL+VJ7+v47WJ9OCVjCeRRyvaAozISCYfdSAi
kSTcYIPj1hZ1MtWn/7B7BumHNqkx1z8Tol7EIlwoW9jDnONuLdnFGeIxtWKmFHi+h7nN2Q5pXAXo
mv4HlYLBB+fJcPAnRZsSN7RlxiLIzTaXaJRI3ZYu+Zglh2cQZ7cF9Nf5bN6+QU1FF0Wbfx44FaeJ
6edPihaVi+zBWASw+TvUoycZ7Oa2H6BH4KEVEYFyf8AenNFYEZqYA2GEYrJE4i2smIJCFGjcoWbm
s207A6iIHMQIZMTyAUDfgrvU61kBeC7MpURZWWGVWeZPGFlC2pHZaBfO0DFVUznp3zcgfmRGfK/h
fAyGODIMIWLSthYtLkY5dozR5zw1juFOULmngN3A8cSM5wBRVzEpZr/PKvu0AZ7+skxCPlSWDvAf
afY/4oQ4IT5PKwdfVn1jQuNnvhHk55zk90yxuLHjnDOwUgpObDLn/gFxR0elmniB+C2ZgrWzOXWP
852Sl+Dz7qflTFuJSbLJx0Vsala5jtvfavRuHUlqfLUpd7GsRdNVjgRoq96KJxlfxNnBT0mytnKT
lU4ZyXlgzzkw4Od6SjUghVZfRRwW7eZFN/cvxGCUI+1/CdIbHbVKDNGE9EJKK9TzMO1eW/Ts7yt2
umE8q/JBLkvL1tvrRU3JxmHZ81ghIAMkVGWVC/1AomXlLH2j7h8Eb+rSDcF6WVyc6Ld+9StMdn91
JgL3I0k4TKroRHLw/oRKcHf20qyZCU1UQ46TzmPizVXR6SgkStZ5t/OxBcuvxeuKp9JM7avTNZUJ
6u0NVMReqvbV75FIuiYj0o6w5mgLOISZ+J22uYUaUBA59nFxO+J9Kc2KOpDvIle0vmdmiun/9ND1
C2i+J9+cQrU4VF2sHGauvUna/rnCyeSyfdI7boEoG/cdkO4DWI6cK6NWAJAPHCO3G4onssqkFRH4
aRCIsJ4FXZ2KHClHrKHqCYF58l07AOAosYVx6j4FUbnOF/bQiTQIuWVD/7anT707dsl5R++GhmXh
1ZHmTkIKuV49fpPxPBT6/h6BGBnwiu2DUQdVZQrF9b4TqncFjuNp0ijZmBUhv7Ikp6/wK26XZgTf
EOyieYRNq6bnk2viCaB2l3EnLK3//YwYbXgqhI2FvrIdFz7rJf+jMkhJyhmyUzecY7+6xKAURdpk
/VSzurJILE4MQWOxc2OmZRWEK2/I1jGY1hX2W5zowmbt0KM+7c3C6IORPNqj5nHfjrB0AV4R+9/q
8lNn3LUAmNvKz6VVPOEOSAk1DKGByzsk+zY/qp8XbcjLJBdwpfZKkGhjYL7D97NbEuLJvGKn1V4L
XYGozaEENO41uTq7H//yANrnmCDrr13eTjCBfgoUBTjhjoyX8xv5SXpSpynf5Bj9ATYhraHAtj8P
6WYh2TjsISj5AblQdnoztvEylIwgzv9CMQNIqSn6DIJZxXO35q+dnQQtxYN5KNmRe7nWvNCwjOFD
bl2vY5lwYbi1SONIOVQl5CsDhWeI/vSlXmeIMBUzF//bhcj/S9ec2iS97O5HxTbVZ8tGGSqBQkXx
BGia9vb68EB0/G0IIUe3FbY8kptu6UZjoUQgeQzTNfs7EzpEiwJDC3p2lNQ1nije/pHQjfhBVHkm
1OSBhY1y0TqInTRW6MQUftvHN/b9588ylRP6L7F/tr/IyH0pRFLrjaXXRRVtZfCclaRLq2yfkbX9
N+mncHM58/hAmsK2gXN3ffs65Ox/Sa3ylHtl1HNi7U/oAqYoi4nqWTofenxApw06KK1OVY1sesH9
UWuFauvA+VLfnMe3lXuZDsw/hU4jQBfGBE93XfqWAFQZ4T2jf3G65z6msoJfjV/CpjrDlsSk6UP6
3ue6YoAU1WcswoHDcU+cZwaUwqAccP0+BeDsJsMNxMiMw1aRwH1p6vyE+zsYA3Ah7cq/FyWlLJO5
l20jrQOmOEONjv8O/TBJfDX/rlOHpgkAwPVw47V/LDmTfG/1bXcilN0q8neHmV1AQyE1B97sbsc5
gVhasbJ5E6c+M1djYdRpXg2mQVuGBWjT4ORoPDty2/HS/k7UreF5zmc2ajHcVdI/tewP23nGY7jq
fobXVsUOWJvJRYAT9U53ABE+c431aK+Po7YLVdZz7TogO6aeQ2HmhC+DcZiq4s8MTPZxWvNVt3qa
vXAmkVEB4sjEuAfA38xc5q4vQcPWlMbcsWaTkzzjPTrAyFNs8bKyrOSIcrUWPjkuI8JjyaVX+MMq
5fvoPM+BZxTwEBv/DMVOpmMCAQqX+TuVjh5MTgst0B1UL7L9+tBePqLcdMA3JahLf7s1zXWqDR6g
NORPtpAhEXPt+8BtF6HiVDVQoZNEyTVUp0igp93SeTdv2J2jtySfOo5Mm58v4SSQUhzrfmEeDLuh
/qhmNC4IuhD+fxR+4lCqXgReP1LixZn9DENuZNl4VhswuS6sjjfkUfCMQTzIL8tEMluUGLxj+z5p
TrJ/CfB3Ja+8FXC/Wy+b5f9EV+VQ73HnO8o2JofVKLX0q7OD+6vm964hXiXIlrXrzh1HOUn0E3pN
CwoTLm6v4qAqkWgtQk53XDGRt/gl9ts3lKyy9BR7+OwsSU4nMR8dqgYFzTPycsym5Gn15OgyoMtY
mrKFtGdIzn/une2lx2mO5lX7LtQRXDLLaNEgjnh2ENZvJaNb5/0pKm3pzgqMQQpBqCmYIWy4hVL/
MKVVPVtwUXwGSwHjYmSupSLvSC/uFIWykraGSZ3LqKLmEKkIpAQvYzW1dys+tqFrAKWgw9HD6Bw/
Vi2DO1mxxL51YK0VxbM/lkGCe7zvuIRSh2xr9hBQNWFS90rdOQNL16OCvhbGDMwP41wNOeJtMNSI
ORY/Yp4Ck3UVM1ZOOwi53VvTJtp35sxd+k/xg/zkOM9x4DvvIVAVfWBBWzlwTNGBTN1dHAMOsQFU
XsqA+6kHmf6OI+R9mjHG6s6fclTW6c+tCbe9NA4p/q0TKXqHa5TdRCj7et2OrmmXlvyEDvB8BeSM
yGZykzGsnNg3NlDq7VGlV+Mv8xM0qkke4a/DNHmGixjv1fsZ4dLwYnaPZ7BJX+sHLx7iYdu+SZsH
NM8uuiqbcujJWdUK+5Koe8zJW82aoS1J1OJ0GBqyZUid7zNx01Q2q98XoJzEO0sbAz83BrmkJiKM
dSW8fEokTdYKVPbIrhQ5Cw3+0rD7X1Py2b/CjkAZtojJRecHiUnx+yvdXUsscVm5yWr2KZoRm/ar
W3jpy0PanVSJJUVyHlbwnCoUOrVdHfPm3s60tuc/qCQzrvgn6dSNN/OymI+ACQBn54ZOTA2AnX0r
MK1zTCdyJtd4UWzBj8dRiTq+RFuJfJtWFDPVQt5YowXcUF+LU7/ErAZ43jjlw1Ah3HItaEGSaPCh
TN1nd5SVjLtQCUFoHi4sqjWW9mvrNGZ4IuYmERNg3LiOYNrsrWTJNQBdp/9CUhUONJ2vc+5ZeLdW
vMxLI1pmQ8jrJOOg8ZheMhCmXJaIk6Y5NJdh+k4Udkl8oBrLsrHSk/zlo6fFRZLJzZDrnMatVZss
ESi72loehBpDeXPZfzbPaIaxWG1lx1PB2tiGgAh/R7aQh/5e7khBwh/9kXNYUXwZ0YmvZPEfdvN7
Rxx5huraGWUU8FatW6C2hBdSMJG+MZPyqYDGNmhv8xcfsJULmViL1eCtMP20Xg25gIu3iAcVvS7P
NLqYiVijmX7CkxhvxJv6dz4qn7YzVFqk9p7k0wEhIYDCBzjFAeZbdN3cngUXqncHvxO+46tVxzzc
QN21q4J3VPDseXQdUQIDHUOGwGXRmERbwRphYhc5xxrLrTe+0F2ibB7Rbu1fbBv6KIwCuT/hD2az
xc5pDrlESKII26Tn8GtRFkaM93IbbrZlDMBPJ5KLzTSo8Xh1YqaHeSNid2vvMQcSMzbYzbtHHQDb
HFNb9CC2x6EfgQP1nJtkqoK6EVp7CsnmhhlprLshkzarChooLbZo0mm8nFnVqvcRzXpphiLFQjj5
LjkUs5ozGeDjctVDEKnc4JV22+mNj3PJYpBXz6fICAuj1edevo3ogSj+9J0U2WCIebCydCn59/hc
V9p3zF3++QxdnDEFOQ2lLwZVX8nPoniBBBvU8XWThgEuUQfX7FQ26aGhQeZAFJ5kPB4fkLFsbIQY
QXl5p4eUkvqewRBX/5nkYTvlE/DPCD2M/fYQWQEV0byGSR9UZMn/VBmaGjXySUJCaTkiUJUsSttW
/fIR42piWAkNG/Qa0n1UdMqyEJ4Bwt+Ln9/8iNMtE7/+8bLT+RaTg5CnT2fOXcTAIsS6BnQk0S9h
nUDxUEAn3XghcXb/5V4Q8k57Lav51E4Jou0ezol4ZSPeYWvDP3D74DjG0E4gvE0MuEmnV3O00e+2
hzp7Wcb+8ySA16wxHktvZ7P/UCWzCGY4xVVDQ/a8pcBBg8meRskGeQ+BSGEW94FT1/GNkTFcyLCN
KciaYZHT2cjVvPEROOqKPh6fICEAbEKf7srWn76gpw2xRlj79xTmu/X//QnHNwxuJ18hqIGr0gtf
ZUwg3bZh0RMis3puua5O/+PzFWAMp364TEdRkgNhgVVZz675BVjaBn9py84KnWJXoSl9MWdRBcC6
ylJhG5okNQeYl3eAmnAfSH+UtYK5Pmwvx+Et3Mo7FwJDopGUXuNZwzBLtZvwCI5+9VK4Qn7DpIPU
ld7D1ufhZ57TlBS6cQjgo0cJkWNOWnS4RvzxdUYCI9V45936QNIXdziOTaNP2Dst+ozK8W2OXbJ/
cr5KAp/1MOQmyWbXP5f9oyuWO9C2ZuFg+ysN0P7QwurObTvGgXq6tJEwPW6aJ6Ip83CoWSt7cS9z
7EmMiyZehGd0He0AG0auTfdaLwGkg4rGE2wXCPH9MdQxA6o2uOYFi7jrOOar7/5ler/ZQTARtR30
SbBRkddBwCDYf/4Vq/XWBy/EOqtA5Fbltfq1GA3GlksTQs3ZS0EvT7ax0HDYdrTQ7r8n8dlJa+oW
tRAqILNlGUWnVpHh7AQwbiMj33xFUJEa3EWczSE0D9VHnuJ6I2ZrNaethBxMr/P800aNsqUHmIHZ
fBdMgYOTOWiki6/oL3nOISx9XWD4fELLl5q8IbLAm9XGrSzCvEV2NnLqqn3Qo4OGYnwJvagdAhy5
MxzPqMw5O0s3L6qWP7V6nWrtnud4VZDCeBZ3wMF12CPyGFugm8sjhHRT1jRQnQB6uXggxlXV5Evm
gK4XWE5vHohGg7HWqM2Mz9bfIig3YhND8rWIgynSvNCsiOA4yBIhePUA6zKZC6Jr9c295LBdPg2P
V/mw1o6F/lzv0egcmccGOgh96MXqRpX25tcshgM+kX6OlIJ4TjcsRqZkS4xC/5uEYJaV/uuz8dJk
STCPXT8p4TanXCfFvyfj8OnSbeMSSdNesFZTaoYPxOSNUADLsi4UsUhrhkQF3WlQH/j73+q3qgms
VXI10HUvDH9yUtJycezApGmTMJFImdwpaTuGMkoBLZyKxOzqmMj5onIxBd2h941Rm2BUqxewuEPt
tSHEU7/I7Q/hixJQNw9KdhKOciTVfG19+47FXNWWbJcQiL7M/6lE8ey6XNfiPDlvISmeiVmpPb/s
gkezzREwRW4TXaCb3+4nLGHCR7OBWo3BWdmeYjlw5kPNbjTOPaOMd00/IC8BUU0tL+PS2qTE2cKY
bTWJhxMfrcku/XAe1W2o7OtYu2/MIIDFmgsU8T0XqK1+509srZl83LofM2smYmEITPBNoSx3VCKy
s7CaSCRAsPJZlNuA5stjZahxGmuN/oX9IGwkRTkBNVs6yecZfFUtKEkD6FEJxLaSmmKf8ZHC0GBK
reDf3t9qLTZXt2Viv0ZKrAsZEARidp/MBy5mCYGImWSfI7YRCpN/soWpop+w6RZiI3UYmvTwOxfQ
64Ln8iFtUrRHdSzMjBqJpyKUc5xUAIsNm7y8eRU5DIlCdhhO2CIGokN8kbwieOgDjjjyobA+tu0x
6J+r2l3eGj8u35pq1RWB4nOqwrg6x0H1aElC6Y+Jk0iS3oGLhM6e7FSS2NODFiTMuiYH+eqEx6g3
ihTH+0+P5SNbAxAYSmaQk5hf5dNKi+io/n8B2U8=
`protect end_protected
