��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3���K�U�h�/��������6���0H��ŀ�N+
�\M�=!�*J盝�l�eQ��Tws�94�m;�>�4�eONG�!�ĕ[�\@��X���P��G�n��K����o%�{�f-a�E� ;���1}>����*#XQ�V.�E��h߷��4 ]Lw\��+o?kì���),5BG]�G/� j:g0��,�����a�]�'+��)��9���T+���wwXcV��c�w�A�F@G��*6'�G��1~A�C��v��a1 ���XI ���$���n/�1��� ����Ã�o��yk#N���wCHIB��G���s�4�����#(�K��|yS��)J*{�ݴ��}���iq�h#��
̄7��|����QY�ϵX���[���3�&�Fhwd��� .ɨмW��`�C��4� {7���k�9� 7�*@�Ki-�eބ����c���*���-g�CHCl�U�E�ד�Sr �ؒ1~!E�T���O��Ж��X�KI��f�S��J�V#萾;������uC����x��rdo�>�f���c��@m�\�_�-�wQ\e?�LbMv(�o7˛|O�g����"��R��P���(��r�Q����J͠��7��9=�Q�A��h�����爰�FiO�lX����H��0�u2����^�����vA:�r�5YZ!FV^7z�xT�C�Z�@�[چ'MR��͙�H���. �0������we���4}��X�A$fg�Mf�S{Ia4G ��3>g�L۴:�D!����99����^�S�T�\�PR$���q�dZ��S�Չғ�A�	��ϡ���p:��Vl���ȖK�ׂ�m�����p^R�[p��CH�̆��|@?��PAb��G��kbrwas�q�|,<����ADl�{��q,���~������i����F@����>�7ߑ䅷CgcAvK���&_�q��>��Cì�`H���>��3OA>+y��^>���>��袹v�љ��WP�ަU��X¤���i�r��~�����n�SaY���t��Z���E��sA[�-��z���.�$���/���e���}|�&p��w{��<�d�;��aȏ����\�}�|��d�{�\_��³4'�0jZ��U��5�.��Z��~l�42�����¤y��k=Y�˝ }��~f*`�>�ĒzA(=�/�����I�tp��ک�y��Ԁ	��󇈕�,��k�؝�qP���6_2(�;�CȜ��݁ Z���!L��1K��?_�dS��/�i)���Alhx�r/N�|^�F$F>#�}���wC����P���3F�A/j�t�:�`�v�gP�'���,�E����l:�kH�Q����R�q�	��E��G��J��z�'H�B�4\`�B���K:@��%�)�gJ7"��m�{��<��)܊�=� ��|%!����\��CI �)U�P4v�$ؙ�?e��ni�W��un3Ѣ�B;\Su}��
��:�K�τ�N��⛼��J�L-
ٖO�Y�d��@a�k���=j<ۯ����O�~Q,�9��D���E�T�5���(O�w~�� !M���(�~���s)۹�\<�HPF��~�l��f@7��6��]�� ��VQ�C��!=X���.c�I�N��+��'9α�'��%�7��,U,2���i�r!y�c$I(ۣ���ki�&Q֯Q��SJ>��9�G�v�Ӱ2d//j�P���������X3�K�qOW�"�Ub��� ��F�����	���e5s�d��5����-����Ψ�R�]go�#�w�^�q$vI�c?s4���8dm�⳦�����u˝Y=s��Д?	��6�ܼ�ɱm&�h���uP����P1
�,���Sj���N�ͬ �����v�q�H�4��݇�Y/����<!fݚ�~S�%��i98��m�L8��hU*�f���-R���)�w#��7��·+Xt���=�X�.RO��%�'�MR�U��c�����Z:��&�̈S�~��;�.�b��[о�R¦(�15~�زLO�yg��	�:�"������7b�TW��ȄĦU��idz�b�*��K��5�Ɯ��>Jg�hpv%�7��Wv�;��[3H ���*��!�y�KַY�,?���d������h{T�4 4])������1~{Vᝯ[�-V�GKp����k5�	x���[O��4��_�ʚ�n�\p2HDr�ǃ� 4�����'�u��#˥��8N�* 	�7"����Pv2bW5��@�
3�n����p�����/(�~R��x�1f)D���������21�H��p@�����`嗹�+�'��2��M��_��4�/�Fesb��e9oXq��� ��$�zKK�����*̓�7I/�8�滉�X+���*?V�2	x�h�ٍ�1�z�]��N˜�]���V9F�Dm�w��wn�f䴴�Ż|�4mف��򩠋Ac'�T^��JtR�y�kax��C�o�q�k�9�m�m4���/������׋� ������5�����Tl�k�}�n1����C��H/�d���U ⴄU}%����N3�=د9�1D��\��� ������Q�A��~�₲L�̻�nf�
.��p��/�� �{�=pL� m�=��^��9b����!���X�2,�qQ��܉�N���*.�Pcm�zІ�? Xo6�qls��*�κ�y{�����9�)NV㩋e�g�X�	g,�*�B�ܧ��ڽ��zl�O
����~M�����A�k��M���x��)���K�����B̎�k{U�L��!<æ�8?������=�>9�-�R�Si��<Y�q+���Ba�S��sL<��x/M�zD��+x��G���x�]BE2��ެ�}�kj�;͓�K��-�A����#�����j�.F�X�=��wA�d�$��"�R��q�tá_����Br��x��1�&j������Bn9�6kŰ��¹���i#��i���hOJ��c_����'�*`m�(r�3��Y=Y��*>Cˈ?��� �~N�EA��5?�3m�g�5w-�L�ؕ%U�B�nSX��[���o�1�g�wN���-�g��A&	i0��NiJ��?~_sꬒhu�hH�-�f� <A�CT�����p��FҚ��]-���C����)IuӶ�6�� ��m�]����B��ZM���̓�K/�A���v���}�sdY���I^���'fEmmi{7g$6�<Ț�A��)�{J�G=��Ԥr� ���a
!�_LE_�9��b籤��P�6K32,��U_�#" kD�`G��&n��ڹ��.a����.C"hX*GeB*}�ʌ֤n6�S:F���b΋���3�#<⟌���(�z:�Cd�kРvѢ��x���D���y\�g؁
�� '�����!LF���ͱ�w}-[Z}��D���"�ikK�|��j(k#��^�z�s�/�0e�Z��}��N;&���N1���_����Ė�Cy�9�-� ���&%�Ԡ
,�ى��j�55N�)�c�Rhe�2��� n���j	��a��$�vڵ����U����k8Jc��V�9|����4����9 Tƒ�g\A���	�ٜ{[�mFx\����J���h~��t4-�j��3�q�Ҕ9�)����1&���������D���~�G~�P꿸�y�5^���!���у������gt�F�,�,v�!GҦ� �!�֎���2��j�!Dﶿ�>,8X��m.��}�&C!Z��t��7��Jb����ɩ^��]�$Y����1ent����?��l2Wx�~W+Lp���O`=C74z)1�~Gj
�����Nٶz����v��:_���Z�L1_C7]��Y���Z���~mI�z��s�k�Ob@�TM��=
�94K@6z��0�ے����((OxP[˚xԄ^�W���e��o���^�6�G5� ,<������d�j�w�McH�ZG����A����^%&M��Y�������.w]���\��iD�6�F��p���[�*�8��5r���r{/�
�@�lR�I	�|��~���"P]$��r�Ơl�f>��&H`(.86�4�7.m7�#T^r� ��"U����n���+`��4�Oda~?Q�j�1L,����Bd9p��PG�B�$!r� ����n�[6��)x�_�b�o%q&)y�H�M��ޡ��~H��ŏWo��l�־����A�d����r��D�h�m��W4���-��x�J(̫i�ט5��f��z�R�(rr��������7�~.�����̫1���	����	sI�,��zrm���_�X nt�B��I(�H��MC'{�KE4���N��D�6@�&���ū�諞�1Z�7�;��:�+Tc�I2�~��~P�b.��ޘJ��ܫ9���~��|�3��'։��	�����.D1��S���ſ#�,V�La���E��ӡ�!��������мK����O�R�]�WR^FG���6���U���e��A8͘y�e{�:QN���2��]�5������y�Vp��{k{���K��W�z�JE�-5m�Q�������v��j��{Ϗ;�������M*�"���F�dˁ���ߴ�T��W�Ԫ:��L��wX}\�-ɕU��r��@��+]�ӴQo{g�t�h$25�>X��7�����z ��k���OW�@��&C9�>=�j�[>s��4�����K�yl�r�ޢ� ��,s�do2��ű�=��j`$���|�Rs`V;��� ��eA�Y��|,�:hPF��b��W�s9iJ�:+�`�p/�����=�	,(�Bj���Xz��x��S.Hȗ�౵���>��;ڕD� ��~!�#o�q#í��6���ۅ�^H���I��K�}����YO3�NN�b���=�w���z}��ʙ��B���JJ�R�J��\��T�g�&���dQ酜�];�c7��	I2���W��6a.G�إZ��}Q'�gG'5�V���M�/,�=w����VoY6$��|��=����>��[R��H{�v��H��&�:9��+�Z��z^�M׈ J��q�"G��d��F��)�
Nڨ�jut�P�t�SɅd��RH�(OWv_��3N���[�;$���9�(�x.0�e:{����^��7Q��K�W���J7��\edg�pj�^�Rt�U2�{�����e����M���?&��V:�cK���/]	̉D,Q��m�����Җ�n�ى��y�X0"nyu����I)(&[��UMQ=��U]�8�"�OEl�蹌�;V�O��@L7s�����~E}ƔA|t��}�0��#flp��������f���?�gK��h�`�!o������:���������~έc�����& P��6�o�QOc`����}p<�E�݇vg��(���Vl��*���Hī>l}�+'��/s
��tK�7��յ6���h��5��aU+�T��|nw��֜)
�+�6��$�65�C=����t����8 �}�ڰ��� �<�rˏKK.�ܷ�s���Vp�'K2zG���%������ˁ�6���kW�O�O*b�sUI\��7wse͈���5ݧ��y�ؾ�pպu�ռL��W�H���������J���V����?"'p�`SE���m��&���h�Ε��m�̼���篚��/M/�}�+3�W�����_l�E(�+��ɼd�f<�ru;�?¥�n����׾��1�R9�O@��/	u�"�)�Z���J/x6jRR�
�җ�4���7�	#�0f�D c��b���Ѽ u��d�:,�S�r^�>��l��/K��ӹ���b;ʉ\�9���$���}-�������E�?��<�+A�ƗS?  �i���"�1�����d���M����6߱�TN���ȸ��U����`���y�*/ᤪD� �pS�t��%�j#j�n	Cj�9H�ڟ��1�٘A��t{8��=+^c��5B|��2���S5�w=�#�ח�7�Z�1�m&e��!�-�	V'��C|�6��P������
����|Go���1�w��*qw�Ȅ��6^/�%�s<�U�I�#X�K|��8_tl&-x��z�0jUk��)����e��Ғ4J��s�gT��K�oZ�X�ɾR,j\��li��y�5\Զ����.]]��ȶ���̥�,�\�EN���fR���:����Q���zoo���!8�.rvi�u(�nE��ݮ�Hrf��P�a��n�R5�Y�G��T�\���+��i!���Q%E!��N�M��߳�T+roye�Ҧ�S��e>q�]�̌����o�6��RN1�>��o[��\�H7����`/@8�ӄ7l�]DKN��_U������Lmw�c0��t�"
amU�X�#�٦|t��_�~t
7c����옕\%b;#�/瘈�T9bHz�kڄq����?��-�ߝs�ecKѠ8����QƊ�ÎPQ��AO~$][�࡙z��6��$�rG�(�GD	&�%de F�����N�ٜ�]��؏d1�[���$���N9��<��o�����ˏ����*�So�%��sk�f _DKɠ��������QgT�rY�	��I&�&�ͷс�?ȳS�(�[��מv3���v_�nђ��d���]�����v��eM�� �Z�r���L9Yd��̡���CQ#�u��:7:��O��ХS�z�)I�EwH��H���%2���g� }
2~���lpHP6��tEJ}�X'�P�@�j�����=n�1������������1�[��(����^:#E�u2
���W����	��+U�B�B�j�<����i�4J:�U��}�|��F�2D 5���H�Oz����1�@�_�Jm��R4ږ'��$ތڄ��[iE���=2����[*�&�ʵD�=ѶK��4X�tH�Ԟ�{�#����3*EPZq��ͧS�&7��,J3��FŌ�K9V�x�&�vk�f]0���~����.Q�H����H���;Vߗr$Ȩ�,Rj ���餛�����h���6��m����"U�]����Y,Ef�4��g�U�1���@Sj5�6����H A@�D�J� ��37 �c��.HxSB����Z��7���#��)�\�Z LKY�����\�lI��4oEm.�-h��,�l�I������PaaҴ��:��0.3Ku�{��%�锳�?��8/BOsm���x��H��g���~�G��{�_��'jh�N\�Q��A��B Q��4�A�i��V�7���0�W�O3oi�h�j�W�CA
�@�������[J�?�����I�eb����c6�'~t��zc�*8�b� ��m��۟�<��r�i�/{?b�&��o��Թ5nPhL�}���u���p�RչQP���jף��Н >�Xk�W���2�n��Ո�g�\"��*zѕԳ�Tlo��{
{'��5�
>�
�<��~s�կ��m2�TY~Xc7gTY�9�i�_P��Q���F�#���a�_�0�#��`�v�Ɉ���ɾ?�m(ˮ�N�[�.��QQ�-�����c�sե[���qǲ���!8��P�b���鬺n��a`d�l����b����CCu%����*��M�Zٝ�-㧥�&�"ԗ���>�Z�U��3��?Y�j�V�����9�9�E#�T/�^Ȕ�ߥ)@���5̋�xӚ�ѫR�&��k�RTq�?�5~����䔤��W�Y��ku4+��Z+�Ċ���cԑL��0��$MW�Sܜ����s�7�����@�[��MKA�iVE
�@�V�\��cgs`^aB>�&oj2��l>E/��:ED,�l��u5���!_Nċj���l�ɿ1�YYN8k�T��^����0���6��u���W0}��or��/��h�Xѧ'9��\��x�}�$�(����Tq^6?O�	�>�sPg�G��;~.f?����9o������a���!90Wu��.о�g����z W�M!�7�F%�1�Hc���틣��l�����[NE9���R�;K
+���z��,�%ye��+�?:��2u�A���4��0O�%1��	��Z���er���ٌ���Ğ>�\� X^�4�}�P���Q�_C� Ĉ�N��$/b�eжҰ�;`P���7O��~Ē�z40�u�+����",��^�:��x�*�Rc�]�@n� ��ޱ^�QS���5��W�:�<�)`��n�׺�ȝ���hAI��C��w���aV���۬�?��(c��#>Lx�Jq���qi���  �t��H���{��te��'��h�����\67yv���-�ʘ5�!�^V�/
��N��VT��h!��єD��v_2���/	֙�A_w��-����j�a��H��f q;�vD������/�Z,̈́�)FW�:S�3�����F~�/���M�*3�bn�n��P+$t�۪m��VСH��_�S ;��Ƃ#�/��N,M�T5��~kw�iw�M@�<X.!��6�Me���J[��I%�{�h'��J��Q�;��s;�I�8��Sr'}?��C�,��3H<n�j��|WMm�H�&+{��\��B<3�ų���v$)���H��i��0�PR;�=L�������L���}xV�of��Gy\8\�t�M�2��(�Qs� �Bb��$�r���W�,���VT�~_�zS>0�)�Ct��b��s��8�2߸���5BZ�d�0�U:�'9��W���)B@7a��b\��MQ���I�gZ(�R�]�M�����з���h��+vF�0����Xd���fwX�{?���D�"��\}��A�����f��,g��$��G�߮�-�%��¦*<L�Yዣ7{�`�4�m�٦�"�.j���>�gG0����S��E/h�W��̺ùy�.0�*Ip]J�"�u;ѕ�<s�����=�F��{�}Iwt�X�70tl�;����Z�Z8۩��xnu>���u#�Q����y8�ߒȩD��	vJ_;�M��hS��@��dɉ0�{��N�?�9X�Tq�A*�m�?�ܧ5h�Y�*XݒV�i*�쬣��@�K���S��F��k����L�3��+��;�����\eD��O[d�~�Jj=G��D'^��hrXCQ�����tY���ǩ�a�
	��
Ɇ��_ې��CE `�ӭ����Z�z�A8��#��Th�$�ᕀ����RO�c��4%�8��
�Ǵ(���B�������Ȃ5s�������,嶺v��$汃�B�r<%�㙨V�NP�x	���#���Z�	gtō#�}�S����Џf� ]�m<0F�ꆂ�m�`����O���M!��&Ҵ�&���~3 ��f�g{�o��dp��v�W�l��^��m���r�!�M)�>NJ���@O?"���з�� ��Q�A�Y�`�����M�B�;�q�۾�e+p��J��+z��S��7�Կ2+$C�S*��������b��#����wW-CG��M�
��n��~�~~�.-���I�9l8z(������+-�qԨR�����' BK�	Z,�:|��Y��ž���n(�
蔻ȱe@��9��k|�`0�4X��E�/�fm��mx6ū�NG^=�μ��ٍ3�J&���}(�$�{B�>л�x$2yK�P����6���nA{��o���H����pkF~m�z�`��#gJ<޽��c.� c���3�F���������?�}�Ө�^�lKWm�ͼ+D��v'�p�)��9ɗE O��ٮNn墕��b5�Z�T�{�yj�`���yl��O�=l]<�7�I���xs�Ak��Z��������m����tЏ��=}3�ڸ[��e��,3z��o%��[�a�5T������
�W��QI����y��ъ)��$��!�\���~���)�c�-�s�E�k
�8�r��u�/1�7�ݭߎ�(����������B�,B^RÚ�hدB��y��#Q���P����It��$3�_�7��Ƭv�)΋4���v�[���ʦ>�8��~������{)J7<�?r�`��z�x��moǤT���e&�rܡ�6��iN^���r�j��:�	�����U�"&@6�����s�BȢ4Tz
�m~4��8�*��煐�@-�A��+?Ar;W�����Z�h��d|pg,T-�ͦ�����!��g��hq�U�E_�<�S�t@j<�ӛb�2LJa�sݭZU"�U}�` �l��96fgqD�ؾ��$)1k���D��v�b��OX���S����(�.8�:�n�U�I�e>�0��f���ǟ{�6��$,�?J%�ƏTg���uX1_����W��sK��3��;�����ۣ<�'�[L�<����ZKη`VD�w��`��-�����P4�AW9$��c�L��7�+r�-)����4v�EQ�S�x�����W�����y�Ϥb[�w&�N��X%o�?�b��u�q��.��=Ѥu(΀ؼ��0��r��Az�Q����y �Hك��P����Jn��I,+ c
�9+0�����xvT�l��V��`u�2$���Alqa���N@�mѣ���б�=E��)����l�����Wc��5�0���L���RCWT~�����C�K.]���e7�±=���.��6�;�6wƠ�ҟ�|��n
1�TI�r?���W&��:�&���W̕v|N���'��9PC���N���&��`h���
+�	�F��~c���Ŧ�39�$o����@H��iUSyց%=�f�/,���I]����m�a[W��I{$��T�DsÅe2�턊}ଆz��`�)q�b���ڪ$)�)�P�l��]n~ʗ@V�=�Ў���T�yJ-;~U	�tVz^	���cB�MH�Y���O�O PH6�<mv�*0�����������3�Y	�;���9iU~���y�ዅ�V�˺�OF��Wa�q�?�B�)�G��*J�y��p�{j��5ʎ�}��Tt��ǆ��_�L��h�+����b�\Q�����V8�L�"�%�Ԓt<�i�1�_�5-� Yl���&I$�m�P�f��Y��b%wn�Q1ƪ�p+j��:X��^��P
����(�Y���aj-�	榻�٧e��dO5�?.n*q�Ir�������粍����IQp�)E�U����Cf%�����4��B��=g��p+wf�{�e�㪸��L��[f���t<�I�����Fi��9J�Q(�1C���Ɛ�.�F-�p���4�{ Ux��y����
`�ҌQ���f7�����\��Yض�^n����D5�9]Ă�'ۥNi�#b��w����0	9]PC�Oqp��1�3�t��t���N�t6�I<"N���/+W�!jbX踕��vQ'�oK���#�uJ�z��$�O�~l*���������cKW�-d���u��,[a(���#S���2ǵ�x�ժCj���QJD�����C����-��er�#�b�^�^]��F�^��k����΁D��N�ݘ�	dژ�tbw�B�a���8�Y*�H`������CNG�����2kj���nc����j�q?9�Qǯ��SY/�->w�Q|J�p8��;@Hc`	y�zb�A��}�Um�P���G�u�տ�*,#�e~܄�dh��H���KAp�Y�9<������'�,��E�7�G+��.���}8�ڷ�mVm{4�w�uܬ�q��B�<�[0�����f[壳�Ѧ���=�605�$poa��+��?��d3��ҝ�Z�V�z�cZ!���+Ƞ��H�P* �e��ş;p<e]�
��T3�.�4ċs�x�����nTf���3ɰǚI��k�1c��f��Pg��j;Tez�)���{trN@z���C���i4��v���A�xܛ��������[s��0��A�����@�le�@����Ң�Y�o���gM�?������)�1,�_7ʰ7b�a�MV�4R�7WqA����DUS�s�i�o�/��'�2�3-!�ey�[C����m(�@F^o���(8Ĵ��ǃkT�:xA.���7��O�muW�4!{�h������l�Q9n�Q��-|�Y�*�9;6����	[�)�x6�Q;>4�mģo>A��+�~��T�R���<xa^��,w�7�E�T��� n�
�\E,
�QЬJ I�t�#��]�MXрp�<ۣu��J�S�؋2��u���	{L��fN�{F[U昨�.�J��c#edS٬6�<L�<'N����_��r�����%�(}���j�\*�x�3C!��X입��KF��Ț�>h�4B�Rz#��4+,h@�G�
p�HN΍�r+��	��/�/F����q@�0��A��9���k:8g��YP��3wӽ�뇮�M�����3��X	�0w_�"FFܧ�����e��g��F��"���K\��lt��<4@��/!�M I7�))��ļ��f�v���%N����`4zӏ"1��"�0��U�\B���s�6{��Kb���3�U�S��j�h �d�bثȧ~l�S��F���c"��PU(�H'��Р��"�Y�e��{�P�TxՇc�j�!�؅?��OF��쇡�[��,
��IzpiaJ��C�k����� r� V�?�53ϙ&&�	��:}�l�F���I����)8<y�5�E*��׆,�d�)����5�k?�My�L5�X���o8u]�-o�~�ԟ�x���F�1NB��ȃ���Ob�+!]A]��=�Ӌ�O�;/PKpIi�ˋ6?y�Z���D+��3+��G: +$�2�a7�O���sVj6:87�Q>����ٍñ�F?��d���ăZ�dxP��f�2���.�NKS&�����G^#�w
��_fK�HJiG�.+�
$��:�%�2�a��h^/x�4TN��G%�Q����<3��N�!�Jx>�U��=�mu.�@�U4�\s��G��q�h#���4b~����ž�7��n�	WML��MM� M�[3����7�'���MiG��FK6 ���\o���t{I3�8��|�(+RAcvjM��Z����X"|P��f�U�:};�%j���� r��Ǉר ���Br��LJT���7k�h:k�+�V0���M��Iv��M^��V.u�fZ���	*V�9yR���-H(����Ƙ#�S�J#�~�p� _�異�S�*�7���f�@�I�(��X`��1�r�c�v�x�60��re����C���@��`|��L�Ӕz�Q�g�냘WD���N��1�	���@M:`��VPZ��Kԝ�ȼ�@��$N��B�9�9<%���q�/�c����n��~̉�!<���B�LK7%4�����F���#�Ȇ���X���))v2pwա�Vǳ��z�1""=�bҦx���n�?? �/�X�ni��l~�w�7��:��l��sͩ����K�6�\tl�nX�c�k�$r�?�$u�(Ƣ��v��v����t�q[͖��Q�"j7>���#�JTO��D����. {�y@���� d%�HH�6@��s�����Q����?���y9	�Qs�Yz���C���鞅rL��Y�s�~3+;����٩Et��e�7��gG�ŋGs?����L�n����W�t:j�Dɦ�e�ۺ�Xw�'Qx����7_�A�h�l`�_�ւ���me[Z�yը�E��܉���'��N�������7��7)�<#Mr��v����.}�Å2����)�Wd�b1��y�†n��A�S�ߋ�F2e�a��1A�h�;a����� n��K.�v�@�#���Z���8��bf��C�LHm��K�!�i��Zp���R^�2L�FZ)O��'b	ڹ|r�i���vg�RC��;t�6Y����©�?�����{+SK�Rr6��=�Q(-��n��L\����_�T��d.��4�Q�PΛ�Z	6q��+
��[M5���x�
G�{
�qZ�Pڏ2�9���t-�saa쐅����QI��i
���C����E�<�F�Gh�ϟ�bP�I�%���b��pm9��zJ+J������^ܹ8��#!��^jbm����]P��{��IǴw?�&�4���v|����%(M�Ϯ��m�c��Ѵ�0�a�2'*���!��7���� � "SeCC�UW���ci����@��������݁[	�;3.��W�x$Ȯ� �0��.����ek/�n�7� �ӊ���)K��h��5a�R�?\@0�����Z�#�W&��x�/��CR֙��\����zxEF�6}ΆK��,o��+�T���q.n	�������9M`Z +�73f<���!U	����!�BF>��哇b��
N!Bm+.��8XS��X�"�Q��n�L &��ş�+��U=~C�c ���5Ng8���䯍��wf䋌�|f�+��<3Ω�C-��M5
�PՉ��D�j���B��O�W,ʻ{ v�����
W�g۱�}���fի�Je�!H+�t ��JBM�㖀
 �_l�<�C����
�]�Dg���A�I��|+ͪÉO�K��P��;�Bb�~����y��̾:�U]�J\�� ����dB�:D�E9��\ͷb������kM����;.���=��/"Nt^K���r�3�U���������2���!��Z�Z�p*��!ۭO����OJ�q���e�l��,q�t��:$wR܀��.���^]�x<�f�:D�'M*�`�ּ��#c�M�����xg\QQ�8�e��O������~%�e��qb�GfcT�4<��34�i�cl��#r!*��T�Q\�M�G� 	�5�W���p���Q�j��cՎl�5�Y��Y�b��::Ge�P�cu�O�ϓ�����ސ��`�(���O&��+�I�w�(���E'Pq5�?H�ysC��fM�B��
��i%�CT': ��_���S1�F�@m�
��-��ߙi�`;.ApPӢ`���� rZ-��|	��I+��8$���FEf�M���ȷ9�V�ľ��J�����
��vP�|�D���v��o%e�?�b�u9"C���0MK�!9ƶw����J�xt��|��ǹ���.�do�������.�.��ڱ�c��T�ku,;1qg�+G�d����"�{�I��gu�(�Δ.���8ΐv[��W@��,h�[��I�P���՜)��-R��Ͼ���L��ts)@j���
q�i(X��V�A;��7����sV\�{��^,�[�żj&���Z�Cs��Q�kkE^q�e��W�o+ k� ��N�xj������,}��k1�������#t��.۟�w��`�5���[P7�yp�\:!Z�)m\a��8sv��elw�`�/�T=�yu��P��ye�lTI�'^3D�q����a�~<�uu�Ho΀�����ҔP����5�{l�$�Ww�K����		�ͬ�tt>�_�u0�|JQ����Z������l�p�4���=�'Sz������sִ���q|$����.k��3\z֐[2��|*�}�A�7�څ�W"��-�{�|זM���J2�Cj��e6I��� �+��#��Mٽv�E�_���q�6��>h�`�.>���)��Tt��D�
A���	%����Z-JZ�<�
"�!YQJz*�-[�2��5�Q�8fjA'9��㻝rM��o�d���<�M�jm㐿��n�#*��0Kѹ�N��� �lJAW�dk�	��ÎA�]<h�v��#����?	ßn�iϨZz����W��9x�z���ɃI��;�S�nn^��8?��4�_�7� ����˕Q�8m���`72��Vй��~�`,;�;�(����Ӛqn�Q�	S�����ww�N�;�W��-���j&K��y���}2A�����*rՎ��	�����A_�M�+�Q��S[B�t� _�ɶ�I9ʕ�0��3ڃ~�.�ѣ�9���>��>!�Ҟ��6!~ KoP$�;� w���3M��u ���M4l'��p R�A�S8�Y��U�lc�>'�B�y��d�|U��a�W���A5bfȶ yO%�F�p&�̞G\py&iv% CUd ��Y�7^��D���t�:c���	cJ<���kN�e�+����y��<!|څ�kr�豯u݉����-Q���E�Bo��	*U����w��8����������J�֑��2a���{:3��w�=H��l�Ό��@RL �~U�d��ba�$�^�����AE�[����I��h��xF�� E�q.
�Q��Z�����'t<��V�cd�7z��Ķм�&�||����ܧ�ʰ��ܲع��zՎ��/^� �_d�?�xг� U��e�5L�Ց��;��%�S��h�-����!�8�ɉ��H į#g���E�±t�.kV�!e�r�k�&(�v�� Mw�zpu$>�A�J��;��Ή�s|����T� ��j��.�ѱ ������4�����%�Y����򌵘���
��� �G��&��+wf17�����_�P�*��ߑ�;#ļD��Mf�q-�ia�B��	���ֿ^���M�}��Z�V�_x�x�&����I�)i<��K��> ��.Oy̙�]�-�/5�U����bS����_����"���_s���R�Q�|}���SjD�"�
�;�8q�GM:��o��pr�)�8 ��W ��]��^��)"�P}Ű����lE[�6�RGϾ�� We ��a
�;���l�Q_�jr���.�.8g��	�6E�p���,�+	�e�U�O÷*�,���d_Y�����=҉�ٰ�7fm�<��`�K0�;�W��Pb��z�o��3���V��������Si�`�VqU����l�!h��F��54�bą%����dC���e�#�vx�h"�Vo��1�H�#�<s�)���rY������kh���y�l`�R_Z�d�����4`)�۰���PŴZ�Lz�a��`��Q�v������l3=7CF�;�!ߛEP+���/<�F��'�?:��m�֨ܦ"g$�+o+�)�p�L)Q  �v#�z*�x��cMo��C���Xbd wB~�-ă9A�c�9�,��F��V~�-#k"��m[<=	�>We�RR^+��յ�v��[ W��!���n����E{�-���.:m^SP��^��e��!0:.#����$���8Z�W�HvRN�+dG���N��B��Z~g~��&Z����u�kd����sN ��mۼ-wy��*��Ԛ'�4u��)>�$�r�&�%	W9;�Q�A@H��"=W�Ў5�:~[җ�4�jo�q� 	����|<,7	9S�����P$��c��"��S��?+w�/ռK� NJ#���{b���:�X�űu~�@���
��!����lx�n*S����!L�p^�&K0���5f7�ʓN�_��诲��s�	���~L�kp����s0
h`̈́f|�}�m��
ȷ	O�����=�������G��|?<y:w�\��!(�^ف�g��OP��Ilgﬡ[�R����0	2g�Y�M)/��v&u�NCIN��(9��_R�Q�/6&S0�_�p"D�x��~;��P��０��W�U�RB'��D>�7��N�x�p(�Ht�5�(d��a��0w�s��G�!���b;h�χ��(����7_+� E/���.R,�1lYC���(b�?�5���&ĉ숸$���d_9��8|�؛��5�e�(�
�tv�휣-.߇*ڹ��N �C�'O�șx.
�c��y0W�W����z>�,��E~�*ɤ���q����7�&'O�u�2������za�1��ϙ�ֈ��a����wn��#��g��3$<w���;A�� ���&s�Z7DAzLRWD�@[Lp�т�v�P���S�����S7��A�!oy1�L��b�S_<	^�2Q���O�#0���
AHc�>B~_��ʇ���_<�W�@7{,�*M�f��|4@9^�����^�F~� @~O�L,�~N��Q�<!Q2�ǽ� �ַ�q��l�.����ר޻خ�X��~b쳉�t� �ܶb��<ݘ`.5��6���^�K����*�y�Ni�f�L{ܳ�&�8i��y�,��>ey�&�j�}�7��H��gO^@�ml$b��
4k9y�v��]�r᧛���b{0���H���p6dĻz���nD�[��@A�
$�`:�%]�1['ӊ��_f&qo��0:��ըJ��o��?�)�5 �N}��w��� ���C�d����=��%q���
��Q��?�d�|�W����9�8�v����3?^�S������}?nD�.�B
�*���}�Ǹ3y�n7, w��Ŕ3DR����ER�k?.�i���a�ЏF%�M��S琵 ��wX[ʦ�o��B"^]=eG���ý~3˽�8�uج�����-�/#�R��Y[0BGK5H
��=+DЫ�����Δ��2����#���;`�vN�؍aZ/O1��*P����h8��l^������+��(E���b?�iV��K���R��I�Pe��D�O��|�1��I`^Ju�a|���#�B�F(g�@TN�b�d���'��w����OT܇����+8��27��i�M��J����x�9������G��y��=�T�s��q�o�v�"/�_g����c+,�/�R���u�H(��K�v����L���$(j����2�Ĝ 򝤆�J���O��R������SW���rǜ��?���4Ǯ�k�[� �����]t"��H���A�@�z~m�7�Ч�e��[e���D2�Zw!���1q�w�Wnc�;�`>�P<m���!�u�k���}>{�&�͂�R����b0�U��?gwy�pjb���\9%8�wmw�:M��Wu�2�����2��H�)U�86�(�!
(D������Ƿ���L�����g@�}�+�C�"27gP{g/���m}F�m#`#x�m�fzAM�뜗�M��٧q�訃R�x�|���'��Ph�� d1,�,ӨPs '��R4�&��>���~���-�k ;��L5k:�w;M���� �H5� �F�<E�v�Z5�M
u���J`�(尾�/u�/Ak���x2"�
��ݙȜ�* ��lV�N�a&��E�$2�eS�Im�zz������m*���X ��� �!9=��t4���yT4G[̒+��J��یAt	@�pO��'W)�6��eĎmǌ��\����xL��o�N���g���eK-�"Hp���&�{L@�ɽ��=�׃-�(��S�����>��0���������[^���o��aiC)"ŪJŤ��r_K��06���I��\��T����+bt��w�^�����20��9|�cc���J����|�&¾���嗚T�^9����׏�[���[�S�]0��5H`��
}y� l̠�
(�PԞ!o֌+��EQ\��yAfy��;U�y@��� ����q���������%&�ܓ�E@�����w���o&]fy`��l��1�=���F�t�|��e�#a�͜��EKo)�0NU8�=�ҡ�����L���A>�?�k��"u���w��*�ml�֎���\�g͒±G��;W[��ͤF�����+����۾��
���`�=����q�!$�Aa�<�2V��Ou�����V|Q
)�)�uҟ���u�	UI���l	�E\�ъ[ա�����0�K8_1��&�}�KӷЎ[�LL3�� ��Go�]��K�d�I�`A5hb|�iJ�$��rA?ջq��i�H�����f4����X^od��fs�&�!	I�̭�n^��N1`
���-�k&^���Y������l�"U��v�
d���Ok���uԇX�ŵ'TZl���Ba%�����/���md�ɇt���UI|��C>vhN�DX����j�2���6�����d�߄��o�$ �j�u�[���ї�}��@!'�;Җ@F��A��e�"p���L�̬���7�ysF����r��Z���!tn6�- ����J�_\�8���V�a��{)��̕���6G�`ؙ�
r�e���q���+�3|Z�2	�S�v�(��^��7�+�/ =�ͺ��OՃ���.���R9�*���z�b�z�F���OΉn�)6/�r9]2�a����wlWq�H���hxxW���^���؞��2�k�by��� [XG4*�s��[�����!��͔R�+�C���'֐o�����AIpa��^�TV}��"��<*���!#�wd�[����r<X�"����#jJ ��۰7�FTef}]8�D[���x�q���D�K�d���qn������I��Fb�h�O�Z�tB/��ܾc�]��x��	���f�$�.��h��f�OR
FD���j��2Q0��'J�iI��
�	�m���꟟b�۾�`P3�IG��(��okGo��U�< ��X���W�D�:���E�� q���8X����$*V��i?%�H���X���{2Z6���Ȍ_L�����ız/9���ӣ����qJ�ٲ�BԔ@f+�y�r����ˆ'������G��qqO�i+˲�����fF1�3*����u�5wm�
�RR
�AO�>I��Q�TW����3y�Գ����[���[k�ػ��OH���/pa�"�v��n��-�L��!lt%�lt�}���c�c�����t��
R
�<d��`��,��k�h�s�D��(��'��t�k�2ft�A�4�
N������@~����$������5����Y��Du�@����s�>k�����v��8�ˤ�A�%��r�2n�������[e�k\{������y��M�
f� 8ɖ���"�)��a�did��M�ӑ����~B�J�Ee��X������H̰H+�"?\o%($��Z>�(ȍ奀�L��=�]�*h�"A�o��g��8b9�4��vO�����N����-����!B8���wi�Z�$'�A�%5M�4���O�HFx�^�a���������$ �Ua����ྛ3�f:;�x�(�~Uy�=��-���E �o�=�x�L�_�I�|��*d����eX%Ģ�qIT
��i����A����y[>�eL.���H:�P0D���u=�Нz#:��qB�.�z��Z\{ ̨����sG����S��*9O���~Ung�< ��^*y��_��
:.z�����v��ޡd些_�/p�(���ȡD㒛������TNd3�ʣK ����C�� �j[�""�_А��q��_Qi7�SQ
K)2���[M�-�&E��|TŃdM��B �=���;V&.3\����4ИP�M��{lSa4e_�F۳a���H��1�M�����w��}`̱ԅ������|ݽD��	3T�w�':�9V2�e�Y��������A��9�KvX%à_�i�r�|�أ�
$���4�����~�GG�+�\&6AW�/���CK��Dt�M�(�x��;������:����Fa�b�t�K"qr��,���%z�a���=��ƪ2��S��
 �����$ȡ���=��iN1ё�_k�E��!LY�+^�J?i[ۓ���D3O*�ZA�{��t-��lAƧt��� �2�	���
!��t1��� �X�k�B�ҝ��� Gg���}cP8�~2$��Gۘ(X��`TkχŦ�_.��w�H�/�Rf��k���zk@urh���X��������,�*�S�>C~�7�k�{���x���i���9�V�/��Ȑ6��M�y���
Y���6��w����\N�*M����t�2���}�Rs�I��A�$���V�_r]��^��Vm@�����w���6�DFV!B�{|���ʆ�)�.��ڢ�����ָ���u:-ȳD����kf8a+e�@�/,�G��j�P'�� �r�V�CP��$2� �Ѿ�5&��Thg����N~���)�s���Z����)��2�@0�߸o`6:���e_���?�fO�*,7]��`��3�d�Jt7r2;�z&��{WO�R.B	 ��-r����e��;B%�.4:���O��OHQ5���y����������݇+O[���Lx�ͪ�J'`cT��S�����U��
��U��[�����W�(Ha|�8���J�� sR���:��^��jk|�������� 4?hH�|-cͫH~K�	CAyڒ���S�ioN�|~���ʒ�m�~�����eK�i��t�P�d��@�)+3��<��u�[F^�@L)=$&�<�*O1/���-�E|\�<�o�������%������,_�WPh�$�]dY��}�vĲ��f�7�q�4��G�J!�,Hq��U����V���D�J���"됇f�ଽ׵5�s���U@��I�@�G�t7N�ÀX��NfT��xc7(�w���ף���=�+�/�W���p��)XzBTM)��HÛ� 񵡩�9&�1�J��o@���fdP&��2#��¥�ů��M��:�w���^��4�H8�.P�V��$��p$F�G��J��P{���Ճ{Ky��2��&��$���1�Z���Ɨ�řg4��Bp~k��W}�QΆH�B�
[������ᬧ�fu  N��c�j��Eb�=�e��*���r1}�ҩ8��\�Hs�)`>!$+ꨙ\��N=�lB�߱{����x�M�}�@����D7��m
�5��]��p SF4\	�9����[	}]�ܱ&�@l���HoŴ�$O�'�o��$ &���9P��J�)�
R�ԝZx�'VM�@s�u(L8���:r�s�Bq����b��	�{�J ����3U��qxy8��A>�!k�(����L�_ j٫aSw�^n�hMY����Ԁ�t�����4"Y�-��rsZ�G�����s� #���W!�T���T���YY��;엕s��Qe��K80Z���=|�U*И���'=���Z`��1dfv��w��PI��'l]4Sn�Dlݟ����od���N8�N[�Q�ލ�^� T(ݹ��4����@H��ȳʟu)ͻ��Z�Ø�g��;K�.e~~A���?]A�N���4|1�kU����_���O������Yhzv���u}ZK�����?���u��`ա��W*��k�ܯ��찷y3�Q�$���������w��dA�gq��V2}7,�ķ���zBDP&����F�Ǆ>0Wi�9<F�a�{��ǁ1찢�+�)Y�B�J������*��Uӿ��vA�(�e���+���v$�M��q�}�����$��oш�*S�J�ʎ�!�2,��\�uܼ֚VU>��~�����*IY�A��6��;��%q�㛝��a_*���C��=w�����m�Mm����~T��Uf�?��vCwfH��F2S�m}P�~,��8��v�>���O�򴍧���<O��7�(�����K���L�M�i�SvR��7��w
�Ǖ�JD�N�y�t��0��We�V������9�R`+::���?v�UKڛzL���7��`oisy6 L�|(�?5���0���$��Zd1�n�
j��Z���X�-�-"�Bs��A����҉y�y��XF�@�dā��m���\nnAl�oj�5���u��W��:䓕h
?��ه��������Aal�PھH�~�厠r�?�5�g�Ň�N�o�>O	����n7*�kOp&�$�'*O{�wNw��cuF��;^>%�>.����?�dF��"NA�X1*�pL�Ɵ��'A�ΔJ˜�@�ذur�J�G�^ADp��#:P�&Y_�jƭ=��/>��UH#93	Ěİ5ݹ��^Q�T�0�.d Eh�(;������l�����JѶA������7z��cQz_Oh3@HՔm�x��C�x�d)93���ҁӸ��2���t�2��/9�P$��|�h'S6t���N����~�����M�x�����/pIQ�x`�0�Hl'��_Q�G�� ���P�=��<�Ӻ{���k�/=�M�a��p�E�[����}\�j�r�6����!5�D��vk'�!3w8I�l��3��B0�4_ۥ!��t�C5}Bt{Z�}�HRL�������I���(u�>� %�O;W�#�_�>q��Ⰷ���-���lUb\����H2�6��Z~�s!_I��Jr��Xc*�c~Z�>X���w�[��|v�xj�vƘ��|HE�_ԅL<�S���K�Q���%�ݤf��z����� $�V�a��/u(�@د�)*cb��8��c~G���V1�1�̨�cz_����.�5�@p^彰^�0�kŖ��Ӽue��\Z�:��S����B��v��!6��uM����'�ꩥ�w<�}���Q�@8��e1�s�r�(a����c������YH�u������|�tդ�x���W3��#y�ξH�[,�z�@iR���Ig�X���P���@�},7v4�g�$R��g?v2ޤ�Q�@Y�{0�\ygHcGz£CC�� >�裦�ۧ�LR�Y��s9����C��5��U���{����'�� �F��5����18ɢ��6b�b����8�/W+�B<�ŷ"�SU+3��rmX j+F���K�_�@�K�1���wJ���	�E���&�ׇ���Z���z�)�a~��n��NU�2� �+�.�Rv?��Ƒ-W\[��+m�X1M#�9�����/��(�IT�-���5Bu�\ʩ�{A�<ĊqD�R#�7�)t����A/�/�����S��-e�m� ;��p�̠�	Y�ٌ؁�_Ħu���Pg^�N Ry7��^%@k9O>^�8�q��]ܢ�0q�~��g��M,�Ȅ$"~�
��zF<�ڕ��5�#�������d��9�"�%�i)����f������Y�S��6@J!��5e�]�`nJ��@��jThTP��]��Q��[iҒ�|�)t���s�2��$�Di	-v���eE*��o���lW[<��5���2�.�lڙiFZ���"-������[�՛��9C����j3�w�a�d�^�k�qw��ᓢ���=A9�(��I�Ֆ�4�1ą�,��f`#wf3�A��S"�$��;�V���~�E="%����G�F�)�6�����&�K���f�?�q����T��@�֢cҙ��/�>�J���(�eK+�3�B�3��"M���i��7��g���w�2R@�FB�>n�r`:�3�ʭN��kf߫Z/N���l#���.�#�tԖ9g#j~ܼt�[+^s
�}FI����E�w՛4y��pi(��쒘��j���+�{<W�lsT�"z&���XD��Q��)L��z�g�r��/����
�xi�z2��I8�c�k��������2�~C��w����^UO�Fʵ�+��UYT�D��X�Sޏ��i�8zX����kA>*��Owk:�v�ul�/U���I$j�?�0#�kR�(y��[�-�[K����}EEi��.iw���Xk��OqzD�jv� -Q�u]ȦM_N͑�4����>�z�˶��9@��j�ӎl-yGNZ���?6g���v�^��+n����������WĿ��m�T�A\���<YB��H��Y����w	k�V�R߰E�C�Fp�r�kH�d�WGM��Ǖu��� �&0e�5��b� ������O��U�q悓~Z��)�T�D'��͉������77��b�$�y�M/`�آR4l�iJ����W�`"�%��p  ���	ux�x��eN)|�?{i��B�:�T���B��㋝����@�?Q��nWo0jY��zh��9�v���<�)&6:�h�R��ܜ����S}h�4�:@ZK���m�N���k|o���6l�p#ń\oF9V~G+f�F�Y�A� �b:��,u�n�ŁA����4<Q� nÈv��|�K���mORQhε����LE�.�H1�MD��u�xӲ��G�dF���q�-�I�j�E)� 1x'4=,����$r�a�� ��1T�n!�k�p!��@vʇ���ض�%\\|�0��%w�����2�#��ġ6E��~�bd�U��&���0�~�k��͋��� E��ѹ�0��P��2���E�"���M��V�C�i|�x����~Q��Q8�t��Ja8��۾k®4���L�<tx�����T���1�G�c�+�/��2V�'u`�|���)�a�F۪�:�gc���J$���xjHF�Ek�[�4���k�ꁑ�}A���?; !ʙ�2؏���>�t�x��A$�u�#�>����ٻ��?t�H-i�F�)/.o+��ST��v�Pͷ_����c�\j4ۧ-O�-Po�럮�ྚ�(�l?Wn(�d�lz��fu��hc�"�G.p�g)�"���j�}�D��#=\Ԓ<���l v]��'��/�q"P�hN@�Ʊ�W(���`�a
�+9���\;n� [�5���&f�M4��#����e��`�a8�A�:TH�#{�`�P�/�1�9�c8�KE�4�$���!���Sc����X��b��O4Q$Z�cYf�cF��S���D_�(Wm�ߝ������G��q���޿F�>ԀJ�~|ԍ+��:��u:§ᚐ�8*��C�AZ��6?\�)�#�ˢ��7U�@@�t��̌�-ּz�n)�*�εx�ӑ���CqT\oVG�.��@F\���KL�ȷ~���'\s�"�Tx�GC����]�cDٞ��P�a��n�H�a�*��s�Um���n\A��&� �,�2o�^h�g&�vΉ�˔�:�栥h���4���j�e�ߝ(��n|CY��(,�#�J��f���I:39�6�)�œ���;8E����A�w���W5rh�@tw�ew|[�����VcY���X���ڙH�5�~����u�j�����	)�]t��Ū��@У�0T������ DE��^	��}���.t�������p;ɾ�+̡�Z�5��u|���ޛ]>eL�;./��t[x`�)a=�{��4UL���)�$�4L�xT��7�e�㎔�ɨG�G��1np�固8�$`���$��v��,Wk�~���1#�^�L1�p
v��.?7k���s�BL%뺯피)�'}(�k�M,���FW�|�����ͪ�j��XV�],���U[����f>��9�H�9b��d��Nܸ����\	A�$���@c�q��Ŀ]
�iZz�?n��ㅒ��z�Y���"�A-�f��R�'�ݞ�����;Ғل�M���Ƞ�;�oV/�ګF5��2i�}Ё'�)*�L� ��Vt�%,��X�� ՘�c��.���,]e�DOɚ�&�D���M8��j���6�Yi�Xò�����	<9X�z^�~<��߇
��S��~2WJc�[gߜ��|��4�@I���u�x��j_V3��r9�y�o�XLg���ӹq��"�Ӊ�Tv�Tow��[X��=K9�
�o�7�u�ݫo���>�.�V���	��C�o���$�w�2\���q��~�X���t�Kal�Grw?
ʕ����6I�V,ʹKc��I(�	�ğ�2�O�g+d�Q3��|���z%��+���>�.����z���6��3i�b��D�a��5&D<�-�r\�>d.�M������w�I�`��V���,�-����g�b���r�S/�Nn��Hc�<}�����.oJnOڊ���+�QgG��0ZU�G��,�AB�&����]l�h�ŞD���8����?�Ў�4��i:nVl<�y~/�/�v�+'��F��|�[>K�~ۦ>;� �#]8_"Dߔ�;o�M��#��[(aԀR6��i��zz�%0`@�v	�O*G5��t�&P� �V:xB���8�6x��V"e�w�X<��
s��_��Œ%�����dՕq���I�"g:5c���5������`�l��Zcp�ŧ�g�>���kV-�l��Ծ%4��hؘ�>MDN54�7>��Ն氏
��z�p^�P�鵗nZ��Q����:4qbG�5?p@��o.A��e����c�����HRȘ�v�����@�<B��\��r$.�)���l�V	��t��Œ�gk��0cC�ˈD�Eؔ-i;&�/�:v�f{�b�����|`��39��*x4�s�6@�S��Pc����O)�p��)NI���#0�ť��(�"�fV>yB�4�V[sԖ	Oߕ�����	`���ȫ����C� G�I�M�Kns� JګUJx^��7�ߧ0��P`
(F.�s2ß�%0hS�V�a
�Xm��<8��yƵ��$3j) �Sڌ�D9P��Q�����0��!���3��
"�ϤE�'f�y/}3���/2�y�m#5x!����"RZx���TǺr�<r��M����ۗ���N�l*���@�C�1K�8��8�i=1���ayG��B���!�������h�?�=]�L=���C�a-x��R����ib��W�W��G^�2N�<��d�V�F�o� |���x72���W�*�:pw[�
5R��� �LD!��H�UH:�mAy3�B��B��p���k�nȥ\�Z{�O�4��ح��
�<���9	�=\X��5�:��2�d�K<1�La�|���ԪD?�Ƀ���b���%�v�9<�άT�z?4�ź=��ڇ+Hh�{Ɵ�b-������{�����Ǘ�<z�T��j?���?��$�ĉở��3D���?��>�Q��%S��,�`�,������,˟2�{?��� �ab��ОsD
o'�R�)
P�B� ȕ���M�+�ǁąt\�h9��8W�V����m"��%�?ezX���X��Z|�����/z��)�"��5��+����:p3.1�2���҇��2%�'��I�Ȏ����#ξ���!�a�ޏ���FDS���D�[�ߑ�,��35�E���<�f��o6��Ϳ��r[h֕��>��U����^ ��=��1j:��[ҢhK�K�"d�T۳�]������?�Ec�`$f�����ɩ�����}�943)&�E�_��Aj�<�҅�<Àp��I1� ���Y`��'Z(�yK8[V���
NQ�u�^���/���a�
���ΔsM�'~���X�{a��EɡiH]�ke37y2+2��n��<�h��2��_'54QlWNh�����]۱UT��i#|���^χe�j f���,���M���-v�}-P{��J�a��oF��=N���%� X)+�qȆ�1���}%;\ukd�R�tҷ����"*f�b���Y%�3ӈ�V��WD�:��Z���,�h�	WȝZ(�����y I��e:�r�H�0�� ��[�JK���?ܮy��eVp�e��|pAe!.�	U3���w,ԃ5�&���D�]hB	)�)n�����;}|���fJZܣ<��?{�sX+��,Q�L�o���m��-�K�4��Cf��]�����E����%��F���P��f4l!��Y��¯���H��+qu�d�G(ԋ��w!3�4��#���i:����������$K�?+9Y*{����$Z� ���e�x����Ց����tW�n>�T�G��xp4h�H�̚h<FS�|�A���*��o?�,�c �n�Ӳ��_5��l��͜�@�G�[�s��G������R�~�!Kxa2U&�|�B�K3�q��M������S��E��n+r�����`�r�ܦt ���?H�������i�oK�Á�ք����BɌ��([����_���X|��H��
�b�I":�Cl.���'Pf�-����N�����a���'TuȢ������h�N|%e�Ս	�T[b����-P�9~Կ���&>MV�!�ř5H�NTO~�1���.�t�a��K^N���˲�'M�2#�P���^Z�q�x1t�D;r�Sm 5W`�S
�����/��C��Nw@��mno���F/���	�+ja�XȎ�B�#��U\MkK�ޔ!��)�%!U�dw�5@Ƭ>livW��`
x���Dh�j�����/���	�:�C�br��}��)���9o�͑f�ѡZMFY3�`��9b���f�!�f܆���[�������7$g7���'xׁrÙ��+��3x?y4m�Ŕ���ׇ3��B��+��nTwb@9��n8L�*��%��P�S��n|��74.-�˻���Y�Φ'V��nU4����jVă��o+�B˸z$GWj��vtl6�k�"=�?p��F�3Hɝ۝k���\��N�\8ZK�}K��ɘ/#�2�/��d��tO}�Ef��{\&b�Vo��>=��W><]>j�h	��ˈ$�Т(I��b��l>נ�LIi"��*aa��%�|�����fA��� Ga�V>V�#�8�6xt�m�N@���~v�@N�ϡ��bdѦ����n{��"�����2 �8;cN���!������[�Y�5��2�����Y�������x�YS<n	7>����^�����ɧ㾹kCC�C1���K�$LeT�wUybҢqx�=�`#���r�1��q�ʌ�h�:�p�]O�*rS1���3��m��$�����We��EGe���Z��&��E4<B�U:�۱ǋ��R��C��*^f5�-& ��e������l����:6����c�v����X���c�^���Z�i�g�7��I�
+��,��R`�A�m�v��]W��0=��=�J��?l�t�6�O����� ���Q�6a�,%�iF���!.�:v`!'ٜ莶�p�'��9
�e�b�Q�w�P�ڕ��tD�檓�>�Ш)�ox��n1]M�׽p�C��V�Y�v)�� k:!�S�=	2�vrp&�}e2���x�~$�s��h+����"��y���G���~7ۻKE8���$P�B��j:vH�r*���\������'��2ճ�@@��m�w`d0��)��	�3sm�<1�5��c{U�շ݀�\p��/�Y��Kg��J8m8�É������OhZzn�AN[�%|��<N��>��F1��-��L1�+ǵ �4b����ܖ���T_x�d���z�f�p04Z9�/>�1{���q�eo�I�6b�CP,��WGZ���/ͮAFrv:9����IکG5*�� ��MsL�;>��7��}}b�H��H�J��Lɼ��Dk��N��ȚE0y�\�&��@�[�%\����R-��iJ�U�C:MU_e����<ktz����fִ�5�h
���vw��M��WG#�J)t��GyBX����߫�^�m�7��uG�?�{A���|���,VRp��]E�O��lE+�K0�bM����y��Fj��(_�h_���B8Rqa�`k��.qO�^��E�Z�����[�Rz�p�ί�H��e�\�?X�����`�+�HÑ��?c��Ə�Rǥ�ں,T�}.���pF���Y�����*L��hj����k��Se�k-�ڍr�ʃ�*�I6��z>{bP��H`���ܡ*p���`U9Q����hXx��0�H��zÏG�7�o�^[���|k�O=��'�`��4k"� ��qH!i�����1��Y�-�$H��+��5f�j>@\�ͳA&	�{���SRu�[8��bo��`�'Ӭ!9ܕ��l��&�a�u��<%м(uP��Y�7=�箆�z���y^�Q�0�܌�e#ֶٷ��M>�A._�t7� ����&��Bw�H�#��Jn9�Z_�-��X�N��_��X*��ݓ>Vz���x\�NP����I�$�T�d>�ؿg�G�$�T����q����P`M�R-쐳NbjyEB1�zg��y������X����[��C�����y}gg�e7�6�~�SR	y��p&v�@�Ң6u�ac��9H}���W/��D�#�X(g�
�UX&��J2�DЗ#�]��xp
��zSL�����<5���͋�SU?�K8�V�wB�&�r����R��y��D�a-I� �7+61��-�Yo�'�ȉ����(����*���ri�-��R���m���9��/��VO��U�i�إ.�Ə��S3և�_ _hĺt���g��sd�Ց�W�8M��*HoC� �?6'�q���:���R+�eP
�vJ&K]�&Sk�	���_X�\�8��p\Р*!�Bb[z��]���!n���*����^�.}��	���l�+��Ehtg��S�[;�&Ώ@k�%��wo��Ӽ���D��d�Pc�)JC7#j&C�i�Q#��G����G�Fb�ȶ0y�3`	U�������̣���1��3�_=`�Rq̌Re�V�v��f��]��,���	H%��'�M�Ȣ����:� 6-Q��<\�+�JC
X���9��诚�;'�w�l����*j���sYZ6j�_Z���G��kJ ��,��՚�����(�w�MnJ3}�MP���_]�ԂR���"��gύ�<�:2KJ���¸{c1:*�R~t�P�o3���E%��Y��[����&�t�j4���=�������M�	�f����;����T�f�����3G����:�s���>�$��LI�{�yT6�� �G������ӈ����D>8�w�d6f���	c�d�s��a`�ۦ�� �4/d�?Wߺ�������K2�������l���n���ɸ"8���Rpb!Ad* ���I��d,���ā�����iC'�O�b)0���G����(��"O��N�H�F��R0 QQ�h�uQa�.z���z3#��LS������Zh0�X�){\�I0�Ee���aiy��M_�%
�Y3��-���j˒y��C��4�? ���%>�VF���sucɪ�+�A7P}���G4��ZyA@�a��ul>Է0��v�o���`?[�/Q�D��`�Ȣ�
R�L���P�%�
o�_E�1:V�lI�I��3�Js|~4c9)LG[fW��f#*��o
�������1��[b�.��k�W�ԋ���j��_���(K�e%.`���_��ʊ�zn��[*Yq��摜�E�-�Vm:_��'*"4�����<��? �:c�nu�� ����nʭ��\���2�h?�Q�	s�6G��<���]�N��k�`դ���۔�uͦ�#/!3(�T9�[0M�p}���J���_O.��(AR�e@+�"`��7��B=��@��W�p�0��o�3iB�!f֬���\;U��T.ʃ��ְt��R-��g`L��6cC(����A�~[�9����>Dw���A������������R�;����?TWT���#C�=@�#V��c�e�F� ���nX�r�$^A�Pd=�2V�6��Y#�܌.yε�{���{��tTij��@C$}����==�)H��f��V��x�TҬEL�G���5űr��܋�P[�UI^v���GQwk�W����z��)���!��T�! Oo�)mJ�CӔ��ݺ�V(L�b�����K��)�w��!���[��9p%Xi�AA#��m�Ѕ�2Z��~�\�� :���ٛ�MO�v݋<�mkfє�U�A���}M��ܛPۘ��	��q4 /Q��u*��&��]]���6t E_�Gq(]��\/6�!IÕ��y������m7l�\B$q���%�ʙ�d��2��e��RrK�1=�������1�~�xG�j���ޞZX�gB;|���3<\�l�ϕ��; �X�ͫ�?����)���x���x����,�YQ#�^�,�M8:<�'���@���T�|���v.�J���!���g�_�b������cMl�@;�_���a�	7�%γ�^B�!��s��ڻF�H6+Ć��?v����
�aVK&���ɾ��>��4�]�1���'â��n������!�fU��u��;J5��*�,�V���>A�ґ�	ߪ'���f]2��nΕ�,�T+�U�#���ǡy/�N�c���$��\;�4�������<]���Y[aO���:<ri��(~S�LR��X{����~臒n`&����R��\�}��gR8Иnr(���rx\�3��dIf'� 9����+v_A8�v�����b� ��/ bE~%_�'��LJ-7�bN��OB�L�����`7���jD ъi���r�Q�=A��NW_����"}��Y7	�+�M��"��A��!0b���^�3d-�Og��p��K�y��c��w�0�-���B�Ԅ���gF$�=G��l�U;�;K�CS8���-_\�\OwF�J��a|S�U�w˼i��t�Y�3��e����N��ם�t�%3�kt��[��ͨ[�S�_/�78�G>|���"�~Ű*f޸\ʽ�6q[��ʛU�i0M9�$�0&�`	q,�} M5I��0���v��ά���¹�U�V�?�ͺ"��K*���,zp��!�t��@��0�"u�y�����2�:ޥ����e�@:h��&Źvj���瑏�7 �.1s�!=��uy'�;W��bƾ�mzȐ[΄(�0�^ߔ�H���1�&@|~x�N�i�~0E�A2¼?����2
̴ ���/�zuL�=������kf^�:c����Ϧ��m,��x��s�p�l%�O.3k~���n��@��g�I��br�K<F'3�bS��,��z�`ˀ��5��Y ����,`���J�'z.�Y�I�(.��L����Պd-_���rfN�mh�iD����E�����v���0x�z^�};���Hl�J�P���7�����˂���	(��-�?�#(U������O���=�&�������+�^�����=�Huak~�΂=�~A�����#"�+OL����B��g%
h�:lm����[x�Y�?Ҍ���k
���ctX*��W!����`6|A�v͂Q�T�VI�i��?I>�!���a:M�=���ް��/w,S�����N"���.�񣚡X�  U]���P��0P�qi��x/Ǆ֤��2��Ɍ�'&�kMD��3y�v>�05Ryb��%{x�x*��%����>S�r�hTJT��Do^Y.[��mzDȐ� h�Ftם ����pN�y�U�(�R�ps=�S�Pf�#lq����@�������O��t	}�����K
b�'��f��f��l����\#�O1���(�����8
�I�_?�=\�!��d���]˟�`�8+����t�0K6����5��#FM|g+9d�>����84���Xr�IZ�+ז�^8Y��I�k+��e)�eY��Ex�I�m
G]aL�3k��F�2�++סS�aN� �ӈ��sM%Qx��6ЫI�R�MEk�<���Ëz�y/W�p�y�vq鵶��b�)D��}��n'Ma���Dr�h�B��,���
l#�])�U_<�����jG�)T��O �M4�=��G;q'<�]��pp��G�<�������{~ɣs��s@9C��M��Di��L/l�_��c�7@u
t٧de1���D�3�.���M߃�O�pٓpi6g�}������})��ȷaC�\�)�b#�y/#��&�a�QYZ�$��ĭ�t�Kyf���Z2���g
�]�u�p�����B��.��!鱻�0�u�'���ɎQa�%D-���W��*��v�����h˦��}f��L�Zt"RdV>_#6�����X����ܮ�[��ܰ"m���m�z ���g��(WdP�,��ߜ���$��[eqn4Y���5/�������V�Ғ>_�`p�(X]k���'�kߙ�%�6q��qUX��3���CPj���#�F[����s�PK�r��iFQi��u�T��mى��@��^��;�X��(Q�.�u�ad�h�&��26b����aC���Y��-�0�����9����fo�9�-_P��v~��Z�Z�M)��O����������� �s3d�*}ֳ�xd��;��^r����n�aΣ��܌��I/��NO���n��s"��.U쑨�P�mY���	$S��.c6���Z�Z�&���P��g5��� �q���?����k�tv���^T�ћV;�����n�
j#��Υ��
j����񎚸�ne�<��r���3uև��T
1%Z��ж�V]�3��Q��fa�L*���bE���<�c������iN��h�{�txL�1]F
]U̙��_�5ō�`����J���
��c(�p�[�%-�4��ya�5E˓{�|ȥ%e<��h�`��R&b3չ8�2��}FY��j̫���>aCwlW&�v���~��ig%Pg�p0�[랇�S.�g���)S� �N�$^$�z�q�wS��G.����	��{������Hi��o��d) ��s?@��3\o#]kI�B�B�t����7�n���Ҭ:CԐ��;�N�9�R�D�ah}5e�^���`_8{����Bp�ĘW�1;?^\s�u�m�������|s Q`s�qIgZLL��J�Ε���~�":WV ��l�o��{�t�<����K��ه ϔ-����]��g�A��q���_�B�K�B��A���|������M���}�e)�a�WV,��-�GC\�G�5A�|"ӻާ�
���N`��W�9�N,�L=��1�Cw2x`�vy�y��U�ׇf�F�������=���q��m�a��Eg585g�[*nbm�`�;�`�8�k�-7���kdD�£c�"�{jh?ct^�ԡT�����\vޙ��n�Ny�c��NDW�kv������J;���+�������t��lK��MKO��o%Р�^�����>�j�0�FOǣc�oՆ!\YN��)?���G�G�������7�KT�A��GbP�L�������h��[�4�M�m/���}��\��;W��x�#�ݸ��ဩ�
���ȭ���{h�:�7ӟDؔ��=v�n~�cfkN����1���kZ�EY6�Z�����r� 7t#2p? �@���{G��L�8��wC ܰ��s�$5A���d��_@=�$���/��٨C�a�v@���BuYث����//<�z�� ��ȃ��4��<^�i��������?eqa�}���b����u�]&�7x�%JSd�/�9��[j1��W�'�粼{���s�TeRUkD�_I���6�	H�Z�V֣3c¬�ɪ42�Ay����֫l�J�����x����.s�h/-������܅l9L���
���G�2����GG�����L�o�HV��a�Ń�ӹO�;���͠�]��Z��S����|��v>'0C�e��?���T4�����x#��6���9�v�
ָ��vMd)sj�*M�����pS��n�!)P�c���l��'8���1̀!����T""��lG#\�w�ԭ�z��x� /Q!P7�|8!x��׼���~u���1_Gw�ڻ`}�q�R��=�F�u�EZkш��3���J��C�2G����mu���e�
�	b��n�$-�0S��(�̐�r䇚�)����D��_���]%� �7#q���/�4P;IN��&�=z<LBM!ĎD֞"iDݐM}{Є��x�����|u���'+�g��H�.��mr� ��蔦s�TyiRc~(�u�zB4o�N[��'�,[�w��Q0��oRG��G|o^�VU�m��ŏC�jm���^�4sGnOY-5��,�s�GcPR�_�q1�&KR�Q�t��3aE���j�|{��C�&\0|��`��e����}ՈBu�Vi�`)��~.���M�?%�I&z�k )d��0�=rK���Ë�K���\@92S�O8%�]*_ĳ@�$�A>�|��!��r��R���s�9#ej��oW��D�Q0��'q���d�zIf��K�_\6���4MK��1 �6|'���Xm��|��a��y�ۢ�X��꾚�������-+��l6����P�i�	P�D�n����>����Q�*@���#6
����=�L2B	�Y.x4�N�Qkd�O&\08Sk2�n��L*6�V�c+�-�@���J=�w+m���q�?l��Z��Lû��?h�ȵd\����}>N
N<d*T1���̌�f#@����ꏅU`����0l}#e�����9?g=tRf�H��IDQ
�m`ΫD��zGS����iч�{��4*C�6i?v��Z� 	��3�m�h���X`[a�A������*�M�Η0�/��Ȼ��_�p��ٓ�u��|]p:�������ߦWd���8����oL�)����hZ��̛tFxp�	.W?�q�r��x����l��
��ｈţ��)S��է�8š4�.��.�p�0�\�A�Ek�֭t��$���;ܔ��V�(����N���^p_��c��6�V�c��ױ�|A��y�̓��a���ҷ��W�b	@�Sr[�{h�*����h��"��qxĝ�n|�
*"m=T�/nEf�����(M��:�ʢ3����wN]O.���֡�����Ma^x�QP�\~��Bma]۔�1���]D�ji�_^|傀�(��v���Z=�J�߭��Ӓa��w���J��c�ӗ�w7{Hm�+j�[��}^���ݡw���޹����q��c�&˳���7i(����S(��/11�!��`D�F/EW��'�ֈ�ç�E_����S���H)�a���Dά���TەEP��_�:��v!!0�V���X�#���f���y]�t�u�.�-kQʟ�Q�E��h��_ \+�Sq�	�>��-��^�EP�U�n���87}�,� �T�ب��vdB���B�b��ڪ�6�:�g|��E�$ћ��W�;�*�X%�Py�$#�֛�=���Y�X�g�{�b�9	�
��95+l�se�q�%�&���)�JtX��Ox�,Sc��G̊�[0�d��;.F�F� ��z���Ё�(�^��%p�;<���7�y���@��^9��ߚ�w/�� �$�P�Bl��B/�ⶮ'�@{zbK�f[?�|��I����ʽu�G��^��/:~)�g.��k)V���U��W�E��Rs�f;��<܊N��؇��6�s�=�����V����y�2%e��Ǻ���x�����ǈ�h�?�˘W���s�����d7�"M;D�� B�Q�T}���������D����m8�d��X�$%�\ZXJ9]���>���܀֦��*(����eW_��p̴��m[Y�6j���]�Vn���
q��;�:K�C�'�2m������B7I�"�Y����n� gOj-=��kS�K�CUiW>l4Q�='P(r��_@��â��a����6�Z�[��Ch:����X�?٪�d&��!��3]�|��ȇ�?��X^��@tP˗/��h��oI��s���*�_'%q��^�nQ�b�a�s-�#�i��V�?�5f:�#�`NX��*�%�r���ɻ�WxRW[�|!����@pu��l��`����2���y��l��Y�p��s��"�&*���D7cKw���V�W�%18%��'�ҧ����F�5��<t!���r��t1����w,Sz&�]PX�ۖ������"�O�=`����'(��E�{��\�ls��{��G'���p}pV<%����X:���ȁ�̖�Un}�����!r޴�ߋ�:y���#h��3�6v����NZ fx��h73�rb7Bt��VH�Ha�޲��m&e0x;�ъ8�4����Q*�p��,���f��|� ������qδ4�u7���:�H�gm�(�������iO� 6�������,�7�d���1�m��*�{�TE��z��)Qq����j�d��D�/���*�Z����ְ1m��܋	m����Z�w�|�9d��Lt4��~-�ۡ*�f��rZ��`v�nB��aǚ��a�Ƙ	����`��ԱLc��~s�\��"��q,F��HsR07�3���G����.�:Ci9X��B�+��L	��.�1RO[�3���*c;�m���;�C��^����k붲=Mi���$��uy˟kV#�P-;۠��[�� "��-S��A�s��d�~?���ֲ_�9�P;�3��c��s��?{�a�N�����"#�ב{ʘ���*�������xw�o]ޒ5D-�nI��>'��2�$�*ܳ���)	��z^�[N|F/W �P
���]��&Øt�~�0Y�A�8�Ƕ��ɼ�w�ͥ5f�
D�' ����e�J^��eB+�G���m�:%�H��'����.�I	�Ƅ�B���s�)jq��nl��E5J�VBAFNU�M��e���t�t���Ĺ���⍯�q�Wj��EA��w�Цp��R+A���(�ҲL��K��O��L1�mYj�l�!pՓM���T����w���v	�z%��y��&�AY�c�����u���MoN�;l�r5|�M�F�\��e�x��ק:��D�4�Ѣ5\�97 �'/ ���;+��Ɲ�ɺ?qгU�/0�^v#�QЯ����.��KF������P}�s��A��6(l�w�@�r�cyt'8L��w]���GA
���'ÖJ���d��c��`�y��E����rc3�@��5���}��=	�
�'���1���o+ʣ����Bd�n@DS�Pe�9�|����Z���cPi��{,��4z���� �-�j*.�{���#�������P����d�ܘ�q��&/��
$
W�`�j�;xB��$��J���(g-�9xo������!�b
��6����v1G�o�"�$aW47|�T�n�N��Q�3�R�u]�焜�P�L�_�
�����򇈏����]�������Ǌz���LU�Oc�!@��6��p�"@�mP2�p��'�g�G����2�N+2뱱�(]5��t]`.-N�2\'�H.iۆL�P���P�
E�C�v8�
0��)iI�{Q�W1C���Nwg��k�q&�O[��Es�A7lک̦���K�l��{��F���(h�:6�6�����B�7�����{�F�o�%�s�"m5N��)�ԊzD�Ɖ���">�K�$2*��tb����jC���®CVa����þ�jT� CMӖ�aqN�����;�+<�~v:�}�	}������%zȗ	�������`��w�=�ڿ����>7[n��hw�=�pO\x����6#E2�K˛�Ѐ)�j���)k�5C5F��zE��yȤL�mޭ���9FJՁ5I�ф��D|�� \��0��؛ e�q�D�i	�W��1�Im �4X\QS��R:�<!�JZO�I��t�����Y3Hdp��Ѯ�l��W� �e��RakQ��,	�s��e������;�2��UP�*Oj�P�0��=m��o�{I!e
�Ԕ0�<���R�	bk�7wv��V�]�p�p3��T�^`�6*�~&ו�u!��m�|��F9R�T�ӸI��TX_��^�v]�3�A�	W4s�Hrj����r�[~ԏ�6TS�4aJ|Qq�w�������6�����x_�1�1U9_��w�TݝU�|:U�1����Yҷ���ȱm]���$̼��Z��_8������n�d�Oke�c�3x!ß��p�h4��}\Z�s#�D�l,�Mξ�<|+U�p�v�Z=�I3;(go�5���9�=5���C�}�.��;9����+�e�\����uP�]�'�b�uYq �}�^�SH�v�^�{����}qiF�ǄK7wLM�%;�I[L�{�B9-r9I�{��U3!�h-կzū{f3`.j�K�E��� �}�_v�]��0뛎�4:�M�$�fX�QXK��n�+���^yY@���a���#O��=<lٕ#�З@���&�u�&��F!7_��T0���4���s�!�O��_tL��O)��P���L+w�=�aIl��ͦ
r�N�7�dV�ڄ!�0��>�d��I�@�c��e�X49@q�@BD���.<MN{f�l6��
j�ur�����-�L:BC�lNF��r� ��Y\)�K���!��?M_=v��߃��e������:���b�H�����@�����`�#���"Ǯ��?>�֬aR�*�"h�|�AõO��RV�lrB9��Z�9z�����9�o�σ�l����a�@�mvzޏ M�����L��8͛R��H����s�7��Oj.�a�?���x��[���jh�*_x�)G�M�Jd�:Ei����Ԅ�C��!YQ9'(PÐ}Ԁe�|���ra���@����)='��$���P�ѝK���l|q�shJu�"	�~l�ͨ�8+sê�y��_�E57^W�5��54K��V �H.ˌ,� ٿ��2`�bk�BQ�Yw��3�i�?��b�m1�ܯ0F�{���&����s�}��p�>w/�mRP'ӧY@��£�`x%W��K�I���sÉӲ|>�T�{8P-��Ww)_��젆���]�|�n%&In������D]W��/7������{�0�K�@ɽ���ۼw���O)HL��얉A��D���[ �f�B�fU���J�w'%�qg��Y
*acAI+HG��,����>�Q2�$Yf#��~��YI�Q���z6*�d��a�O�����`�)sB���N~��Y���H)(�'���AEL���~��t�h�����#.�Ġ���DJ�Y(�����1uaB��8��+{�!���T�-�%�O�"�5A��ɣ����X�����X����Q���ه�"�X**��"���@�y�� }x�aq�泐sA�"�N���)��Y�g�����S�X��DtA��_w�	��W8�'xm��,�޶�R��W3~�[diGU��K~!V#�Xr��O� ȒX��*-��D�S����f	�@*�D��f{���F[�Z�b�k*?o�h%#�KjU�}�����/�����2��d���kd��v}����g���-��H�-�cJ~aI���̓JK��;�O�,�_��<r
pD;=6#t�QpI���`k�H$����n���k$�Ȫ�fY��(-'�.:���OZ�4��bx0�ئ��/Ǽ54�Q�#�,�/K�'� ��>Ǻ,��2�Y�޹�?��Hӿ�����q ���a�1�B�8��K��������i��1�+�s�,���g��{�$�_����~L06T���ō�m�
���dЕ,��XuZ3�Ʀ�� ��d�*"�{�0M[=	|h �)K��2�4�/{��k�J���K.��<���0�o�����k��<���0�㫩��y��w���]\O;��$}������\�ڂԄi'�Sc���sxq���|�9����OC�7���6Ǉ�Y�	'��nn{$�.ڈ��ʮ�@��R�{���SՎ���5��h�{Y6��,��O����Q�p�ٶKD�����?^�����h�,���Gb�:0�QWHf�1��*���� �]}E�+pUg���r�8��îب���㩎�1����|~0
R�d�r#�(�q�&��7�Z� ��|�K齄�*�W�
V1St��������W�bxN���v�M�rN�aܶ�b##X@�64x�K��a�|!0��(��R�F�_�[;m����j��#v�5�p
��!)�Mȉ
Q75����m&��^�j��zC���ĳ�#�<�s��E�m��~�Ȁ�1Z@I�Z�t�
}O�~3�蒍�!�{/���ow#�o��.	*R��_������"b+�3�8�*J����X���՝k#kTQ�P��j<��~�?uO!n;%��͐<���������	��C�CE�\q�n�*sW#m�r$Zu����X����L��,�nXd(��x<.�������4zّ��)mc�n��<��:�\y$�����h����ύڱN3X�N�[��g2(����r������_�FB�Ŋ7}�!�1q ����JY	䉸%�����E��q�i�&U�m�Ub8)E��0����@�l�����4�"<�3ٵ�p6}�yj�+	Ɩ�*�L����W�}^��4$xs��>�V���GK�74*U��q��u�Q}#h�n,>�re����lW��d��؏J�Z��C��/�<���t��@�M��m�uk��	�"�UJΨǌ�cw�1@���c�]B�h�b	kc�%e3Ȑ�!9�Ѹ֨�f����c6k�>j��w��3kIT��^�(�m�ݜ�L��vU�m��&��X1>��/��K���C=��();^���S�Id��u��Ej���3�>���
��X�S�d^i]��H����[�jq����!�"��Z貮:�&:�D�2�é�G1Ӳ�����>��f�pC�$�#�(:~JH�I�ڀ�c�1�IQ$s�tقv����ZY��́K��p	�5���jM���E�~DÐ�eq�J��A���h`���(fתR9&	[X7Pk�,	�U�a-I���ҟ]M��M��*��c���`�A�M�l�E���_��S?N�����5S����F�䟆����7Ú!��~tX/+��O�?�C�6:3M�b`-��:�J2-�+�:Nب#ꠎ��O�yܦ!Qf	`ϫ$8�0)ЂXN�Jg[�W�	��B��l�a�;"�k�l�E-\Jb��c�ϊ/��!�J�u��o2���S]�'�ft�V��4��\�&ǁ���?�q�]z�[����f��t�6�3:�[�uL�s�Ejg7�ا���Q��7�n��Yo��B�TZQZ6-2���U�v�[���B�ҪgY� Q]����㒼���0z�����	�J��� ?E�p����!O[�[�����Cǥ"G�JzQ�/E"�@(3dt�ZȒ;��F�N}C�-���x�����m��(	+��k���,!cq?��Z&�>�"\�s�c�9F̸��av
�D��o�A����!�Hc�`�?C^��!���&��jW�����B8'���f�:��M��a�^K�`�ZmN�n����x�K�^�q-�ހ�����ɔ�c��x|=ӭ��ڮQ��3�e/_�A�
Q���l�]���_j��	������`�qu�#*�Úm���ݧT0i
~����D���6"�	Π���a�K4��3�n�i���4��ɐ�n��H��'�"S����u�
�{�Dj�ɠ,��+�8ާ$��KD=gB�h��FD�'�&o�@��0���,KE���'��/�R�x���
��֍h��K��ɉň��z���:�ϹB������ѝH�u�'x
�m���3e{6q�")�v%N���>0�Y���V�3R���;��E""E"��W��{�(�8Q~u��Loˮ
Y>B>�v&�������1�d;����!��Vh;�#v��ٱ��l
�%0���m�T���p9?$��^�P������g5�Tr�n�s�W��B�����P��\�h�K8�r'�n�	ch���r��J��P�9־�E��oٶ���t/��5��n9On�|���<�|�U��ʌWC��9����)i��������\V]��Ko�$�rO�^U�2�/�P���cd����@m��}�ϛ!S��c����H�ˉ%����LX"�㩸l��jP/��.����L�\��h	�Ҋ�ɲD�A$W���w<��1�@�9��'���ڒ��`K�D,�i�v�mr��,2��1���f�$�����t|��V�0�h�(��%�2P+M�TY�������x��ӫf*�Ծ~���ῡ��2�kr��L�5�A���
��n��M���6�vU؏jeVԸ�&#�3VY�P�����C��;�r�8�]���\�Z����{
"�&����Y>�F�cp�EPz��ν��c�҈	������I/m�0z�i>��"��)��xJZ��m�4*��K?Bu�|CK�O��vs�#� З���1������-���)ki/��f:�K=�q.�p�?M����-�H͙%�O4[�nsɵ�>�D�ZLzD�*j Yn�G7�� ��9��Yf��O�p�6��t�:���-�͹�������_�~��Ϊ��ue���5k(�j���)���4i�0U�-�'=�o�W>>[
".���*e���h��=GJ�/���Vt�>�3@?j��Fb�����+����$B�����u"�")���V_���/�H�k6�&(v��N�.O��� g�n�_��� C6�5#( 0@S*��c(q
F��0���U�+!�����)�N�ڎ�:Zt��'H,`��V�9qgόj!}�FjRk��dَ#�O�5,
�KG.JZ�ޡ��X� %;ӑ`�D�-�5��h��t|�ݡ�A��r:�&v�I�IFq��]=��]��YR�M}�*��ǆ��xyfOa#����.���v|b��r/� k`�H�&6��ޗ�v2����{�Fl�}�5s��IH�$�ǁi��Ȕh��%'iض8}]��Ҍ��
W�[�ؾ2e�$���"�����}[\j���@
���������\
 Q���N���b��nAR�%i�#|P�>�}�Ƀn��i=���sy��n�ҹ�$"�*I�Sl��&UN�B���C�-ˬ�+�[y!�RM�u,@�`¯�7�
�IM��$�n>D����;yx��\��.T�s�,�m�k�����!�i���Ψ�7��g���)A���)��	(v�Rۑ�ŭ6,Kă�)M�
௛a��Oo$�N�&��;g�6���;9*?e
���5Y�4�����ȔI/�l�I��bZ
�Q�~���ľ
G�A�i�)g�,3X�6.)�����l��ݑR��nAPfBo�׮Vl+��v{iI���/��NT�^L9�몁}/��nx��'-�Z�D/{'��ݢ[�-�F���(��f�p��KW�Fq���d���VJ�%}��)��m�湷U��D�"9�]�j?��*���v�N�%3�w���P����n�����V>���J^8j%e�Qj)|�g�DmQ�'S� �:Df� ��%��U�5V��3��xYWM&�:[�cF�3�ݧ��$i1Py6n���\ؖ�`�9	��5$���K.s���CYKŚ$���#g�_-��M�{�͛���k�gB����<��z:�D軣�έ�++��\�lw��Xk矎�=L�/��譁�9A�f�y�Xق���6�^@�	�oF0�]���{��o�������-?�+K�Z�/��Ol�->�=&(x�ZZ�>�S ZF��c�"׉�=iv�F���>(t�p�9u�֍|D��(=�!�E{1T.�D�D��%�l��/-�r�f|;����ph"�_k���X��$�;5�{�"��P�LLd8*(�|8���1�#a���Ȝ󷐿�+2n�CƷ�6A�6&�H�\�S����^��B��9 ^�0D�=��#�>#��@�}��`�����ghؕNt�Y�)��SNX��1�I�*�����5�$/����
dwLi�ّ�;���ۑD���k��V���^/J�m�p�N'��y��לwAiA��u����w�+�{��f0c-/n�+��J�PO����FM�榚8+]�bp.��(M�^o�u&�ln+=�}��8��p~1ʵ�Ђ7�uA�8�������/�q�lM����#�䰦�o����X��J���k�w��=X�D���U�(��w��r+ ��4v�d�
�RR V��Ч�_��=l�'(_����b�����3�k
k1�6��A�;�"u�ԓ4qK2���<�6��Q��>׺���څJNEݣ��!\ҩ��}WGl��"?0��kJ�O���R�K?D I��}�s^C�v6>���&�^O�G\8c���v|��+������h>J]s6���1Ϛ��o��Y�pJ%A�<��$Tp���"ȝ�H��z������n�Jʥ�7%�U�-I�e-s�@�mn��ʇ�O��c�7	\ni�Od�>�A�vt�䊑v���"�u0p;|��<r�"-����6+�(=y(�����Ĵ4&4n8�P�J[�xEo�R���z/}SM`�T$�U=Z�|`�0���<O�v�ĳ����@Y��֮��ب�|Y\]�s�D����:��:<@��̻ׄd9.\��G��9J&�. 7(O���܎ЋY���_��IaG۪�Y��+���=���*.Ǎ�������c�<�,Q`R4_��Q����S�9�}��$�!�h''G!�&+i"�P^$���}L�
x¦���!O_�@������C���/mBF�Ȃ�v4�)�7a\D��Z�ML��9��f��܋��r`��c9/!�jp)�I3�bTK+d��e�P���t�kV3&���L�$O�'�� +x�ᛦ<�AO���`���,� )�l����
�����7-�׫���UCE����\.�Bn�t+�V�yCq��"�iBۋT��o�:����tl޺>�|��I�Ȯx��}@��+U��QA���j�Q�%�(3��� $ꝩ�t��4˰Qɵ�s�����.�'����@�N5gj���z�Seʔ�U�0O�=Q״u_�Θ��R�C�3}A�z"��BK���n��А;i�:�Y��n�ʗ� �Mށ~gVh���=U�#R�(�W��D*��"�;3-SV��p
T�rL\��̈́e��OXpͻ=IӍ�:2W�^�y�1���j��.���C������T Bx��C�#�3��������*Q�֛NUɥa������Db�;�ǫ�E��BK|F����v�B6m�v�(�K皟*$6=ĐOS�i�o����h�8{��ٺL����t���E�\z���_+��ǥ	t �x��
�}�3���8N�r�;���xt�]�Ο�Έ	'`xzZ��G��4<�}LF�4��@65�m�$��p5y���
��@����49�n�U�vi��?�"�+��Xi4����Y�������ѐ�e����:9~��}w�׋k�+R0�+b��7L��,�\cqL�n�gD�g���/PX� �� &�]�gI@��Dw�`�(Ǫj���r�RB+s��)S'ئ�β�-���~��FP��5��ാ���U����~uo�q�Mf�w���u���~�}Ͳ�l��%-HB�=u�t�7��p�4#��m;z����`f���d�9���*�ne�M���,�����5Z����fM�(9k�HE�e�F�X��gq40��L9OҢ��59&!xM#A�p�snq���c�I4ں��4͙$Wf����:�V=d��Y�Q�a�=q˃W{d{n5q�ܑ,]7�`��Fm�-����\���^ʊY���?����9�/�~+ Lj�4�mѫƈ�����ĹF�݄Q=:�f3]�^���S����ܴ)M+�qO�ײ�@���VlJ8�y���y��>��i��͆A}���#3�?���>�W[K&�����e{Z5?�i���W{:����|K X8�Tد���1��{Q�:��ٸm��j�4?��}e:���]D;��o��Ϊ�M4(���K�+x�Z$�`i��aj�@F�V7¡*p�G�Q �\�R���H�q�i��}|�Z+���l���/�gc۪n?�Hw��khO�[�z;~	�o�vq��	�|�RT~>�tn�GKL�'�M��]^ ��,jRg2*������Ɲ�: FG��[�(����Y]y���l���u�P�ŷ=����a&q^���s~�\w(60�q�º�Kx������ą �~�gA� s�9�+�h\6� �V�!ί�w�DO�8k�JWt�\�䖶1���l��v㩩�v��q>��G�D��Y����48�M�8I'2)�{����"t�� B��r(�wMM��>����9�k����'@A]B�%��+\��v^�R���:ק�<�.�|��K5� �7�k�7`�?��쌓ԏ*Ѡ:G=�:���w�$C���w�*j�Ѷ`��ћ^Y�/��5�M�:�l��ЕS!�����?����RYoZ���A�P�U$�N���Zk������n����7)�%�G^�z�	���Q|���{����`�h���	�'�(� %���n������xC>{8j���6�CWXe)��>��@R����`E�'0Q�����^JE��>��q���S� ��5O+��I��r��-?��PM�nl�����9�f*��C��`�SΘ�T�@�vzɅ<pC��A�u/wOd'�ž��a�L�ӑ�_(Ȏ�Gc��
�+�T�UҢ�B�e}# �� ̽sv �M���&Ҭ�����+ɡs�!�	+��~l��F�I�c�o�^�(��Vi܏%���/L,R����05��~���\�<4��,w�d��f����:�,/������Y�"c��=�֯X ص�c!���=��KJ�7����o.D��\zi��Az�� sY�cKM|jG���``uR���٣�kҋ6��D��ʨ�z�c�f��〵 �H��. ���~d��Yx��Sd �m�����Po�f����+���,Y"�0�~���u�C����^�3��f��.\����Кy9�#�����Z���R@������V�[D�E|��/Z���Y'�ݮ��v4o�-@���J�FX*�3�z.,��7��kH�.HԠ��\��x�߸$�=���s� ,XK�5��hjX�,��|�-�ίm�.x�FG&�mY����iv���o;k�)��R�+��n��A��F@�{9�� �qvr���$j�*�q��B��0��(�2"ս�Fj��1�/a�/F����%Q��4s���q.5�*'���q�cII.J���G��y��X,�&���ϗ���%��Q�y���f3�ә���)Y������`7 �?������D*|魷���?�`��	ڄ��d�;���q
��9\��CQV�(e��<�zB��8�w��/7�tI5�^�j/��g���P盧���ᔑ���9�bYR#B��
-ں�E�hP�UFme�\2Oظ�c��;/}�}P�Q<��Gt �֍Iƅ�\���j��Pڪԑl�܄��}�P?�xX��\�Oy嫼�(R6Tߢ�= ��5jJX��9�}��2���r�(�E��ix�IiDJ����������W��Y���/B���L�w�����jtg��N[(��D�M�����3�҄
H #&62K�Oj00��M�U��5y���'�ʝ��<�e�{����=X�ݗ�-ϱ�E��ꏆ{]$��{�[�*3�蛿>&"�Ha��/���EQY�Pw���!rrE�����mvb�&G?r�@ww2^�cK�"Y�/�^Z��ا����+'�a�?z~��3e12����k-���X�TL�}���S}3�����j��*�7¾��0=�T>4H��Ě�!gI��&��W������F��1'���&����(�,�,�/�垟��F��� [��C�����m�틂�J�,�t��=��"i��j���?�pe��x?��+�$����K��	�&�����)�{9�ʭ�:��7�ڱ��z9��w��u�L��0RS|�BB�������c*b@N!��@�W�'"C�_�I{�{��.�\m'���R�ǳ�f��,���ߣ�)�߷�I6ėp`�Т�g�o2r��j��Q"V����O=��mP����Jp^ ��N������$y�.!�M9E_�ZbE�H4m��ˣ��x������1�3f����?�|)r�D+j�M��g�p �.��#o{�,"�Y#i?�-/�s$*���b���_3�Dրc�ۜ����u	�=�>�~{Sv"tVe M���,>-Ym����P�64G����z�7�=l�v���:CLw�2��Cg��v�ד7�t��#�㋸�Öe�-��"������4����cu�`?�FGl��A��˥�{fI��K�5Z>��!!$�P�u�-�����0�����A;T�7����6zy
�J�Nv����~"%�\~َ����Eq���' X:�pwZz� ��ϫ����_O��JΦf�+�@P��)�v��rkR�5����oB�мk�eE�x0[2�3�nH�k�ؼ����=�G ܴ:����a�it�qܤ���M(� %,��l)U
���i��R�mAuq��Z �h��[}����;BU�Wg�D7.U�X�
�{u��	#�~�mO�5�(|F�/ΐW�����aNU� +��y5b,�܅-ٱ�#7$*���,]��R��:�al�V����-�:	!ۓ���ڦ>�������dW������ח�\tvԃӐ�9��>+��iW��r���ؤǖ������!�$�'d���X�|W4*�I-!m��5�������_�����E��
����V�'!"h���	!�<B_��<']�N�D�oX��%�k��ٿ�����r�3La	��2�O%9z���vRL�:a)���hHRfA��]6�ص���b�M�+3��Y���T��:�|o�3_�����EEOv�|z�'߲��S���d9|C�imJb;��Ώ�	,�.�	^U7ż�Pd	&h0��F��3[��U妶k�$@�N��̹6����^Xr��+����i"��P��F��V��̽��zSA��Ǝ��ю]�Y��y(��U��}�ʗ�����������v4�
e=��%=aEU��*Z���n��-�vg��m�HH/�:�bx�G�����5l��1�(Srj���r�C}�:t~	[F�-�%�ts�;sE�Zݵ���ZI�`j���$��D��@��~^^�ޭ�ϰaa�蟈�D�ف�Hp��I:�5B@�u�J�;��Y�6��Vq-.wD56I��iS��co�Mr*M	�".K\��5��q��A�b|���ރ��$��#2tܩ�O�r��3��z�������[NuU|1F!Eܿ��y��P���.,�E�r�DNp{R�	�]�~�5ٚ_���E6��y~X��p��yЧ�;Q,{��*��:��?sCX���cX�O�d|)�@��;Gt��p+��=�>�1i��Zm�ID����7Xs�N}��#d�W�����f���4 ����9�6'�R���f��glY�ʾ����P�A�.��_����R��t/P�����G��V��Pdԝ�/H��n1���!�$�>��1l@���	��@n�S=oeF�K��Dn�v���E@4�-��6UWS�q-Qs���+�@R��\�rq�Opa�S����ތh$K��KqJ��J��v�����V�����(���(���Ǡ���_V�~Q{�����U����d�� ���iy��v9��G3��j�mU_�V��	���\wɧ�"d�5����]�Yx��))[�jKT���.�q���Unx��A�X<Ef�Fq�PR�	�~Iŏ�n�z�=28�0�x5���;!rZ�Q(�~?��I�K^ӻ�6����|����$��&�.n��X��y{'c��H\����O���L���20wZ͍�SP.'w��]��N'^\�{q�����r3�����R8;_j�ZgJq���8��蓨���Lm0�p�V/(40�I,���X��8t��@")[͕9�I��k�!n����_+�ȩ-��SЇ<�����#�MƦ�}U&�ݻ^hpv-oz��X&����r�7n�#���V����v����&�J�;9�	��E��9qr��T]����QE{o�v��9C�:�(���,�%�(7����na��C�Qp2���B�e����k �^�'D�L����m�d^C��g�A���N�a�d`�^�H����I�Y+��V]�����Ģr)����h/ ��a@���YBN>�Qv���n�y����E]#N!]���1(}�m�mL(t���WXC�	�����K5���z�r��6��6{�}$fp�t�ni�,�$!�sPls��/�qK�e}v��O�.�I�TA0�y��o�,�D7�@��\.?��_1ƣ��K���
i�\dqZ=�:�4�̮�b�?
��>�qOs{`�E�p���L2�*�*<�ef��H����(�IC��P���	�u炚B�K�11^�:,����,��9��ֹ��+�	K��)t�0������<���'�� �(r�qPY6�m�*۸�ޙ.8����[������SK5�w�k�T���t/q����l���gM*o�
=fW�_��Bk�M]�������!�3�k)�x���*&p*`�����/P"�͐�O��X����-5��4fLX�]�3+iQ�2I�eM=���,�|*���f멻c�wA����X�קw�rۯ�JNh�;�͘�ۥ�\�,/B��A�֡X�
,�3>�(J��!iw���I�zJ�&�O��;�ӱ��Y���!}1�1��G\�� ��;H�I z�\R$.Hf�-��R%��H�A�q����x�0���zb��VU�����TOk��PK�ǣ�hj�?��a�#;�i��ȏrء�6���(�։�U9���ԺEA(�31����,Z���g87�&v����d9=��,YP���'�	��<P�������.%������)|s�9i�/f�.��-&?�dx�F?��Gs�U��f?������TMGu�U^+�1�­�)��W=�&�D����
��V�����7��M&S@\B��~[r;���yx�e�����WZw�";�]����ˮ�W�]��܋	�#nN|��C�I��6)F����-\�H����nԋd�E�����M�̀�N#��e��w�q��I|\�aGRs��f>�{���@�|���?�[?��o�9�� �NT�{�^J ��7 ��aS�P���Ѣ���Ǳ�M�7�x��%qc�ǔTQ��	Mh�"��c~3��	��N�p�-�a~�]�o94%��;K|J��m����BP����>�Ő|��I�F��ᡔ��M4m�G���`㯶����0����C&�J!��;K�J�_,���GԄ?�Y�	}G�J����ghra�m!H1�PdBP��Kk���j���iq�S0f�
���T9-Ҁ�:�����cT�������$m\�#L�d�|,��6��K����N^b�7�i�(<3�J&9�T�ۿ�=p����k	��%�#��G�	�U����恖�(Wz��C�i�9�=���8���~���_��?D��������rپ|g<{�(c���&�����l_��X�Q��%�e<>�k*m��n\ZՖJ��4=����8M�77꼹 b3�GGBM��77�?_�+/��8؂�C��58�mVBVd��;=�h�%k&�������������3�!	�ޒƼ��6�k�o��s��V��>���-}1��{_�p�x�_̏+^dO��-��!�m	\���q��o����'S��]�yۖuv��ك^M�sgz�i���WfsBe.X��!%���Z�c��v[d�W��޵R�\����*��(�2g�R�ш��c�I��6��b⩕	z���G�������5�ő^I�p���v�a���6�0?�+�t��9K�l�HeCՋZ�V4��ü{�c�u�n>�4 �dږ^�/�5�eU*�&�˻���(�3���4ٮ�,�Hz�d4j�b��]�Q��������K;����i�PO��vV�� zU5�g5�e�ެJ�
ԛLo���B��'�`'��ql7d>�G^7���*)�+-X�l��H���Hu� F3�Yy8@�e,�fgS&+�˓v�$������}g+�D��ex�9{�J`�#p�/i�����+�T�䲥��=���z*!#v�����.~���A"�37p�F��P^�꫗��={�di�$���wm�.����0��'l��Pfo)+`G9�:I�k��w_~5����B������¢�����NZ,�f`n��E\ј�_�'�3�&�\�sH;���!M�_ԉ�Z!k����N���&XlX��r�`j{���"��.)�-�B�<A�����vD�~���SӢ.z'J�r�F��䔳��ABu�6�z|i=��훌T	%2��%4Z��>N.M�V�JLg�b���ȼ���ӣ6�ׇ�\eU��ѣ�����򧏨,��bB9n?�`�r���Pl	i
�m�����&�<f&> ���p-�(���(�Z}\5�@�!�¿äh���78a̛�Kӛ���ɂ�Doz����΃`���]))tp�{ݩ��-��ļ�sk�8��9��Ҏ�IG���k���:�$����~h���D�V��_��'A˶5㖶�}ĖD�M��"��M�C�����^_���>o1}���a�a�O�.�|�ē�P�w�4:2����!C�e��������eF��uwZ�I���ﾗ����7s ���*���`�)�*�#��(�Z.-���� �n�t��#�{���%�2�]��Q��]�
�,�,��X2e�5�ua쁄u<ۼ4M�W��T�,��	q#bW�l~�2��*��J�� �3����Ï�4IO)UL���uy�0�YeC���'W;�d/~'a�Y�?���h9��Op@�7kע�uL,�u'@ fvI �	uu�1�k#9��+{�V!�kw�:�><v�$0^�z'�I�����|�*�	4�.<_�uZgx�f��a��8$=��{�*VC73��B'�է�����Ť|��mo�儙#�Yh�9b
��QA(�-��&K���O�Aq԰T=�	C��,�-X�'q��`�k�8�N e+0��s�j�T�[��\�l�_M��¶@�fKw���Z�*1�=�/O��N���Y�2 a�k���.¢?����lH��f&P��d&i��p�E똕?4��^%�uY��V� ck�����,�5�*@i��l��PO�K
y�S�XV�`�����2?潥�S����0t�Ke4�
�Z7�,.��9[Տ6��wv!�C� ���Q��m�M���A�I���1��R��oi=��;d�(Ve���za�K�e'�:��7�0_$��¨k5^&5����(��o���k����*��-�Jߋf����_F���a�z�V�ﯳl.��V(Lj"|K�?C})G-A��Y�\K=��㼐1�M�[.=�ˑ�;}�}γ��+Hw�@.Ύ���͇�ϋ1=I`Q7U�y�a��Xg>m���G��q�Q>_`�Y���űD�L�jy�Qv���Ea.D2I!΄�P^��Kĭ{�yǑVN�܀��ip�eR�L������׾�IG�v���.�ZGB�$3˛�����pR���@ �z�x�=FfJ>,��F�����C�@	��9���FM:a &���9"�{(��PM�(��öY�C����Ծ%�Դ�D#]� �*K�C�ZЪV�6��9pb�t�?���<�
i�d�,�<��u��gb�剈%)�� o0[�gځB�e";Z-��GɌ�o�3}/%��1�-�X�"��#��nmX2��U��ڸ�@�!+@Ⱦ���YI�eL�3��$U"bx�J��RxR���N>Ihh�s�,��2rKS�z������ҕE˷�,%
&si�Q���J^ڠ�8�N���	S1��@��q�x��'�����6��=�L��ۇ�nJ�%.����P����?�O�t<���0.��xY����Z�N證D�M��	�=t�s�{�ײ�Y/�g���ʭ�F�C-5�Ť���BH��r;F<�x�
�
s�_�8�C�,6Ӏ"��b�_Y`.���k�#��V�#$,�fB�fW�8t��$�R���B9;��|�'{>K�W���\��̮���.��?K�`�)Ki� v6Pv<e15"pRe�֧��lD!A��:��#��q��|r��f�Nn�>oؒ3p8����x+�x�oS�e%0���G���W����;jmD�U����_���F�Sy̡A/�,tc�M��������{�7r50�$�;�T��n���I��;��'ru#;�6ޫ��驇%UO@*�����Uu`I���ڒV�]���ℑ�y�,s�N�(y9����~�$���/�X�����,O>�n�m��[m'qAR,��w���p������<�s��j�����#��z�^������E�������+��*p���kI�.���I�i�����CUy�5�$n�F��˚�o���z�j�-��1W
m������1��>��y�Xyڎ��r���_F�[���Ҁ����-�Q��i�V>��HXnD�-����^~�o�h4+�x,�/p^�9@�5���&�Zom�x�0:k���v��6
�v���-��H� &���؟C�ә�$�P���5�T��犨�#^?�3�ۙ}�=���u�Y3R+?ߙe)�We�>g�G�{S��|K�e{�V����dv�NP�*��Q�7��92oȣ{��J�f�SꪠsX�)�1=����~�s~�<"lpV���(�vJ�]2�ϩ��ҭVt<i��P�WP0�Du� �R��~���1��Ɩ3,$~JP&�g*�<�M�vD����Z03 իG[I���g�z$V��̩����J��^z!#�Z�8׵e�Z:���oT}2���wr�j���B#�geU�t�$ޟ=y=0��u����G�9�Q�aa�B��2�RμC�����!�!�_���ld�AdZ��n����\�a��l�4�������J�f���Y~WK��K���\i9�T;��5�ZH��� ��O1bE��S�zƬ���E�A�S��3�'A���5ڮ3l۹��J����{i��>��������oL2&�7���_��,(��,;��?P6k3^��я�W�p�!vV_���֫��>��j��?�%���9
?9�՛�yҸ�㋣^�#K�s��
���~d4~�>�����aޥ)?X��w��GK*Tu��uȅؐ�,��dR5\�D�n�+N�=��$�Y��,gp�x���Vc��Mt/�%�N\��p�����|ﴤ�o��n���[�¨ď�eӿ{,�_gHh�kS�5R� �N��9���U:���!f�i�٠�C�	I�d`<�p*E{|6��'X�������xs��q��Qf�7@�O�H�!�Ѕ����6&h]_P���T��Y�����܆�;����i�@~���p����Ǵ�y��7�o�x-��>�J<c�ZA��{�[��:��V165�P��]�F6iwJ���*�s�O�wjF��nއM��]�X��9�n�r�N1地1�����2~Xd�]��n#�J_��s9s���\�ؤ�N�3�ƻ>
�8��҄�	"�ǻև���M��T���v��(I���@ ]���u�:ϳ��{~�+�;:�|���QR7��zA�jyut�b^dĎ��q��h���@^�6�[� � c�ry4���Q;�=�o�+E���|�mߨ�����<���>@���]9qn�g�}̚r9^A2�6�UG����R~|N|7,�9�?��8C����*����خ :5*/ιý)q��PWмZ5.ߐ!�10��	j��i��w8i#�U�d�:Wk����}]�;\��=���l	e�
6?c5KI�S����� 7����f���Ue�6.(3,���0�6_[�r�(;�@v;fĀ��q�.�������-�/9����܄_%��>�%+(�yb$EY,���p;��r�̈́�C�"��LF����ݚh����UG�����_��Ui{i�����b% S��w��s�u�^b���^�p"�a7u7�W�b��nA�.����F��ZLd:�P�]���#,��h�F~"�%Z^��P�LV�~''Q�
���� �=���X�T@�U�6�	��(k�����������ϊ@'^��9��OGS�F(Sn��Aj��
�|�&$��e�)�z�z�	��}SEԮ�C�k��t{��b�VfCD:�'�W�3�S^�V�vŚ���4�4���׀+�7b͗���E�_�قH��U@�c����տ"}�bCj����M����"������J0|���G�vY�!�)�I�Y9ڬXq��I������=B���T�K�r��Ct� |4��@�n��OZm,�)A3C����c���ʎl���٫޶A����f*l�Q���v�ҥr��S$�x���o?�b���_��	3�K�;�)4�贌����������ehӿ��q���V^Кq�H���	_����\	@+6.>����-))!yb%���]&}\��s2=>����oK��o6�ڟ�v�r�[��q�SK</oގ6���Y����f�}�tO��EZ|pp6=m����&�9T���/�z�G�}��+��O|~S��Gi䑨a́�\�Z�����`r�f`�#у�3�����[����µ{ѮL:�z���EXY�\S�U�n�K����!v6lF�����<q�(�^��_�7��򗎿A�SU���@ϲ6�.ib2����ᕙ.`[�C�
�KP����,R,�ʛ���m �nA b�#&�̕Q{�4�C��6�n}U�å��-M�y!"C#�\ǥ���)|���jܴG��7M挩�æ�z�@�ƶ�ENov���Vi����v��Z�=PH���Ƒ�i����Z9���fVX�ç2��(����W�<fk��ﳋf9>�q��K�̈MEdf�#yD��>j즥��c\���Hq���ܲFy�2靓�
�,p�]��^PRg lz���ۨ2fIxo(�Ę��Du-X�8d/�~r��E!�xa(���,�l �zF�����K�� �7k�`�������4xú��h0U���e�JV8�n�g��MJ5?ğ#�KMFn$���c`�Wl�S���K'���ן�/���p놞y��|}�5�:)e��HQ����X��?X�Ԣ
X*��o�8��R(�U� Z��}��N����'�
P�Բ�mUQɊ����Wy�n�$�2��㒓���D��o�;�
��s�!g��J�5�0)���\qJpBL��PGnN�4m��n��]~��;�<�Ơ��<�>k=�d�5�X����ȳ�R��}!�5� ��A5���:SN춒����3�%���̗w�L�ݮ�<���E�aoVԿd���	wDy	X����x�圄BKU���/�<��ۋd���1tI�9�q�'����{�`��ގcI�#4�Q5�}Mu_`�c�V�Y;zn_������mM�ȶ������tz$K��aqs��aC�4q./l&)9��gі���-��n����^�At;�~�ω���K��$L�0�&Y��oWY�x��;�r�7Nǝ-Ú)���	���>����ɉ[��ݷ�L�.1�+ٹ!*�'�ˍE��Y�(l"+$�-���}(����&�M���������_��P��<�-t<� jx�ʎ t��U�a�J�}�-EN]3��B{��u"�z-R�P�l��v�cP��L;M���&/e��hi�ٴ
����S�$۔4���5���-��a1f3���. ll�����&&��^�$����W������3�a�o_��E.u-بI*�v��Lıy�Yf@o�h��=����x���F9��g7|���I���� s�}���U:��oJ}�w��UUES
m�uHKGhyN�BԴ=��T�O&I�4S<�hN��3h��lՅ�N_Z�Vh4��XM�Fq�FQ�.��r��r5�ݿ(���t_C���EůJ"Ϳ}��4�kt����~�E�*IX�7�CRw��"����h2hi�]t��gn˴䃹q]�T��Q"0�vo�s��Z��r�Z��h�%��聾(�^uN]Yb֨�t��q���&�����:f���F,k���~l\>�e�α+�ӹ�x�e��X������y���w���G�馯��M c���E$lYa�Xaq0��BRz	47?8�TG��P	ٕ3�o,�ue2�?#c�Uܻ�B�_z�1(�~C��[p	�s>�?>��`��Tw��]�(8A����PHk�4�e_J=l��+������ ��" ��W�`��r-���E(��]J�����:l��:q�L�(���G �>����F�����h�3V0s;�>��YSĹ*��!#'�x϶b��o��ƙ���ڤ��r6�{-V�vb*~��`���%�T��y��Ы���<aQ�%B�m��88j�� �(6�~���<5���9{�����<�@��
G��lO0��$������"�%�Q��EG��T�U��o���!�L��Y������Sd��J� �Edw��۾<O��'�2ȟu3�6�����T�O�fS��|�~q�W��e�W��e$�̀%�_���(9�m�¯���m�e$^_*�>���=b탬�$�,�0@���w}&r
�3��GZx��"����?�Q��HW8�)�F���8��Ԟ �v{��F�D���gW��Թ@�&:�`z�z�U5#:P�a/k�l�Tc���ނ6+iv��±�2Iv��C��j4��$EE�:s�$ȸ�[���1�<�����
�
��i�8�����Cڣa��Wn~0�f(e����� �e��Սp[�a$=�Z��h���\�R �1��"
�גe�!3~�ꦖ�s���H%z��F7 ��	-"�ٯbp�<�m�H&��\�r���}�L�ơtA2H��T�:����ˠ���g��Hʬ,�D��%*l�4�0��NT+�T+���Ђp��^�W��o��膋���#d�α���n*��T��0�h����i��* /h�Mk�ӗ3x��U��Mc��jaF̏k9�\(��Y�)ު����Ff7y+R{��/*����y�@.e��r������d[,��7�ɺ�^t��˴\���^���F�	��7��LZ�	����~`�ư��(�w�(�)���pN���~)�y�r�B�����h��a�o�ٟ\�ٮZ�yb������	��W�kk��[&X:�o�&�O����G��/H�O�W�i���H�����YBw�RF�^ԫ.�}��i;7�F<�}/�I2��{�j��0ꮭ�Ԑ=���^jE�'�p�WBI�CܗTs�t�d.'r����!;�vꯌ�E���l<�ד�@�V�沪r&
��p\�cL�e�|1�q���|���|�@X�g�!���B�P�u���p�CFT�堢0�V�{��p8X0n? 4�=�02*�~�����ѧ��[��A�D��}�!�5
�h����OT'�����1+ъ��F3?�ֆ~��O������Ǌ�ϡ���%2JOZf�����	7��ש��� ���R�Q��o�����D�"
�g��e���{�����pW��k�w�j�:��(�Sh�qz�|7%�����t�sg�O�uO���x��i�����k��7J�}�ƴ�Kh�M���ia�?+�#g�9~Z1�**rQ2��r|:	{]�����~C��O�}@�s�� %\�yA�3Q��P�:������a&�~B�(���U�L!�� sQ�� �9"s���;�Ґ�'���cŏOn��6�^7�":�������+�[���*�鴈0��w��IM�[FG�3U���P!g�������ť���-�Ae�W�Ｌ��H!q�F
��M:$N	���)U8��P�c�,Jo��z9UQ��aD0��|<�#D�9��&U�|�Qu��$�K��!�|tV�o�G��Co3Ǟ��Hi)���Y��,,�Y�qR߮�ba�7{刢���ak6Z���b�b�B4�`kԿs||7J�&]�p�Fv��KC$6��:f���s���h�FC�<�N���#�
,}ؿ4�%%:�g���^b�蔈~�c����$9�D[MP&�ɛ�&e����R�S�2]9|�c��A*��L���Ѕ����}f��?�vI�є�V�a}��K��'0����]�s�H�����T��
�nӝ4�5�;�Ed��֧�3��2Q���i�uxG�
	+E(���\Y�^×��a��ΪY��Aܤ2�T�Х������Әv)��G��2>���	�>}�[�<:�(I�)H�p��H6���'w�4ڭ%+��r̊�3�� c R�L�l�G��7���ߢ3�o��K3����m�������� ����K��Z����;�K�rd�U�2"ˏǶ^n",�֐�5��I�3���0��Cl�Z��*�to0hךt2F;�'p�;a��T��V���2�j�Xa�YV�����/ ��=�s�Ϝ�^��2�|+��.?N> w��=���q���$�
E�rӴc-�j[*���jl<�8����]6����|���;�{�âx���]Ґ��9�T$��B�&�0L�S����@���=86�'N�n�IX�Z<��/���:F0,��1H���՝NG��؁M\>�\�ۉX.H���,��G�1���]��)����4������U_�$�w
���J�~ъ�Š�r�}=�b�l=9P�㛧��խ�&;�(5hP�S�T��@Tb��-��ڑ�$��q���� �,�R�X���t7��;���r���'�f"1%��&-f��'��[��k������e|�Ϸ��gvB��n�����Y�.V
��Q^͛K�r�\�Q ��YT�X�{�K��+eR�ϰa�߆�������ض��}��3qѭ�����F�f�Dp!M��۝��l��ce��Y<��M(~��m*�eQ�A ��t�z?/���L�<
�^�ͩ������B��\�F�<x�+۹,è��%=�B�frK\مi{��9~`��Z<,)���y��Y����/E�wx �!2�>�)�#���*�{��+T?Ӄ����.��{��-h�X����� ~�ta|�Q����>]�S:�1	��|�!l3@�8(E$�߅&+�<"4����D��(%��:��d��p;YQc;��P�u^�=���kLX�.�P+i���ZQ����bV���׋f�^�Mg����*��cz>d&|�����U�.���I�d��lb��������2N��Vr��:_ּ^���q#�慻** >K�b��{�'��S�t[���>����|��G�M��%�[�
>]�Kt�����<ߌ%Z��Ģ�"�7�a�{�[ ��ss��q������s
-]��7<��p����?̪�|,�<�Y�v�:!����r����,��&�w]��)�ɳL�O1,:m
ͬ��I�_juš*��y��nX\lm�p5�LN=@N_Զ� �y�g$�1��-g�����>�r�R|ߜj�&�KUSghj�#�F&��)�D]S_^9�\@��,�J����bm�r�N��i���S���7�N�9�$÷��9Fa�h�_�,�J��lI���-R��?�S^�E~ʿ��i�{��aq���,��Y.id��U��w��2��¿���u���4�k.��K��S���jp��_Bݱ�<�~�nПȜ2�r��2WC��t:���ɫQ�_E���.��L����=%h|�.�ÁHÊ����jA���;�����:�Ȇ/g��EU�C�6+h���]7b�$j�����=�^W~~���b�z������y�8�z�=��_��B�R�K/%�_�мё�/��"Nrɡy)�PƓ5��D�+��	:��D��8�E	�1�7�`�N�#���O&I�ۨ�\�s��睢db��糁�f�㨿����G+Ya�NU�RP�T�F �/��ْZ|>|T�����1�HH�����h��:��&�3(�3`�~��Q�:.r��*�_>�����|G�2R�9^t��9�Mc��ZS@��k<_�4�8��"���2�q8��td�`=����F��zE�+�X��fs�HqTP)�"Nԁ���݈��y��j������l�OG���t��ܒ�� m �9u�;B��i�I|��=+R�;G<HE�bSh�!"l�v���keR���hJ��b!�iKD�\w7�fXl���sO��ӈcV�&Ύ5 9�j���,:��!���ȓ�����rgѷ��_\ZI#?2H6��R״���O�ps��1P5V
�^�x??$+�|��R'�}&�ߛD~���"֔��h +����~��Ffy�>�#?�ȴ�a�1��X��A�t��4 >�S�˞*�@����·.w�L�r��KX[�dN'(�"lV=1�=�j���l���~UxA�h�8h�FP�Yg���j:�w �vy>�#IVr�M��R��Ӈ�˜o���	#*��aڒN���0c��P7 [R|Wz>��ݭmSt1�����7�:MT�oj�ä�X1�,`y8��8�>J�����렍�r�w|��q 3�y��a�@(�1
�S�#I��[��8��$&���H~U|�?���ÇM)i�д�Ԉ��80MW��@JT��cwlFѯ����Ay(YY#��j_��x��7�p�5Z�G�Zd�:�V����W�B��n�؛�&�cUNhi���ޜ��[0T�[]��O�R]3Ę����G<$���\�h/,���\��� $�j�`�߇"�3�J�	�.���qO8�j�JA �~Ā��z���޸��?���.j&N۝�� J�O�"��R��!��}%<��1=N������5d.�J��iΏU��5շl�������O\���Ae_x��<p.�Yy@=Es�?M����6�l��\��x�E�U�m�����3j� �'�b��̖�ub�Pzݲ�S��� rE� \��P�ܽ�Z����V���hM5�v���?�pп��U�:7M8ۚ`**���x`���id�]�-�����p�%@g6�8���tV�>k�a��O���K{pي"ֈ �� ��dX��a7ޣu�5x��
eZ��:>�@�N���uY�W.F�����CG��(�ێ�-WA*���\]iR��l�R�X9��Y�ܧDsE>�Әy�eKBq�o����.Ԝ{ڛ	$"k��e���3��l�0�n�P��JZ15�-P;�K�뙺O߾��͕�85��=E�5Q@{� �	dܭR�ޅ$��s5�	��͝�?�+Y���A�xa�A�<�R.�D�y{�#+*C<�e�M2����>��M��d}\ks|�U��ߖ<�&���Ե���ا2�����١H��N�Xee��t�w"-ο�J�<Y�v���D�>�M^�N�6�������F{�זf4!�ɣ��(�rq����I����߮�!#��"�����DLe�8s_"l����[O|C/�2AJ�0zF����&E��m�SݔhV�������Z�K��cW�d4R&�n&��⭲��9X�&r
�3X�����SPpF'���Q�C���v��I��TS�e�M�|�q�ɉ�Hp��:h��CM�s]���l̴j��O���q�ִ4  3�^�Z(�@����x��f�q�}�)6��1�T�\��OK�xwL��-��6;8Ň�b�s��WH��8��r�i^��Y��a��%R���ÅB�D��F���d����L�Y�1��B	"���G�#��]��W.p6H8Wp�������_GL]��6�0�ε�|@���v0#y{aڱ?�=�7��������׵�� b7�M�����T�b>��jR��͗��Hm���D���
���Gu��rIp�3�E�)f� �IE�$��h�TΡP����ԟ[+-��,E��x�|hΩ�FR��Ɩѱ�;�[h凫�2�`���#~$�An�՘\���l�_�6;`޷���(O>�x���[-zڋ���*�_�k)0E��Z>�,Ƒ��f���� `2�^�v�j�\R�D{o�v�,.�H�S�x,o?��2����?����E�~�wnJ�v�!fWB�2}�l�����0��O�=٘�a���C�����7o*S����ћ��5���$�~1[���K��Fe
\SMT��S͐l�X�E��e�v�݉X�oI*;�m��IO�D'�H��[��Rh��*C/x>g�T!�~Rd������X�ԧ�-���Q�l�w9i�t��jzx�p+j����E�x�E�U����WY2O�WqD�֤)2���ا5]�Ay�[�&��Ǚ�Վ	[� =�ԇ�.���O��pI�;6M�R�}�U�:����V/ƺ�,�h�C�O���0Ϥ&���Mf�{G*�x�
�&�T{�!	�7i�zL���>p�GP��ǌel15�	T�|�2�`���a�`MK�D��le�&�h��I�FAC;���pu���^�Fwi/Dײ��n'���ֈ�yI8����Y�E9ʸ���T!�oUǳ�u���лj���ٳ�#>�`�ܳ�����^��V=G����W�:x���7STqE�rb*$�#q_�.t�ժ��8hQ1�� ���0��-�%�)�?��B�;N�r�����%������cj+c?���g��*Ȼn�N߰��X���t��%��_[WC�)�~ +�J�Da���r�kG���x�*�~�  �2�K�`^z�Z�]��L���y�m���ݾ��}��gsS���(3����1��j��J5L�,�Zdc�� �0�lvא��EM\��_�;%6O�E�Gm����1t��g9�u��pc���&�1UX("��C�eH+�Ƨ�Cp���-첌y^«�r�r3���������\�$`^	�62�Z	�m�&0�r+%�= l]N` V�6�-�D����A�zf�	���K,X��;���rȑx%BX��6X4��\�u����,��F���®�[�v{[�F���  [D/�23�{���kS�Q����v�됓��4��&�6�G.��(!`�aK�ֲ5��B�L/��Ʒ}��-�����^1���T|K�)�`�nF1������vi:~U�s�	��:v��`3k/D�T����H_ዖ��)o���,������<$:�qgD>�=H���[�z;>
C�@@T�ZG����W�.�M%�p&��cO��sY�h����ޙxh�
l3j�Ď�8Zr�H�N$�r>����mj�]@H�{�,[�3����\ �eB�u2d�ŇȠ�/����xu����O��Y����c|C�q7J=��Uy��\95���g�s���~z0�P��1���zm�Q��,��)OV��>g4� j{��F�W�l��¸�,ʽ{l�{���g0�4�x������;_:8�E�m?��%����{��~�
������[&������ˎ���72�o�ȇ��,aGA��z��c�JȘmҳ!���w�0c�%��6�iXE/5}��̴V/=���̤];`:��&�<	��O�hT�6��5E��Pp�%��������h̖����X!cF�ꍤVy����p�f�������
'!��V��ݬ.�U�zD��Z�:����̖��e�X��d&@59�$ڑ���:�Gk����\�XF��CL���k��WN��q`�[��T0%U�i?�`%�"�;,Ȅ�����O:��D���N��I2W!/����ص2+�����^��ۍ���$�ZL���l�ĝ(��~^��"N��N{��<P�󠾲�W�}K��¨@4�����1�v��rYoYig�N�
8��.a�y$�-�é�ݼ��j��Ҩ2������pb��N�Juwpbc0� �����R�c�@C��RRg�w���m*�s��Oa�]�gXz�3����@��]��G^s+%�-�A�>ez��M-u.��H!�m�皝{�����X��&�@F�xg	q�ֆa�烈O�]�=Gp׼xFV@5v��iuBcrZ����ꝲ9��8�����w�P1�A��t6iXˉD�+�+�"��F
���T��e֭j���~�lB��l�RV
bP��Ց����"y�2E�~��L����?��#k��b4Km$*ThGr��Kq�Xǹ�*�}���ȑ�"X`���i�t�/��}�|{�^�P&���!q���#G���������V�@:���	�4�(����a����>s�#:�l��k}��G/V�qYß���;�����*^,A6)��D�.}OY�ݎ��&:{>�����Q�{�;�B��}���x ���goýA�T�@���PF�$���,��ړ�e=8��ە�7��i�	m�%t�_���!{�3��I2�+j$��w�@֒���\�\��~�F��P�o
ܥ0�_g�P�1i�kͷ��v��(�u0�����G?u])�u�DѪ51��z����df��أ7��0�A��1��O?p
ǔ����^"��]�7}��M��E;(�G�pu�< )O:۟�B�Tf�ai�����1��M��}�Z�D�O��k��P���y�$�����@�����}�H"�/"b!����
�8��S���.��?�m5D����_���n��\��ްD�}�;���#�Y��%;�bC������}���J���ؤS�Wv/ �h��HG�	u{���Md��1�@������$���I\rjq���.M��|�ܛ�w����w�ݢ�� DvY��a���
A���~�M�)H�~ix]y/���5����?:�y��#".�.��_�+�O�!g��o%\5�gV���2n�N����ux� �'��v�� 3�	d��ou;����·�.�C������E摟	�:ήbDt��&�j��#l� $��u1���%�O�o۶oW5����>���#����cF�NW�!��{�u��3 �/��)�'�t����ÓOp�\�ٜ�@�"�5�nA0I���~���0��5�w�R�@��)c"*y�����Ac.�5"�~g���+i���?�u���_8.��8Ҽ��@�&D�c:��2���f�٨�N܂��r��/ ��X��:!7�m�E�N��a�蝣e�[B3�t�`B��Q��Ȇ�<�:5��,�mu�c���x�l�Ɋ����$b%Y^I��'��Tt�9���+np$��^�-&n����3�u�;�;�ⵂ��,�jl�V�<z��265��({�����=i�L]'�/f!e�;E:+������`T<�����Κ�䞼��E���a��g�3�?��(m$c�F$Z��[�q���*��0���q���zI�S3�S�&��B���n �&�]��[�t�NA6�8�QIv	�h�S��͹I�UD�r0�P��^#�NҖG���n?@qͼ�.���~���~�0�վ�y��mv�����ُ��^m�ۂ4�fq!�S�-G5ǲ�&�	���[�V]=y�a�A�᷆�*3��-���(�f)Һ�O�A�ĥ�䪠�iR�$`�i���XTL���ÌB�@�M��LU�M����*$�W"=��<5�H�]S�v�(� )��#�i������M�~,5���D}RFi�kɢ��e=Ov�q`�K����ӜB�mh��`VXA�48�7T��M��F�:;v�qDj�sY^.u%[Ob��x�=8�N/F_���T>� _����qs��gCۍ�%3��K���e��_㽴'�㣱���,��vD�451�-�Tܑ����R��8F�pH�{�iv���a���m��y��c���L`��H�H�?Z=$�:p�S�<U�ue+G�F� զ�� Sz�1�����j�Tz�]J��.�(��m��u��QT�WE
"#*As�ǐ��,B���M(a�c��U����(��Kև�^��l�{��B�8QȠ��B�_����O��ۇ2����=��I�U���v��A�:k��l6�������
���.C�̼>��òfO P9�����]�%�?��8^f�`6pF�T��[���)66<##��yvݕlӘNˎ����C��Syv!�}���X�Ғ�Jvz0"[��i��/�4 ���fɘ)Q��Np,&f���Pڥ����6������3V���1��&F�f�`	��~����;J�3��Zrۣ~Ɠ���Z~��f0�6��>rv����w;^h�)�B0;��~�뉾
�$N�f0h�����I17߻�.� �Ou�I�\3y��!�b�xvW�z�[C��� � �ӯ��o��[��[:�2�TV�����QW�Z�ft�������鲏�o��)&VsjKt��5v�](;�VtU�<t�;�3�'T�p�R-��>$�Ra����ꩽ	Qh#�cR��|C@��q����m�����Y��,Ţ	5'��y���%vǺ� Pq��>V�UW]���I��������-�+�������8L���+2̞4YI������'|5Tmm��N�#`_��5���I|ߪ�eɢ9�I+��I�~�+��N�e��s�mM(����Y6�ɨc=5���|v�ܩ���J��������Z<+{�d��-#��P�R�C:�*$LC��5&D�_W�nX8�@��i�)q�B���߄��x������ސ�i)���v�(�p ��h��T'�p3�,:�kW_6��5!]�oab��s�B$�U��ن1�����$�y�x'^᱊��˶�d}�D3�@�����20v�w��ϵ�k;�@l��O��������W�b�~�co�/v��)v���D��[��|�l�So�qW�yO�m�|��_�I�����/����}���-�[��G�`mCȍ�ۺu+���Cp&�L� �D�s�ѵ�x�7�EEQ������ޛu '�"���{T����0r�j@��
����J�A�Yq�?�����(��
�����k������+��j�	SZ���e�M��4	K��0A��Zjѕ��7Y�c��P,U&��?�9��P
t/�:��=�`K�����R"��4�E:�Z�h�߾_)�>�X6��[[#��>��)v�f�B��P��c���	��G�X���]���>&�JGEl�������k��(I(��_T�rMw�ʍE;(�'�|)�V�o�����Z9�A8����(?#J���%w���!�ח���_;eʘ�C��e�Õ ��"����'��Zْe��]�U�<���sӴY���㭗9l�!5���覬�|��YB�ݗ�y�i�:�b�pE�4ۖS�Y\�(y�L�P�>��F�L�΅�[G��ɇ�s�����;�g���`Rg�uD_����Z�����w^č�3}���:'+���#s9YL�T栭�0黬����s٫���aw�3"F�/��G�\�ZL�����)oi��u>nv[_qf�'o��v��(���Jo���i�.�G�Wx�>�Z2�)EM	��c&�ZhV�6^�ʢ�!��P���nh��rB��
���4?�ڡ��.|�ؓ��6s���d�ܭ^��e�/�s�̥xyH��">9�<P�|\*�����E6X�+����Uk!A���n��g-��ubr�� 7�6���j�o����è� ĕ8�s�bJ`6��xoh٬�dV5!5�}���^Y0������<Xxx;�
�^%F&��t�	���G���h�?mǦ��3x�b�����M�;����d^�}7��ب,ʆi�|�x����'� �wۻ���(�T��Ś��Ы��
���ρ���:��PQ�H|���G'��G�M/�{[A����B���W���s�Y�t�ڝ)6���iV�a�ro2p�]�BW�?�D=* ��J��K�|ȼ�ok�6(��o�������+��pud{2e��X�i��{�QB���P�+C����0��eB�R��Y*�NM~�',	d�?b�)�3�#�k�P.�p��D��g�E���=���w>�ۡ�+i�ю�Tڻ�E!Y�d�vB�c��T�	ٸ�;�Dn���c����t	��84U�N@,G���b ���8��M�S����'ɜ)�#�i��	)�k��5���������x�͢�$`��,�64o?��Hr�Ȧ~��5������l"~�ϷZ@h��x�8~Z�rA�$�>M�p⥴��M7�o��h\���'���N���X���Pc5�����D�_7�uq����sU7Ģ�c�7	���n;H�n�op˰�� ���J������D?���F��^�v$��s��g�Kא򛖺�y�	�$a���7a�RK}+����ΐڀ�"xv��p��W�C������"޻��p׾�
J���.�1I���*J�@L�FT�I���Ce�����o'��|���]�U��_������/��~M�<�i�=~�H�ė��1�i��ȕiV��M��gA�M�|���/l�F^gsu�\����D�'P6x@�����O�}�S%?L��c���c����ˎ����ߴ�	�L����T&%���|�h	nf�I�$����ۣ���_��|7��N1��݃J|4�Jx�����\r��C8��|w����T��누C5�"2�f;ڄ�B�N�s:V��"�r�m�V��s����� d����>�ԣ��e���s (��&P4\��l~׏\<J�t��vFB5e�A�����U�\1J�ϭ*2�To��lx�;�*�g��SV�Mݟ�5��9<_
9(��B����Z��G$���û]�B;2H3A�`�twR�
��ƞt�`���K�,	�&�q/L��(�#��v_og|�!w�_��[�C�)�Q֊��N���o�IE���a���&S�i��6�B���89u�޳���W�ay�)?eN�zKW��7Qz��Iv!����ώ�c�����{<���+QJ�*�dLm �p� V��gNu��[�pt�Y�_�`���}9����֊��J�  (J�HF�!(9���?3� |�7vIǡ�"	��!���AL�6�v�e��=-X�7�L�/��6���3RQR�HWL���X�����ի]n��qT�,�ҔR���ǒ����+\�{b�l�?+E.�2c�.`�
�m'�l����	�ԝ�~�I�[7
�R@M,�/���FR1���4ԧxLCZ�f���E؎���b�ES��Yc?U��Us��h���{��
����P���+z������ESkQ�ՙ-�:��ODT��My�[��*��k��i<G��vF<�)��{@،
+�2�Ki�fm|���(�K�C��n��m��y�/��Jx��NW��-�Br�;��}/�3B=_��u��`��]��qf+�L�G�xv;�@�-�]��zV��)�5A�������B@<��c���zk��ꉙl�N.M�a� �4�h�=�������x�` ���P;�#L�Z��- �"��u��F��mL[��w���>:�52?�TX�n86�1'��缷L������।)0]M/�^�9!�$�iwr�ֹ��g�Y��i��4����
�I��g�],ؠ������`'�_V�^N5�	�>D����֜�gk����9t�3FP� ��)]����S4��`����jMt͈D*�m��{Ք[�Yʭ*�t�K��������Du��Σ�fn�Ƀ��ul�~7_%�S���gN&�p��~����&�u'Y��QCʡ���ת��K7�-�E���E�:�`��lf����nY���k��|�rN���hF���������l��'�%c�=�k2�SS���mdG�h���Y���t�6{x��X�R�
�+��~�gou�6NA���)Ʉ�[������������j�kk7� �}��5��Ӆ2�}�Ŭ�6�����		e:?��D<) �R���%達ʹ�w��X�HpE�i��z��Qt}B(w����w��,��	��U����6NY�K����S�g��7��-�z��?8�Ɣ�q��U0�BK"p��S� �p��>hg:"��Ҧ&�qq&�>��@@ť�M-��4�BB���ef����U�"8��-Uc#�;���MH4�$������?��;���w���Z���'��>@Z+ɾm���ό)18�.��|�m�� �E��2���e��Ig��Y����*�~f�Z"��C* � 8rUPM�P=}��{�_aAW^�'7 n�nr��i>׺��q�G1�qq^��f8]�I�v�C�����a<�႔�岋-[��b�{�D�bd[�=��)�gLT�Xa��ٸ
�I���#�W$��52p��Ku���z�yx���c�־�m�ݲ���0�B0��³U��bL�c0�6/����d����p��'�������cTq����x���h�(�0XV��B<��1�p)`A;J�����A����%˙mB�) 4f"�������)J7N��7�<�5�J�ca_&K����2ǝ ���a���K�-���p�\��,D8h����F�.\ǬO(����[�?����l�s%ͅ�\n��ts�y�r��[�H��K���gh�jlj���a\�L���C4�g�1�����̊Ok�F���= Ƽf*����e�>k_�Q�R���j�ظ��S�%�`ʈ��S����u���F�K���Q@k3�#�Ly�<�����D��Bd��_dlSf4!>�|z
�WI.��I��7�uS�_W��:'��y���˝��_o����0f�:�w��߇�l���DK�k�Y��Pjjw0m�8�Tpa�����#.��J���.b_58)�k��V	�G�	�ȟ�<u��$�Y\�e)��ﲐא����"ef����Ʀ�ݪ�a(�ɿ�ݜ&f��C��Lr�wU�	Y$.W3*��&.�s���m=�}�����D�9&��L��5�e�XR�� |uk��?�Za��F�=cI�RX?�5����!��+vT/{����$>����ˎ!�OI:��p��DwEK�讂�"y�ی�z��{|��(��|f��$w��S'�@�U��/R��o�	 �H���2��������"�����답X��͢�\	u��xx�9	@�5"�� ^��P5�:�=4�Jk}�$:zG�>L�M6�a����ͮ3Ro��|��]�m�es�X�TO�Q�}5���k���{i�����,�e8��lT�U��J�,�r�ڮ�clBK����oh�Mt�H򰟉��0J_��Bq�Di쓞L�(1���8;
`�M�I��v�n��2�v�4�6-�d�����r.}�)���L���{����[�mv����,zv5u�^����8-m����Э=�]F�P�]癣TU]��Q��H��e,��:@��+"xƓ�(��]Ć:��.��q���Up��V�]�'D�}s�<޻ `�7˪(@b��O���nP��vS4z�|޵ve���ޖ�g�`xj�o��0C�^���CuG!��I剶�Pl\a�E�&k�kM�+�������u�~ H`]�%��P��c;ѳ7��0�An���*?���y{�)-�Y�="?���4'��OwL9��h��9rF�J��P|��Y/�t�3�%�lz�cU ��}����1Q����V����T����v�k��|3�)��`';M�Ȕ����n�V��F�B�8�c����F���oR�qv,��݇�L�A�Rug!��J�M�n�#e_��Ϙ��-p�+3���K�f��K��u�8�'Gjk���Q���KK*��&������Q���U?�
�S̑��aJ��q���0�7��.���ڢ�����h�Ֆ@����Mp:�s:����=�]��
a��r�ۻ�$C�l.w�r7�	����8�#q�)��EB��"���Y���s4�"��>� D-ح����#Ff��b�W|�,!����2)�Dpo�E�>}�GV*��n��p���h ��&߶d�Q�dʐ}����,y��2x<Ț�1��B�j�)Ţ��yH��yT�L�.�<W��Ou:x�䓼K9ǉ�C ߴ�a%2Do�C�ٰ�G�.��ʫe���3�Q|E5":[O�B a_�����0��^��θ{�b�3o2�|:��ўd<<�Rs��N��l��������B�r����-i�����mD��G�6'���3b����%��0p��ؘj��M|��\4�G?��g�C�ɵ�>������2|����j�K�5���ӛ�A��Cx�φg]�o���ӭ���*��� P4�LQɫ�	�lV.'yNH���S��Xj����?���a%�\n�Qf8�s��<9�.ܠ.�*bo�mtw��L��{��c���%�v�Z�Z�KT����g[D�"��WN���Q�F���'���=��3�-�`nƉ;�l�n<�5H)�I���:�J��Y��
 �͜L�R��}�9�Nȵ\"k�%�s�
��쑳�����K8D��[�b��,B�voU��o�T��d-m@OPxe��$jѬ��mj��AՀx�1/���s���m���2Xz�Y�i����>�fI����'�S3�I����Ȭ�?a���f+���n�O��*P+Kp�8�[.^�87]��萰�2���f��
��1�'��svP��X�����>����⫊q��?��q%�	<_����ј
�z��:<�G
!	L�>A�mq��� ��ƒ赠(��vjP��$�rf�X^���72�#�Aׅb�C�xQ%{^������V9U��ГT��;)�)�E�á��u�A����խ\[�J�kH�Y	�:�>||
���]6�Ȋ���Ӛ��9�Ҝ���`��:�>��C��,m0��'盡�c����=CC���������25%m'Ub`�� �}�Ņp�ݦ�J Q�L��h��{mo��]?�'I1�s&%����l��U뼶F��.b�a�E��R$�#UQ�:]cs��;�BZ��GKy�����_���Zb ���y6?VP �xN�a����iu"���\��Sv*N��W�^��w���;�u*d�����:�ld�܈��e�����V>`��2���(��c%hP
H ����p���JC�h�S��$��Ao)42��]���0*Z��I�S��$�W���caM�� �d�ܩW��b�������$G��68��l����7Z���[ ��~%�������-S�#l��[@rG�]8�f���� ��9��#����he�#gP;}�� �\#wt�;(���jP�m���}���c�$ְ."����x�{�	��ּ��Ř��
HPr;���dmo>�J�Z�������dD~y�� �T���5�s���Q�Bt�b^FЖ $ќ��o���`
�@-+�)����m6�##B̨�y�T���j`��g��Ǒ���!� ����L�,RaXo���W�7��+L<���E������D���gWa�m���Ls��=0�G�z��(y�oD@w��Q8.�Z����M��V���o��fE��)C�ރg��Ǯ�� ����j�+@���������b�퐜=}/�O+����Ev���
�ב�H��d�����D�V{,mU6-�x�Fj�ȝ�%�N�������+�B�K����Կ� ���w�l��/��	��3�9g��
��
��#���0�]S��D��=L����ke��qyNMԳ�؇��"���)6�l�������\��
$�2q����W�X�-a��t��U]���L�<��jR���QH^]$,;�ᑹFm>6Des1���Lm����]v;G��r�U�������Xj����+��],)mI��'\3����a�Sg�dϢ.5��(���ыvʦH��P�ǒ���#��^���!��+|z��OX�1�|���=��PͯajF�[je���׭�1&�Au���!݅��F��T�3�j6Jf�2���,5��ؚ�g-�@�o�ٽ����P��v��e���SU@�L�<��T�y���`������ɼ3����%ڷ�(+�����|�T��3�g����U��h�P�#ͻc�s��S˱Z����ڷ�>q���}��K�ͪ3u�^�sFtL�Pw�NS�X=����	�����l��REL��#*�PsBDS�tP�������bI{f4��[�>I}�J�䚊�Ut����
��H�9�J�hD8v�`�ut"�!3a ,�zհ���AX���z�V���Ԅ2j��_jqc�f��/5B�V,X�I|��G�ݐW�H���?*��d$��F;�K�݂���ᣘ�k�1�xyo��{��{Q4�R{�rp�f��að���c��w�tk�o J��˝7R��M%aR�߲�-��*s���Ql���ِ�R`�YC�3�������eg����@%�y-"8�2ޞD��M���j)�����Z��F�y`T�n�鳬�
rpi7��(��tʘ���GN�ɡ����&k��D�J��_(q�Ԡ��N-a$�����f���eG��k�I���uӼ$D�����������g��b=]�#rS�̭��&vG�w&(ݡ���wZ�ؖ9���S�\q���Zg7��k��ϱf�YG"�>���Z��Tq#-�bc=n�9�� ���p\�b����g��[���*r�)a#��d��xU�'?�^���e�����m�4��z��|���ˑ���&���'�K��8ϧ3�YN��8��jWf�'+y�a1Q~�W��-W�h1�����/`U�Z��=r�������ba#����od��FB��z�����=��l\/̒��s�9x�,�Q�p2� ?�H��`�cdO%XT�K�cyf7X�*�,�?��^r �&g�X�3�:��45�b��R.{��F�� �:(��l�I��E����E�~�7��\��[Cz�Ft	�kl?J�3��9!I4��B����(ZeC�M4�E�A�٫��j�I$�����Rp�s;T������m��v�A��C�-�	�CY����h�LK�5~��gU�_,i�v_uă\�&l���e��h~��6����^ځ�%�"��Y����,��<���]�n$��'O
�x�Y
�l�y9��v�}.���������$��,��.�9uĮ���Aml�\��ɉ�9:���!{EGM_+�I���?��{:�\f��\�;���Q�e]J?U�&i.��5��[0ޝ�� Y��u�!e������4���x�t&���	�fy,���Mn��/o����Z����ox������Nw�0������Ss�9�Ζ+Y*}���6ҋR�2k�^�z��ڗ�![R��9���2zF�t�43��
�y���đ��B]�ɢ���X��U�=��z�;S&� �~$�uݖ���r0q��Md�!�:h�5Xk�|�Ⱥ&��*vy�I��[���`c��gZ�� �J����9�~b��#-A��_���H>�A`�-kfȆ]3���2�S�T�=����H9��|��(�'�Q����<����LW�џ=H����}~���Q s���U��YCކ����(���a
0���6H�5����P�ĥ��!9����+Ԃ?ޕ,5�-�,�OQBYRϘ��F[�l�u<>�VKx䣱��x��v�������8�n�6D�7@�C%��;��}@�,��k�_[�7���z�1�.���/.#"����4 :���2�O!5�����J�D]3���z|���}%�'����.3�l���+�Z�X��D�_PG���IN���N�qNHr��H�+��.�c| Agߦ�%���wmڸ�um��\0��9� ?�C�gG�\��� 2��x#�#��C@���<��f�\Ϲe�ae�z�#��r�����|�9�0C��c[�&5�>G!�p)���;��Z���� ��������-��&ԧ4��t����Ag������$5,���BEi8�A�$��"t���Z+JL��Vٻ=kVk*���b�Q�]mft����x����C
+�����>���(Ki�O�ƨL�����q֨��9�"���3}���#VK�{H��G@z-�)�:)1g
�y$�|���h��+n�U��E�������x���r����>�k:MW{�T+��F�>��IP�����խg�`�����zb�'n"U���%��4�}�#�f�	]�
Ԑ��M���)4�Ǌ��J6 �N'�م����I���.�p�S0\��w�Z�=|����y�ڠ6��T�D��"4��l &tMFqX���v����نiM��R�j<��(/*+ �N����:����5�p��s�!-�1Jj��9M����_v��{��U���S�k7�r���ّ���s�m-��I-�l�q�`�����|NU�Y%**��aYK�z�D!�X�����`�+]����莳��7]���]*�с�@E)�ʛ0
�»�_SS�@�Uw�7X��`��wN6�0���rM�OS�*ӳO�G��ط��3��;q���19o ɢ9I�Jc$�A�{���+<u�Ͽ;J��������|qT2;�{�q��0ea6XJ)wSSX=	��]+��DS��j�U{��勍%�����.4J.�߀`:��p�a�X7��Nnt�����,��@.L_��hl.b�P�ߛx�b:�	OmdX��>3��  �2��Ve[����q�~+7�􍽋N�G��?$v�c�Z�g$�o������9\&&Q�F=$ax��A�6�5��"4�"�N�XF{hw+�:��ǔ|����ʏ�p�O`�J�4,q��Hi�O����7�%�Pb��M��Tӌ�=JU_������F3��f4����C�$9r�!��bu�l�~v��e��3-�nԍ�wf�<*50�����`�0�ChrVɟ��,<a���KYC�y}[����q6����^3�ǵ�ha�&��:�7�JO�t3r���mR��ŧ��ke]B*�i����XYy�M���(�C/���D��)�����#<s���a�a��3~$�M��ٻ�������}�!�c5��;���<������#|���7?�~��&�a�T�e}*�J���̙�������|�9�z�$_���N�z;+��P�E�<�G���#S�[#����C�`��
�
;Z0��	���Ls�L����.����97�\);V�uZ�����d_Hh��(>�_�����7�ø	�;�]�z��|Ӏ�z����xWUM�G��������@�Ԃ3����O�ퟪl..9S�q��~�����)��j�$Ϟ�A����ג��Å�z,�C�#��)�e���n����#rD
�p_綎
��
���3�3)`bN����?��Qb?�Ҭ�g�މ�&L�����+�pN���?J�����+����^M'J��	�޸ХN�g�&TQ�"���2g��YT�R��8��m�s��! ��(��(�>�6��T�k~���Kckp�zyH|�CU��3_�f$l̎N̒q�����/�Z��'�.�t��(�xҸ9ɾ=�}F�� GK��s�`�gSY/�*h܋��~��с�wρ�RSάF���bίo2:m�c#���`����#h���D ^@7[|ا�J^�(q��px��1e�)���T�d|� w$�pgc�1�MqGivd�u�׆�Ĺ��Hha)|&�c�iMҐ~d��UG<MR_����'�qꩽ2ē�({���-<A�a^�U�n��3jW0��T��)��Vt Cd�����'lt������o#�>u?4����$�i���ʵ�^���(�(E$F3a�*���G���$5��m��<�ҟ_��7��i�L�a�=��+�B/��y�p���A�z-�)���+Z�wU��g��E�zb�8{��A�F?Fkԅ��F�jv5�_����S�Ԇ�@�<�Q�$�{�r��t+v+4:�_�6T�	�.9��]����Rneaf������;^���Ga���\�Bة������ �a~,Ι�3A�`2���7�S���J�^��#5&:��؜.�jS�d"t7���a�@9d�G5@���K��^�a,���]9Ɩm4"������A��Z��	��e{����r�������z)7B�q{�=ZrR�4���������$�Jzﺾ�x�P�%Oi�_���]��&��K8�a�?�g
��Bi��(ќŢԓ���ǅkr��`{ ��M�y����j��3Y�r�`�p���}H<�kg�5�Z��(i��)6H��P�����&��u�{��>�M��w����6�Sz\�]�#������Wܐ�U~�k䅮����$�F�Ҙ;�i��ҭ%��9��E�s�F�b��I)�(�Ƣx�ׯ��ԦsIcg��ww����B��s�ަ��T]��%�o�+�*T�����2��_f��s�̟�{�t�șM�������l�dȭ�J`��)8;�(��UK���a{#�\&t|kퟨ�P�~�W��C�	�����k�>�H����--�!Gsq�d}���7�G��"sUь<�/Z�.�Wh��һ}*À�]s��( �f(%6|m���]��V�(�6��f!%uU}��\1G���/�iU�1��0w��L�m4�F{���F��3D��C�8;�K�W�w�X��h!8�*����DN_�}t��=��@p|��+h7�#?�q[�%"sU�[�58Dir��Hp�b���t����d_�5�^��@l��&H�.Gu*K�k����P69����56:�K��D�.�~
��Te�b��(�]��櫾�&B�ӹ`ᐴVr��]�T$��u���[��w�=Xh5#�Kb��<y=+vG.>���!\姇0N!Pqh��P��t�w�V���z&��^�j�Ş,
c��j�X����;�A�� g�LB'�uonX^.-{eW�;�Lk�����@g`�J-�\��9"}�1n����T\F��F����)v��m�8G���=��h�t+f#� p���P�_��vWGn&�8�D�<��Dc�&�_'��D-������O�ٷI�������ʉ��^�;m6R���~�2��qyWގ��w}ݰq:�.}g#h��{��L��]�C�����5w�+
�?υv�Τ��	�V[�/��>5�1���%펾O�̇bHon�5��z*���v�zm���a\��r�2�-�3��W��1���S*��7�
�B�Z^>T�E�3Q�l.f{��n�����LU�l��������ͼb,�LMT[�'6;&[����k��0�ƒ�1�1h��P���]#z/�5�E� �`��|޴~dN>A���J�iݻ�̧���=��'~�%�=����M��0?������?�* O��8zK�"�dul-c�������-��88 <g���3Tͽ��v2|xߴ�J�X�&�
�8I�UL�5�J����n�����fYr���(����	a�8��}��U��s��˥������H���݆�y�٥�ߐ$)��x0�bP����)-���+A�R[� �p 2{�>�Rp�~fi��Yȯ�-��x��\���Ek>bH����n��������P-����c "�35Gj��R� ��(�/m<����|��6z�)�欖�����L=��J��֍h;�4���90BJ~ea�ߝ�u7��G	Lews��.���:j�'1�Rׁ�֗~o�=XMw�� ������z�z;ƯK�G*@�'�^�1����Iǔ ���d2A`����S)��F�]\�:�.���9������DČ��<*=��Y����E^{e�<���L�G*~��ȅ[*0f�����V�tUF�(�ܲ~JX�t�lѴ��K�m6���W�)}�*����B&��
㽘� Uࣔ�tѲ���������8О�0_	�4Ɂ��v��o�̜�(_ h���4gꀟ�Q�C&S�⍇�ܪ)a\L�2��x�����j���>h\�j���<�+�������dM� Na�f~��1h�}�.>e�_,|I.��j�V��AJ~�10�}i�+b���������,�n�@e�r�ۄ�����L{�w���a;	���<=[�d"�.䆖2�Ñ���@iɷ����O�Z���Lj#i��-č��盌f�eq[M:}���W����F���^0�����^�-����@w�b��w�eo������]�� ��&�CwZ��L'�@r
k�)s��C��^��=�n���ה]��)1�!*����D��) 
�v�B�#�-ӜDa'��n�g����X>5���o �6�x���=qbU���&GGgl��!1�����C�h��gPq���������'��-"�M���:=���/j��(QvT}e=|����Y����A[F�4��{��
��� �S�ƽF5�*I���EC��.��TW%�A� b���E�}l�9���	W���OH/#� �x��@��ٽ�k��H� ��9�6>��i����i�e�⹧G��+���,\t�z�|\o��J��@[]�*~6�����8���}��\��W~��{b�1MR��<Mx"uF��٩��*�3��cO��S�]�iN����XYwv��J��F��2۾Kf8������o��p�M�w
�����A�U���A�2�Gn��8�|�$:���h��V��0]�\������}������Qm�e��չ���N~�?��D@s��Z�Ma�#�_��Փ(�?��Pq�K���%�C�þ("Qu���q�����:{���Cj��3���#?W���e�U�Ϲ=���JN�>lɅb��2��Q5��� @�lU|�|���-�daL�R�>�	JD��R[��W�h��41����ʞ@�'���WB£���D���m���q��;�Y����uwB$�������\�9�/?~�&�ǜ<R�q5J��{5B���ʘ����5]��֙eIs���v�uk$�b�G-T.C��$��p+��/d�
��2]b��s�9_���Y���D�܆/l2J:�{e�u��.�8]1ã(�[v�ڐ�c���:�>��S�`��~��uL���FL�S�kRM5�m;�_«<����`ˁ@~"�T9˱��-�h z�8���v*�xa�����yP�^��	�ֿfZ��\�w4neXN��(�R+{f!��Yѯ�� SR��6W��t*�O|"ҴO�L.�H�j�"�D�ۮ���LV��Rv��9c��eٜ-�����r��iR4�|�Z9�6��%��$믮	D
h9�oIDM��$�� �|����$�_W-�E�o�z��eM�gz��O�,I��i��x��v�p�'m&�	S��ܽ�\jȄ�%4�S���-�U�����2�C��|��u��W`mk�z��M��Ü��ƟcX�����­F��/�ߠ�?���j63�Q�g ���X�m0�=���A�p�mMG�Pa��?9���۳nU�'YDa0+2�DK}�H�r���n�T7ѩ_���ۮE9���򷽍�$]g��?$Y��opM�6ъ���8d��!��o��TZ�S��,��\��3ҿ` �(L�A��S�� �X^{��S�O���߻�1BQˎ��H
QvSm�����!��K��|���;N���_�|�ʟ����⺉��陪�@)�~�(T w"�KQ���i5��1E��Y�,����I���,n(����5���m`�2����f�y�[A\wOs��`=qX��LX"�����̢���}�˳pPhC����i�lW��$|����j���^�g�5m+Y��i��5<1�������7*�e�bh9�^���KZI�/t�2\���^D~%���F�#�EE�{H��ʔ�6�Ą?k0�;-/U�v��ef�D�H�R=�|�c6.���1��	0�!�� ū������N�O��7�z4�U�q�d�ITcW)l�Z4����@=bU���J8S�¹:5M�z���!�XW�p6z��/�K��;l��%pR�� [�xҡev0�[NX^���
h>�!=�<����kl �j=jN�nC�q�̋cm�g�98=�c6����7Ro�d����i���w�Zs"�Ƚ\���뗻�$I�XV�X��~@\J�en��3%�U@<ԡv��I#j�*�����u��0����pPg3�:;�D����C��[]r��-��W�#�a����,�~��HXU�	�u^��!�S�:��4��}O��D�Z����8ǩ)6>D���{)֫0��$]>�^�r��\G����TSB�|�yWds�A(p!�����`ڳ��?���gg=�7u~�Z�y�gf����D�pK��F���_��45̙��G���8�'��(bI��9�ES��NX�=l��) ��3C��٫�3��u�jS<Pw���(�]cr����	Q����qdN���vr��IH�z��ާ�xc��Q��8��unA'z�f	3p�D^L�RS��_2~�x�D@����$��XL��i��+3�],�:X�m����) �p�yx�Ή�i��krc2p�-F�۰{�$d[���J��}�jcJu-�2K�΋����II��s5�dI7'�~�|
��ԟݯ���LX�E�r�,7Y�nf�ݽQj�V[�}��L4W����v�q�5!�I6g�٧PO��6N֣��̹Xi�?WW�c�������2>pP� �7�e�G&_�3���8D�@s�����\+7(���IQ�f���gW��%c�#��z�?<�鏭�����ה���{�1H뙀������ElO/$&������.��@0���*�i�J�aI������懎5'Ξ��8r�Z=ɨ����/洸d��1'kk"d!��t�r<<J)��kҎ�R��:e��r�����J҂�N���-n�����<F5���k//�*�ѐ&P�L*@`�j��V���],|)��ÏR,Ux�[>��TI��KA��-��m���@��#���9L1�����u}𛸇�w[T�,��p��BL�[�d#K#��"+(�O#iD�����|�Y�b�R
ca��;v����U@0f�8�����Ε�ZP�5۲HL�:�{�tpoB� �{�gｱl�`������`oE��e�#��V��ǩ�BC�| ���)�q��=��R'�b�Q�1��9vj�Dz��kɃ�S��*K�cϽ(uE�_j�b%Ëıl�TB>���B��퐄�s��J��vu��	��'q���2�:{�!W-�d�ľsY)Fˏ�p�i�%�o�N9��2�!�?��=z�£�|�#��"�����(�=��}�u��J6��#ϣ=FnS9s�L@��%�o=����%��ńT�)�a�L�V�vkK�z�����/�RI��"�
n����P��dU4��6�1 LCu�I$��dJ?>� �~��[`�v�L7w���d8�$Ì� -�Ǔ�#$;{נ �Z�$�����Ia ��o|}��3u#�ykW�E�67cᤉp��`��z���{VT�NP3��^�pvY��i��vR�yJ��!�.��:���W~��~��s��B��mʌ�W���v�&v�3D�ߝ����ͨD�$�V}�<��Ŝ*I��MvM�)��E$ί��{�z�but-�<
4�܎H���؍O�.ZG�.�w4�P������؝7^�|�S�بR��&�����/-���ΦΥj��K>�uH�����PKo����=���ĶM�-��YAu��T�v�������I�zA�z���1�J��]���R�p��R�@4�u�J��J{��A��$�- 9�U�1Ơ3�@��ؿ�����B�2@�0���!��5ݤ��3j��=��&��A�@C{ሾD���?�MG�{�dē�"�r���6�b��֛��^Pb���!�N�nlc�?���']��˩(]ES�fÎ4����MQF���B�
���.�i=y#�ۗJf2띗1a�)՚�D[���a�73Q��حL�|�e���s��.�0�E�2�"7�Y�"��Z�
��{'Z⼩�`� ���|���H6@p��
>N�N�S����l��j.�$���J|D�Uk]n\e1&�s��ң��|��'�'|VQ�I����χ�ھ��ʌn���_|�E3� �S�e�u��-�'��[�G HDu�K�����a�W{@�3M����j�b@[4?�̖��A���h���sK�E頳�n"�kph@x���'eY���ϔ�D�*7:���H�=R��ğ$����ܼ�S���vY��=4A�@�5��)�c��J��3�\��t�4X���DJX��kꀨ���Z��	�����'z�ro�t���h5T�C��2�p���T@�>�Z�b7o��_
�m�)��f
}=K��e-��Ў�����e���^�V���8B�k`>u�xV!8<�7Z�:�"�2�����yE�L�&�cgh��O�p�T0Wy=����S��]z�L��JL���ĥ�����K� �����B��B������=���#%X#c�lq�4YS��v���fͼ���`�/�/��&����\r��[�D �l�Z#	�����:i�½vm�S�� a5<�$�b�R�+��K�1��tX�,�Bs<����f]�q�ʳJ8?_\�� ��(�ڶ?q��G����D���"��уVB�+_k��c�H������^��Im��\���Ǵ�VG~8qѺ�=�Bg����=�=P��i�HdF��]J~��E�AK�.A$AX^C��ҝ<Ҝ�Z♊��0W�[1;��?KQ�c��]��L#��D�>X֨�Yg����c�űuI����>U����c��bQUѼ	yŖ�?�<��^��*U�~��Wt���쟙RGO�csT���@H�����fh�L'�@ o���:��1�-bP�Q�Ji
�)�DR�uO$�A��/�|q���;�?I��I���'���4y-���2���A
��������َ;����;x��9�^mq\��| ����$h R�h:�X�8��^�xP�`e��Z	����Mzt��l�]{-C��K�L��N�Mp��.
_�s������}�H�.�q��J;���@(A`2������M���}%�g�$+K���ڮ j���|Y���V����m�F��Aߜ��(_n��;�wy��u��n9"�0޴���@��H_J�a��99��A[]���
�8�$��6wE�2�ݵ�1>14o�ƹ��%`���_�����e��d�R:n��p2�8�_��ޏ(`4�Y�jh�OI��>3�{���lB���2��q���>��w�fX7%w�ȶտ�?�Q䭙uS��2�-�9��?k���e6
4�R\ā��I��C�����͇���hsZ����f[�	h�x6&�pG�7D�f�����<ywH���!�����G�����=�ٷH�u�#�	v���ɞM�w�2"+�5�+HP�B��+i�)�Y�����.]L�u6��6s���(o��(W����&p>����E,��$��,;�����ۘ�,G��nE�>պ���L�7f7���*4"� ���0��x7!�`�cyS8<�g��d�b��9�ӥx�Wl#�л0l$���T�d��6*�(	{`�Y�l�75(ig�dml�cK�X*��b�hL(ۆ��>RZx&��իX���Ɖf�R��	`M��If��T~6������M�b�9���٣��ݿv:xa�Վ)�|���Dk@ȑ���`�[��4��V�b�PߎxA�-)_�/��&�zH�����@�8`{v(e�l7x,gh���g��u�׾k0���U���E�������:��NF�&�e���5�t(�i:c��I2�0�X��Rʀ�R�;�C���Z�b��J���9��jo�Ae�&Ŏ��i&)�_q@I�S����rJo��A������������4�*�ӊ��x��eŋkm{��7���3���zq����fƾO�{���_7�����y ��Q߈r83��n:e�f�;�9��/Ұm(qP�-���'�KV!S͎`xY�(#�%��yl��CmK��Qڣ&%����@�������Z��{��xGJ{����4f��Ռ��نH(X>�(�yTJ*Ut`�M�]C�)I�<ȇ�^�ǃ}uS�W�y�,���������]�I��"#�CU�x��"�o$����ܪ��`|V2�a9ڽ�ԯވ�O��c����W�U�-@�Y�s�q�[,6�WR���&�;�k.ڥ%�a4.�R�O�o93N�=~f�t����4�Ap�.���8vUȎ0 �����E�B������?���n�%x'\K��Iõ�g���G��J����Ƌ2v]WK
]�)�ங����l�DJ�n}��65ZaW�m�.D�U�� ��M����m��:I��Fj ?�#��[@��rH'6�|8�P��#Z7|0��d�[*4$@��Ba�@yڎ��W�d�r˥��I�'X2֪yD���3ɺ��~�/or��ü�� ������>�d>���E�)��G%g�:��,��R�v�qFں
+P�B�N�K!������{���y����BTF�_��a�l�<w��޸\:�~<m�V�BHަ�(*��4�h]�5@�Tm����\�*'~JOx3�+,�	({ZI�Pc�'�%�|b�䷼�-�WQ��hT�1P4�`}6\N�Cp���A�,�����S&��(W��{����U D����L!߸�����aI�	���|�%�}E��-�3'wo����P^H�>�{�$`��@�Mq:z�|3Z�`#�7��bJ&���E�'�_bP�2O%���
�����nJ4&j���a��S���*�m������b?*�q���ݰ���Mh��E������!=J����3j����.�I��A���D�jY힘���{1`xb2<�p;�^.�T���^��+�kW�\U�>�[r���X��ֲ/�%�mo��݉�0�]��P���^��ѽ�B�
_��?k�t��`Y�����nUD�ɸ�|-d��Õ�����Dm����-����Z�de|G�t_h��y�.�Yc�l ��?	���Ŵ�y	b��/�CѢd2z������я�5e#8�H��F�f�zzq�9�D�T2�Ϗ��J���'�v���+USp�XV�6ꀔ�L[Q� �qa��He
�=W]�r�L=v�)��ʕnn�Gfv��)d��E�8�1X��	
)�~N\�^�?.�C�A������ʞR�*.90�$���RC'�u���~g8D���9h��G[&�:��'3
�\����8Ͱ��c�̒9p,F��4oo�gk�j%?<>@mx��%նm�YX��1F��[�MEFB���Ϛ�^=:�S~��u�g*$U�%��ߟ���\)Ϧ/8(�+�{s%_�7�Jg�^&���f�.W�&���(���9�r��}�q�*{���Qj���"�2ı{,QU� �z�?R�u�$B���x+��H����
�݇M��`�m������ �Q@��?^!�ʅ���[�c��[Ē](��z�*��GX�-��~gy�b4��7��B���j�r�:Ux�2-�TQ��`��L�a$}r�H��#�俔͸�G���<�W�Z���ޡ���C*6����A���Q�wX�l�����x{Q O2��H�WVi������R�tJ����^B�ߙa�hc�wR��(|���0�����d�*��o<�=N��;@���0!A~j,=��,S�r������C7�JL����%���Z&�D����{ ���䡢����ك�����"���vB~���z��YN	���\Y{����u��qc�;G�2a�X\��k	�ۓ�M����?U�xj^q�?��
q��-��tt��ޡp���B�e\v	L�@V�{�Z�ܰ�W �K��{7��iy�e�.�6L]�y��]PC��Hzd^��%�^d}/���+�%���rЏݴ�OWC���{� |{p��������f�z�U�$�����f>�8�gIU�ob�)��h֠���nao��I[�0�j���>�h��j`���u4Y�^A-^Y��JI���]+��!��m�+�h�~S���1A��W�+ �G��#���e�lL���Z&�k���WFL�Cֽ[�J?�����i�t�@��#����O1�K���z�BQ������� G7�6 �T)=A�*́� �m��9�S�H�����x��4��}@�k�!�J���Iì:!9r����5����Xw�^B�M�"_뉓;�/���͂�5��)S���%S���&��j8I���:�u����J�QFɈ
��ߏ((-��a8߇�#A����M�8 ����T ���z�C7����4�W��e(�*�v1�k/6Pݍ?Q�1|Qf�=�����%�3�$�Vu���E��\��t���Y��>⿍=��V����O����:}�n~9,[�q.�<�2�<�뢅���7�Xɐ�`� @��n������ �s���Џ�z��]yi{Q'���_����3_��#��qs?�q����'�kF�Hu��h�E,� �.�˧a�{�L�l�*�\�q}|��e�+&pΦۓ+zO��AMF�A�3V2����t�UP�E��Q�C[֮���K¡ �$�8k��bz����U�i �I����\�P ɚ3=��*쪐o��r�j����u?�ĉ��^���u�;?ܻ(iR�U����H�L�1)�$���C�E��c����Ƣ��2]->�.Y��ٔv��^/�s$Qp�61C�E[�(>5��@��K�*ۮ�}h!�m������T�)-�s��Q�}ˤ�E�[�0	(G���Q\U���0����(#�j�� ��0�
��&e�r��}P��nS�Qh���W���;s-X�i�ɋ �� �D��>)v? ��A.6��	:�o�Eۊ�<��,"�κ�5D�
�=4#��&�U�*��Xfu�;.���F�<���0�^b��ٙ����Ay�NVi|�|A��k�j �����8:DfD����7*{s�:���3@T,G���$R��������$�Zc�)��E��Miv���b�I�!3�ZH��5ڪ�d4��6~�t]���ڜ^E�V��*7�(�� �G�[� d���2ĕ[�U���'���@�	@?lB�ka��^��r����i~Q��B}^���Q���Щ9#ۤ�<�j㚝�֫Y�3�� �Fl���>M���#��/�蠩�0�d(��|���*D�$E�Լpr����I�1)��U!���@��8^�kq�گ�sj��I��V'5�9��m�M����r�&�i�\��(7�4��a��隄�fjMӿ�2L_����-g��������|�d{U��xg0����H!�@4��y&W&Z2����8.�g������B���&�J�`xy�=�3���
FC��ʎ�wG�t79r���T�1��GJ��dk9t7r-i$�Lu�ǫ/<�s7�z̸!��,\`@���7_���5�V#q��m�N/�~��T֜�D,�fe����%v)�7Հ�;�H*⪰��<$B�`,%^)O;$�Z�Ï�q�g7ς��!ᠻ�ذ��3Y�$���<>q��K����$��k(F�*�����<��ghz���W�o�X՝\���Ѹ�bb��8���N�0��f��*8iN��G�}�_Z�zT�|]I��j�@e@�Yޕ��F1X�_�Ra�#�����l��WL!�Ţo�k�q��cAt���k�2ɱ��u��{�o�9�	���0�T��m��I���pr��*���|d��2�RX��ȬT]8T�ͨ�L E:$H]+�MF��"���`�r($�"�q`���[Y��3#g]��	�8[^{v������l��f/��I����$��h#7�@}����7Ƙ\��ј�7�j���<$���#O��`��������,��~�2(��+��7��:��4�5�_��� ��͓+�w�}͸�p=,���9��_�x�����C<��ktN�Wf���P�83�D5���ҡ���U����.5�
�	��:�h�!=<>��2^�q�Pr� �P'��@o���>���7_r�o��(�p��i�M���,��#�ݸ~D+�ղ��s�̆��'���A������?���z��t���bs�����l,]9b)���۶��$�:�@	Ɉv	���=��N��O�����Ҝ�e��߲O���%e��Y�mup�e�����y��ۃ�w�<8ݜ�ۄ�#C�ɱ"�W����yG�`�_?.XġG�gWD;�|�E��BP_%˗�
��7'�I��M�J�93�a+C0o�Z��[	��B*ea�Z��)���о��f�_Cw��~��^-�,�F���y?����7PbV� �D�OmB#�`V��O�@�h���#@�XN��^]��_��F7OW�wW� ��<���;�on�Mw..}����S���"W=��l8�@_y,-�G��Z�W�I�gj��3�B���؀��d��9�-$ɲ���Wjі�P������{�}�?P���%5M+f�N(�K�8ұ���������X{kz���Z��T����#Z$?�sy\M�sc���R@�Ǎ<��2��� G�b�� g,�"DX�a�8Q�Y���DS�L�0���L�Ō-_�NH�'[ğX��#�C���ź��N��ʏl���H~ m^O����eˈW��ɼ��n�;������wC�nn���C��14��Xv&.	O-��M�^A�D4/#�=��F������T6ح�Y;|+�g簀�5
�m�<]��	���0�G���	�k)���]+ba�{�)S�$J�8��Q{�ܰ�\l7E��?��dJ�S�p��\AU�}�9��ޣjg��z��m��v���S�f-�;��|�Vw�·�˵[�3Q.�B�~_W�!ۚ%�D�3�l|C�+|O5Yڌ�vC�+ЌU+������X�(�� ��a��Nx�K��fZ��aL�k��˜��ؕ�P�e5�[*h�C;�7������g���Ki�E`㝎��694E�����Ɛ����:���uKY8�2*Rώe8����j�$7I�3����y�����C�u�te�O'q��
�ëUˋY%��E.�R+w/�g-P=P��t�Xߺ_@*髫����"�|�N����Rm�l�B��_��J5�O7k^��Z;���C\�S��q���+���Ɇ��	!n����h��:b����uz���3���O�K�v�_��.L$��he'u���@����[_���[Dl�헖�Զ���ҨQ�>Է=��t�=���a_�{�IonՀ��K��(�%-r����r���&�dOp�sA�������u>D49�h����'Xu�Et��@R����V��٫u1[��C�jA[��)K;eM�'�b�5	Vd��=��c僈e����q����#��e�����[�B܎�A�=�J����{�����)f�26�p����?�b��L0d[�|��'�M�i�M��q�V�Z[�g��ڲ!H�_������X�q�8�����%����z�H�����yKF�X:�:aw�D��5gv�5)�l<y�)�Z}Z|s���,�ّ��Ӿ�!�=���v`�ۈ:���_�;�A��k��M��ү}���b����j�ݻ�3Q����V��R�*݋�5�I����'�`�13�0`t���<W����H#� Vj.@&	{���+Bb�6E>7|���K���:w��ƮSn�L�����ă��XȈ��s���b��4<�b t�\X��YS�����?eMn8~�w�D:G2˫H10�&8I0,H�E�?Ί�(iT�}hA����F/ضe��_���Ș���Ψc
1�qǇ�c
���)���&Uݲ0T�\		3���m	jjLE\��n5����o�n�m7��`��8bNm�xM��������/����gH�p��vF�'�Jk0�wVlέz���:�O��	�x��@g��zs��]����n;	�/�Y�ǣ�/��?=v�G� !�7�g!Q�L�����d�����/>�>)��K��sAgޢ�<�j2\�[z6�N��1����!TLq@�u��a'������f��z�h��C�q4��PG��|Kr$�wO�A�\><��!8q����[� D+H�����b���Q_�������%���}n�����a���e��V��ٙs*��˟p�����e>�r�{��o�.+B��A�|a�6�ze���z!��
$�ӕ�Cղ��|��ޢ#�3g2�\7��&B2�����=�����Z�oʡGvS��u��|����Gg�*��]�!+B<���������R�ƃ���X�>��Y�D-hM>� i�S��y]�����&�����3��]RBzQ����+��#2����J}��=��!�3x�����@�GI�b ��8X�?5-�h=��2H!4w��f��<8�}��*л�3�ǃf�O�+��eHq��-I�/����TJ�_a�k��e��5�0�n��%<m��0���U���Ex���4{k�[��&�__Ia߿�w\�`�f�*�Λr��Q�>�;`e4�t��2��̡�j�`������=H+xS]̉��vX5p㘲��!�x��<SEz� ]S:x��=sH�"��\t�"��w tёXGFl��ZdA�x��[1Rb����h�bϣ[��on��{A��*GH��i�]OK��r-�K:��NA��]Ñ� ����}ߏ��m:�������R4}��S��F�/Y�z���.*�	�B=�?C��JQNs�x���`xyG }�=س�\���ej��y��ߌ����@�mɗ�6�f$�?��8��-�q2%I�;���G.fP�w���sC{�Ek�l��εg�%4��-�c-]p����������;�Sd���6h��������|�m�(���F��2���1�/�1�u�Ҹ���(o���3�p��p<G+xen47�t����/�����sH��Cc���z��#\�_��	�k�Mc芧�8�n�f���Bo�B`�,/d���n����q�@Z�����r�s�Qw�r�5�8Y*b�ؙ���6�vU�?|y����	���f�A��vܕm��;-���{��B��KN�>�E����� �xeq�x��.���C�s�z�wi��Q��Y����f�X��}Q����;'���yXS�)�dW}�OD��Dgu[!�v����g�Z��>��M,t�c��{������A�M]֧�F�#q3+yh�r��(�?6�=�3hO�@��1��,y�ȯE�5����Q�Z>P]����iذ�'�Yɨ�uR�	��� ��g��f'sͷ���
�<��cR�q��2��b�pͅ����qz=���ݹ��K�������QGUR�v� ���`��;Ee���yu�F>�*ϑ#�&Yr�9HY��T�ߜ�g�l�N	a�.�I�F��y&]	�*W��)ϯs��4��e84i�x(�-9��Zf��p�?�<txP�Η��*����!�/6�׋�>M��+K���b��dh �vOv�fa��M�C��@6PWv1_�o�aV��C�;X�I�U��3�	n���i��Is5����s�(]�w�f�G�@NF�l9�e��am��++F���Ȧ?�e�0�=U�WLO��߁|���C_5�6H��@xQ�ɂ�inUPU|W���Gle[I�(��x�c1⽜sR�f�n���������^���F+i7���r�JPl�bʽb��|d���%��)z�e���#�_��ry@�.~���li`ŵYk]�������8s/�(�S�ښ��y�v�j����o��UV�C��1��\����r���Rj��=}cʕ��$w ����0���� o�,Kj��$��@��=�.��0?U)��Ӌ�d��<d��*�aj�� ��}�-w,����M15�)��ϭ�o}��$w��,@�'����/IZ���탪�Ί�8�UhU�}D���55�F����2�x:��p�ݑUP[������&�RJL���i"��sUz,���n��s�R�}i5׵:(�P>���8����^{�������}{����T����U%O������ёg��	Vr��he_��?01>>�;���\��Nm�&��?�pqP�����ͫh:3�S>e��|�D<�1Qro!�`�EpF�}\%f��kPduG����o���iV�t�-Q�k1����=��9�3�Nk�b��_�!�V�"3rQZ��yY� ���4��Y ��J@��u5�N�"�!a�P�5�H�+&��xK��g8�ǉ��b���Ϊ��GhJi��:/�72��V���D�~�f�q�i���1�{Ʋ�m51�	�����c,$��
�����F.K�����I1�.�U�ɒP9ky���vL�F��##�'�o�c2�R`���?{�j �
�Bt�1�4�� �R}]���eݛ�<vP����.;��c|�F��4�*���y6/1���N� |_��-��b�d�n����;�-��.��$�٭p�O��윙4�)��Ma���>/��T0Ɂ��BI� 5�/\�����S�le��{��-�]��,s�����ƛ��y22�@Z�fi�����~�������?���=���ى�(��Lu�y�H�iqݞ��!`�t����64T�B<ԌE��HGZ��~��L2�H"|��5��x��n�ި�,<]OP�!��	�������3�q��*�ڭ�&�*{���o�S��3u;C̩Ҩ��c������lZ��~�a�F&1�M��3�S�3^�ޡM_ǉ#�o��V��vJX	3�+�NG3_�U���T�����{�*x�ԝt�)1v��p8o�-L�"�R��?����v�.0wy�Z�E{�0ٕvލIW�VЇy��t�n�Q�����q��L��T�Ep����xY@�H~�##�3�-zt
B��{w�k�~(x�BBh%;�JpŶ6�fx�8���#�k*��]Π�w4��LwWH�
8�)�o�� X����t�.�|��^� �4��*8ؤ���%&E7s��oA�<-�I���M<)V7
��-�v�����#�T� /c�'��M6�N|�Y����}��x�a�K��K܉�6�[K]�9VG�w(�3����Z����w���9	*�dn3��A2>���U�(}�����YDI�'.g�p�'��G��B8���d�������h@��ȫ�?t��E��&�B�[L�(G"����ͻ��دF�έ�z��ҘnX�j4�q��ئPF�U4�cܴN��=s7Ih�ŝ�r�$�u��}4P��^d5ߪ��g7�&�q|!	��7�%�6�n��7./k�sc�C�	co0�����b;�^nb)s�G��m���ĕv�9o�i�]%�@@V�M/���Z��q�������E�����ឮ�D ���u����^�&<�;��>���	In\�^�(K�.��&!�O��LTrU9/T�p㙞+����O�Q��S�ɥ��+�uu>��6�\u�!=����k{2��|�:A���ǳ4?�^>k�=k����V8Æ�4nJ,�q�0˲�Dj��Z��N>w�J�"sy�$�@)!1��wϏV�)VОc�gȃx����e�$8��u����yF��N1���v'������9�J�(��Z�[�Ƅ?��P6w�@$��c�bSB��C��\:���b��~^���"��q��T��ibfv�Y�􄍉�� k[���2J�$?9EÕ{���"��\x��]`��pˆͶ)�&�?�'��� ��|[/Fo����O48��[,e5׫8��_��,�ʤ����_q�X6��U�*�6��Lq��=��/F��t`�x�[%Փ�:ƃZ�x�}@N~,P�_��	�B��Q1µ��h�i�?ح��$"O���W<B�mK��:�j^k6����&e��5��ӡ�v�jQZ���o;���L7Cl�S1����!���g�r~�U��æ�`E�\��iv�,I9��0}2���W�1����L+?Y��le�tSkǻ�L~c���kյ���[w�Ш�e�S�_�fS����{L5�m:�&�2�t7�
�f���S�MrQ82�R������νV�зh��B��aû,`d�V��`�"���13Z�ci�|,8����"���ojb��N���=�`�t5ɔ���Y0Bk-��<YPZxo_������u8������Td�|V����_�9�g6�����Z��Kac��M?h>uF.6\���,����|�`��w����8�/�(��$����u����W/D��VJ=ܹ%�c�(�~�b�G���ʕf�\-/Q�Wg�M'�տ����3�����!p�bzǧ4��_�-�>L�y���־uD����C�ThY��&�$�w�vL[����\B��M�nB���\��^>����P:�l���������)f�,KQ��ã�E���>z?ݪ7�oA��Wk��TS����N-ٗ�=�=���G_�R��e�Dy����rN�Rz��RC����>ސG��`x�d�1�1rlk��C���4"5���n��]�%����0PiȒ��u���?m-l?��u`�i?^>����o����4���PͧѬ�PE�/����@+�;e�}�������T�,]��g1F��8�f�:X��+���@e'��L��*Vڰ'`}mh�ؙ�T��ã|���Ư�Ҳ�5)�S�d�u��N+3�QP<5�D{�
2\���["��rܐ;��vI�yi�Js�h��=~���rp\��1D#���UG�<I���P��/�B����kSW����+#�g;<K���Q��ҁ)���=bD{0 ��y-�sǘV�*�iQ��ӓ_�
�����&��g���l��u&���\HP��<�;!�~�_��8�T��N�����+�W�}��5ɧ�I�J��T#?�^8�]���!�Մ���a���r����2�s�iy\�YQǄ��raQ�MA�J���rIm���ٓ��G��9�,6�Q['��<��2*�Ji�Y��]�N��{��LKd�@���I;��.P: ���6���`\�����^�|�6%�2�<[�<|O�C����S�&�Bj�����SɁ=������֥�|]Q�JY�yG�1�ڭ��h�8�iWC5�є��u�rDr�7�2D`~����Zi+�k�qcRm�ީ]g�'Wz;��=|�SZt�z1���M�5���^�{��^�]�nj�s)BF\7�?&9{k�I�X4p�__�g�mD��63÷v�VC���3��j����Bs��B�����TK�7�I�>Ɍn��L�P�/0<z$��/��,�w�-e� ���\��[�.�Ѫu��{�
�x��o\K���X��\�\@�u�8§t�M.��p��H2v\80"_я>&��ͼ�� �P���=$˃N>�v@M����Wi" bc�D���{9+��>��^��Q-]�ӈ�x�ƈaL�BA���`��2��3��T��H���N�t�̎�u���Aȯ�Hc�r,�;[J2V�[�G�߷=7m�>�|�����5��{2IHG�>�E�z���0�e�8~��֧��������>�}������+@̥1���dO*��c`����߿�	�
��N�>�+&��ߓS_�Kz/�����v���'O����t>��A<8��a����^�M���;�6���8���UX_��2�Q���7a�c�;T� �
�>��=x�&Jm����e�C��V`���Q*�p!T=lG��Kԕ$��
��b�oR�A�ڀ���T�}w6�B�}�ޯ�c]S�������%�wNq�U0o�y��ʙ,�ĺ���!�� ӡ!%5�S,v����:Ld-�����F��+�ͯT�V�n~pp����������Y9g��1��ր�M��]?�8����]4o��~9�����U��7��'�I7�'G#ŗלּ2��W�E����t�W%�sDj]��$�P�����T��x*�_��n�=��/���,�Y3�D5yd|#��/��|��sbk���rC��\�s��͓|�L!�
��q1�	`R�v'z֘)�?�ؼ�X:&бG�[:��I�ݒ�ŵR��Ժ���������W=+_�J%� 1%�{M�'��d�ª��h�������׏��b��ޭ�a��h0���]���i�Q_�t��;�мC>ܾ�_��|Sl�b9v��S��߉+SX�L�g/+�IpAx{�U�l,Z~�vcD�©��;8H�`���F_	�@S�R+ h�3yײ�+M��3]b�M�����(��zL��ɝ�3��B٤GP~�v�N%_bQ,��x�+r�ȭ�|��(_��@5-\���7��r(�'pT+(#BD��BWBLG[	����ϧ������M~��]<�z0�9����a��W=�̥ݭ�K��؄���R�>A��/����tC�p�w�h�������V��:��3��/	纃�����i�����������C�c�լV~����3x���4꽺�cl��������Y����f�@�2�g����p�^���Gq��1��˯�D��H>'�|�yi��
�+9�}E����_X��]�d�: ��jiթQ��;��$hbIB�ih�Z% s�'�����ι�PI�=7��Tn��N�P�s��&�W73����9o����qZY7�*�[�h��Ä}B� |>�J���7�+��`=3ӏ�og�!�H��KL�Hz��k��-��63;��xmcņI�0jьSc�`+��hE�� -j�}�A�
�U8��hX�䰂�q�!?��G�9,��<%�hU�������@��[�N`�'�2ed��@����7�B�y�e���v��L�����*��՚��<@�f�g�x۩�P�[�R�~�4]D)���+I~�hzi�v�?@(V�g|��V��D��wdq�f��&)��_��r�Z{�VF@&�L���$7���:l�*�Y��:�wT`tQJ��[r/\�q���DI-QD��&;�(�ܝ�.�)�$W��'��0��+(ZC`��`G�\D��4Ӈ�ig�e�ž�)-=�rf�l�I_�cK6�C�B��YKg>4�S�[����Ð:�*�X�η�OEP�L�D.�����K�����*D��d$���ASs@�+e��a�9�&xH-���c�X:����4i#c'3���Z̆*�I/�3�c7�f�І4�ި۹O ,���޽/r�i��<�6{�Ū����|�F5�*@3�j���6�Xn]�|Qߞ���)&V�,D�X z�C�����r%,6�5W�7��A�
?o:���b���_�H�L=��ǭo� ��֋I�-�*��ܐ��k/��s�Lb��_s5�oYpw����c@�s��A/�sfKZT��{$��h�������;���Þ����un�VxϿ�ڔ8�0WJ�����I��|���6�Ka}dG�gg<�4W�ا�%:��s]} �ޥ�نW*�ս�ֹsJ߹���2�'��r*٥��*P�;$���H�X�X�I���y��#(����J|Ż�Ȧ �n��2�7ʬ�����
ð�*`�@���W*��F��5�}"��pG�W}�	b>
��>7"�%~$G�L��~Y�
2��v ��;m[!��&�A� f�Fr-}�Wm�C�oO˄0��
RV�0�LF�X��q6՝L���ѩV�b_�E�f����wx�)28���1eX4���=�Y���	f�9N1ZU�i'�~Hd��|�&����:�K��߰mv+z*�S1��\����=h}�U�s<ޏ�3s��9AbЕ�ҧ��	W��<̍����{���A,�V��N�I�b1�z��ڋ�b���#Pu�:ǹ*s��Ȧ�$���m�(>�&	u�����9]\�*�8��T1��<U��}��
�B�Bd`�d�x4��+l.��+U��8����S�3p�r�pG�K�i Y�x'��� �ҁ�a 2��i1X�Y�/k;Xr�)�7$���}7�<@�a����;t��Bt��dfE�jZ���{� o�x�=�9^����YF���ߊ]�{ڷY�톕�Bd�<�tM�
�W�SF5��خ&#M��`p�"�I�?�St.L/~���K�6Z��!�[�e�2�$��PȚb��Y����v�1p�u�&b 8E���M�*IKj��q���g�n7������i2��b�\�:PV�z���-Z�h�g�AIBb���fD��	���_*�-�_k��t���/�X��� �?���`-�\�\���1�:��~@ �t"_���xh0�	�B�g����6�}ޤa3�ba��	���V�dGj�[̖���>hȮ���A���9�	RL��T�Fh���Gop2�&�PĿ��X��p��zB	a���9*mx �]�śn���O�$�/T�u��n�ayvt�A_"ֺ �˚�M�7��ofE�v��_f�҈e �&��h)��N [}��ݷ�ȼ��,úa�*0i���s:F�^�	�8�ęl��}�d��C��a���3��2��ε[��z�d����y<[����i!��uÉ�q:������������^�-G9c(-��$#�/Lu�qR@�$y���7��M�|w�6h�NZ8���>Xџ�"�Wb�m�3�YA�.�ǵ��!L��m�:Ճ6`U1���X�Ú������S[�����y�[;`�Kx~O�k��\���*;�x@ �Ta�,���>��O�M��^��<�3޳�7��a(���L|�6�u^�Ъ�(*���P}���p� ��/�J�6&�N�O9����t�R���+��̇���h���(t�T�Zs
$��� �"#Y(�/��zX ��`wJ#����&�����������y(�ǽ��֮D�ʬ<�n:�A���AyBUL%�l>ʤ��t���AR'������ky�](WVRn����j}��Pj�HƐr�����x&%{��8�̕���2i<�i��l[B^]᲋ON:o��l+s�.�k7G���Z�@\A��c�Ȓ�E�����k���Y�7tN�{�2h����øZi�2<�)/�����G]\��_�L���e}<��Z��P_;����x�������R�V�Ew���CHQ�^(|,�o} >`��)�����jd�[;fS�~���#1�Ƒ�bR#����jK��x^/R!�Z�NN�
'���h	��UT�f��665�����}�Q��%3�����UH��n��|i�H�앙�6>���>,+�"�ZY��>B�NK8�et�1�'�=�x9�%��J�*tȜ�"�y��"��#'�s�*���n������%:�
Gs�w_ΰ�D��h	�U�*��M�&W���)��$�g.�@�E�i���3-�~c�sp���h]֝���V[�XL̿�D��B�9_8��5�f�OD?Jvm$�@Nb�1��j��,-����{K��|�)n�Z�8�/K0�ժ�;�g�qW� �*<Rb��<@6�֘����	�W�`3�4��ZEY���F�ؾ�K��@ӆN$��$Nq�84�S��-M}*:[8�c�y��x�p�J���H-��٢�����C�x&߭�,u��M4W����l�w5���{��psY�z�0R(�m�2���xM�ofTi��V����4[ߍͲ��2ט�
��N 3j+
.�Rc�H�9\��!%�W�q��7�A,��̬I�Ո�ڸ0m��Wδ*���B�n�舻��t'�+�6
F��f~<W0�RO���eX��K&$�����I5=�-�#�U�7�	�
Ș^1,f���C������B�X���j�@�� �L��H��l�(�1��S?��"�7c�GU\��n��Q�v*��<<��$Lq.�K8�+�_�m�Yr����8;� \J�s�^8"�G�Ԏd9;	Q`��
��}̍Sd6D)fߙ�,>.t��~H�����|��&�ʎ�H@-�����8[�ks`�r�J��2��D.}���͉z�#o��Ö�`��6�I<V�BT�~���Q�,76q8�l��[��?�؉�P�s�M�W��~c�"-}�j_�p��>+-rY��ܙ�,bW'٫�~_�u�,ᒥ;)O���X]^��&ߢw�a�Ro���XU��O��#BG�yTo#n�lg�Y��W������(�� !����� Os�{rD�[�?*EPD�1�5[�