-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mKVqwy+9j+Xm7erd/SOfQCns++YtDhjoHMNUoU9Ly7XFklDDfRE+V8KRwDlcxNFIp+CNVi8DNHk9
0lySyGrj0DdV7BRvbgwfFsPnxyMzfy9j5Rsa7jKFA0xUa01rK4ugRjHwISr1lXDzOlrMHxJiaab7
xhtRv69ys4w8ksvB2n9uMauekjZgu1sfqHgaeBtkGQBO3cR2Xeg1E0DKjIaiGqYaxhcw5uwAKpvM
IcSfNYSycaD/lxZXcJREwg2ne9GtGiG/m/8pC11YlFFuBDt2ltGDR2ap19RLJ5kbxcyUMhqkNv8e
bMC+wXCLH4J6U45UljORxA5FUd0KF5zD1H8z9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
Nc6NEcbkkQPWd/mvmwU5M/mQdi+K3RdGozTYdQZwj0i8k3FbQMouu2ynZBIfa6uICV7VR1jEjiR8
WzUwR0AG6RGAnW8fNlN4BDEyjp8AeEWn8OwpoEesm/HSEpwYrcQqfCxvQWy72w/B0ewkhtO4NORF
7IBKFxKeVdcu314rNsxAFsA1/R9+a2q/CDSIj/csVoZ90d7rNNXdNVmPHVRiipl2XxR7wrFw2mE2
hoX2akiZ7C8u7qJdLyse132jtoSEm68GTfJpgNyu9PGOHi6zzuSCpV/Gu+XPz8wrve7I15tizDVH
NM7xI/7Ghc0t3QqEveO7CFD13srBo7zBsBI19aa+bwcIdex/nNxKfFoGHpRorwafEV1TfUCcjWvI
B9iTL/HmP6ud9P/opwVjNWsU+lLKHO/rJ6WQaM+w2c6PiFVtPz4DPpeWXvCbUtMmaNxYEXA/Reuj
yY8W3U7T8pcGPOg3dnwqPfPBgPdTz/z13hnPh2DUIY+oD/+Se0jLLjYg9+fiwtHh463ndiy/0dpY
U1M2IiJ7JAJbr4hwaTQ6OG4/g7lw59Umj3nfWcSnr74kO7ZcBV8gdskga7f2MGs9j9fS8kdqCmL2
hPsCiHDBqO0sJ7fUNi0l1Onf7N1NNGScnzATjhfZvzA4rUmPdferFKUEVfoTAqlQfxYJPUSWH14a
yhBKyUTT+oxtitvmU+nmQPe4ir0w6Rtoq8JpeunEP3hrRu+D8MsNSOWx+izr4RIYlniTz6kItxV1
oGxGCl5XDJdyxE1vLPlrWnUggiOmeUTSxCvvcrz2Rinj988gekdgd7eSU4UBvysOqOX+WJTFztZF
2cCk9fnZMX23o8bXFoMRpH6KCvlTsNzxutBS7X3YKYa4CtaHaVS8n1Q+UE2xc5wpOHTxDqFJ1DQS
MStA4KnBydKSKB8lYYHRfq343QGwONS/0yowokiObdZ+KBA0XOE0OFm1Wlr9RVAkzJ0iRsQKS+a6
08mo83lIoJPWKkcs3oaNbvyp8F1Qy3KKs9K+SWtxXFhzPdNe6P+2w6RD9VYFW6j/jhLFl1RoB3Ug
Leh5KbNW1qkjbJnq+ZaOvBrHRsyxILikZzdaoIATldB9Ar15UjZ9B0y1IDXGgK4fKsu9O2Yh3UWK
ydC7NeYgWh+oFhuFj3V4rz7Pe4vebSxsVJnFNN3dPQ4rRAZMtHbmTWg1PR3M8oeKzhjsL1n7Aa2l
CPvkhngbFFtUguHNnDBl/6PlORMAhjF/XVUU6xTqZwRUXxrHD+rdJgYSLoYR2gmwFRBkrszRT/3O
jLkftMjPZsOkERBuLUX0qf5GnYPL2QbREdw169AtbThvI3YyTMK4Uu5oYa33S6UgFeb3PzUFDSf5
UNS3lnwSdzdLZ1/5ymSEfOk6UeTmjFms3UHpANoBDAYd3zxTIW9Qixu5zf/GO8IUom2NKIkUZ6eo
mUOHxts9Zorcu3F5iFnqPHNAnNstadAGUqCJQrVhC9bCQCYbY3Xexw6cuZd8kNZjga1J7RxM5P07
vp9dat9J3tu6qLCb31QfNIrEPr7h65+VaTP15NXgOVkG2xJUCEIgXMgDoILh9H2ZnsmCUeCfUrPv
qjr+lorcn0tfepVf0bCN8cl/x41Xfq1TEZEQEkE5d/iWnHNtVSHN49osyZn866IMXp/o0DKqXxDz
/ENZ4q7ADM6WieVSJk3jllThlHCdKiIw8xayqCQbcXwuIGGVrF6nEqa4gXX/q4gb1VpOAq3B9Buy
8FMNAUFNOwBI2VaStX/ML2f4lfI1pJnJJ1cgCQgmizIezzPoKyVfuMnRR1Aq7sATlVRcq05MF36M
FpHVJ1fOTNZV+TyURFZdRnqPOkVPOXq55uMc4eTRuYKMZV+MvVYphtt/J14lLrGFDEFzZoHGFERh
zU8vZas+CcF5PJUFKh+nACFpJnDfKyu5yFRPwqdtXhUNagk+VH+uDNo0pXvgl//3Sr7A/2n/6TKE
pS+Hpq6YuG74JUjkiyz2Td+HEnuppgOSDQYLRfBb7tYWlU52Blo3sxavTjTwFCKSZ/zkyeglotb8
X2Hpr9agEum1dJDrSicvZBzNTCLhyWf3hFVdErZ/lP07eMHvcMUNdnUwZT7QJ4BtWzM4SoD02Psl
t2zf9WskSRzkZkmT1m7GLMlpbDu74Tsq29R5kv19rhyoSldZVhGZK6qWlMySs5Ku7kFZZ7oBwxqQ
ZElpyn27UWYC4Z/1eX5w+5cFcOasyvwZZ/x2x2D96m3iTAqj4EIA7P6Yb0LtQhtaRYmrUaspTHPO
3tJ1paaFadYEng6hZNmER/LePeMK5DB/o8y6TkN7M1n4NsnMhHbJbq5EriTQ1iscyZkTBmSBsohV
9TpNDZpcR4/1SajbMGyCerXae5F5BUPZrInsjLdWzErRu2S9aA9d9V9KjJ90UJ9DJ0PZa0xRWsfB
f0thBeWw3SkDlgvv5jWX/DaDVn1Q7P9+fFxBzJIaZ4kVDBwv5XC07hWcmfl2rgiEYR5sWHG8AqP7
R4rJ/nmEBYrJQhBSzcmo+oWSqMV5mFwVsePI3F/ZyB7/BnQYcOcnawb9rG9wukQ9VnZme9IGnZSX
2y1qKtPr0MguEbLD3VnaoKpiC8dk4MzNXl4BBgsyjwqGMcVfpIY7jfP5F/z3ZYn0JGLO/Q6ObiOt
dYYb2GaO2ZA4PEuM0LqeF7U+zCJfxTzNCim0p57k4nq/OGZJ1d71hA5zH2h+F97ocVi7861kQytl
FkSW1DfH1+xiHDz6EqWOaLSi30Zdeq6ipOzwg3XVVWUFI8WyiXChYVN2CFwQ3jtxlLQ7XHJpONz2
FSNH6nJfadxM0PlfNn1ip4IeNOskxR2aQhBmoMrkV0j2mIbmSPNjma9jCinImI+Re6AWgFPO5lAh
jrG0gmCQ+xRVaeT7Zh8YKIWqlvKs4jfdte+oWCdZVGzTs4xk2Gc8K1ctfwMrUY0cGhoxEaiX+Hhq
h1/UUyAsX9nzFqHFADooxWr7w/WvtyDHt9JWHle7TFrKGl5PTH+qY3kEo29sX7izWBo5gY/PKwhj
Qi5vIF85KSamFmWUI/NUGdgPeRAZSikjnEjnTVOIt+s5qscX2U2p8HQVDxgFin8IiuQIZvwCLcUi
xdNUoC5BsQv5OFP071iiSK00jDluIbShUS8CPQTjS8uQ5RtsOXRMjBKga4T0rcOvbpU0UQrQXQfo
5AvbBxA0IAuelYrWNykHqCSAU98x8hDIETnf8XrJHzGYyyYteqbC9ALz92f9zGts8jbGlsKZw2Xy
zWJX6/98NRAAk/s623PiEjV65x/a8DLEqVKKOyaF3gaI4VIF8JB5P2+8ZikTQ3NAafWYoQw2gU8i
QYIjWThRbqywI/su22NA9M4kIybNoHJOWZWHP6e+/Qsqm5iYRq8tIqf4FcIY+23qA5nJ04FqlCHH
DGFAcuCHsOdYBmMKnvsCGtjb4vmogaNPNSGCQH1qqfgX+lC6iKI2JZWMoly5M40tucRcfDRLreGa
lOCGZImxyc8Y7aQR8LDC7oa6Dc6w91UMoG8fvFYyqi6tvJ+zzqhTq1t8k0fldSnR/mMQpoh8lwmU
fdCzahf1EPqbS2NxKYIvt3QI3vAjq8BBpPCB6VUzfzmfH4lij04SwsdWTqR85qLiZBwZVNuOxktQ
LZUmppMEeiRcn/K6crIiOXZLihc5lYxMGHLwNllT4U+iIKqsc/XLHHMYuc9VGqTMmT59vtW91EHQ
a4zpQxNnTGOB3TBQAfHDqCZ339Md8sEhKWeVdJFFS53nMEH/X9ZY/Z1WXhpe7XvSO0A8pK3xRhK1
ebBPVqMXp0JH7X//4iSQq3IlwC+LFOkPWU2tZHXc9Ga9qBrJRQJpGTuY5OLdtBR6zA69eAUjhp3F
b+4aaAI/IcDW8CtnhNNZFKPuS1u6TqBZpfX9u7lNRiTkk4dUMu1PJjen+rGaAwRy5P3FL13ksK8a
J/F5cZHkDYS3Maurkl9G9ndKDesx8hBbmtiBdipVPwFkvJP+Gk1+TOzF1mOa0asnjdJrT8AdSO6b
/UpClSMDzLcTyVN5b+rXCbkMgnec6HRBwyPdSaPNMQTXoxLkvSD6arEss24lCXtAHRfIcboYl1es
PKhW7kXvPL4Zd0ioLToWjVfEbtUdzXyzTUmfiZet58wjxuJvmZn0s4lfulY0K3VdJyMvP+jZnu9s
EZnWRk6k4QAAWOXiXqaPOIAgY61yPuXxlcCnwq0us6mUbXejuSTyc6kT4B3VG8ldexuCwyDKU/zH
6wuSudcCZgr413exuYxjr+OW3BygnV7IJS+dj7uWklJU1PllStrIJ1hYIH4SCA8StgfQQK+dl9WW
grIaqszA8/O65csG+CYI7jsX3e0SROi55CNhvSLj/xUqbT6YtFt9pblk+Po9Ii0EoUqVF5mKet/m
M/m+ofcb7dR6FBkJHojQQ4ggV+B+QfENrDkpK5efN/mzNyGKkvxR+A7ZSRPAqHQozkbJoODbZ/eC
1YfAGYRrR5buAezZBkd0lx9+cY0Ps9RZY5neqvnT2iZVyuQea+86IsQz6Wgf8nXgY/FjARkiNoep
cHrO2vavAxh3IyEPlLuEf0wzjRAt+bSBHMfDUNlk22PbW8pn2svDNsDsabChZo1Y9YNQBOZ7lkwV
6uZUcDwgzS9DiVZqtvD7ONq/VOkB0GMPYZ0/wKNHfCUSkXwfjo7m4pD6CcqPZF/59kbdplQQM7yM
qMoeQNBAwoC6cd6pPZOB4o4QgGsfmpBZuJM4Ii+JWKOy0xU6zlSoG8nZ5TdQ36lP02WUJ03QB+3C
bR7XPkGBvzsIqG6+FFP2H+YTI82TWY5+PYz/vY9lwEvX7bPloEkB/7Gbd/pgpzPU52mzWC6TICmo
tGEmUiWcO5F80CxFAmoMvluHAVlYhRs3DWSVAZuZ8PJY9mTR/ehfErSgfulsglFI6GNcMxpitAPF
F5jTq5fNmXDY9KA2qEPEprm4ixtgWEMsJ8wSuVIz4cAD6fkOopX+EkZm6xWMNp1TNZduW/y2o6Ce
l4333+8hRkZ4BmIZtvyOmzYetBKvaaTLzuNrDUuiQvUP72V1smJxkkENg8MYxduPR9g12XDu+Aln
t5itF9fCeqcNZ1lkXq1wtnTjSazqfdUVGAlBh1tUmeyACk8XGmLJ98DlG4hoVWTXRPddGOKT6707
wk4gIlH6KcbRTBoaFmWiQo0nlc9pjxtEy9m6FcYPWpYdbFYN3PszA7cgD471sYO3DXEtYP921E6t
+3piGi5EZ4EcZoTc9XnvpqsZnKnZz8o6BivMOJujfMBXLARp8omRTn5GL1VewdFAS7N0DMc3/kzo
JtQ1ZR0gCBsfe0VCC6YH1mnFd7JJk3pJaX+WJTzbT67ysTJdqzsNtVAt5zZitkR0ays5TgNrAWwH
s8KI5Bm+46zl2Q3WplIOUrYT5slSRmCGKmj5utT/dXVPnXCSCCBb+ldBzIttpdWku3K10T5acjfx
Gcn/uPgVbQHn/hx72qU8rKs8hzDmTK+8K5NXlAOZH0Vg+W9s/fwWh8Zafkq7NyDTyKWPSc7xwoAm
r7BKlBz4cEPIoalj8YRq1BrKDL2oYMII1Rj1WL617MnD0Zewu5IrQMTCTr2NFPQWMJw6/ghB0FAi
6gxDzJE8GZNlME+ERiGovbl5WMccZ/x+PPxtvVDM0Bg1OshCPuLTq88KOBGTqtz+U4Ccf+qFUJjB
UFtu7s5Ps6yRNjcrslOAzxDZYeoRp74B4NNgnbT7LUGw0CXEOL1uOyA6FSqEw3EEJjgg/w+C48hb
rHh44o+lVmfEM1DqYKdHhy09xqNd1xtdpneNK/r5nJZonHBDExhHjY1r4zWOVFZoQgZk2PV4qGY5
+VfWr9t7MrZzRvGr8g7lRZAh9gy/HsaILaL24b6QSIhuC/Gr9cyT6qrHOgijt+6XTOdRui6vUiqZ
KCoejn+KHP9MCkJz0736jc+LOoYGX/D4XRFiUNW3ncP6zwjV6wfOnQNdi5AVMksTEzIMRrzK6/Wg
47yHS9fsw246jQ4w79ybBe8B8STDE9hap3YlGndpTBtnxJ76wh5rUgTq4/N9dKNN3zqZfII2fNfI
2MUvf7TTJkGbD6mymoxnJZ6R6/AFw4+2aGf3zw6OJh3BrBG9Vvg3iFnsuxjWlMBX93eP3gYXvXU+
s3NurE7CgGXa3z9OZsRl8M5kDI7bVDYKdxwtS/01UvbrglzVc7Vju38BXIY9bnbARdE6wWpuGq6K
yGZNGZqOi69fItng80L1VTwOgU9YFhfGG9rjSmkTXfAVmP42Y8+svUNZniLLCzKeRYmF3MNh0OYu
VPrFCAm1I8OUeGdfT8hw7HlqQSf4zsOK1hybZxUlRqW0ljZxxDJ+DcwAxBXcjP/hBUfo9sJC8NTO
7j43j6cW7PfTgcLAD9oW1FZ5t9shuRg0OMpIWzJGmCPyaiuJHW+lliSvo1Gq8S0567sX51m/cdpv
TV3wpY7bgJlFgIwuZC4pNM98elGrxt0kJId5RuCMJ5xlRAspGDKQ0XBN39Z3lTIq6hZXFu/w913h
5MElTjxGbPTSmKTmFJ3lvPXs+RTLOtgcEGdl6TaJjc9Z/1L/A5GgZhqzIMZ7rHHa5zcxJnaAnEaL
khKbQb7KZqyt1j5KYPdmfT9xAFgYoB94OEKd4MrA/Rwxm7FedO9F1+J7ZqSMIPLGjBdiGK70oh/G
7lbEsub6Uq9rHHBqYDjGn+ndWiTi8XLMVzpLBphVgJzkWzrAgenxVXKsbJPZg4QsJOh1illsnhVs
uwD4zMxnGznG8SkpfYwIT7dC9oR9pCMG8NT8L1tHqx6jGOozLL9UlMFLqFh8Am0fRlg14QD/62v4
Ksi0vcq6LdYlQ3EiDbAsjUfiOT20rm9GR/AwdrZ7RABPdJBJbrYiShU2xW1SpbgOafKHVxA9cnCO
HgwFL8he1S9oz8jseDaC2paMEM0/TwklHOmGBTOyXmkJHBhf8CaYFGVZdy3qeYk9IU/pSCaDExKI
K0og6pxF30jXxPPZA98yRYSkRYsabOg9TveYS6/GRtHJjItwyq4Mn7Wl1LBV2doKf4jUv+cRGvJV
iP+gOQZQjLMtyRH0uVnZ5FbkBPG5tRUu3VebEi/EUnBQXANyzMx6K8WuraDiCMtFDUq17yq3nFso
dLlxOf6SUOnNFIBoHp/+fo6OEiVvPH8oyEMKPsC/uiPoXcy8b/JqK3cBXnYxIWrPfbzqb6SDmOoe
NJQ5WJweGbZGrLS8Jnkb7pO6owqW0sYoWvICq7UvWS/YlS2j98mtYH3/vXLenedZaqardf1Jj3Td
8cXNCektBFYnf7tgcN4Q4vRZA/BFxErVf7uatC7bDCRVDRbWLdFcbrkcRKCIguIo+jXXFggVhV9S
VF9HnSHB3DuIk0Ih0FYgtdws/0AJ9MZ2ekwwtHpU95oXRg5nGGGW76xg/GA3M6APngmSUFjPL2/p
KQiNiFJG3bq9eFzgoEbKW7jMtyoFMqQLCauCkaJgXKVfdJ+Smo6gxHt9POXhZbxyMcZptXeXqwCq
oLUK/jcOpmzBEX/mDEFWSNpQgMjabkWoNcHFDhZqqxtOCs/ldwTyPlooFsy1zjLuHQ2pstvtFgIw
lkJY5V2b0N2BX++HbU83plvHpkN5EVjzRyMewLrT4fTP6U6HialhBzZoumy/XHQWkNalwb5IBiGT
1Td2CsrbNezI1gVI8lQbPP1lSFlmGtAt9W4dn+4lfXinaPVyT/AkM9g5Yu5wn5zZhd4JsJveXlJX
ju+X7pkey7lXuGMlJ318/QOg+RcJYwwKD+LMbrVcLblxUZwXYpjDnNeuelGdi3YN9bYg1iDytEfe
ZCbM1W2vWteFhc+4sJ9d8IRGKwZ3Pp3JE4pdTUwV1vqKTNgkC+AUWvxD93eo3ZKv+aCnQH2Iq7Wz
+MkJwfwzCmrRrQqu9z3g6ncvJlYr0/E0DPzXvjvEetmZ55iRUT8rZv6l3OGkRD5lcgr/j3w0rqV4
2PGqBxOVvqjsBG0MgXMuIB8mqxtBrwC5w9xXd9SObj7bwkVyG1BoURZhMlYP7Ek2LQGnAxMujNpo
WPww9v/2Gs4bY2Ti8gEql54yn7rmtdyaHi77pTDkXQi1gr+yUaiIiG+YnVVWVpv+CBfaosej1RRI
erUvMJXmcKv9htokyUmFXApbGnJl/X6zfWbC7OSeF6ERW3H+rCpjUAM9EL9Aga5qSE4yNZUNhktV
3O6DITUOy8+lij7C9te342aNFxv1aZRB3kq5eovpXlH32KV1Zn/Nj7Z39kUIPxMJTltxtjWay1UJ
h93Nq0TzHVaj4qRrdTeUQcKnmfKVYMaPuUJMAXFI98qWlRTUMl0BeARpZ9pUA7pqvZr1sYJKDUz4
UeEG34uQL9lMd+a84hQMLBA7pt+mQLjwkv1SNQmKfvc4klx12gDy9ZCXsVDLlRw3bXu+K3UO6PaC
390Wbxdin9U3ZckNjink5nHBX7AIEfJXeJBo3QeaqxNNI99r0BwO9afADxLgSqVcvTzCnjEdo1Z7
amGoergWGJWLt0zRwisi3/ZoqefRI7C0o6MfXIgUzSH8aiT5d+Q1j+bqnAlLHLmCtn7sTgsBI17R
3KlyJpP2UjH9lpekeoK4FRXHw/ItQBYa0tWodxDYFLKoROHj6OT7GyJEaN14euHjvq7O63xWk8Dz
11hN+ieNl39q7k7ETK1ewa0M3kTJN6ru10RqYzLF0UcPjSM7ulk9msE3687plgwRN6L1PxfG7yKG
ldwj7nBB99BHNbrBJ1I0FXvWOjMMjpiw6jRo1Bp4JkjWpNhEytJKcVVQ6M8j8vtzquF0kKstJvjE
QQ2NZvhR+0Hf/+Y9nSRgcE67d0WjqJ/Pjk0xn169it+uMtrCv9Jj8pT64wyb5xIlTmTQ7QjGGLDc
QTcFdTs0F9NsY7sBo/4Y92YTRANwbSlCLgeENDx53rWiEf1/rk27I6BImHUS23f2FugUdqw6iHvO
EdOLcbw4tRuZYN4jrEg9vdbqRcu11y66j3FJvnTFvKQODKK8fFedP1mm3bhX+gTiF6ajoXKMOYEp
G1iq4LDglxl9NNzyq62IVejrc0RaqvarsJn9dSqlSBfMHiXe44VBGYHX9YPMfZlijcpiq0Zu0HYF
X/8ohLGALKA3ouXIh9K6cZmkXe1NNunQd54KcDgYqIpkrIFtYnyoHIMBP/x/mUsa0f07KjokoIen
0g4vJ48Hq+gZJZQS5Shl3p7VaB/BL3wdzCcoCAk2r+06kgcuypTeWxH3wTTEK7MkIQt5Yrfap4vj
0gU56OZ+QHPxZXqb+0q9pQMTgmFTXnspgufdG7H8aqanj1t07EOm8NH5JRmNzKzVif1YcPXvAOLz
q4Lt307zutiI4CTYN0MnwbSMlpn6uGbXCPvrtajRSosn5f7rLz+iKyaNEFbZmF6SNscRVdW3IFUZ
IEDVvaeaGuYZSgmhE+Fv1hBis+7rguCp0QxAcDPuoW4dFXOC0irGPA/EaxqO6ybyjULvX7au+ES7
8FF67EsUzq2k3kan0b8W2+Z/vUNSmYr9Vjtmtx8DLYh+ZzU+vSvrhKxzF7GKYPc1vtxI+81/Re3h
RYKt/e2Jq/VmfyetHE5yynckdj4cBR+cUXZxL5iOb5SpzgCJQq88v87ExegO17bwmBbIjFzmK4ft
YEtESbNteb37HSvPwQ1wSuLhcLK+Hxt+FKy0W7NG2GADzzP474G65W6/EEvcGndp+dnbZxcCY+tb
Do5wb8NpRVGMhf94873vAXUZsCEDIpnjfoZcrhKI3/x+KMtCFaaIkYN5JL5CZIBuF3y7dY1IQdFr
R51hME9Z9Rw4wV5cPzD0VGhgfAmEv9S6eg/BcV8GSjGkwUeK3NDDDFCkqyrfoeaGjiftuJyRpWZR
BJTXuQ83D5oBTIiO6nTlznjijyFXf7xF6hCNebOEDxaKayD926enkq8Kga/k0HyUTM1dRco10KjN
X1cZorInZQBTZ/Et5JMwjxsNBK2ag2WBMor3uJ41tWgvybMIWMJd6liXudxExwoKtIuRN9RUvloE
ABsGfYFzI9v9QNqBSypOkUNtyBD6qqX6gD4fcFQIyu/QbS2n4GmBoJD9bQqXqQNPYpgt0UK7LSFW
J4kv3qct2UEz0ahAOiujsquyMT8D4DOwJeghsJy16w2xDZUVF0Ofm+0KEns3+sgz2KrosT4rQ+49
I8Tyc81/e108gXhdOGJvjSLyiVMSsld27Wyru2gITSyrjbwD8tBuTFK7yb65aOKpyppLSH0hmY05
eB3D7lv5lFmDU0NrL1Pcu0Aq5TRO1tde8fR2C/30DOMkKTlyrG5ZRVYs/Mq8J02IJ0O8l0QUoJl5
o0wF4w5MIUGBJGMyfN8cAfncOC8ZxczMele2eDAzSrPFArG4iK2BhcQxwXK35awH0ji9RnR0Y8Rl
L2o6U5zFoMpu1CNSwct55u33XRAKGtSOBXYzJ50sylgftJMIkC413raLHT6gp2Gk8c2HUEbw82Ho
PxwPzmzX1bpwCTkiC1/gHIIaUo0q6D+wOzrNHci0jZhound3p+Cz7SD5a1Rp//w8fLiyB7mwpzGM
Ps/C8tmBKVViXpzCu7JmOTO6BHYOmygi0vGghtgM8oNHdIJ+q5S1sIX3szyBM9IDyPfs+7IvYlqF
UOz7P/+09yL7Ww82c26/3Le7axUiLXqndsdnDxJwM35OgBtykUVbQPc6TUQ37fw+QZzI7JxTtmNl
E2K9PMtsrwbyPN8ws+gOxM6WEIjcLGz2UvJpTKj9NxHNac1Q4NKC/3qVwcn9L0TyBJ6jStQMhIzt
20sP2gdS3hXoAQQ8kbAfZ8KnQO+vlNX860ZprnSCTk3zn+x1WVx1/aJL39Ll06YvOsriAcT8iSkZ
eoa3YSne57rnqi9jYDeq+EE0p5YnE1+5AUFRD+z0ZqlZHUeICYP0t72YoOUFbZGKDFVtQy2rzzMw
ldwDcY5gig1CFn14JTQizp7KtrtWQ6QgGpQWBGS1x4xG8CHrksKFEyEFz7jM8CiuqPOCJ0xnu0YC
RWTwSs3lsvfX0wbzkJhMZhdBjLT+x9cdlnIweSdIwCVlXhwYhw1800pC5tYCZxNcJ01TYoCX2rH2
6dtXYbLyWL1hawGkW8ZQqs4nIXu9nNSANWdphyQeSwhnjP/ZDVCRskKXv2Sf1oNOrPuXnMVL2+EK
+Hn93RFqDO5iCiXamQIGKYhc7ZhgzMT8fZ62fruhTzngahiluDkcNYovru/g5VERy+HZdkbFPaK2
joSO6Yb+YVY04ooCSLQZB+5/U/MnUS3XK7YGhF2mbVpC97Lpdd1mc1ATT0BqBuVWdjxSgZqApiVo
LzNsSjT6gHPdjiFa8UzGrroq9e/dwdHjg6g2+MTKMzzCTiC/3FHAdIJKkGIc8Q9XSKl1bndgx5xK
sHq78KT7uHL0brEoBNkJXvd2mzNgdBtH5bsywCBw2WaVNEImRk3FywDzyRuo37i2gP2fcWdtHAOy
F3qdjjkdKexkY+XKJogGkvaKXvL1Fw08jpOlfw2jgsOFZrgLv8VfY68qmksnXG7imUovkNP+yJdl
HZXh8Zef0mAZomV2Ms80CMfPxf6QpmWwhvXtLOTt3mI5/1V1WlksdX2UOFVm9OwWhjSCnWa4oFgG
TXVNboTGqT2betOYDC4EheXnPJuD1YVL/Sz1VcEdvAaEntYV8LfKjCiheRmWClvAichpcwRnLBzb
7kYtoFjeD/TmFUJbm5sKHvS2y6BaM6pyQILL6sbkE0SFCEN8kr4Bj6czsVYHNwevtKe1bTbggq3W
dApD/EG7OW3QJC1mx6oDNbFYfhMQGlMLuCWc1whhiIeQIuGs+qVIpIwfMVa9tbFHjqHfC8NkmH98
jLmWL5OsQnIGjDb85YSiM0A2udl5LrzGMDyH0BnHDXOWGRa/ZwoYn228anBBJooXST65OWnK13/t
ZkeGT0Cf5siD9kO/EzfcgqdOOb7kaTdW6DGEWWAqa+vHBcceoMhFcvSTj1/nsfF6cPA+bQL7L/h2
VT/r/B1/MQ1uACRP8OYHxvZ+oFxJUIfI+HFE6UbzmcvoZ19IXvzTmgss6iotVLXNyqMPMp6Bpru8
8O6a+YWBxyBO6JK2vxZ4QzT1yub1RCOaiCwkFTqOchKeQm3IB0w3ONFSSCA1eDN7Wo+nVN+/NXZQ
rmoh6fpsz9/KLxPgfKTpURIlYwM48gULRkndDJBhFK9PUVio7sgBHb7GtDZqm1yV0yLe9IMGDh/G
tNX0AApDesGD/ce+TYcTrMkJzqhGAHNzXdfvlxD7i4utprV1w9FCdy2er7pkGIYBgOellR9S09kr
75MqYa+Y2Bzb8qu98jaJFOC0PQXRs6kiwAR4GlKeuhR2+GdYgTYW55iXSci2MRHeIw9eFDFw0BXo
+V9ro9l1pa53TuaX1bHPIEFX+kbqf0oUUEGrAZukFXRIZuR4c5w0ERb0ghlyOmK0BQ8+YjLMGVEu
e8kPxX0hHfF3r/XL7cW3Dkh3W9QS5s3ArpJOC1OwxrU+KeeA+ovD9RISyrmy0o8iuCELqZumGYO4
hUr6o9AVJ+UcTlwrE0hTjXaaJTpPaw8I7A4RLWoTvAizOGxvAVtjIWZgDKyxiN3d1J7uBr/YURWp
nFQUqqUj/bxoDsKQCi0Ksr2iqexvkFT9mcNWeFqMHQYjxBogeYUjtNybTftDD7Pd+4LvLnjA+VWV
Od9vOQgigU9P9UfkIaoy3wEt+Mgcg+3I9rpRpqM8jNIj/TM21We8QuvhV5qishKGI9xLkFOqRPWa
HQVz3D5gnjokJ3oUvP56a1M3BpwglerbDSn1X0/KsXVmFX3Rx09LTGStxWU70OYngjLWzVLx4LNB
tsiODfySNy5p/y7JI8Fu/QmuzgBhtL0zdBzPclHyR5cu3E6BBWJKg1kRPAeLd5E7KA1VAan9D2VU
zfKZcdp75MeTaQOP7sBdoGg7MMQGuXDPeh4BjXT6sJ8Tv50GO1CLXFLTP1w/P0A2jKvPPzC6PIMA
lfS6PPJ9kp4uSvSI3BpmbokwyB8MFBCR4APihStBjoVLDMgMWraxpT5+THOjVF+wWkBESKNHb+c+
6Fjl5ovSXb5GZzZG45YG++13L8jEdpIEe40VTDZzRawdoyNwgaggkO8CVuZBg3p6C7v41K7T1AK+
xZscVyI4Rg4ORBQ+Tqd5cqii+y92RcLPWFpFa90meaPA/6qSYUDwr6XrJZG4cImOIcRWEsaPf+Ax
ixedRpnOITs0HCBkMZaEOmr22uZAGG/Hg8m8vViz9p9n+B48YjBwG2ZEBE7LAHMbuur6WxA3faBh
sg6+jCwKxBh7DU0mwZwZ6l9pc0ENh31CooLBoa9qVMlT8k/lU5UszsJl2rt+TlsAz3Rb2vZX2npp
6g98dsqU5GbSbuuYzScWBP5g86HJAEL5BRcnVsqLklTTL53KjsUXcMETimoxDY2+7nuzI8vlw4Sj
U/wAj4bKlUbUm6gk0IpiMNuiDxNnGrvRjzF1v8wb+W4XxZUbAEuRIS3NMvGkLzDAkAMkI/tgUtEN
dmoGeVZnDiLYyRS5sUz2iKLvwfsNZQDl8QESbWYOC5ms+pLpqfZC1nWuyWt2WA66CbvFKlQq0DZd
ajYU+aBDMssSawwJX1P9UTs2h14U+qsE+AOIyn5ycp9uacgKPyFant+X+4VcYDg+AfQ4DMAAHwaS
4Fzz6avmybk6UrLTd7QRarpCYJqibuA+a+1K34cAbi7jiuxV93kN1xjfbz7Ik8PSt5oz4uSXaEtw
OFjFQI5S8MkW3wAMkzlk4A/dygU1zvUzvST6ucSE+Ccc8iuWxNH/jI6WJ6qpZky2wDVsJaQbqDx8
bTXB/5b383AUOZruAPyaoOOaqJf5imY+L47ooBGr0E96DRmzd8EQ4bNdcg4Nzusb1RGsTu6iJP9u
TldDL25v2+rEJdJY4w1UCVjhxNyCck7myZ4h7EpPF23BinDL0kFv0OK1zqKRx2gYglbJ1aE7NPte
qbS4JG0Ii2pFUDs68/YdlixWPW0ansU+/k1qfACmvuDJEH3UQVw037fR9FDQXOU3V2fVNLaVfIrJ
wbUA1J7k4+STdgd43Dj5PJoen9Q1fH/mEWzQ4loLreFFgBSLDL0jQbwWLubzvtVln4UOLbSFPPne
KLCjyayHrD8n6+W6g42e64uzJEiRII36MZ3dBVI/EqZzHK7KY13zC086V7FTuwJS2nZXfIdWDHiI
npGokjIR1W9su3L/T47XTsUqBV8Kb6Kv9IFxBiPqct/lL0juSda4n9Z39AcPaAJaclyNTIIYgfkv
0BiEVAe6lIF1a/8wt79uZAV2c8ULLbY5sNV6JyzdCwbdxQ8o0SeXz97H6gCiLo2PVlawf6KK9wUc
mL3mluMnT1XDXaVHRxfjydGVvYTVmsyiXTb3qw6AjGG4tZhawifHPW2mD6EcpdEclv7Nx/9EvGQJ
LJqsEW35C0jnNNKGTx1kAAyC4XnGs29QelzF/jwauyNGWZEjZNW+C9Nz7WijiEgrotDmYDfkkvh3
wwj5HXQDL1AZzJWqz9LuNUxG7JcPkfxZ95MefVWmMTSJLYH/GjN186LHJ389OTwUjq4rB8oXhBEr
6MDNnd1aPB1khK9A6VbW1CsHMUSw6N7/IsjU7HxUbn0KgBtAHMVgPg2MWFNeS3BraPVX4eCfl1mI
5WaFoih/7MLLzUQnUQJAOf8TV6bvbfXsKA9aaMeSM2Rnweo1kMXr1fpaN7IcL75z6x7sLSUMcmGb
OO9lHLCTIAvYtUC0bw72un8prbOYY87jcT0HoRQm1w1po+JDnt0vAF2PIw6tvpJTZtmzPlfWTMru
D313Wr6qxma9k/uWtlSHebwv5zflMBOI1nxcvyjS/efD82dB9Ac5c5vTEsNDIyKCbx8d9waC96+r
XiG6MkppmNwy/aLgwEJqBs9ZBQg1/L2Z0FqDOiA4cUb3un6LJjy6NgjYkLMCBAwiHzctitOKirXH
zi9mpsDrWjWvUIVnf8CO90xSDQi9YQjDmiahD7mr86RYJhT69dNaX0YuwFx8WWwbUyXN7M6LKRux
yj9kg7u/TtOCjLPNvb+rxdkiWogmJbmWHonVrLc1v9bYvEkSSGF1g4ygvjM/Cxg9yrpz4/E9RjRL
TCOCVBb/ZqyPFNHrf6Xfmh+CVi7TVBUGcBUg3NSeNc2W5HFLjqvrsRzLysISxV7Bj3BnhPv8iBw4
yM8TZPZJdhlT5QXzct89oYtrqEVcHjA+JDvBFOUpaFcX4IDUzjfGIXsXTQ8vnBrCdoIC1/Vi+3Ll
uE2VjxCzu/zn9dhqe+NzhkhHZAPAiaO5DduoEY5Av85NmuKiSyHg7Faso0JaqioVqvRX592PVifK
Hjh0PPKP0xDnyv+bGpioGsauNKXL2vmes7Ftz3OhPVIyX/8t7oEqhg0U5nLMRsGp/ZoIS5ZKWV+x
UDZX6DUtKlLDX6rNZVy4Kufoqp9I7Duyxljbtp9beKhxV1BA3x5UBm+mDu/9XBYvah9Q6biRBFdh
LwS8LnNXbmdf87tHD4mwbLb2JWA3xi3KNzOK+FIuDv7anu5lcLVB9nJPNxJLhpt/R6Xm2bz+IesC
HfPsRIvMkk2GlOOpXljC2eLz4Nc+FnSuRR+0kBcbhygO2yHeU3xNMkL5zo2ztYhW8eEjUrcwhw3r
an7axeg5QIj02Qr2x6Qzv0rA+qL9aqr9xu2gj/RQGd6GJWi0DY9h5Dbevmed/J4+1LewAtPsaGRw
jItt1+r/j6JmrQjA9JI9KuKMh2ulwsuODOLP6DwdROkn+m6LX/eCdiVyVO5etLeUZpaN7UGaA8Vq
/sfkavejA3Tlm9htAbtVll5Xdm1lVovVxkb5jzJTG8IDrk6e78X/ZWvTDxwekPXgJsb7sEyoCDak
4z2zk4juqz5+8nKBjZnrGEBkbzooAdJCtk23CSEK0T5yDtrXfBUIjuBkOUcMX4Jky/st4jJwMx8h
iBgi2hBfncJPrrX0/VUEkBtjAoNLkUVba0lmvC3mM1X9vCHn34uEWP67nEWbB4yKmSbN3zZDtoG2
zWoiRKNgltc4Z5Ks6bQya6tDGi7t0ulm2FqF7iZcYxi5EOF7Z5xhU2G5FLIwfuTl2UL9Z8aHdAsk
6amOd/MlYNITzCoEAm+IxsOTZKtS+0PLw3G+vwjkcCSEmrBQJ3r+wkid7BmbCeISSrwAOtjikMbs
3X5W/+gtAva1CV+31TZ/uG1n8Ifh7wgHsxer7Ci780qpHzBE2HXH4DGvZJqK+f77dnnh1RY/vhWv
1Y0tLHlevMhVFQXdANgNna2k6pNA2wjxnbVR2UiABkBHtlIPfzytT70ryCmNqKujZ9nu5PNLPCGd
T0i+GR/VsTwfifCMp1LGFmMmSWGyvQyO76f3bbivZwbNfJp0ofPN4rjqZQWQw5Fi2a8TCTbcOb4B
qgIIkVIL19XDhj8PUJyiPt5+qLbkeUopBwlICR1HqjyZQuczs9Dm28z+hBwngE/kypTyoCMCVotj
OBJsjCULVCdy+XlPDaXphmwU64nL4iVsFBQUFfT5/86N7to2bSyr5Tg2KGqPzYCX91GAVudpecrL
nHyAmLycJP3bslWaYsWwRSxCNO1wDN9WiwCKqdChSc/16jqtO2f+jbuwcO8wyJUaWTTnzaU5Iqpc
3WV9TOV17RW4d7NhiW16OOgQLOW/suR+hj2VwB0cNn9jgnaGP9fAh5wR5AwHI9sxXXhS4IM8C6ea
RWEx+P1biyTo8c7Ns11eLdV4DdRQr71xLvOp5Ju0j7qjcDFKEvJM5iw4QaJXsKcth9pz+YjL9/um
GNnStlFLSOdeZL9cUuFesPVlSCU54WmATxt+aPLapa+A5OJ0+zfR8XrK2Fp4nf8fIAnTxCur+4J7
Fcj8HGtNL4q0ZuIzv4IWQNSN/Z0mjaivkkpLkQSDg5z0BPSLWKpfOSckAwx/S61p2HzTgQLQDZUl
wqx8ZIKGXa7kaLmPHX8jrKOLuOHmqXFRoVRjN+2uG9RyhT6sJgw85Wb66kpuCUtCOhZ3FTHv6rTV
hFWL0jZjp1mDtdzL0T0fTQJfipZr+EuZnKcrwqphkqC8kHnJbG+7WlnhMyQNMkaJQDuSsLXmqBmp
TuP84vPsTxZBAbZISoVwPu0lWv+cZ6S+Gfu2bvUrN0yPf/V3aiwefEFO7wl5dA09CuYqFXUO2y/U
34wiIheX3BlIf2x9EJ0K4HK4MPtFy+GM26ynA9Bkq463cVkQuBM0ayn9AvqZujnd43xCUC8gUESi
poTlXm/7PSNjADna/2MIINuJgBUkqy4zAWlE3xw6purrFZX2KZ7VuUJc+1BPkqRezp8YlaIlgzsR
k0q2SdOePQlPMBPZGoIVH9noiKdx4Bl+sU0V9ylUh+pY7P7UWpqc12782mhe57dBh6GjhXydxCYh
c3wqnwrm1dgfqH0EoFaTieHhBlvJeifnYtP0Zp5FXz4X/grDik7ai+O7RL12wvzeXRZekX4QAgQQ
EaepV3mTJjJP5HTMgrN+Uv6yCr4vNQrpAYxf0snbjH2PP9VPcZbiknaYRJY9PdsVUKQyV6ICbawj
fIujzhPb3q0Zzhq5z1E7R0ZVJ8InaR8QwJ/hidiBiaUN6svZVqyMikfx8Oi/4QKNWF2qScHoewSf
4O1MRtojMtpMCN2VktxJRHWy4gbROZhRTwNA+m6MpwNZndYvXsTSvdU5458UqGV40jdRlhHcxQne
TqLK6UbMNh0fYrWxv/Ud0wTl1TJh6qRzelqPPxYLbc4huEZPUW9+ApM41chI3tA3e0QLXudv6dtE
WYMwe0AMIQFA6L4Bt/e2RvGzTQZsIQSEUk7uBGuvyBFcxJIC+khip2xliNeMzlv6DongMukenROD
pzYkqomDR+LHdbPmaoaVSczc++UdmGIHMmg7NSnL9S69pfqBHZrSNpOFLWXbHcGegP6703eatAaz
SF3Hvea0h8RncRQzD6il8JIMLEarSiaDyjxj/JTIdpy3bht2A2DC5OjS4QobmSj6ypo+JUr3KIhC
ksm1wbnixFG6+zxUTAjBUV8kdstxeweNKD7mD24OVWXoz0c2dQht0VC1kofQp9b4dU4/m4RhCQFJ
+ghlwNMEND68Dvjc4AW7CqE3enYWkX8PIsrLwMWNgObCYhLFYnOIO9dtyIuMj4tVrkpuI8dFlnH9
EeudfW0PXN/wpewIUPq5J73PAmKRyljJMnqud+9HhzeEu+Tc0dcu7aGpFTnEHvZKiDBiUG3ai7sZ
fA4Zj057rXn5vZqXQk0CL3eBW1h3b9WXJPVfz9OSKMWKo2VPl7bYgyDeWZ3wgEoQ9u3tmMA5WgOr
jJGSHsFY+TCL+6Bs8Q0ALnZLCYmRxloxMcyr0VnBUXTxpIkVgnZShImk/LE9zLE/Ymb8sGl4Bqv7
SE0Tm+dqQhgFMIEOjCEXiffrCZlcwl/fq0FMtqQE5U1jchBdyIZBISORmFP+mq0LKLEcs7a7dyWL
pZpVH31gsKkoQhBGj8p32jO4PfR8pA0qMFb47XbLfTg7AIQchtY75imLY7ubsk1tq4khS+8C+O+S
5/9o5WCUBUUE/S24stVTCY1UL7qTzOmgailQTEZnbuQjfyb8nTfokX5CW2PqHdsWwiS+YM1wSqEe
PHrp5K7Qpy7zwK23rFQfu9GFx4toiaxGEH2oWSV7Ol1jcESxE5X0609OH9+vpHogWqH42uoLkuwy
dzUnupbsqs6V4I1nUfFNBw5avnNIs6ahJKXoRS490aBvGdfIXtG/xr/KjQG5NTShm576cEWIreFX
0XNj3jtiZ88nSzVJMnHXkUob0DQyHAN3KhMgH0H4s7CXqBxZ5Cglo1nOCOoYzyWg7+3pwOCwMa80
v4Ai3BGEvfX5/5ifkYn42HVSrtl+aPO7kDGUxLGORXQYlm3uL+DL6OcZbqe3Pfp6JtcpNMdBlmkL
ja/6454vpq71j/covRGndNyBeIqYYttIPq+LZ2htZIYWpb59b27WoKISdW7m87hpb3AnN0pa1+KI
qz0h9kRATO9kuZvyf0PFrCPtiiQZcrQ0kFi4ayJL9GYuW7DwvmWcJ/r/3HTnw71WV/mlRuHVYbtI
SF9Lq2/K1O+5o1lZb80G89UO47DCP5BxqxZEWMbSDKFoVFHyqUKH/pXAj+Y1H9lx07A+k/xe8Dyr
Dh0dMliHiV1iGXHq0JwQ72V7bvJPmyD5VicQ8uwbbI6Sjh+/VQyFwx81P6cYNRphG3Wf9ruE/NbF
Or3tSLwEpEJR7OItjXk32h66McRtpYdkF6vWlEOI6OxEUKaMf8csIFD+49p/X770aFtHlcdte49s
uDmr2vVt4EHt39vxZnG4wFGcVtrUbUGHUqj4tor/TbSE2MgxZlsekZbAQBVGYcL1+VT7/plRSLm4
xAFeF2TBm9YPEL1YkXZCJaTKBGfrCljlYDpybMXKAVpAcUeOgDF9Y2Lck3LD83f9GR0iXTjR1sJh
tQIlBCveJMTiIW2AyX/RX9r/dTqzPO9RB/o1SRZitx90ui7R+h+bjyUbwBemvjq6s1jI2H7Hv9eT
6ulE8gc1ia4EIsiXNlwPlPu7LYR6vGxMaY2RI0zHV6b1dImBFZn0uCMlK3kkEx7+jPp0Wjx/A5dM
3W5WtuPV3ZAU0XcdRTHgfgslRdwFXE71nvdu+EhPJF518QqXDAn/hiQ2JdJdYm4OncD9+j6UBx8f
6/hVyg/feRTChXP1+MqQVQ+i6O5XAisDy/IH29yZIsxQj67qXRWkUf6DpC6w9GQCBXl+Mab3xHPc
55FXbJ0P1EasvLgU6wMYskDSN8knQFwW84VTw107SpX8tYrRjiExmX/k7H++b2n+ko5kj+GijGvA
CA9kuuayEQ0jwp2GwT7y8vf1QZrnxhk20GjUYMtjRRD60MeKlgYFPPYXgIWMTD38f+zFAAujiJpk
jNK4/qg21xQFiG1MmMla4XcSzUfdtvleIrAP7Pfdkqp3NB36TE4vs8cP/CyLZjKSVrNT4+j1Xbo2
ULUMS0eEKK7/1X9BU53ZNlnly3RnRjSJW2M+ihUuS4kevmknE0EV4/Vb11TQPCP5UU6toDW86wP7
IBm6tWa2Tbe0QYNsHcj2ZHFnQuCXU8mK4hXgN+ryJLzUfy/VO4ON7O8wVpRyF2HAnSKlhIuqgS7q
vCJU7BoqbuLnMZIiicw61kfDTrMCN0t4ojZXIIrQGQnck3rabeaXlfEcKSV39ps9p6cxQ1Ypz74D
Ado9+KkSxZINHLeDAvxuehla2CDjnZTsZLyZI1D+jtZRs/xxJgLxMBb+LorwkU7AM29idwFiMH7V
I4S+vXae2Cp0EVbBftwx7x5KcERxPifoio+B63N537Lwvl/yfN+/gzGE9FpeJHiDd+aNVyzebFZK
8DcwrAlmm6oL6Uu7H9Koo7sQAXJD5ETjDhockgXmoqUkXbCCozdcpItJEVPTyINDLsZSMU1zCr5n
rLNfTWhbOBpKViz/c1i2s+B4XxQoxrpjRXu05URCglm4VHkD53upXGLsh1kNdHkEhd8nYPXcH6Z0
bby8YxGf8gRX3XP6kET3oDh+n16C8h4ir+lLNiR4aKpXUHlLGmzQ9nie8GUqElW/H2kw3Z2SZ5Fz
Ay/TC9dQTxOLwuOKOxsaCXICmY6WrfokIPtuvPVuU3vZwnubXH0zV7xGALVeq7ZgP58YPPeNBfbu
qxt4OmaBaZ/WWfpnlWQbUIcyCfZ3qvZKYzBmv4I514e97vVSLMjpfTbb16P5ORwH/3m217v9us7x
Tk/KSoGER5gvpKfwHYMbCNA/3RyWcQif+3O6H9EpMBC8ZdS7Uo1XcY/qkq1CGYISKW9ydUvFO6KJ
YNkP/17vRReETokLjDSnjr/CYpVqOvICNMWtMzGYd73EJseS6bDwDlGbeebrf2m4WM4manEDrII2
Uy9zd8dOGrGl28ThHTdqnRwyJ1coEOO0vkrj3Lzu6cyeVbo1CVLfSqo8VKswCtoaN1c2Aca2uCZC
fy7fiRlwtrtenehYxRphC0gjdyj+VUz4pDfS1xEWuwH0V+orJ4wu+W7CPNYVLY/pBCYW9bytz1pr
FOGWKbiWL6eVFtH2yHrWveJwDtZhuWX8wkxvh0qweWJO1qzEm8b4MqDgAmBudXAUhGwtvEsiPKKO
ZaJPYoKlvzPaxknoYS3IiVpyzE5dGqtdRN3VEjDQQhZlYCYGpu/IlOdt24rAUltEAsY4My9KXLHT
mdgbnaj33ZiVhuMNeixTdNi0xLfCP9AvPGGRN02whgZXEv5kibYg1TtTlrePzGR2hDC8quz4Tk6a
boFvscTfOsfGA2+0jXRp640Z9AKYtb6rOGD8lZFyy9K4kAkV+HxVJ0g/WyNFHpdXcUdGyTRJRFWz
rEVK2iOB0QvRjXJBYuzN8enVVBpKbbcX9I79yf/rNkqtlIDq4PHhsP1pmlT2jptSadJieB6CEuPP
AxRUBVB6B58mRqDRukq/KTjTa/G9miNgfojtJj9PXt2NP0oc9IEy8s0W0cFh858LU3I4Ph0q6g8X
H6A7y7snWSkdISO276NKQ+4TT0tOgH+PxWUBpcwO2HFw2tA8cIrYUY70xbG7lwwxukitT4JaaDkd
pO6dDHfKMnh7iegMMOGChevsK7YBqKMTAT85yBiSo33MdOZRVq0hmaVQM30zCoZfYqH7iOBirGaf
dPs/qx0Wq9ujx1zK2SpstlIIrQr4cTIA9ddH57LZpkwpgIaaFyKR/t7hISexbHsKBEYM6G2YaT8Z
udw7qA/T/rnuuj2VwegBhwUA/5ZL5pZCecWLRE8B2necr+D1oC/vzA1369KfUdLUtjTVEnjFMkG9
+PURb3KLv1jZHdUivSwaiKq6Lf7abaws4mHaiixo3DNVjDDX5grj6fmiZysecY8Q7LG8NvraV/UQ
24/9w3YXvX0CrtA4zkxNyssv4kHJ/FLsLOBxtcL8/wLgPnZTqs+5dVA2t7rAN7ZfWxv1yGuiOYcr
o6cQ6eJeogsV7twt/qXmCcjrQJphKZjT4a5RNxLVVyMyxHAu4HisULd3r9cIhAsWdnIbTu9ZpnKH
V3W4TVuNRRN87gB63fane5nkMMMHBq/XbsCVYTOMeth3txbRpX1tDUKzZwxbkXYeFSpK0iDUM6sN
Kv+jSbq8LtfdOaXDAqgANfcXAjQvUvrZFDBjwGqOcOEjjLcX9Gs4WrSuW0St4/R/NXETbvJDmSyD
zMn2mFq7YEvvY0rJ7/J2r7mpAnM3jflsps541BVxFJ7xRCJ/nV7K2JW2z14OvJzUNI85oEzs1cdZ
5abb+3QK+I7Qq+NJXKySAvXLIBszXPu8Mt9/Pc08ka54ahWCiQicLpBIuXeAR1f43ruckKxGmpJA
rDEaBHDvXc10SWU3ZxMpoxJi/XSXl0m7VCEGdjn4eqjsz9cm6bWMdvncJga6dqGNzTmine5S9T4o
PF1zaBdctwABRA7EkmItWe41S9gCehEH+NHGEJ4uzm5kHCagbXU0YQvkh5q9nnZWeJRr+mZ6Sv4x
UWTFmn537vsOprdjplsl8dtIcrCJLWdxO+vcP/aoydFKkrueLorP503Xu5zrvEzzZ7uzbZqk3O/N
Hog4lRSpa+RmLYYQBebD1rsGhSYPi8dVVLZfPcXvY3i/zr9LvT+BJiPjnzwXnT9IGJd1x5zCLm/A
E7VE2ZbujHFB1oZKB1NSicGK9NvTCCDWNPG0fFWKxrOrFJmuAK9lwBtjMrPoZGpelUAoYg48bkhR
uo7jHEGPkPSr4Dnw5NJ54NapcACvoMvAn7vJnOTxdMqZegfKvqC2Ai8vhHZv3Kh670Q9v/okh1AU
1kBwxkcbUd8oNWLW+W8u+wEZmj9MMtQEhjd3J6LQQM3rtwx22rD5ooF7/M5U3Jlq/FVwhGcebcKS
zb78l/t5LlWpbmdpRU2Wur2UQI2AJB+LH6yFzTkJcIPYovWci5Cy1His7ertZ90OknYA9mBt+Yw7
5/OijRyKLaVWnmJNcE0dI0SncXzwPxZvIyV75fYEaNPK6nTSZU1WLS8yThO46wKrDGOHCc38+Zlu
fgdpB0gJxz39voJQ5XmWFifQj/KJ4oq/B44TUMGGEjRX2JMNk4bw+LuFffXYCvr1jvWAJgKhhjpu
eUqVRmidZA6AmOlJW1VBVDRdUphkWzztKrIizAtyUkoq8x5WotLpLFgXNsUXbyfCG/Jd9Ig8TzuU
N4wXVfbVw6KCupcWLuRSZomzbOXGfQbWvPVAFRuk289nwlj+L/cP83BPPpGDi3n19++D/ODffAqK
0o6Ra/SfUgNwQFKD/1EhspsC6VJRA8r7hMSSL1hOf5zEAKrWUUgTONnZPzJeexqSBm/rrSfO4Du5
RDO15EKpHe2ghaqMSasGq7RRFWXOzZ6T2Z4+CRC8F6CdQoasQT3zKzL5ps02sZtqIMcnDUwYYsGJ
dn9/11NNUMlbIh5ko/eLma6hW/EVKIWABg9YqM8aS3lQuDY5wcxDLlFl3ktPIgaDqQ6dJGeH1dJk
sTGd62toFDJ5tn4A6vpbYoIcZh45czMeBZjSunUc/UNkJ4VxEHuqA4MBC41JK9PB+pvRruAh9rvR
xjiFsPFLjewVy6oQV00XaqLRcwVocDaltZig8Z91BUTP7stRlNMh7eND8fulW94NzmF0CCSAMQI2
2D3nkelx3/yPJW+RBT6RfgIc5zV1X90RyKHeMQOav5u/GHsH1/o0ystfRUqgAJonqq4CAN4JtgHm
24hj6Y/I0OesS9YT0dtsqaCbFmwuoLTRgYEzdE/t6hO0XvCIRecVf/AGEjA/HQheTvLK11XgUrAf
q8VKCnvf2OGCCY+q2PRnr6ANEDanpsmPxcN+1I1TWk7LbVKEAK9Knv3iFn6MN6/duIIxYbE9c0PD
YZcM1jwKLb1gG6N2eGFzKLdhrQGkAx21da+ABscOpQbJXOsTdkbxtVzPnnvYko+j802C/bJ1ucMs
fU3tfGxwaNRV4lHIXtYAAroquj65ADddcet5VmZmQBR+G98Kua3a9kDxnnqMzL0K9zlH2C/VRFIL
iNSSeii2Lc8WvMzhONtdJR8TtQlcoYMs6H+HeKvNS9RjNROTttWmxq8G9O23QmzK0fPz/KSsaviW
sio6JcWOF+WFWzJ/c+RKiR+AvIiIyIDLcJ4D7v4Rk58aatjiKi1qEAkS7BW3O6DS1Vb0gEAFV7Lo
BpGGmUxjDCtzoUqthSsDDlPw5+K/1tSXZkRdKVVUG93kJh0by6yReVczqje+qXZw08fLTW9RY81G
4sw4wHUvtEzxf2MK9UZiUW9/O/K5qnj5k+2F1o1QLBnHMNmf0ydz1BHlRh7+M3WiWyLoENXR3Agx
jww97limptM3HCLUJi4JjxP0QSbs2b5eNUfA2cXX0LCYg6jju2u2m2/GR0jcXZr0xC5U2cwbckdR
6BUQPX2HWfPT2S1+TvSulEG1Zg1wXrEtXpM138fwP2eAuIpzff5K2PWdHN80Ru6GcjX3Fn+wfOa4
pRrbeDY7Le0xGNfGsF4ewR+nx/6j7IBjy5j+MXISG/4Lr734/wxZ5fIim7uoDQD3KdfZIzBfrWEz
th4PxpvAkdn0MTVhdoVI/EQ+7xB15zanO9zIi50B67DR4dl4juB9XZcQDzBKKn7UxhDVMPCbm9I1
o8X/BUZmJr/mP6wgOh66rcPRqyGMiHaBKI5XxE0rOKNzB/esrMNWL9r9SCdKCy9N1dlC0huQoSr1
jSseY3c5LcmNCLDBvK7y1eEwS2ZX3H8qM2CIX3dZeL/ujyKRnLgtkVnHNBqjgor4JrthVQyVjsOV
s3dUTsntn7b5qNgfGLFhSYu0jpbuYgnsEpIxRm1lfcuMJ0Oai3efGxHsU9XlaKCiI3bQoVeXT0Uj
UXNayI2AmFnmMtdK/imlQjogXEUeYm0kntopRDhVah/DfhfGxLna2pD+UNvu2cuwOU6M+B2592rT
0riekPE91p/4/2TZGMNQxJQsSIkBKvCKu7hQWXdR3Y4+VIq+18l6ZcMosm0CQT5Bf1snVzqbWx/J
Cch0C/3aXFEd+2qF3B6bGAFI/RMbY6F9puCJpsViwQM2+zEaYv9PV9VFRpp9oOfCgS0PCgs3qT31
ZwmViC5Bw9Y2cNN/oRCVMvm8jJYdZbULpDxGRuG36fTdlyN0a2ppNfx2SMAWnYHFPG6CHoVoCemq
YjiqVtybCSZWoyYS6AhGLS4aDGAbyxYRLsE4rzgiI/lQ0XjzXUugB98tDEFNl28BFJnuLEyb3Mq7
Q3Cs+emUdHS2VNz/vn3sxd2GlQUq+FEWHvmDAczM2z3hJ/T8ZZEcNTc4VN3Tjq57YRJ2jiPiD9F6
vBvVL8nyZWRubxGZkmsGmekFIX9ob7dPbKz7TbdtnVgy/VhJSXIsCsjg8WWeJbxOxYYnBvYKbW0t
bmKFARsazYxexYgE/uyNznAG/PPb5empX/ybfgFnGTiXmhLGvxC6yRpoz+SHUya+RyIib5ECDVuv
j79i2c1L51EZYnbumKspZ9sU/h0BeVBdEC+BfXLzYycCcEQH/GL9TkimH5yrmzBHP9PQTnNuzDst
by+wDFym19TMbCkgCWGRCsmdIFerODWNVg/5D1SoX/l+zJdxtnis82yWJitOX7RyoF7/3+xNdzCI
M/4CE5wApypLe2tYxvA55JQ0fdVz/Yh3nvqqJaPllaodWxBE057M8RbamKPD5P7UOIqnOMm1T5g8
D1hptIUKNT3psUeNlO+Ku99D6pRRvSfmqQGiCHZHAYlfTAuiKs/KFlS7/zzApD4kPycBuoCYQjR4
A06xPLkEqDKbEyZ6/OpM/H+zhsqbtL9Vjx1Ey+KKX5Uq3X0ifowqoBfBtOX6AYr20901mYlKuI2G
zOjoEGDvRyen600/WdvYz921e/p+IwROqKCjVBj3wPBMSog7L1QRuQbuqmgOTZi6bZRVzZhtwhz8
2ANZJPAkARH1HaRb2KWnQXJofoEpKK3VgStN+9nMAzlcH953NFODudJoF4knrhYF3PaNoI4T6vLs
stOZxyTUDo4l/CTep/chMPUHUI3sJDoCQ3YJE+lqiOfqUBvbFghAfF4WG8GtLcPc4NWZMtDerjA3
/U+1WtJV9n2OeCtzn3qa7FmfsCqdUenwVkm7FQYjuXiEZ1IUC8lBOdul+lQkwhYP3vGKk31Q+Gj/
5VYELoppPyramvRhH+Jn5LQsTFCUEUE3VrcUb2xnrYROQ9DWyK2Q/RvY/0fPShiXwsAT+bvQp2YJ
HYgSZGZC6Ip5AuNXJP5yL2lyJkA8dTd/ixUPIwz8L3aqaWHUEz1yH67IvO1qzFRlNPFm5t/wPs1e
iSK6ExdoBAIYBJ/ARdsGfwFe/Jdipv70wyFc1OoR7XxuyF6hBKrZyY2qDJdDJ7Pmw2VEeXOSTyKy
CRvG3I6I2lu+xPFLoXz/IONWpGPn69iT0u1bRCUVncJSRLqpZc6swNeYGcD+ztW5Ex50HkAZ7ZI0
17dqACIZkIIaoBXNEGxEHgyyyXKDiRKy8SeWdINUg8DuUQiCbusB2xNwUJAFR7rtWZZlEu2yRhCb
uWaIQN6aeMTppDUisNYOVL1pt9ok9LQU70RATXcdD4dtT1V94xALjfP4D3H9JX5QckTwyBkkRn3F
aQbortvLg9/+HXrBA4M7GuS642ox3n+NKtNMx43+ob2T3oj3qAJ9ARbi/K3um5u6S+v9Tgp+d0d2
hpGd1YktUnpoZdxKbrjpFfx9DQNt6LW6nykS9rH2/WAnytrroj2d6qznC3lUtDJkEuX4KIDOWePy
Gy/3JtwGEUPxDO0KnqPx2g89Q3VlwOQYvCrEvPWGaQ1i/LSd0hslOrCfiO603efpT5nhALnPyhDR
NgjdoIJBnPOa38Wm09fsfU6zhZNnTolgRjW9lVHi6/vcYFDMaOk2z0LW1ekOYFmlemO6qchezo0g
hCb25viXy1hK3SJ2h7d4AQM4LG0WwT0IEtmWE5o6tZcBKwGsManjxWZXPzeoie1WxW9q3bwB326L
qsfKYvsjRYrtOoE/O9Lnj5+kEb4mzfWwZkkZUd7cProzgZ/fncgDjhVzqOBDVhkqk59XS04O/kq7
5XMn3rpX3/RK09wlZjAxuyBTm2TFL3Fd8iiWzUl0gUNwkOnZPdJI1iweoSRAw77ibO9cCZ4/GR/A
/AraMWe/P/voWAcV3Cn+CMn6QjNZ9zpLuIK78L1N9bLd/C+OBKc5uXxarESeraYNNCA2V7U4EVGL
RdtEhTYHHX9Eav0iDwU6ZDByi7r1Et6D9KU5yyCqIBJ76eJXu35sZ1xQ+Nej2UN7PGy2UfbeOmuR
hcoR/AqQFa3SYakZUiG5bXVD4u4S4vq/9kVwRa5HalQi7VOeHGGMyZh3uD5J44Mmw29OwQLONbCh
KYt7eRynKWxXZWAOSRMfCfPWOg3085MatG0RnIizQwA3JxYPqCC1JYphg86SLT0zkB/GPWYEUuPh
+9xTuRk5qGh7QbwOF/e/DQkXVtLqYUc+o88REgPQKu4kujmOUXdvsbQR06TaAs8DPEgY1zO2kOKv
LYoOMFC277g604S0fg/rlAqmXbpTJqFor/wyFNtL3i6U4+bq0rAC8I6YTxiMX7C3TFvurAIZ8ATW
VzMvvf2W4lRlFBuJkh8fMJouCXr35KT/IIdiKLN5zT1foVLh5NOxRVxnfsNnw81ddQwEXlE8XMKE
olvh9Zcx+VyxI5ptPuDK49VLMh85MdOMqNftDasCHSfdkNd+uCc3U0jmwCmgQhbpDS2Cd2piyf9z
mmrdgQva+x2bA3Xvd49fCUrZxJEfIdA1GgQSE0QXcoITxmZQVV12400r0PyqU3WCXCBDnbXlz+ai
IdK/SSLXQbVRgHFHiri9jF1Ctf1CKD7yR+KRDwetNyfbJi9gfCW7rvQiwhx7z4uuSBc9wcac0wOf
KQtjBY7F/4V3mNbdLi9uRCQz8e/Y8wGczs683mESj2mJo7Ui+O2wg2ZINBRYtwPut3Nef+vrKQA2
ymDDAJ3I9lNt85DhpmX+duz4az8mieVECmy/up+u1xEzyE5+TSjXrXYjA9EaPvDx9HeDErfOzuFw
LNNZz1Q/hTmqJSXj/1pcQfqp/giUN1sVJH5ZDtQyfg9Wu5U3h0/1VlQwOjsA9Av1Pua5I0Q211Y0
IxIRF2KElH647crFa52ja1Dxh3zpaeDxsvTcU563sTzqWz51NMxDBypxdFZgcsYSfu24Sz4uBgFw
v8vgIVt97+efbCUDM1qkuVDSUBa2bpB5URKMJBR67ysH5BMGBCW8upD12tkv0lmNeUxogWLXwcWO
QhG2pFzoeyg88S67Wzh5BB0+YI47UCJo9IIwSuUzLTHX1GLqCQbBqFUc0xMpZgmoAv7ElJ530SMz
d3kMqf4PVTbiS1MVXGR6I/1EcExqJ0g8MzB3RosnRzWSENmaiGlT5pVNjP2FSoeKt0X9PIf+NZoJ
m1G8wcEJQ2I5+HlHwdTi+til0ZfG3aDwpd19i0x60vD3nhKKnMfLG2HuwSlUltIVpszFRBlpSu5L
Oy6dJ28NbPq3QolGmft6+BXTsgkAboducoUqxJhMaFfVxAbVtCGTNnAAZLx4AtFLCe2dHmaUPgvS
oaWuuT/H8RsG00mMV3z1w1G7sSudqauAhG4a1SHBPlnGoYUU7CH+BQ/CKNPpl7kNehsCVRhIH6Mv
NmYWHVqmFCtHxpcnbRyVGwDAu6SmLCB2o09i3BQiLrM6luvCuLlk0cuJef1PZaItE2kdem685AEL
xpcyVfV6iz3pJl3gG6tp3Ba3487s5TQ3TNzInIzDupuzvWp74taMS9T7UULzZkLiHMN40RE4SHuw
hrdpbSmToknvL49ibAvnsO3A+TjxRn6ZZZThYO8D9yFV/KVfDxtKSSKacrS1QQc0v1826Iwcu9o8
sOxNvsq48v8uIZESA8LCwnu2+Q9ZoBfmF5hoFg7fCRrMTDJ7ffoOIGgI2C8qs1/8QAseZ1tMme8I
a9P7EGNj0hajbphLdEZSuy82zvh+STBMsof1wf3nQurKQSBiFuGAFV3Lf/KEzctqTd6MW1ixzDfZ
6q6wleGoJodOGFnkNQKNeGgNAHtF0JjWIPLbHR0ahINB7pO9LPHcWm+mFicxMU/dzYVr6m/yAi2G
FScE3BBIqwZAjmR33rLiY0H5LYgm2j7qURWEBbaZxuIOXkmk+SDbsg+YKqwRcdTOg6H3S1dC3bZs
D7rRyn8jRuzX51LqGXYagTim8izJo8DHD4ZEno9mwxs06itOgy9XdYZYX4s+jUV8GuI6xyUzwT29
LO/e/IR1vjwGpl+6UiCUdfuc1VslH8Zk2S+607BZnLoQib3fQvRemoi84YzlrBhcNH3l9y0nI1jr
PG7/fSOmNNlT8xUd5oSC4sS0amX+SsLp0l+1nAa3yyagRA/UEnPqUjvMAtiz5HRW2uWlDHPTNCPt
F+x26lJ9isq4RFkOPL2q8GF59CwWoHN3tUIjh2/RrH9Wy4zVbx9jnWRs3S7lAZ/MYpT9BokCdBEt
wopv4Zl7FHlsSSHgrj4AHkiFPg5syla/fpGR6v5ry9HrQc8yUtnidEMUfDERTSb5AwdWTNly5l7M
eQJRVFtf6MxmF9D2q+ZpSxQqSfiCeCT4xBgFiReoWKLMH9CnO7qNmd060WXqBFovVnEkltlBjLyb
r2hpYkF1Y9sb1zF1gVkyQQosmRd5hmdT7XpfQZa5Avr+IKHT0hNHZQ0jghctk98l0haI5i6zXUWb
HX0xh/UDtxhB3xEfywDM+IA2uMJvZ5cemdnVSO/WlRUyxX5ks9Ad0U8ZKVK5Q7NNYYMNrjyqL7Fa
gXyXjjt39EDYziZUKyQXqfZ8OyGyIAVIKjWHm8/U03u6o7sv12bmbELLQ/H2qYlfY8i9rWZqeUZS
SaMBc4BRrtxhaL7E8G6MBCpcP+BtEEAoQyxQTwBIi6zf8KgalpdODQZA0lYdbXPFfWeh5xIN+2j7
XBAR9wsO33tRsJY21ksDX0cmvBkUD0uK+/8xhz9oBiexC9J2J8Cofk2mBMfm9vi/RP66/qGpYk/s
5of61v+zhBQknY735x2bt3pwjvB0jv4E7Ai2n+FgvK+VazJjeXhReo30f6NkiNPFd2O81rjF//R7
2bIJDfD8cnTxhoIgPLwTqwphBkqzPPs+W0PK6fpcvhl3/cB1Gvh3ITfueX1K/AejOn6csmBxl/Wf
Fsf69Q1MjvrtvlmhX3G3lh10IMF7OzdbzNQRY3+y5ogon/6M1oxtwZpsT1L/En+VI8Hs37BKZApI
mGqDOl1G+gCegrng/pme9CbrZt5+y++ZN+CQy1fhkq5kqNf+RjhU9s6yGPLoydRLIM7zFssRVnrG
my2xm+N/K9Z1X0dS+8Fg+eVMpKeek74LqWmNpoYQpHHXUcqRoymPNgxHEpMqfn3VBstFrajSIwpW
fd0wkNkqSpxs9T070l5/UxgwTyRMCNzhlHO/elWBwCJmzOjqYJdLjBatvkg0SGZCYWay9NKi49ag
xzWnxGuKpB5yg/YEGFgpC+4rv4H3wLgHMrVsMKCu1KB9jQyytOJ26g0vdGGpTRA+Zc1sl0nEp6h+
K9UjuxX/C1YC8iHi4WddZ9xd8zlM3nyBnCXsULaef6NHru+ClERbVezt1+Gm9aUyM4ouLwUiS/D/
o0a/tMalAGr3SyBQDYfNyWltqiZjVjMSh1nOfFNQdB/cIsGzXtkTyxU9K66pasGcwAmpE/1R3Q1m
jQBqid2z7tmvQwl3DJliYLxjC7+19b//qxeSGD+1UltP1wB9qavp68M70k7pFeMioX50umW2lSBw
BRQAyhLWJm8+OD0j4L4Lb+EL3XcUYN+Ahpr8Xe30Q2MeKHVy66U03iUcXBgQC+CKq8A3t8hhoSot
0JjOQEuG9x7/GekVd3FcVq4AuIHRwl5LHY/ItdNSYogWNlq4lT10mYQ3KPfLFzuRUvuxNrVg4vIg
+0gt6TpABOSL1gTt9BuncD8P5iMMMwjiujdbTpMQYOjpfYRngxTZNDX1/y2UNldBZEIQmr3tTFYN
sDCGcBMulBbmhGOgB3zyamS/otpLlStTiV0fTTK45aFQqkKvNNDxAUCZDLgu0wG0xyLNpKnWh9mv
QHv4aAJOpQLc+Ov19nGo+2aAVA8gaMZaGrm6KvKtX9C72G5hclZVu5NyAM2umLyWEzWp97dBuHBP
4tUboxpLuYwwb9zWs6o/Pe31vMdmSS+BVIK2cXW7cm4htbxsrQn5nPUukT1cnH1zP2vzcB5kM3HR
QBDzWS8395K6JHzedOCRMW+78OFC4BA3TpkDrWlEZcI06HTLusn/uQRP8Ptp4F0LcgOQ8ozJI6Ab
AZhsemmtP7xF//A8P0zTjIMjzlTg/bm3DZcV4yXqfmYpO3VzeVE6q6j5HhdfsuFGQEyxlTDv7Xj0
6nlIql/A6cssnXVST9u5m59f1Jl5czt/QbmEUy/fgYT7x87tfs0SU+mjabQKly/PzE18h3ASPB5N
L+qXtu6GqVa0d7ezJoQ75v3o8Z4LW5UlTMSVViYYG1iuSAcn+PRS3vUjD4Xj0UTs42WTNyYc7Y+1
Qo25x0EYaBf1cdAiJQ0Skt1fakKI3IhQFJTMCCI/4hcD0fG5wNXpFjftm8ZjSoDtC93qEPvyUMXC
XhWFk5Uwapbuhz0Hmj1jpQweqH2wznzd+w0luGVOowsqBjE/SAi3IlMfN25Qed9KoUD79o/rp0ZQ
lFkmdleCwdMivyL1ZivhtXWWpo91oYSdbJYflrsK+zoO95wWGFaMPb4BZAuOi2XG8KCgdHxb5OHt
N6TZXLLCZpTloO89M7kroG09/oaN3sjw/IN8SOU6ZPfn6VsLX0lo8SMCrmnR/6rGmampXygxTz5K
g0qVb55PD7uVpP3XyTAF2N96M4E5ww1w0hvOOd62xAbfgmXbZTyxC1JGyMjHMTFIM2HOprgYx7QN
1zTkeub6p7rOE1wYm+PNjC3/it6bYfk7pyP92PFwrs+JmRNnf/pMJq92oQGJsoFIwEYCAHOeC0hy
maUO6vEBP0qFk6catne61IvwpHiqcPh7horcXIDd3qyBCBhb3Nssd/bQN5ALc9aBNT0kdqXumUau
donPaGG65BqM0ngEXGRJmQ3iKT8KqsB9isSjPaUe4dhPl4964sZRZZL7QecFudaR4jkTlkS6gbvO
/p2S7EvhckHI9BIj2sF78ACyrPwLIhCgzzVdTg5MVL1jLnLFvnrJwZtlAz1d++sCtXgfY+BwJ9IQ
fz1/O1mgP2zS4XXmOjguq9SGoJ9+fV5xkcjTRPDTyFgwgAE/hHS9q+w5miJpIWLzRRM47mX943nd
UiHBR43ASvPCzr+4hWoLKQAdqdgY9lBPJPt37B63PJ7C9w20wlJXc2RC4uShGP5AOTUMAt7GOj6B
NQnwL8YmGdMY0d9g3zlBLm+OW6swi+2+1bbOCi8rlyvBC/2iAjZ3Lnpi7hkp1MUC0/57NLKGcDCC
yPH39uEbb/23Qxak4wLicxSKd3ZehWssLQhZ0UrjHRpKh1P9WYT3nGrIexDbw5SU6i3rm47bp03B
rMddqCvGIS+2sMHDo5sxl5eLnZGMTSm6ElxOqdfKYTPQKaEVAmjFOq9HtGqH91CbRpOtmuVSdVRD
tI0JBgDtRcBOyPMvWcIJuRyjH5CDcFeSkAqonJ0uBjzckzXxDTtSYrGbfgrUJeHavk/kavZ1CdQA
pZ7CWxbrgRBljf6TnyPnaQd+5ALbKDMESfd4b9ZFlthjd0RtF8i44XOWXhl9A4QdmpicYd+R4blx
YwgClDp2zxqmiil4CyjlJy5rQBQGOGvYMSujaM+5a0vXt4n57Vc0YicLkssK99KtKo1klZCw9Hm6
uPok6acpLTaecgUPt1rAMux2/3TTgcIaGWiwbpVGvEl5yHwl1e9zpIKxdGABu8VrVqwX005uIdU9
v49olKUDieKA74Iy2DXrp/+gHTfZ7q6Vmr8uo+PPLH27DEBrkJiVxmtyAZ2qQ2ZcdC1y5X07iYly
XelHs+rXaE7WkrR5tRO5+SEHHv1dlN9NF8uNmTnJBUp3je/xzHN0jlSNWf98uQFb53H0QwE3vc8c
hhSolRDnON+3TZeW5RE9hSfzljmtBaSOzl/Y8DmfAy5HX1+gFjbs+uta8+HsM/DOvLRh8GoOFT++
oI4tPPBH5Lr6zrbY6YjOugdrCQLkjk4AaCGEbBzHXcE7Osy+uV55PTBmuGKvKAhraL5yJySL/47P
PdTYYfhiX9tbiAooHsc07C31xHeYUrZNQXm8t/1nu8Du4DUJa/RJfKYMWR6QHkqRUYagsaBGsh9J
KYWzqstAVTmTE7r0BfjMNA7Npv27EwSLHcIKg2zEr3r5u5yQsI4mc0M6JSoX2ObjeJMMvaBIescu
6HQCTcHG4P+sFpXzrFupPud7+uhcPnqW8cNynbZZ0zfdkw4cOPIf4T8K3T6oSQqBUaCDBaFX/+Bj
f+yb6sEvl+Tdfx+K/VHJhUfXQ5FJtigYAt5l0yTbOMh+IGWGhbgQsnmeZmrkZfddkpFMAvSEMS6X
V1pyZnr81xYExLOHHdaSGiVP89YEcB4audopHHWM94luLeYFKBRhdI4C4mWTz4dRn70673x0KotG
1Pr1h/lAoi64xQygXSrCNsiOMKJrZSdD52SfcVm3CcUDUIcNiq0Qt+zrMYFrtBm0ZBxLFFJ2fbGK
t/V18KXm+04T1FhthQOK6Uj6mgSz+5WWocTuKKwYJpEKkLdup/x6MK7Oz4PAbc2k4KMCMQUL2VIR
BCS5PVTB+poL7dfkfpjoeuovefsWGXmDwjqtDL41+Wg2OZwYz6SdOTu4nN7UcdQhPblN8t0bIrns
/xscieRsGVKPNyfg1oRtye66RGwEIc12h/kPMG8nSC/TKXnrREtu6da7VM8EAHJvjs0mqrGEbfPo
qZg7Eul7SvwcViBU7ghqa6ZMFVpwLse6qiO5Wsw7MEaBqR4UT8fJ5kdXBXDyUu9Okwj01AXtHg8I
CrK826YU1LAFEqNHBWrGxnj9hYBbtHhZeaIFmcOb49fzltR/vVqJSonmr9csOSn5xGfb5cPVAxg2
uaWQjxF+9e61ABQ3I2+/JAIuLwpMviF+unMeKK8moZVNEWvNxU281fffmfBrKzZYOZGytuFosaOh
ibQncTntgd8hOixNEe/6B+oYKLIqIHnP4GUri7mFt2Tkcehetk11886QBqBXcMWxV5bTtaxFUfpf
B/PcP4RDFa+Htqv9E2zcBlNoDjjEZ/oJMQ90FFQ7BgGL2xuYXXVgDUeEf39M+odgdqe08JHYwOo2
Un1KzKhD5VTbLrG847WeKA5/ySGyBnufReoA7VKbljvlcuh7/hizC0GO1UNPdHtdsdJVb8pEFpNe
Qv3mLfR23pXbyNHANYwGHx52CBOQqHzRHjeTQKZthaHFaIJ7WXo9AA21tq4jijX/TgHbT/sE2a8O
6Nt65a1PwP5sQwRAtij8fVXMeH37QCBx0A3cYNLbvsZxCVTSDhCaTWp4fSQlO5isi2GLHeYUs40N
B8nrXRIrjKmrLKsxO3v7xPJ63JVC6WRNDtKbHJTtFPoedwaesfmaALvuEP0ADI5+xiHv1Kb+Jd3n
NKKmOcVaujYgOEUAZa48v45Pb1DasTAyl0kMCUYFTO4TQyKYqGBtEAG7M+EM+OJOax7oYEDixShV
kIG/kSzwgoY6SMyRMnZtTgx5NxhlrcnJOcFiaqRCfIaZpoRrUeXxmZG2FqaLSovcSkccE0WdHxKS
EXKhDoeGIoxYO7qjABlABGjpm9oPmh054ekZGDHuQvXeAzKYGnyQtlfn7cL4VOZb8RA4lvQjNTe3
Ij/eP/xjEo7pJANpvjih0cCGFRoifWreSswhey2HTG/KnLqXnfHjO5FleA0FKeNyijlBzjrh+Oe6
fTI5RKFUAN73qis7M+0Dm4fblQVuz8N9G5nDz6ND/lJsj7Ddd4zuUwZ3nusVcmou6A0kRuBgGrwt
plF8bcw0H5le5ReCOx36dMuk4cuSbcz9nZbzyDq052/rcLxjvaTULpk1eJngbxgNZZL+OAJednn9
b2EODcx2zvhMjpc+LhqTA00jnRC915FxlisQ48RqgHrA5RjzBFrSEkJvIJ+xWp+yRBNSKjZBlG2U
Lk1eQOgygZBlyD+59BjJrrQjIe0Ne0z72exoPz5RPJpAMbB5SMwTdoQnOwo7Ltls5EmOmn8ZFZm2
LG2dTyL2+VWqBaW90yXbTJcNZG07zqE8BfmjTrE+4BDjKybmEg0Uk6eyPIRh4JA350HKXrLI2Y4P
VmvfUxoTHa/Uj3Bhvc5mYoVPVOxYiDbbEFWfHjbw8BnqYmx4N1JxhudJEfuTUpWaft26SLaOcrwC
hFNUfWiLXlNXnmeKwSnqNeYvaICwSFNIjfoZLc+9txcLWhvZWWg0iONQJweKiqfYnx3dH8a64XMb
vJ3lZJiPp57ndM9N5IupNF/p5J0FypgfWS+3qEJsVRpWu0B4bO5+ZzMfq6SN2UdOwQ1RR/ZrO6pM
cDL3nhZbKVcfME7N9lelV1TWXSNBKZvjG2a7RorYr9Q4V1+FOiRPQnOUIj5Y6dcIaGzqLYmu0cvQ
GVxyYHNJtcgIlaqk/fELkRbJO7jqFe+BrGk/c79MQg/saxo85uBZRPs4p2XS103eDMXr4it/bZJ0
bMvg2Brze7HEvU5yoBjFAIN05K8RKNzZxTJbXSW2tQ3sE5CFK9kM55rqiXAajbHacsuQ7GUIAJzB
Rc17o4qQg+VRE33HDE1yzNGqy8LgX1Dq6Ib2SvxH8sikXRHIvJ+QW0kkuZFKktiE2PY5o5z3v/Lh
l/70SZRRQnfAtHaul7oeQZ1LEelXgeh9uEIlyFk94mSFiU779Z1u/yA00MTUb4Xr8r9z2/bOMnQO
TYv3C7iB3LRqjC8PY+dnuc7RsA/xR4nTqOm1wEI7nX8AoPrGdz66RzLpD8mKYlxjiwL54drK7K/B
3pKlm+D+T+mm6gimZRWT4LlGtXmYqaIm4CdHay4Kw+7POa0pywfBQ+4aYb7TPFfGo8TkGrxeimc0
ulOXDr8RyWyBhSg/LfFMiKkGvrUZl/Bxe+NUPxvw4swM50THZtlOvIcpBGvtPYyE+ykmWIBcohLe
P16ogiqXVSb2pHPHsd4b/PGL0jI3+mYP8O3ZfpIHGXQiOQ9c6zVqIvNfjyEus99mEgBFFzU3prji
+6MFviQs3okLCCppv4Jk/VUkHYt61MbfTCfjZDkX8wWeaP9cKzgnZsURWWHu9xQGdBEJB6tqYcsq
dbxeSKzCfmPwA7QfzCH9dkMGg6N9Vj0rvrpkEPKH5Duyi1M8l+zFp2d8IgZ1MVoO4hWvCGMyn3rz
fsgD+kL9YzM8drf1qMQBDnAoD/13DA1zn+lLCYQnrSgrab75uCCq4+i28joS/qNCuJtLmzuisJgu
rCdjPihYnq0ddNn1yRKZf48EaJPkTkWZTVqv3oYUXFWzTuVxaGqkcXhx/setNNqEAQ0YFNiAJZEL
WgcVJth70QjVV99lBgvNQljG3ngxMB1T9qUxvKOC/Vi56qXpzP6J82zSacjuoUVtGaPbK/jeGy0F
S2DZXxtNBy8sM/4G+iZ9NLdNdKymKaGy2qPI/Fdirrp11P7zKECTpHvepp5fmh3DfeKBkaBJzJBF
r3ZAMAEenrJxTlQvB6jKTCSw161St4T/IVzphiDIOtJ5AhkXeqaYUaRtMIQD7i9tJ/RU5qOO1QD2
r4rIupZeQc4w+UG5bvmCT06d2Wq76Jhl3jVJdPjP/Dnfj0nT42mji9ghrqalShfnlrzRaYNHUVnk
S4ak5cX5K2WeZA1vbUCrEy3fx/fUm+G3XKcXpp3jFuNkMXUO8hGNXl/dxxaQQXHYB3BJ7kRfA8NS
ZIYl1IHGStShOWX1Cy6DXhsFbRdePEmNQ+nk56F04YJ9dnGcHO/OIKOud2ZRKaU+e1skNfN0pw2x
JEi++VMM7bMcKbR8G6Xeq8N74Upc2TLc0du3du4vAo9ab9w0M5+I3wFpx6mWM0J2MqJTLzWR7221
lgV5aEXUybo6K7XsIdscS+4Wdix2PXjwrclCN081nqFK8NSrhHSaUwvPe7YFIjWYIjmrORN+aL+K
4ymeNsJrbM1LHd0LdA+FZfnPgF/K20XpecDgw2TTLOD88glCzte/iNuREQUH2XGxjSWvCNmls7hw
3R2/VUBUwRfblGy7l7lqLGZccqK6U4lmFguMS/ra8Y4HZH1J91uBrFy3FLW15wAJ5EEkZevVVUxT
iMsPPFahMgcsy6k9F4A54PA/do2G7YmEEJYM1XpbCM1I0HwSPqvTY31+cLurLhficGsGz3SDXY88
b9e9odtr/H0bVh56XfPtK+TpfqPOW37YnDvrsa0wxrPeSG5PZl6Em4y1lAIATkJS6CoSPmygYgkU
fGfHOfpwktQvWOHS4odCr1va3l7UtoRNMnp9Playsvx/lG/dnF43mmW2dfBR1jOka1jng4wW7inb
JoslQzTfv73mG9mtkdRCAQ0KAXR22bdK/1nW1ErxzOJJATjlgxO5mQPM0gFKYuKeyQd4CS+HMAYo
UVj2gHOpPBY8kNc6667Vgsoo4gywYmOLBry661ez6Tx4Sj9NxLkpzhg/66cu84L73oqIUBEXWyPP
mGnFcvQFmnJb6syev2KUTMz62yQOM2QH3IVXCq4KGeAbLpW+yfCZSII265/KQmJ8Rpr/5tsXILqf
PTr8ea5LYc25A0Mmc1I76yMxTHRO7TMKRfMSfugKwlH5k8I4ubotXFUAAQIgqCMDrmljdq6moTc7
EH7Y8KJAdp3OdqsaUA5FRLTR6AoxVgalaUi2Ho4FHjea+3Knxe4e0oDL0SrMed4yoG9vfrBbsrQ9
0oO0jgiduQGqtRQchLu6o9tnnSqEr2Xzz2afzGJycWL/QjyGd80SQVVl2G0DTq4FNLcWS7uwDEfY
3A92zVwiKMgAsYLLFaDaH2q678/ZChRzgXJbHEcIIj08QL+KaXluISHsetvc8dcZSSnuf0GzBJw3
467/7fx0qu+dhW0yskQJMaLVI9nUHJVIhcSFRx3Hiz9MEyyeZPtTqUiM9N/jvg3QbqQMgOJqn+oI
IAvUhxlSoiQVCHCK9vP3O1IiYNYQ0Mh8xwdFus2h8NY/rFwyL+TWc1+5Ep82D6SKGDFgLsOFmVyk
InRKuiQ8tDimamASKFNCc46Laj7B+AW+qdUQR6yGBDe3q0umIobPm9jtCzhyj93TJKJ7ML/ar8l7
0Ltl5RdlAV0dPyVn5BQgPprII85mtbfjbTM04ajLkBllIi/JNpUXiqxsCO/oUGZU6tAwrKG/06bl
Syq07iaapEnADaRXWWE1lvU63GBQj9N05pFVskmZPBniAeztsxZ9R4a9FxE6FESZb6AIkiU9a2Sz
eB18cA2lMRNYLbWeZqOEdcdFINFqfO1BNDztchVf9wyzpvpuuCPXgVFjPhOkn3eBIXKIInbHLYMh
q83Nsc6GuZ3Vdq9drFwtt7Nl98tidTYlEkkiE99b26z8fIGkV3JQc4LQaXFveIQwf9ZThVYZR9cu
ZFOrv9fno34LtU6QElA8iLq5lyj4vKy164xvUhgv/1Mbdbfx4qWeJk0iFes6W8q8d940GgcvztI1
Nv9lxm7WLcW7Hb7VaDefVrmAnr74PaC6Dmr5Oj9GLlITyjqlES3NI7r2W5xC2x+XNhsOlxf8SJ8V
PpO6loe3yDrIvW/z17Pp/oNl71QtokMWFJY/Y85sdL/CwjH64V1rYmw1jH/2f90fzkxwJKz9HVSg
w3ozrWdVvOaVgqaN2rVTZc+9Raqpn5rcQZiXnwQTWah//+lyu5s+L9DmGHQByiXTPi4kCMbDV9bH
knsZjEOFv19aSN8E50z5l9S1dkj4WoRLbRinSLPezmKuhb7eeg7JPuqZliEYUJEW1EgY2OYXKSRF
Plg71NABLp3Zs7JYvVk/BakFUALO8t+6Mlw5RKQ79vBVHBHIAx1WtJ9eCb9lVD+IWGHtxHImqppk
wG0++lzX0sToF1/O7vI/DfEgyPoV3PPjscZAs+z3nPpPK7dUsxo7zEX6ukYIf2yHSTcqbUA9xm0T
BwGKgdi4gU+IHdR5wguAwPyBCftP/D/llSxqFVKIeovSJixjJ0B2N46S4exno6AxaOE7hiLjRD2K
6Yaa/38V8zUNyL7uaHOLDsdkEJjJsGVnU7sVmU9nxBgshzpM1vqa9zdM97TCPhK2puSP3MrgCLix
CHtLpFC8+2cOSmRQzGFJPYFAkBoT6HmiDmTxSI6nvDoFMU7G5/AODSGYhXTpnaiGT1DPQZs4+bEY
a99PqykrZVXC1z5XRkXdfWX8C3RxhiEGKpb7sa8XW382k+4VDfunRJ12fmgUcBDxHtImV9hyKxo9
2N5T42HizkfoqzAhwDho6syVu85MaxS4R1oexR0sKC7T25AEHBKWNput2B4QGemWB+8ZqK2qP7/A
vfw68r4xnzwA2VW0m+xPYGiFON5Nn8Pu3dV/c2rSQp2pKuJ6Rpkrtt0n4dIuR0z5uifs9zed+QeQ
+qspUPnanXqNd3eiIEtHacf301c9E57UvgYIzOxasMKpjx8JZZaW1kWsjeRbvnPEcaLfWViLdVWB
5KaR9f0PlfLwatBfvN75XmlhfVidR0IKLv02hx8VZvCkQM+BhlXnwTiAvOt7DNhdFqBzWuJm2GMb
0w054WFoTtQUhh33l/9Bao8L2I+FwybRCEY//fXz0n3u3XbGvCIArxybyV+Bsn5QZSUiJlCEH8dZ
Y9pD7xllDL3wtF4fvgI2hAgqIamW8EUx12KR32V96vg4515Bw5+xig2YLn2309iikk5l4jC1QaZB
1xg8e6i91PDqpbt+tVIzoBXhPvmIZJYU/8IFKGIqW1srMfVhwIWh6q5NBNbZ3h5Wy05mnBlOft83
dDwgnMMtzJOwY+toKY9EmqwhGl9W6e0Dc55Vr2j2XeImrGn/T3Ja7Uw1rj79qsCmxHmGO5QISHTH
kl8MsniQ6IVjh65arYYDK6fVeNNNcFRd/JIy+kdF7HXkmUZFcxSI/k163Mdc4qVD0s479HT5Cu4V
RDVsIdqgrOwPmCvfn81f/ZHdF68SAqXIOX/Z3z8LZrXl4q+vlNrkJbWscqW+qQ/cQbixAFowb9Nr
GZU3Bzp9lAWSORsp/JagPgZe8dUD16q20rY2W4ucBz7cBkTrBcr4t5XBMds2iyVAaPt25xwL5EP7
YGoxN/AKymzDH1s5CTk2q+2Qmx3hZBAQGEmh62L7yycbsAq6WtZY2ez6+569GelodBUqyZlJ4g0r
9wNC3c6oWsJYtF8456IM6cTRjfQ5TnLtcC6NJS2HNDn0QBKnnd/cxxy9zEY6a8Hem1SYXxb4MZ5N
GR2QGVlytVk0JIF7CAKoBQQZGldWWAeCTguUamAJf23ORi21BGqZfbepYTk70iyO2wP3E1qNd54l
zLvKlgnjtNT749wWZ/+9C4M/RXyfbdaiJlvtm0mUBd5hpl248n7RhEFy3zhfrNuo8GUmLhda8f0Q
Y8CwxTML9F+Yu6vLK4/oG/QWAVWKlUhw7OASicbQCNhi7ZQDoIdLBe1CazaLzHVss99/uQkzo0CC
WkmSm6gQnkH2KqUbvpvZwCRXeLMdtnZvxrYDNH4wBi3o2evBspOHgP9iovx1pdzRSwjTFRWBqY4N
H4y4qzPrzx2ESCn7lrZeUk5Uz0TJ0hwZCjzvGKleTjcMLbCCLYj9NXOTtw6gcZU90jlxKFSz7qK9
OtKrZraVjElT9kK5w44a0hpMcofLjctyC7MfVc5YBDEltnjzx2UPll+2rTmoIDv4DrvVA7zq5Vz8
30Aay+zxU1TR82uXIWc790XRc/fXEsR7JvnRdobbt3L0WVPOuYfAC/TFNislrQ6UYE8QACa1FQYf
uavxXCjuwKyyvk4D0QuoFzqcfW/LYH4g4PzK2uWL0n+NPRpKzJjDnfSGEoc4UwH2tAOdMthu0dCs
odJGeaPjoZ7czTCNMa4jv0WO8pyO+aP9T+KCXI5Tz63e3yBADLmAGayN/cdan6R1RszTXy0rLhg5
AoXd06P6IWogwbDJJWBvJFb1mjX5EIAEsCyRCw0/tyxpZDV42l+qStIsnNr0+Hc7grJJ1uJ5eI61
0MiSWVNqASMmvBSKNN9uFniNY0kE8tjDTLNFRt67Ff0lsMKKMzBewPJE+/gRgsMIAA4F0x+Xc6ea
QBMjpSDtfUZGW3pM4XW7ZUzfBzKHGiKE9Rm7wyOAsr1RbGtd0FGJpe4bUB3mOAl9YbWxiazM77AE
OKbPPzQgMHRo/cAwe+EwijbpvgVhLQaFw7wUh8gY2hFIuwVuVOaZhm//kOfA3NN/oLGXQtLwkQJ4
KrwM1UDqQSUPoN/bjcBFZ0Y1/FZjKON+TgFM723A0EqUcBqe++Ask97xbCmcpC/o2gQCWzK+l9ab
Ti7tbCjSbmw7jovwwstZzhjbhVOAX/9+sDQ69dlz+PQ0lovu24hiMGp92YLIojXlNbAVw6CzWm83
U43/ClVGJXo5A9LAwI9AzL/va6LlsH9pAY4+Q0SWz+jw5KASDJvnlOBou/7auLBNRLX8jjFHn0VL
uDqqD0l35jFN+PChq1QHtB2F+NRkJwMz4qqQte/gthqVppaST3gTJxYQH6BeUOWsMvK3TCiPmd6K
H92bvszsYpjapnGUJUMqROhqmi8r87u7m6Ei3Aanqv3jSz4AZJ2Us8Jflk5ato5U014zpcs4KXl+
LB4T/1ZNSvnviv3J/93Fi8b75CjA/Ol2BEhVnssxRt/cfYPgeElfvJQhanzGSpw7vh+219n8PLVf
DKRG0dKHY7xTknmZV+CpSfEpGWvaV1vic9EdeeEA6onXe8RJ3wXywUi7r3AF0na2qKvGGtDAH6dg
xfEDY0MT1aerlt8q+mMNmcYLT77nsD131DCZ+4Rqa15A6nWl/fZetx+dlHU7mAq5XTKa1G5VMXI8
F44a1Tknp0uvHwJTx5IbZbV7GaGWhGOxGao5+QP7tzHCAjaI69pRBdb0ZoAc5FcDU7DbCN+G7kSV
mj8b+1d8GdIQJ0ZBlZVBtfF1NylqHaksl+X+yJ+x9ADki1U6ibtoy1YQDiLMYuc2XBlKw0heWYYn
d87n9p6syBDOjrpRJQBq0PkT/isaPE9PCBZPjkzit/L1SU/ZJ6fLTGqXR5Qi+ij8k0tQFIJpSPZd
VyMOLmXQZXpeqqxzen28Hha/slfyFFcNhHUI3XbSuD5k+RFVh/3TpfnvgC4WqmWdYHFKeFCpAyf7
CLcv+DRCurgnY7SzPsA2XsKBaVQgrbCqK2oyiebXd1NpHssmmEzW32016/rRplSbi6tNE5jKdKes
QKeozzm7KD6Vqhgngl6hD+wZQRyiowsYXjYoAOMfxbFFkGdEu19Ju9aI8ZaXZHUPAHPELtwLS1tf
QS3Z0nkeAbVD8QMYDtScpUeZahLyazC8cTYWltfsIT3iCHHXpLm8ePh4tg6yf9YOSFPG0uCxRWda
ve0QHlvD+O0rZaQJcQjnuiXkRTS4NGZURUkv6B0DBGV8O3BCqQc6mKYJLMfEqyEJ6LHT3XCx26r3
njLo+pGz7xZUTCRgrSeLwYbLTOfQgbVZPxJTOQqP5ZrKkztwn2C4g2g3Y3aoHysAfeA7JZz2fv1r
NJwppCY1o8fuwuNBneQ3jOff7vNrMLkU2TywF4mArONzkfDGckDRlL1uKsnSeub95OQwzg6sqQC5
lNRQ11GEXc6jAKLB96abE5tYa+pyRCj4LsGIMViAqPUytCv5uNC+hORC7TkZa9ODjOS0DkD9XysZ
PZGXnhoLQTwYavmVEHxBa8SddczGQDISTsLb2iZzHUfCQBuBf7HcZs0FW8P0+Lt1BetKUmUQIBls
YMRBpKl26OwbSPok/Veb0/3WpCdL0fDMMvyPypX4p9fyp1ytHu5DGkG87TEQnLYGIVDaV0+Pa2sL
K7C86b2HQmphHHRHkiRVdze+lH86cQ0nNUoRZDzu2SDqikS9n/jajqSMq7H9FEmT6f25cKfPebRZ
9WV60q8piS/UROCtPhIdgjhDmB2OSRUATriHPWJpJzBHojCBEb15Rx6R2V143Mkuo93XS7Y399dj
7PJ3vlRw18PzPb/kRJHn8C/N2cv/tvdpMJsMipk9s5hhSl2fuLqtFvc8jR7YW+ePxZ75vMhvcyK8
VB2HEu48nLxIhSg3UasGjrkX/Wmaw6GrfmyRMz972ZO4QNMY4lVdETasARtXFks3/A98vduhQMeP
LqfAW4Bj1yVWMYcQbv8SALKEovpW9/4UMffn+Hl9LCPmszNG9neD04KULWgHrtyDN0xaSbG2kWO+
NTewZjKglaDu2rKIeRXLRJEXawuI5jvBefsX3Sb/TAjxNUDyHgptJxXf9jjT+kidHSGyEdPVfuRR
E1mSsBuzEd+lkZD0PFFzyRqTc/vxJ8mM9G7BwzWmmzNRoRUoX/5WSxapiOY/m+Xeeyd9venMuzN3
DJqWvr37WZuNr4stIjnpqJ5FKl5IwCYW0ro7ZIG+5kQT0FdSevzhXDVpnEuLgM40KH8GD/4nM0dP
/aCjI7Z1LrgGCkzNELeyK6IDpc3y3klawFOfKiLLFHPy3u1L3LDzpQuF3PBScomSfqRRnPU/Szu4
Jon1VfB4vAn3MhFCsVdRS8MctAMRbtzJkmpMxwJ8VqJ3pHN1sLxAJWR1bUOBfx4RCnW2Hmx0kgLX
/ITe8XhoXpU65z4da7l6aDYTB6I5JVYr1UaVJmG8Oc/tzMTQGf67lJLvTrVQJP06G+mxPHldSGPR
yneYtfDxzRv3pXhllV99An8h994Ic6MbRmlalOOo3zvj8utxAarmgohhT0Lc5B9raYDEtegeqHwh
Cxs2czUvOxqFO6hDxECYeSBopSrnloRIY5HJKln1vazYIvlOFFz7P0rCfc99HIHiuZoe3pBEeJDS
3uJUiKufZndxOi3i139L5zNhc0Ro4tgtb5A5t+oewrSo4+4vo+bhhYBnRGFupmgSVyazxye+C8Qt
wz+nSjfpIjpI9JOayR7fgAqG4DjanWDIoalm5jUk6e3CdLX0xuIeDjMRjeTmeiVFrWJXrPaQtRye
JG6K3MDBJM7PwKcourMdhbbjaq61ZziE6VWz+uHd8rM0U7spJjKg/kYn/UkBeP3582R+MBJNqZjV
155sONXWOUhhrPC6EvwfRl8RJIbaXQeT2pMAk3RVK4DW5dphqApnne94d0U6GhzS7rNMN4j3Lo/3
HyYPuTz0r25w0/I2wBx6DT86DMgdYZ3z35WNPsOyKSndKsyf0KIinMpZJCGs6g8w9l6b2iUqys1J
WIJxXg45J+WNCuHIWfI9Fgo21jMUZ55DftQEknwwEsW7yUnM1vK2n/Wprkq2yTr0uFeqhndCMA65
RBi09/Phe2tRp9pbJkK2RXrKcnpPi/aSWVGgCtNXElQtGUtL9bnfPvCkZNYgoIA70FSjaIpUs0zK
ukME9CnDY+Uq4T5RsTm43xFWptCdSncGS9Cv7TATA3kCPMLj+N53swszeMBVqirlGLik6IYjuUo1
pIDQPQi2TFXdGN6M853yWlo5wR7fq41zoWfZPAXaZZRz6DbhxPB4CNqzQD0Gzv1Zn9BqD7PMUBiH
YlWuHcoCyJLFaIennndRPu1N7g8c/Oo4cwVFL6tNjI98XWbZTbE+ziBOq0nwJuYFKYa7vNVcwuzZ
SW0NGD4U5IY6JnD6ceTkN5EKKcTWjh1dBXSa5NqHZzsOW0SKYjGFqOz/oCd6aKqOIcJu8Ja50j5G
ORbKdO+7s3hTLPqweEo6iIr4nVeNIofirVELPmCzzvyFIzBupGErwcIKPsZC+DrbSPQHL7EHEFCc
aQMpQcDvzlwh9OZFmPwKpHskBWQ2lZt1JH9r4XVqxHzaIoYlGsGoJfimqOvYd2YLaCD5PvvjyhcE
wUbodPIrg3E7w6pXlC5xRJmCFl2IAHiRdV/Ir0KENMmpmsHXCuJCuTXDfmhmVadol3K9qFjxtyWj
iA5TIS6hP+hhrTSkoyF+IEbzAEMy/L6Kfnf0ttzRst5r3R9a53cIHmMIWgtqTden0H5jPHIwSwvM
ZtE52SSv9E7SvW6820cY0CpiB3fR/sovAIHvGIyieb7iredaZJJ/SS5dDZHj43EtFR65eBUainC0
/1lsasH6mKusZnV+5EwlYqRt2U2Zo6adL+vCdmh+Y4JzlroCcnux6dUNl/mweYC2/KIJLPU98q7i
37yGIes4ZTUOvBPuPPpXMaZT8OSqHfPXvbn1I/XA2z3l9lFianQocCRYr6NzhntH5lwlMP2NZePw
ElvLrWf/HjwZhOQWYWMdu++ZI49dR/fnlxuqeypdPewMxazvSh2MMon4a819nzRb2ImFMUFlKdCa
jLa5RjkR/sqORmF1YHdUuPYi/YEYdyn6yo2qKV3fLGJ2nXyzCbnPHY9QdqIT6f6v8WFuBuMKFXvd
y3iR3rtL4hM07MXfJws8+gkxjtyKZAfCVs2tMjXa6PPe9wYRTNra1Q6lrXShxrigld1SGnmj6mk4
ogT2kArTPPgE1pu3pSKVcyhYwM0vF1oLmw8Xi6Fjy2eCdWktIhGlJJUb6BHHO8NI6qdVsnrkHvry
+i2WCZiR91q2tzXLYLnA6HSxBaHdbMk1KPMMe696VlEsqL4wexrDE68qKpO5+Qv0rcLQgNrTMmrt
m2Eir0lhqdl3ucW9GAPpp+D1YH6zJF1hltByYdcqjZLg/L9RTcFNIPUSCevCmjNYU+k9E0qrULDh
8ooI2UfSMfh1RfJXO/bf7ei4RnxoNCWbnzODoIUT3xhmKDQ6rS09HZrktZ5AhIH2dRIAo3OW558X
xZUogqT8k9HdYAYdeLBasrG3bB5FzkCrcFyk6kT5/tLtSqd11awkon8sc1dsu5xzD1JXCPTZ3biF
aU4Js1LUQ4JoDHKSfe8gOg7aTRWTwaE+CYpnsR9lS3XOkt+PHnj3W03TVCWE3aPCfEXx1lo+SKwN
NQFZlyjyBqWNK8KFe4B7Mry/o+q+ILej+Z60R7CQCuXAzfv1q5kwAQqudLADChsYy9+KddJRcpMq
ehpw4Y6YbJGgm6SDYZyEykaFPaO+eoQrauIDiUbxP9gLJ9HgKgfdZXpEC7s1kNx6tTVwKIHG5ERB
HjmX+Fjc92hbUr+cyQ5YDLr0Go4wPJoc5druOGrIhgBgBzP7u7WxJrPskhfUD6z3bgpuzEo2xmzU
o/6qe+73MqRxjxsnLtIMp4kCucl6RNu1oqjwAztEfKGma4UBJUzLoqM+u4rqkfmZ4CrLdyfuoqhE
CoXLIY9wmTPevc5WUL++Ws4Wsbas8QRWOX3YTy6bH5k5lm6pSm8u3KT24ocCw4uLLOCfSmwppk6c
Ad09XJHatRrG92SnLXK07jQyFx5+FJjLT3g64bziAlTjhbhhMBJTODhfffEpBA3SMVgxKisqg71F
sgeWNttA+8rgrcwopd8UC7bfZVLIz0J3qtqtXyI0P+wmjYielbva4BPR8cZoZrEOOfHVVGKFKJyc
wr3VcqRXInVQWbxsStIOqNv8BUDli1HAOUJWxqDd5FO+2g0CXnLQuy7e1IvmWgSeWmn79cTfUOfi
SBWaIkw0Letus5nJ+16F3YdUiNHGhRgc50KrLzkZoh8dJIzcrKOOAAp98Hov9AFig8EHOavsFNm/
XT6wRKXF/SlL88K34zqpQqpc9iWT/JBbss7qO7gVaDjXB7zS+tt3jSX71OoIfjc+2YWtqbm8r5ud
2YOUe62HWQXoEq7DHNDilZ1ZMr/UW+pVdZV+qD/s/tzSUUAe7qyqjCWK3i6VK1rcZcRwUoKsG8S6
V253EYrFKoRFMGwn9mm8IJBMv9wUH7kTDW8p3lRcISYArIyWrxAq2Gw04IM9llrlrHvN+5Hzcw1T
YNeoN4RIKc+SzVnTGYTKNjOYxRollJLdZarzlV32Eab99/mFhLHsLYW4e8G2e9eb6LF1zpmZJZ61
jcJE0QBN9BX5JaQQRAt7UXdJHU74+Q5CnlvWoDCEs2D60kXBPQECAAY8+Gew3pjRY64Kl4QMJmKs
XlisWBUznQpnHm68d+VgIa4qLCDOelcqMSKxchqtcj9g0m/YTKbR5pyLAwFQEbGEhpL0RZ2gEkhP
LepsSMAPfSaFudrnJCL4L8RWh4zGCwI3Kv7o0XQMaIqLmmm9/szmfNXGPg2C4CwQF90ZRVGsIV3I
FAWr0rR4put2eaQz2fjg8uaHiBRIsfSTZTdd6So8/4HtyEArvySRAHRE0qGo2dmZ1fldhpNWlnis
0hKb5fOt9GZlF4IE7SUEypSUF6IMLWw8o7qx8OpwpPGv+3V4Zss2sLYlq8CMTMkZlHcknDRbHssb
2W8XQpK3o5XSEA5GtDfkKAf8lLbVv1pGrJrUjrbmDmyS1+v9BkeZ9AGq6FqkKOuodHqQzRlm9W56
F8STgjrk91YUZdauwJ4gA48uIOnPyS2+U8MUNZdkFOQPsKotkRMdwAZ1jqUVyDJ71CEoErB5ruzR
fYIOa/+M+8jPq333sIUSrMbJE+9mXkOCz/mc9KL+n532JWG1DP0oqI+iEQMwY0NuHhGfAwP5GXw2
1vu3cPFn50GDz3rixwcx4IgvhqscFps8xo8EHUbY5OFmKwjy8Le5NIzKj3NVmDbjCWaprdP8i9FQ
2IVG9p3w2QdvgLn0t7QAeoR10t7RQYWK+NZPvIb9u1yPqWQhiWjGSHNetJIZaQCx9Kpy/iJpxMZV
z011oZYx1KTX0TRtqOhvEmhyT0+6Kb/TzEF+/qn7qwkI+fSm3XFCnEQ+w7jvFiULsR9qT/r84YrO
GHccPpRq8O4kLhX/LhOcG886JoZZwGifbDrhqAfSriM3z0LhidUsWrABitNbzW5QBboA+cs0ABcz
+NOB8qHPT7QK0chvUJQP8Niee8AQr/YiBqdL9fGKdtLi6rFj1oLgdn3+p2ytRN0ynMTUdjN2qEG5
2OjP0Izg/gAjuQcz9vPdR+QEGxe+TXmKVSC5ru/OaBZbkmL2HMWEW8fNFVv4UMbwojlld5t8HIhP
RxEdjk/TzHv0unr/ZN8Qj2wJ66EgwAGi2GwMdnMfk7RcddX9IwWG4QxqYYuigt4ja/7vK7L8fOfC
l/7UPK5cgnvXKtGKeDv4BTNVVcQoZwIr2OVo9a38ANn+Vg9xl3LM56w9TdgwJNLBX5ZA3eusilSW
fC/Yy4Sd19IvcBdtikbSvdXZUoqU9PnwKjckHj1XLQbDCBH9AddovrJO56v5lnBIHfO3Angwkxu5
4da53Ji+mgSOqKuVYa09pWVBmsiOgj2jzWDo7h+4EF3wss1Lt0dUqI4YFWVtF7/ome6r67WLxrR7
h5A30MULdR5QF65RApIv70eIU6LbzEIcbiD8+H76MwAztO3bKdPOWsw8xquIG6V6iQ5SQgIw2Dpn
iVUd3uiwWjvVXQ+rG5UUWmangcjODDwTM60REyfIypBo7leVHmfeRwtJMwJ/pb+L6GmIq7SNmkLw
c0W+p0X8aGoViO+bkhq0/R14d9gB4jIRTG2rRDglMeCI+vZ5asnvVjvxlyzLltRkddFgelE2kp9x
iwb5sMLTqNwddil19rnz4EqfpXpHBkXWP/qn4/Qpl609q6yyIofdFKmMPCBz/PBBP0xBvVcLFJi2
HuabKbITuWLvve0ZsoqPL/C1JkWiB9TtM2B4y4swYsSjBZzMqgHlDELN56z9FY20bUIELfG4RquS
JSrofwQjn/lSzFS6cLXWy+CM/EmCcamJXD8LEMu9WYGqpUVjoqS1cBDbevixURy+Boqo4RWb+8fr
DJLwD9I3EP0Bh3IuGqZWecNMGs6QsZBjtg0hCYKFxg7KAc9emMBT6VXyI1As+d0CNoQnsKkAaJ0U
6ig+PANNHq9VMHo/z9ofKwUa+5rS3BMrZ9VdTO/Ckx9drW6HyT4je6L8pjbu4Vcg8WHI45AfVZg3
+mKQZVAv3Yj/011mtIn9m8ttWE2YdcpzoXHwwLFJQBAKCRqJui+hayWs9r9ZHPBNwzhg4gAFiZO8
hzjoYCgK1XIOzWzrmsM7Rs/uy1E+4ZDpDdIAHbS3A7JRuZ3AlxFhKcvW58thLx/mFnEYKGz7D+8e
iUfOV2fUbMolzf7cP316FPRll/8U6u0ilvFM7KuEJp6J3NPOlLEF1xRfflOhbYAmcPVChzODJmB8
+4l1hmYXBTzKw73pKuQQNfBule5U3d5QxZyVI/fnWssIJEYEtT7OTc1Y2IUZuyPAxh8FfG0z5vFO
CQm8i/saJdM2MutmRQM83mClfbHr0OYpFIF9d8pRlFH67K/J6CzmFGimyV5MDLVOpgdYcEXyifBq
E99fDIh7ZAjpfQausy7GnBy/8Y651ax3U2F0MaMV71noOUG8/iOt+cxyGH3iI2lvHDrj4z6qgnXX
ItWhLDnPtiJYDPsZE6fwjJfa41mTN6GnNJqn1BdD5KErY5rXw1y4pNYJQek3cPyYe3vfefh4Qjbv
HELXcKGFQFkU0CHNJht+re1NKhu0rLEP8NSMrqsyIjVQE0lU2Qntb7kvzi1zcUQDBV+sJUDBiMrG
cLsDVwK31DfAvcgWXJhGxoLufBAPZsCUTR8LqCJyEsZmiOZcVC8iW9Z2zOCvu/+9Hf/EwIjqAcgP
AYWs2YKkSoKtvIiWGoL41uMNi3wXcHAuGlqdJBDYDorb9hZDzG+NVJSVd9B8lELPGRjrHXjzzpUH
KhzCh6t8dPcrVa8jdQSviRgPXgIhsNdIPNA1DE9GreNxKImd7D2qw4u58XOcNp47an4XDN1r5yZG
7QmxGAHZNnP2zT981pe1PG2WcAmJyqoMDvcwFpFAS2BV9plzFxpegctKAQjYrBgK0psVXGA62ney
nXTdxuA+ml5qIKJVUKO5X6vYVJypQ6Ulpod8W1M4c2RKjlPQ9/Gejslen4D6lZOMbGlLL4HaWWRA
NiuiJAgV8sxCVjbqRyjLWAP5xf0Aa+3Rk9pgbveECOhiGKO/3kJ3wAftJOgwdWRz1Wd5X+KCJuLM
NoeyOi6UoJ1LS5vxBffsUOilPuKiO91HlXEwh24mnA54Gp/o5yqP0TxxxKgZ+0DvylmMydS8IBJ6
Pze19hoC84m5nRUZGsX1A5xzq/XjtHgMpvszgGhqP5VzpMqL/AXQmr6AV2nChfmzgr2WM/87bhlR
wjru1TNiukeQmSlzXOFg6CF06DCNNtfQH7opbgV9sTI2xLv6vL3bLRITs6KvrKz1emsSTgq3JLJT
vQ5FF/gxOFQ4Gq3Vqe4AqO6PPRXECV/UaeyvFg8go99McXxh9YxkvwxUpJGgPd5NELyR5c7snM78
Inujy96J0umi4UD1TmDflPUh9n+cZV6hW0sw9G856QTCd+sOTcvlTPF58VktH07THS2X8JH+ZXvj
d803n2nIs/EPK+RqQ/iT81VX50StexcGJzUQxc6+MjNF8pXyiUUa+hnMpNrcuCa11j+bOGiqBA6F
TksUhl+3lGM3vznrBO22c9NiFsF4EbkPw1UMf/RtlI+JXvT+A7IfrQgUqRjlfwCIuerROdo4aDUS
6TT/F0iB78O/QEIJM39KRBm3CGq5omsG58OFP7rm1BGe0HBzca+VrovQraagWUktyqB5xhK1R1pa
8l+oLU4RbmvJNJ8NvGqk29AGYy+tRjtd06ZbeBYkJU2bM6bEgjFn8dUKGOdXH2piyZQoGHYdt1YJ
bbCIAlViT5vWr9fHR+K3sKIl0WyUKf8aUPoeEEAhXNpawpbCgMJOJqSqVanXDOP2DnateXi2G9ZO
7HfpnVCJtrkzP4+JNHxdQ6Tab+W7JJNGGMW1ZIJzs610ijLhF8sx4WzoU2iux8SbdNFqflDH57AM
Gutfb4TM3Ge/vvg12Jb9A2VucU1HcOL78G1RVcJvZhRGajHMrrgMbrEWtKFGbVEtLxmN0fqV30xo
qSbTUuRlU/ZD5bkfMB7F4WOqVaQpXlJ6jXgVdAQHDIUBSC+YUNaMt+s/iF/AZGPbWcP8e8+iPr/n
NyZkhTiac5VdiUgg17LTr2MDq/yjdXAezASERsnX0CLvoaHVpvhx7t1Hj+4RENuhRbYiwySRxu8W
ddKUWJV/ouL1h79Yax2PAQOWONzxxU9eOcb8cX8HEbmxrREeYUsWkLIHLMD6g7Q3Z4XIkIE7gsPb
Z0KD2zsO83gEjdVBOpj5ty5j5OmXd3G0nYZq1Aq0jG1RPGMNKbIReGx9MDYz/1eay71BkGrWUwKZ
jpBXWgGVf9mZki/bGoSZExNijj0mJqQ9tqsEuV5fwdyakF5i2E3cQIUWpynF+dEN1FMTYwP6ktNC
Vu5v4zKShuRSspJcejOa816nhtgXj4BlwGfbHviGMV9K5nvbf6KPeJ2blelf4lve7kEpmClL1K6g
z4V4SDCJBnNZq6nL+Eg57Wult/ezmjuqkakAPrwl9glw0+mzfeQtwXgwIxLVOKKqKr66zhbIPxx3
5F8GMOpa22HBzy/pHiP6nniuAk1Juu8qxa9Wce+LExjIZZvt9EdqsqkBmfKRgWZ149NtUb/XLyxA
RKE2Vftt20UpkRpcjtbe9rxtqDyzpMo0ivS1tAJLc6g6C7I7lS25P2DZWRV3q8mNxItQJHKlOE3Q
IaBe2IgKIQuG3vyjPtAjNW3EQXw+/YDG3OEU7wjqEDnUdryemobjVlc9Hi+Bb6ocanq5aD0SLq0T
XthWlXZWySHD0euZ3hqoaI1KfaFkSsJlfpZ1P+Xa1KWxcm3tZ0UkEh1Hw/s+0LuaGiZDxaxO4MfU
nSGp0q/a+hwSENR3XemBq/MebfzHBZxe8fB+7ufxSyfji98alsxlAVgWq4OSLCEsXycg77etIsYP
yGOBFF5OFzeiIyPsxlKe8ymyUrSwg/uq666yOnRwVbHddlboK+foRyp4YGHbfNo7LE70PGcZwdNg
Ifq4F45NTJKk99s/msu0ySi14xSBOHd5R/g4hZrRxuIJ6u6f4RO41OWJFCegd0OUAg5uZ5oXpcT6
k1gODd+avYV4L2yuNgt4zfFMcrU66bPqkpvqNsAuWjvLneXgFGYM2BgTHMTOK/rjzg843hd25WJv
zKb3ZiGKK/6JvVSXN8aUF8cxJeTNEPTD35qm6h/ztgsjIXRkBH1F4l58JrPLRLiW2WgzxZGS3kVG
YiC/GhFaav9t/Oom77ruSclf+FooMtcuhdBft9+Xcnv8MKwcMZiMfs+LWjuYUsaNjOG5nVUnapLR
ZVmjKoTIWVR2nalG1ha/esrUeRg9BrNuVe7dMWwJwoYr8vAotfZF0XZINajszMruiRUPmVteGywT
RSvDhDd/JRGmMPsXxL4ee19TJO4PuiZFFoYxtgScjdyS0iU+lSt0OTidfCS34TjoeYZ/iHYlofF6
dHfU6XoskByYs9U62Ccqc07xAjcgxq8zdqvNpf9TZKxMv1pzQqmMGn90+dtF2Akq2wfgv6/6vz8Q
2Gw/CyQLYEtICeFgHfTqDOjL/Yq9dO2vGLtmYyBzwqdr8SnGDCkcsGfM5Y7y6qT2A2zxD8BqOzwF
G8MHcp+ZOQKbPLEYRg4fkZkmUF1YlHMWQji7CT/mI3xdfiakREFKf+WNT6fqiFzL/iS877AflEye
twitCPDiPttT67sC0FOUM9MXx3UgheS0Hva+3C+acHitPUCSS0dKARgbl++4d7XsAQB0jG4NxBL8
Qc2v+w/7xC1dk+SlI6CiY6zHvHJDXFmTBCF8aGRh1rS/8Mj/vlgXEptNpnx6O+uldqJbG7RKyWUG
23cly65s6X4g5ZhsmXL2auSD6RLZSfvP4Ph56ieSlBNipWU2HoyDS0oPFNtoxsewXSmZCv77FX2w
JTrxa92ut9o0Wh5VPz8/J/gwrMha4YyseGBH/gNa9+AQ7ffBRw/0nFDFJrRL17NDg1pOVCgaY7Cg
ponpX/Tp/Cn9Z2PHMSLK4opiwmFVws7MhWAkpqfYtLgpRRCREBfE0QqlB5PXMTbqThQjOOS05OhU
4GIHwo7W7rUEnwykAyjnUoq2TTOrbxOd8f0QeirLpN8/QrfEeAZyfdoESyTYupA4vuykcfsrIyQ1
Vn+i7ONDU3ktynYKLgstpfFk9is826bYYOGcIprl54IPu5sy9tQyuT3lqCHg+WMgo1VFVr49Fkoh
l3Cm4/MFYNTRvEe1hLtm4w7Z3vq2HpnzK2pUy6b542eU1GjsSk64SlOP5Zt4nLKaePYOz8C7iB4H
siW/fzaeZK5p1bUXuk2G45iaXlWEGlRnetq9WFUdliYIWc7RWMEZaFoJybPtCpaeIiVyQB928QvY
BrhX4YADrx0hs75l06sQu/dVUqi/XrjTA2p35hDEKx3HcZ5Z3oAeHHDcaXmYHxquuk5e0LlZGExZ
0usOA6h51nJ4URoY3jvt2hoSxmZzPM3aHlEvoozG5HISLu9xrJ1uI7QmkENqfjIYv0UdNODff3ZP
X0B54khtdhPBcsCQEUFsUq9PHxUzTJuC/KS5qcvHPNwgW57M/sW0o1xMFxOseLKqlFpEa67Chit2
gamwfCPrQD/yRdUhYnNoGrxV0cjJxUu0KzSOgS61voQqWHk6Xb8/Eo20fEaPqi/ZoI0tFoTbSmBi
4RpQaWuHnY5Mz9c0HmJB7+/tGyhpWduZ/2WJT337CB+C3VW+Tk4IYGjm17jFoiymGdbmK1xr3k6p
qAn+CPRMiyKGU/DBlVwp3rJwnpvyVN1XGtBdXI+tT8765M/KKBvYEGNxOb2W/gYK6vLp9aIX3mj+
BSkNukJNO0wUG0Y3yuMXN2BqykA3Bq0iehUBYa0+NYqi1ov64CSjqx/JtFMW6TjE4GPDJIcQUP81
6ogDUBqAdQXKDbtxU+FmX+UNV6ingDiopqPtRBpLBQTwvbUM1QRjLVbFJhn0Lpikn+mKMUKefoP4
Txa3dqwD6drzK4y82Pu2oUxUc/P8C5UegcSmPqdI34cqKFVf3Rjko3zCvnAlotnENkRyTj6TQFdG
s+cY1bXjCMxFUs4mKAqAOkRdg4gyPyi7ZVx8EIHghRCwJC5BsxmKHiIa7ZWtDAcRNOQog/K4gFYS
jiJdBEUafdws+aw6q5UVQsbPuTn6WNA6BPTY6bzLEwD3qZezUd/mZQCHSfU7qJ34UzrDarB4Wcs7
3fJus/xc+uNMQe3JsVciP+ePgewPl+JabUytCH3ZJP/C6WRLt4suAjIOJU+7m3p9LBk6ax6Dx12X
jgoWGo+MhXdOYt1YrjskAJ0ersfRp/Htr+DeQdYcxh/vap2CBW3ghRNuDmW1rrH4ZHX2jaJsvg7b
6N2dK9kUP0vhXNmx5r3JaO3OtG/90+BMsTuKkFNmgh+Oq5bJPoo75TLNnI6t3nZAOdbjc1qf4buq
qbh0DEQM3k81k6qZ69KER5osAmrbX+YPxhZZbz4FvjG3x+lP8OgAWrdNyNnOOFCDAAtx48VwXucB
OMJ5n9BuEsJIPre7Yt/yaVNiwCLLPrU1oaiNuhql8CXxkGKgZnd6MoPSn1azR/xTg16/LwA7/wSP
7cKTKYoy++UWmRDdjH5PsFKJAyzjfldyOiarf7Knsx+zIBZmStaRhqNp38DPxIIdYE2DLCibVtiE
KzKS7NMcrP7AAOWvqg47HNTlKs8r48ga8nqX62VEUo+zrIxHKy2te6Ta8zDMUzYC2Ac4nIryZSjP
mHLZujH7Am5bs78D/nfnHM7mTBQ+0wDyikXov/4djPlcH+bPF9OoZ21d96xgf+xXr3kEQsyyP5ME
DUAD9sbBhlDefq1tdu25MMHufM8vJCfYYxrEQzImhHkZqsDkteuyx7GXW14eLOSVdw1wpCc0pLqQ
37HQiJaaOnrb4fDMoNCo71AESYPiGhYSTNJ4IqToyO0Xmq92eJ0wt0lmQDPncqX3pPEIapu8MqAL
LeYTTqTQYs+qhWMVNWi4sOPGgnGlqS8Lc27yKhnvAZkXwb19qXeOUHiTNWcHFrAdMg6KG7ZyP0Jy
ZFueiASugxaufTCSoCi8itzUs033s0GOMjCaDc6Lp/g9JTxQBXhRbsl697hggBNSEKXtesQZwhvh
T3LAK8Or21Xo4u+2lTqB/geD0Ep+VGPcm3BRjpceOBRp1pZPVjFKpk4+eQamGkWGOwpDivJKS+15
bL499OhBvLSRIpySEkp5cm6E65W0MuJlinAs04zFBh/szuGiH/x6Y/bmmQc6h9hVZbfwvB9Otucq
P2GPkW/ny+f+A6wegZ7p9A32jsGA+Bzu2lbyb4/0322dSrDUCrBMNWl2afqFYAwj0GlEHXDs0th8
CsVOMmf/dn4BFuwCV4U6YEGJ3tEvci7J0QGQ4hp24Q7t1jetokVZBHk1/Sb7wn6TaecGIR+sSZRw
ouICNjGYy7/SoxgdCcY8QgI6k1ZQykzjNR/PE3Y58l59msCqsnNbQdz22gqQpDABpaAUp4Iqf5St
Yjr3pePI3vqk623DR6Rx6YKWrO0YQWK4EKv3mF+ksW9SsbmYuiVxAxLRb7M1gJeS/cB0Wg92+VFv
gjk/mTJ4687DfZ7XII0TmzxTMp4p7t3Lrsl9cP2Dz+b/MzHsNdKhkEGS8VfQZ2h5G3GKft0ruK6q
xce/S9TwrK2Qa0pxozoDjyvMp01LYVD6KyBOuJlfbL8UNHH6WMW1l/WwbZbgzVOUDcQ7j3/YwQLs
WiMTK6Scp6jfFQ5abU9efIlNi3Uo3I4cpPZ6DhlJe1c5SYdJwA39UFX6L8Q7Bm619b8+yE+17vvI
6hZhTAVtnSEJC+f4SHLuB9Vi+peHZWsTSiO2RJ9IwX5hmaFN5LpqCbYzKFuCwRGDV4hxHw6o06Zx
H+LDyei9sKKsSWlgv3T9mh5h5/n8Ao8SdUIaso3Oga661teunkFpCkyDVnitp19MOIIftZof5uhD
zXrm7Y2He02eqtBGSCrvCht8QVeEH2EURFOnIHnqPK0A0GuWkbod9hn/9GFFv40YhgYoZIvwUxcm
5qqKIDen15fjzYO1YnNuGd4PMPmLd+NZEti5lmbBGxcOtCOzuWyBZqKgWeHU9q2KmnM/gDAVB6fZ
1E491R5ejSjbnVTLKARuYPNb1WdC0wSzcnbWAC2HoL8Y3SNJEKUK7DudaFFz7CvPAJZMU4gKrdhy
CR7fPISBZFz6qTYOATOoMLDaguYCul4hfpR7j6N9PnH3vGFaAi/FzRBN4MqiRSHKrZn+ewO0ATw0
VUWJddRD6Dip8SgSsGShPMY551ymStXdZ5WUsXOa9xSfm6Fvp9Xh5HOFKwfiFZRjnRTmLTecDSe/
/PMhaOJ2Y5y48Lk6wEuEwCg0d2p26Ljwy0D5hd/v8dPZydlQqktj1zoi/wO5mOV1GctRvO0gferO
gW5cK51l8RYatGngHp/GOBCMvFi+oQ8KyP0Hp3U+DiN3rZrSaLf/XhVkp6hsKEZ4/J4ipSN8JcoN
d/WiWa3K+tfNpCZmKmwEXg2y2KbFk2qR4ovegpOdjcZsf5C1lPRzEUY30hd4Gkfg5KJyguQ0TsnV
sE6QRQ79Hu4h75ipO+cgL0MFYitGYYyiRrwD6elVKqqcE6rvaU8rV9hIiVAlcUsdT/HKLVCHy/lE
4ISNmBtN789GRoc3gPU5U3khObh7wUr1scSZT9CnSYRztZacbDTcdL1c5m5Jmf2J6BV32K9pdyyC
9efkGreAzc4aHIpuJLjIFTr1QYRq1Ys7Mw5DgjPoPX3fy1mr4STMaxEtTHG3Qmi+tvip/6d5mV26
3wZfyoeJ9zlcpVnLDhTWWdvlRwxjofBT79w/m1HNCPJxYvFzB2g7YqjON7aEt7gE74jNZdNC9567
XQWZlhf75kUlF+el0ECU2M/3xlyLmQ4OvFOc4ZNoFrSh7Hw5Rg47jBrOoFQC+QUe49RVSshWAaoh
eeCOvaMLmfHb7lCBfeTy/OFkeoT/xvx75YNAC4JIRNcoCBVRMzRwF5Kq9NVhF336WEnEDlgU2Oiz
hi9SxM5VT9I4//ZbB2BK+748Ktb+lB17Au0VuUKn3QvESf/T6t3T4EwgRR2MNOQA0IY+26KSqNom
U7OCBc4EhsWN7cvzZeYRmnCQxvrUb7H1/jkX9dDgTweStwbWkVpzI/xLATzdDzQ8MXDd8ys3kkX8
bkdpac61zqOg3EjMmKmxrSoU3YW6yVaGYf01Kbb0xICo2NQR3f/7TXr1R1tLPmpgTQPIoVb78qhp
k7Cc6Brn0p+d2sFBxZ99nvEbWip5nWm6XVNPCFFhBx4SZsr/zDoc3hVSNvISsOJpIP0DVktcAfW7
S1qCFWPX4DR9Eg8ryqWCDqi/ix6YlHbjOTSl83wIIVe0ehUUUt1EhFwBFHZKKzP+v8OyfCLkh0VU
vnf+qZV5T2W25NhlaBCC6JTa4JBhkO7Jax5MCqEUBOAIFujkAY4zAUmZIhPj/6exKveTZ6p54QBU
SEe4h+zTsyUvUTsvIn085ncTKOOxSnwY06dolOGIsJRXXlGZH5v2F1MuXL28ZSKj7GhRfm2tm1xE
EIFMZC1PskOxQ0iXsdDXJnhoE8BjoQ/Ks+N5psBxsKjyZWxXwS+u6d8HTdq7mij1DS2h0GiTA632
jfrwDdyuKdwEshyJcbPloa2kmguDTtsZIFJ6lULVPaZ0PsUDb5cr0rAHATaLogue2A5wtfuh5481
/MTTgnXyyUqD/zRUXYAfgV6Oe0rtp9Qh9NQpEm6XfOnP57LzHJdD02cCVFXJNYijwbgZQguASTCO
Du/OaTnPBglrHXrpVNjfteeK0zAww/odR72lOXLfnruvhGx+cl3LLukpfaAa+LxKhtQ4j0Pivkhn
8jM+3+20XXiwI5mfRJ9rvb8BinihHP2wO/9Ca2qisrSyAM76gAyPKjojNzY0/j1tv8jU9nuAScvI
FaibhR9YLjMx2nOrcjSCHaXKI/hss10T03un8EQ9kAOmHI5BheWns9oPk3yipzEdz2rQTtpIDU5w
sYQcOxTg7f2EZVQTM/6HL0qQE2LVopy0O4ATRqdL6UUUB/Nu1AQJ/hYGKDxPKcULjam3Fm1DGwco
O5+adcr8L3/qX6xUO4tN7D1a0hgG+HKKit0B+Rz4G9PcYAfZ0dJ56cDYvManONmswYbiQucsXfz2
TqlBKUQ5jnOMAJSfwoXa0YdLvwIoJVUug+UdZJ8oyKcj4Oll77U61bK0CzVzbMoumXGlQ6dJqkiv
YGB0yHpNfrc6vhixvy/XSsPWeZ5SRAq+rv8nzSzz0KJ9qr0PV8tL3HzoZrcUbMRqQ/bIWFFRGYmP
bsxxpW1M1hhyAoSdVjrNVz2ExER50SYUpvBA9H7IWlGNR11R0wf+inCSRKgxXHvexeQUbFX0C1V2
6iaqkWYnN7KyUWaM8OKRSGlMoGX79NAIprg6MMYEP79Q3cL3INNgef1tfM4Iv1d+AqWlK2+Gcp2+
hYIKaw8+jEep5N1BqvM2I/lR/BUOrV/6caVZ76XsUiAuJXRTpx/Bh6coctoOZ152xkbGscdQxAVx
qThRHHBdXXQrdSou8nKQHzZ70TdlY/GVelMt4qzc3dwlbVnKwO+5+qEATsUBJba87AYVDLYZ385h
6kR6Q2fD17QU+jLLwht2HhEPYFfaiznjWUtNO2NxxFvMa0JfjVAakpYvq6JabEnTisTujNqxIIRy
drNT4TA4rA77yOfemKvVc1qh30SnaF4LaX0fQBUGEOch9JpljIQ7zBhliZrDRnzOejXc2fAxZtzd
KRQYe/a64IGF+WibWZoUmjvMNvcqVWhdSoxJwZAbLgJq68L7YbtE7iSPRt5DlA5dxEaOW+SMcnWB
a8/VSpPNlFy+Jqq4mU9DOvKOcmFc1o8ml/Hkx+Mag95VFQ7SCw8pJTLgj9GvIVqu6+Uoa9PXIo+R
Zm9LUsdxTUmh+8Spj44nNo8sydNRX1OcUXez1Y2xCT8ZVXAwZkRT+Fr4VWzS3FHfSSMTAvOKxMBQ
sfA/USLNWL9PC2xDGOGZ9YkK5tqlGIbkEvDTaIBz7Oe7gUaXPPtxB3L1HoTbpOHVYS0Fkg1Ke/SR
eb7z109vNbkud21o91qzyRUnu5jL+LWVjKSXaZasf3Z8tcT2+q3zQ8gJgPUezdFpgdjlqNah6bW2
KojVqze1+FCDCplX3cxXeOUIweJ3tlEGVEWtjUv2n4d7ZFDSvhJr8u7BEuBhV+ri3ePm+LnfXtlu
xpCwJydY6+GLvzJPiR8IPBsF3Jwgqc5AWN1sZIYxJeN5U5Ed4svV2q4Uv9ir5HQ+2NU+pOjczika
kiOEzYO+9TGzhLSSWKFcOYJlEp+dSLc5S3+FcEu73kr30V5Lbauex21LxKRNQGJY1Yi1bG3WaQGW
y2ic4QRzkRBuUK3C9DT5it3ud9WydhunJbm57vXn0+DbCZxVTSEobMnVi1JowDSq0L3WVODOiz76
AbH+IS5UxBD1/RP1bXzMweqAxXwweZKyMHC85aOAIZWDw875bAnvgusPV5RRlL3AyTqse5K1DlBI
LAN7gCIVePv4JhMehMS0dcr/Fh9qLOLvFAM/GKVGZdQRf71SyAu52kiUg+u+dNcrqBkdAnVFtJcK
ERp2Sh3Po6TvjxOfFPVxzPo1n4f2EqmEHVAmZ9+HghidwjxjCHX+l/YHpNmPTsaIvK6f3aWvHmyD
w3CotM2q7pIVP28ESFRHS750u8LMlSbsRa2dOUjJxzQzDcfmKcQb1/mqi8MPZXAAqrLoC3PqNJ0u
62lGvjWudN1U7MexkdTk83rv/qjF49mLNDvh1WK0bsU0I9BpjWB+sczDVm9Zaklnktl9uo1+v+sS
OuJyIltzbQ2aaDk+ZcdtOTGWH/1FSKEuKVNFsVJ3iVBuCtVMGGdP/bNxvkm7/ghK3ksLnuC7kh4S
sGmalBV6wOToQqwwxW3LzGSTKbggYI1sllLTI0Ik6mwPaL0SMjrC6/0ZYGmAfiKRZVGP81HjqYQt
XECn98nqbEXfUGoFBANa1iTlUYlsT7XlzceOkhKWgfAHo6DddQOGh2Z6iMryW/GjWsNHgKIv6LM8
6JQ8lmCuZXUEMKWa+o5Lpexz0m8yP8ozRSdjXOtrxJyhmV5X37+imTxpsN7HW1Bfh5/ABNDMNEyB
VPun8TaOOCzNMKci+2QWNzqk3r49GA49qGyqBwMr+HjpqDuKHMQB3mIzS2xykdnKkzhvcB/w2892
U0ROTzICeMgG5tqWu0EkyaNhFwb1SUA1Fv3H0s6sZZQWzCaegJX+lqW6OGubpGEuGBaPV159XXss
e6dpSqEMsc5zryU0DIebHRhKcvVVD1c6T16Vf/DybYmexaR9HGEjyETROc+vCpb8QWf1ZXYzJ89s
paY+ndVlN9gihJ+dtjcnXD51PzKwX2yxEhqy+ElOWnwhatYLn/vAQM449MOv6lVq1ECTxDsjt1pC
xFrvaDtZAPh2RcfucdBlN/SPfYJ+NFk8JRJqe4DMMmdSJBBoplAQObmelUu/Z0AoPzxKMfu6OY3M
mhgx91M7KZDnHYfJUZSFpbbWeWfUrjywuOjQ4HpZFt3CJSpkeSwKZc6aztJqm5R5r8BYifm8cIGg
YTM2OUrJ8TwJ1sMK/99jWylAiFRz8SWAHQ9H0kz4+KUc+IBdM30UggJFfFwC92oXBxvMLY4nRmTj
axKsazLOkQdp8QVAL1VSp/RTFj7FQq0+QHURqberOxvRA1WPlNsuDoLnOFy7GG4T2W3G5BaaKWZt
pwVEd+pQ+zH39o9RqiHV6MKklkGhmOfvng1/eTMtD4ltIHlC7AZtQ9SIGyCfwi0Lo5Hzlj2Na4z3
uZKwa9iPGJa1yiAaR5kv1nnOlix5kMCvkON6cBuTB7yH8+vN4GA3zHIvx9jfJ2kgM7Mb78lLH5px
OVxJCmFoDMFw+Se5CdFSV3QVL8xNnkYBFkXF9FoasPLFdkpgna9flR3YT5Bh6JUfpbkgrfORb8e7
9kB9uVU93rsj0Lgn6VbHQ4YJwOLLBMGkokY3BYb7lD9jbZLYX5W2EXAPtHJ3hbg8yx2tsuM+b2ug
g4OSQOwxfSPHaAWdKfHYf0jfF7bnezVg24qzFQlyO/0EpsoiU000VxrIIRBA20uwwh9TsL/La0Do
gIDmfdLLIUINpBqOe111mGqo2ZBHpVhT6FgnWoEF62f1kl8q1fifWnmPn8gLYeoUJguOBVGbmQ+K
KYjoLZ2v9P+EfX2j7k/fw7rScPzCZdcRL5EN6yTA4Vf4JUrZY4lIIaTbhrqfZ7fGhe2sN3344qfP
iro3ZRUdcUL2uiSZ3I1cjBOb6goG/rvfFfXKj4qXB2iGJ/ixftDDY4oSf6kuBcwvcz7bkHq/5AUH
JRvK/qp9Z+sBObt+CTnh1/3tnz4HDCpTgTX/sVEk/4nkff2BCqJ8nVIW7HAcSNp7ClJTUrgsizbd
JYTksgJ1nFNnsXrcrA+/IrYYkInefhx3yLNhix5o5QoFVccba76YeOaB+JCYdmdqov/i8hWVuRkn
W4pwJR6QCnLtkFt9l4GEq1BwWp6758gDmxPkXZ4jPvyyYcvOkRSOVeA7H+aeeTeCJFFMvPvjJX7T
zBpvca+PT4TbnjOZmcTIBPIHUhpMgWJShMtVskmEKLC20KN6WdfUJFyf1C7fKF4dDonunbVtO+7l
5sZ7KajbU9wp+bHhiM9O58PK8PlPcW0nceuO57OVgbxV9t7F5xXv7N3ikCo/RoEoTANyZMTqGpJn
XJbcTYLzo8Qf8egu+2/24OV7IlxTSZaK7riegSWv9+GMqsoKXGJQ8ngvRctd9b/dFP1+YmvJwcrr
99sSnReOyYFUcZ4/mNF2bGm9HZsLVynJ+b+TVM85c4EOceSvdcE4ePI3ak5AEUOfc1BozovDaE55
bi54TMWFAwDAaGuNbzaXVtvbx6/FITrRL618yM2vidfPN8gvLL8l3i+0F0BzzLNlXWu4sQUCuoy3
E0F5dAZ6Or5B1VUfRs/byIkCqrYUm6qAxfkU8DMN1W0wI1Rd3KCQOV+CrMW4cTCIBWC/bZ9SmhJD
aJB58hZv7XPKhfQ4kq080qfK7L/++012TYI0ujb6azjZnOvSvt6mFRTZ8hklvgyjHy31iOGhwSE/
3Lvh3t2NLb7Qq3YHPAzMLP0PsCe5gtMJlCgSKVZs8WC5LYBeQ2bG8F2gqxg9T3KUFc+supF7frFj
ktqT3O9s4N5ZXw8GxkV+6iic1hN5eS4RlZPMtcvgVtji3/R/TR0VkqyRs/dAzvKtlDuflaYT0joA
bXBFvcbQ+7Qx/vIqxu0Npr6fBLcjnkGREL8YD9CnbebhHxf+6Jsdf9IIimbCeCnFurSMpGp/hCp+
qY3uIAiEE/bOfg4n+zqMrOr/bBenirvVXxi5DOYGmiaxuXjbwtonNDHSpOxhIlNbNRlAG2QLVSMT
2saGDBRvOjkpAHCeAzU6xR7YQJO5omeA1Ops02qt67/MAdfBxD8Fuifr1aC9NItKbKc+QnrRLfmI
GuvqhNItPkK7D6qkkzY4FiWiWtJfOmiHF2x4p3E15kf1cL8HCFhXswq9gHzeMEiemXKlMpb7rn8s
Z0f9KaQFT56pNi2LA7A2NYdIwUAcZuhdsjckHNm0lx/efF13BIXneja2F11FhXsNYpSoNyjEA7Bv
Bu+0s23VsV+figmP+gCYCZCAkjdVl3R5NQRYJ5ANbOuskpHiYhKGNBKZZ5gj1t/m4vt5zh2I+08w
C+uNG9/SZnVeEE2DyXHVJlsGGqUmzAS6hPDc7ECyn0+AKZNI1OtTZFTS2sntYuBgqkPAP1tJO/TI
TLen8FMltFNHjjsvAPmIH8x7dhFpz2QO0DkLUx5P/j2dVcYB81pa37LZ3C0rn00d2Lcsxy6AtsKk
hYIpXU7lpq1Ny8wEXGfxcz1yzt6hMJFwRCP7WEibBfRLfzsN3rQKDlui3t1KEoe6f4mzvcf5
`protect end_protected
