-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aVzem5StMIw6OzvNkIP3qSZbC2+vwsRnXXwcANfUHiC6XnXrppDVhM/XAg6oJQfo4UNirEjKRm9k
SILv/er6KWv2zsYxYL1/Ib7pLnzyTmcQYnchVDuWXC28z51ms4Zk2/7d38PeNmuntHCaauyReBV6
E/O+F05RjSnTHjuJunxtVNmNDc32OS2OwGbQ89CWQwJC9Rtyt5S3GbV9fCxBDf0rO15/yANHm7KD
uNyojJCV8Nd3fNE5LbSEJAYznckE4ZzhM6PluvSIT5unnCxsQhRBtvl6A9AeCZgplp4mqPR7Zf+N
nAHohY+uW8qfvbNcFfnTfq3pUTaE2BDNXr0irg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
kJZQNMgopNnUes4/xX0xaYnHbr6EDNx0KRnRzk0NAUzABHX19thNQoYm6UdFJTb9Q5yOgW+x4x2M
+OfQ2KeeWatSzOojzg2f5XipGMSsUYz2CdCv9l1AAJcNjsoJmuQWtUZU7dhH3QDif2TwaV9tuJD6
wfWeQAu/IzWlSrEz/e5ci6145AsYZJq/2InndU136yWdWrqXjO04r24C0pcwk+mLlYrkewe16FWj
h2If/rtm6P95ipimxzNbCPGB9K604Ou1AOciYnxUszMDO0yplN5RmpiC583fCyYmQoAFwOuyXwaV
oFMY+NfaH0RwahKN3l9Wgb3cxOxvtqqIFrSwHLu/nGrQ0yBqbE47VpWKFljOfB4cISM13nFNL9Cp
gklFGRzkLkAds8D8POwxfMK3F10Pp1Ri2MSjYNlZy4lTwqeDFKzoyr98ZKnsQx2uZUNjTY3M8ZQ1
FhX959z+fwfW7hY99MYgByyH3PQWIkgPoPEnmVd3TScQaukeUS6VfyJqfbSAohC42nRAH4zTp1VY
Z96nyasqgRX+S897RHyKH23oRT7hqOVpBJWcZx6ZMXndfccNKm0kcMqA1WscfNeAxZw9tWy8Kxbe
qyXjCITWxp/w0WrtRg5HloSePlbvPb5wzWEOnHieSvXSCxOeDsRZDOPD5D0CdCyNF0BxXUFJW0Hr
ojPu8VctTlggmi0ECK7AkcBte+UCI2hm7S7zZLTSwOJzt04W/55r4xx1oRRXuE1LcVxdH2U3b+bd
WDJ0AcIrFPqV2Zd2IjTez5abiiWHalGyvxvkXw/Qj2XAylj5tWHTT+ZRlshNebgyO0PnlJEohEtd
w7pFX9A+p6HOeAQBdZG1WqsI3FmOzEEskTDvOexWhSCeAuqgqZB75Ocsa7EJ1aojFCer7PMSxRPU
YZyW4Kw+Sf5hblV2fDZ/DwIvw1CpHcJqsmENbnAOa25qCU++J2OvwE1zfsQHIJNr/n18IHTeZ53x
CdSw43EQrqaRAiolfZhSy9zkByUKs2pLY9KM22Xh00CnGA7l/nE+0qbUy4FTt/FuJm326LU77SGC
8tZfPJe5aOiyXIcztF4z+Fd+rfxMWV19SCDjv8sUxsot65Rqqh4sJLbeRpOxPd0hSUGvNkTwK2EE
hcOqpP5L3cjZ9SRL8PlQjuL5ieLD2UJtYbb2fQwsw3vwy4yAh4U9gjJAbxRWKjsx9ocncGGKNqhM
0Dw9TkcoVHSS1AimIVMgU+qEADxZnRMH7QwA3XnWqtMJEeGTEu1AJPPM0qFZOnNbtI1cMfMidKkj
f5JUkuxJa00Eju+U5n8IIXqPCNjonBMX0GCpyK30zgxjj+SbHYuuF70QumDsxC9OKtZLSy/5xqSu
JaJZYM2w2Cx5gqUWFhZ7d+uZboub8jXcGlVjn7Fvq11yVVGGoVRYAgPr7k+om3C+rAIXTNGc0xII
jdnWaoraGzcb1FysDGdnlGFik4OAfy/pWNTrXswaV+jYrNOeVsl6pc/tfI74p+yTiD9VDgmsbvfX
ifUJzweA17iApql3HyiQZDycUosVQm6ANUJUGEr8+kdiDtCLaNHSxXdTElbrFGrDgRAK2xIX9j5L
T89T2nCM22I0d/3AP17G3Yi8D1eh5SmucBt8TTJsYARa/iZ3buqPah3+6+oYewX43lfbxEZn80GI
GJ28iwckJKLFHSkjq5KgLUqAg7Jcq29lKk9cg8rlFwbm3XKuEiQt8776nYd5nOPCMoJqArkivRdW
THaZUVZ3xLDMcFWnM/JvwWZHnqKY64puMIFmPElcOf/P0eqAnYaEdsdJMjN/2LaKfS2XAVEHHv+N
naYw+a1vtkRVMa7DGBWKO6QjLqdwvYSYxStOrlZJKL7xrdI2heBws0NWiPsAF5aWZCrjczzocmiI
r0RKzEyDq29Kgd1nSMuHryLiSXp9+U2vuhmQezPZ5KO4/NhCWgTMK2p4/Mz0PYBLM5ppGLPSc0Fg
0+E94ojFDRlaSYQUIciMR8qS0P7Ginr+xY97PAethuLk5qSP2ol5Czg2yvreJXW8nH3pMLmQ0cNF
YKnbtLLdgh2VYFIFkT5vgKD13TAS0KOYrGkTNwmVWCtErGD2cWItFGw4uOCrD7PSRgiESCW8Qpyh
hAvAsE/3wwBaLO4OzKN6xHIxJIkolTMKXWoNRYYg+S3BY0IUZOU2MUR4VD6F/tU9BmTBdzs4cVRD
OwsSCbleUOGOp30cv1m7nhsIyL0jVQQmGRYF82UwO8QmrvYeWGph3M4CSccZi1nhQY9vdKzvigo4
vqnKSBVo3mcIYUBFkd3AVQKdB9fe0gzAyWnOqfZ7BfmIN/Su2YgmHVbuLmnD2hMYgBd9wTRtdibA
0cY/S2xVtRtXz6LBuYfOmriEgdno7jExMgpk8IBpOrqD5thN/v0q2pvdQdfc98QMcR8A+mZWxXBk
LvX3Q0wCXKq4C+D5XwPCJrwpl7hutsm2r++KGwiYcZfIZ83xBOs9WEzhOHKoWkdGe15LvarlRLGb
wdAMDJJrIXSpryqxX0+2d3Aq609R8wntRg7qBDxHuvWQu/kAzmtOUe54pS+1cxkYGLQMLt0MsKY0
9ncFSBaUjD0obgZgA5vWhAPipy9477QcbgO0Hi1uNxNQZmMjVJO+51aOzuWgM7KdbV8evGKEO60S
UhjWojlWZPX/SsJRlPsAX2UUfMosSlJ4PkJh9lHoHnq/CfwKoH3bR2KU7tIpO2Q/nX1Q+cqPOUod
w58wwLfuuR1MfN4Gg9FGQwyrsQzZXzmatn35mBExsq0lM28bdb45hBBitPsO4dqwrVVn0x/uv05G
bWRVhsejculDZSYtJP+p2mqeQCsA15Q6+xo0gZG5hpj5DOwiEm8N9FP/l2/6x8+jKKEvvXh1uKBd
R2/G4Im5Nl41oPnp0g6i3oIqzjPdcXkEDqWc4oZCkN4T0NhYjU7qHuhCd9lcpeM7n/OM98kH0iHd
rWZGMSy6w9WaSESfOFCZn+Zq2CAp9x5y6CJUhG0tYL15upRhwPmimpuQ39XMEQFRywSVGI11i1sf
I0BxxU7hoxbfk8Dxb+2C/GfVxJ+fTBhFm3rkqP2jWJ2Fzx4qPfqJ4VHvcm3ZGkgGwgOuJ9V7LyYh
9FJIgwXrWd8qKgN5DzVJ9izD+fqecmnSoQdgKQoz79sB3jKtxEtp6OaarMg4zclfHx/MB1xQsnlE
AJqzPhQEFVfK3zpaqX7tPcDwmfpSzbtv85vmACFhbfK7hZriWsFJEzyaw15bINvjThA3JeApJGCn
CFRKkHPnzfvtDoZYxOUYa3BoXv4QzmCbLvbaxp/lkPUt9xKYKJm8qntm6NJayS2lVgLEmuvatp+A
Qqp6Sl6G+yurjaXbXPVIx1cYFvyAd0DDU3v3LwRrH4nJnOXjk6coKPYmOMwiwTTF9yqDHTAEWYao
TvSUwP7WH4ZHfwyCzMNgz1ptdGmFPsdKzGOv7HMIQMYuMR/C9qpr1k+GBVmxD3Ba6yl3QijT8BpQ
NOjRgXDZAzNRMU7Aw0mjmzxwNXBWPD+yf2X0G2KJUMJzaWgZy1Qo9WpmG8Gc/4ud4IAJ/b+z3uPB
L0nTD6MY7h7Yb0Y/Y2gmb6XvzQFRPbPsgLXBqMilNi0CBicDMMOa2ju0oGkvQUsaOge4f4L6XQXM
G6G13CL8Aajnl6AuZWqa4zt/DtEVDucHV09JELn3yb57BbxZV/VnoT+G76IUOHUW3Ckj7VpMhug7
t48xjs5robjioWBkrMLzM0lJsIrK39uC2xIkZIfF/MiIwrbyCH0eF7UXlXQ6XX4iEhpfEsnm3fWS
8VeLQdAfPRR7Th6GDNmUw2rCCGAmarjmFK4FBTOE9ZHy88Sh7/19aCGg+edN8QvoNuDyMdFjzyKj
1oE7fYq9xCHExyKYQJS/DRfLu3GEnCJUmWzf6CzUNVWLDWpULk7I9IWk1c6TlZXPh6ebzGEqYLcr
EiRbTFFKKQHqK4/GIa7L4U1Te3RNVVIgEtprquw1S1kEDNjHGbuGLbjCFHfvilwrFKxV38Cbz5A0
gIodBYcwtioC+sCh+9VkE/rVYj+Q/DkflUTfIy35Z2FJC3vWfoGTurFjf6eH37zAO0kVeaz7N5Pk
OGpdhDtC70h2mteaGSCpj5B4TQM+Fvzm3ikYhAIULeAM50YObqmBAhrzuMUG/+F6fILUIL+9fZSz
B1hw9VZPMqxGo67uaGEky4ns/oNzRBqIwgRy9korKqaY3OCZxuadGxsB1ZUP/nMMRB5L1lQ/ltIC
RwvJVfyZxSFKRVE5EnjQ7zHgCf5DY13yXtnQkjTUJVKK/GE6JINbVsYUqQguUEcROITxjkL1nEIB
mQEGY2up+BWD/p68BlP76PpOLYSJX96vp2Ik8p4PPbtaWWEXt7RljO/mFVSXdAE45CZOka0KtcRb
nKpO/jt+S600qkv71eHVkRXxx6y9KWB/flea8eoMwc9wPrH4NB5uWXkvj62eAyS+q2jbkkQkp93m
oJig6VC0fsAntXn2KU2L3ybV6OuLwvU1VujHm+A5GPoMzUn1e60v1x1/Va4hcHOaSgO/MXUpyJAh
LEs7SRAJ4cDbgfoRhY1GR0rPMv6ho7QcfOoY+j1MnophemCtZSGkObn76F9Xvo6qQ+o/3NqjQ+qh
M5OfShhlnaI6OhyIexZnrfBpGqnmtL8HAdY1fylIqN9EVatIb5pd/0zGExDQVs9Y0UlVjlDGSyOR
POjxOnLe40GPw1fzYpYlRRtC0U2GLZQQArcEgKS7//VEq0t1//WWOZ9KQG6hDuttujUDvjCR1KxO
NE9EJ09hykPW46JbKKlGIk+kvn2/wnG0xsVRV9UhFPRlrjH6lNJInjyx5cwN0RBmToJ9W2oODbOE
qC/743Sg/Q8nzz0Ac8OssdfFHPx6XiZEMe4/JJIAZ+lcxRh2GxaeIrB0nLnLUbo6DMoLmcGjcOay
ARGtXWZX9BOSD5PHyB5E/9qbPTnfK/pwf9+NKIEQGyYk7vHnNjTlUHTD8a47BJiZDaW9DJIVX0tk
uLlw3raHHbGJqa41gIllhJDAxcPc4CqKvn58/eeorDNQm8ZMlATiX3xfor4iZfzRMh0uDJptbwpf
rD1jBDJw+/PySO5CL2JcWqbktK31sygpxift2vnR3bLcWv2AzkCTUcxz6cKZfXzdU7kyrQAbIkUn
XdJbhsJUnwWKjRwMGtvW2r76pumzr4EpaQX0AsdWXkSsbPdwbUglM4yV7s9A2aZnaGEQSa/DGwBP
bcyYviDFQ1ft2bRJx+y54t5dOF/owgri5IIYjBhTCMKLguGvsPc4h8iV8gzaY+CD9HKu+ZfC4hw2
Nyx9xGVGjbPlf5Pgr3thyngWctCxSEYCs3T2X5KaNyoTIdAOyDKK0efNL+P65kZ5nA+MBT/YjW2m
9AFzN72Gmtupu/CF8BqdqCwgcrfG/7ao5kUJ3LTA9z88SmvrVVIl8j1H+EPB0R/RwlI1rNLvt2CX
KzNZiUAp2r1Dv0e+am8c0KT2z6m7xO/dOZPPu/IUR+8CUbHRRfYU5ArheaBSt2fozO+8192KglXd
2o/PL6B5mrtVobjVk0rqfisNzP50WaWD4UBhRAjqXPmjoQ7nLcrsP2+QcAYrwis2yvfpKm1Vqqn2
5dtZlge6TcJ/qkOwyU0q5URSGmBcYjF0kYgWb0Hf0liDOGnhax8B/Ac3RsJhgh8DMxYmZ5prK84A
yStRL66kIVGvAmxKAN98ZE+NzXBfH1cAuNPjSW4oIK2duhnilqFesGtCoFrFhoizyptPoDqtUFgC
PEucT0Oy2EPoOvOFx2C7bUSoYnviyEq9WQ6g2u+J7F5Pgq7X53CgcjHa4ihQJl//+xMfdfaBCtaF
EZEGxk9u2YK+nvhaQeRwcBTj8VU2II7Y8GOVMmfbF4rL/zLdI6C5eCguKsOWyY4QtH3XuHpqYOo0
rHa91AKBOeRVvc+G5h/kfRmdhPqAQ5ovmDKXH9K+PoXn9LFC5L6lK7zwVTsob/iY6qsjz/XKFRu/
eXHfUW02iTCyh+/JkRzp5PPWVGUD696gjDJOi2/20WOBI/wX8N+S3FjUUmRcTjjerbPaCUPE1SkK
nJl+JoBPdDpT8k8ZqkiXF37OnSYrFu3T6uQSe9MMmNe70g+GAoNaBrAoRL+e1iAg5jqtbBTA17ED
FpHp3tIo/EM+fxc/6w+ck3UY8x9ciihbOHUU4MD8kbpGGjwHgr8Oz9QCM5muIe1w6tNDtyil4nMZ
8kZRDEi+mCAuABIaei5KKtUrrH84gJREndTo8gPrO392cKq/Lo/uExYUc0jG99p89/Ze42UfJSoH
MJ/2zrFsCQ/a4ye/94ge1tuGdoilPe/0luKauboUqoBNcdWoWxVrEQMj3DWQ5Z62FCh2m9+eVxLz
Q0tWfn5/Gearse6udnm/yS7DTen9uFIwLdpQgS3L6ZztNaN96xElb0WTN8pHGb/U26QwsLDIh8+f
FmrE55SEx6IwfD0dx4moEyrjbmYUrUzZ8JcEST0Bis8qB3PyJiwldbrwvEpooo7bEFSOXeRRfZ8K
VaEySp8Sqwh9YES8Y/ai1KQF73E+cbKluYUIxZP+T6nD3A2qbPpq1VsSgeNGTU2EjyMb/XAMbGhc
5raImSmz/ubFakATBM7eJ4oJnssDUGCFKtSogDzqvk/6+ZJpZOQp1IS2FiKQI/oCvuozOqnx0sqM
0G7bjjLcl5NEai5CBKtWo4oZYnXO2esgWHj/3LWl9lKiCM4Zm2Hs0sVmtInREL4FZdqsGpqA4GyV
BOtCrRKBpr8jf85N96R07YIkrRHpkU2FJZ0LgQFyy6QcdE+PyVIaH2U2DxI7PEnxua10QHLyODYC
zNUJAVXSRYCXIW5WSWJ3gGKXKUgomJFHer/kutvCMc5m1NFYzgeGLdVx8yC/C7AngagXdAtR9jvB
kKt2xVPkfP2734A0bjtGq/OUQbEgKrBOYnbJsPKu2opcdT+WwkhqnSrBxTkhTcPe/AFH3V8u4b7F
5r0b28/RK17Xz457PnKYfFdgfRPGuMiL7PsmVrGG782i9VB0fB/JU+7hvi6HTXpP2pooJTAs+8oF
v+c5Vsj5BNv+7s9FmZQiK+uLe3jEmZ87XISPj7566Xjpn2fADt0Rq3TSCT+71xsx7oJWL5V3dt83
WdABJ5+jX616mNOByyrcWsuylrWHRUyuJYN2F0l0RHe08QhEkZnTPkeVk5fg0k4yQjA2LGlTWejx
dV3KBiFs9wYZfRtffcKLb6qkG2Idr1vFjl97QQmUymXIs5g2ibQmrK9sIejtkJoWwW4GpidHH8BE
QHgmP3oFriuBjDAdt00XlVBJGIjt3c12NjKVcwewImlePhb9tzMWXXdsPtIqu5VspgCfxiTKkd9S
OuQCVh3H2nErvaYdrLXvFrfjoTHj7JIuK2Xy4wZlNb23zwgOv3e4/cID8wFtP1BSZODM2qlnu7zU
A4Gk5RHdTgZikX+70r6JgTUQg2nWIP8SpJ03JJFGJaf9Qmjg4SCwKxtRK4JRWULc/9HlUi9YSq8r
qMhBcKqM5qEomGlOm+f9ei/+Mr/uZLTfgNdUIe7IK3/w2iH47sYW8p0fLrsXbfUZ0vXAN3y6IbSF
omW3WGhQr4qR7JP2HUa+f/tpFqIwZxjqVP3N0jG/eRreHe5ZyQI3p+TpioQNX4IY8OvzQMHgmYS1
ueBvXwq5DpSioKMuBFx3IZHXbBbjSKV8Gy+8TJkklDPEwsdSEC8G59wmyiDmKHz4/nY756QGjvBq
aiGoGZ5s330hQbfMQn2LZaq8Fro3NUqWZL42nA75PdwC3VfhL0RPrHwla3jrQ4K61KrLQkRh3ONw
EqoRU7ptWWp5k6QHgXKw5kzzE2WSTLpURDCqnTHZb1+dUc2uGfXXycJ69tMZ23TrhDTGnjjClrqN
YZjAyRSTYO+FABMy7SLzAWwxz0ymCXqFk9Nl/nosu446VAutd9jsvWuZ2pdinBFjJzwH3BPveTEh
+UPA3g16YafDAqEgV1o9P3wIIXTh6Ym1KVm1moebEFclT6LNQmWm3pnamT9Bv3ZiX9KF51GIZhzC
lK4KIZAy17ahCj/LgVwTFF02bFDvSdiNfbmjSLZh84T4r4lcWqSW5PBo/VtYeocGUT5ra/WOop62
Cb7fTUlFK/QxliUJG2elUhi5tCCRPZvU4juSUJmIPBPgQqxOFoHBBqqu+a12J3d+fQIXrCI+7OSj
/wGU8jTm9MZQp5CF0CElgad8msp9xmjNl9tv6kDs9/IrXuMDaPvOQJIZQce+fXfP1mbj8K7fd6Gv
4DJOa+2/1Q/Ek3cZffrNhmBtgaaa1GbOXETDjL2Z2Von4dhfTPNx56YdVndmJSW/MkDPu0GSOkbI
Zl2abXrwEFp7lfCWhkU5Fpow/Vrq5/YK5bOSchp6JZ/iKttJm3PziJv+u4N28f+4lIahAi1HXVg9
w5v1fMTwriUVdhoOCaSFs6KI8HtzrB6+neL3D/3keyORTc9PiMuVx46qw736nJZ57BlaG1DBIjYT
EQlW4CFvY/K2shBpQKdK23F+ORK2kSSTAnwh2BQoWHHCOmISN03g7FkQ0NskHl/yC2vmO4vaxJ7q
ndfIqtxM/3lYMXpLNMM9YF/tDgEC2SKZIDpew3McUDi6dIHdavZnulDBJ9FTH3k8aVs9BQ3G8kym
DjZW9eLemkBXrzfxD2ulvbn4Mn7dLG5zJGiQGWBJ2NvXfAzji2HgElIMGVRP9hiZmm7aSLvIx5h+
oP3n2SynRAYcQMVvyGuB8DDJHqecQgrYY8R7Ba9QhUkzrGO15T6yLpKj3GjUbLG7LGB/ZTq6RgG1
c9EMLt8xCfhJy2cM7Kbo5dJi5/ShmlP7ns5ZtgUq+e3Prr50FqFKkQKNy81eJmlZuf6q+tWgBCUU
6uAKM5Q/VZVW2BZg1M8/lCq0Mw1tdwDET+3PazV99Sd4RBL3AZxXsc9VGdNFYIXx793lfGjZunjN
QMjSnbRe5l4lMPbsMtXiWYC6hc0ICZKOaErfdEuFJWM49zRIOvzNn1Xo+Ws2aTQsL7uOndBux2F2
vUS656hs6CS7WoZ6LH03MoFGIUP1RhLYJK1OqaJ+KjUvlBIG6iCtvSQxlT74b+j26lnL7TTEvlhS
6cJEV7Q4rGiEcPUFUlGIR0lsdH35zdzSqPAAln8n16N1OFNzRkzhOUJEaJ5qrlnHCWB8F6IZBmDH
PpNfKN3MHeXc3ZXd6RCYiib88L1FPnltfP0n7W2Huv2ZNAO8//JS2nHU060Puy8BwhNwAHHL3Oyr
6il3mNFGJQhd3108NlaMf4pu5YU8zvSMjuYYp7tulNGSl+d1GVK4Pk3c/ugdW98r06wmbPh1uixS
jesmTuj1LkrenhzjlcltM3tzqnfdemo75nbsVdPjLaCz/Wi4YDnOeY24i46YvWp6BjFAffKh7MjY
ewvjtwrLGzBRbCGEnCabeApdEgWoo3GR6qHQEalgsVJHcuNLUfL5JViOvRRXh4xB18muM9O3ivzW
5RNNjMCuAEmpEBFYeN3Obgr4Wu+2u+dN58Nc1j95/7rMxbtWlSIIr82ouAlJrmvQenaU9faX61Oh
DWVnmm6AH3ufirprqIXqhYVRW+dah5zJres3CoiVLDyIiHkLyYMNVz+FR3vHSQuS2vfna8brKYNA
V7vPRxPAVHCdpel9fs9pir7X7YUcKPRZhI8fZFaBQDI5SP4NUe08KTgq6iXPNjxE2Zi+zGwxz65W
nE37VtC1x29I1RdHl3vnoSuVL4tl8RCh6g87MZACJF8Y8XMw/FZMQbxZSfCAXB9GAF/uUAqNXEyY
dAnw6px87eWFBdeck18kSvtUZLg4Z8ASmKYvbB9G7Arl3kB8L96A5tRgcoRXEOwaCSTZIuUpSKnI
KUv11wkOSsgpExzETHBQkYnmO3Gtk2P4hph9YAd87hSIiRLCvMjdeK1aozONAqirINCKss7GMKPN
RLUZzpAQMOjv82/cXc7mvMy94EZVq9ZEmmLWA81RPx2Sp3560q7LHL9lEkYIxlFjnm26UJst2Wdz
K9QsZbfQYz7VQJIkaNYuzmWjhu+gKu7MRVWCyB5KuAkbodIqCKjD/BjXOCq9nNSzs7ARl5sC/ZU9
agqDgmqm+Lj0PZSfvKzZGKu8t9M0NKuKme56ABCTpY9FT2sZI7fLfspZl0dTsAOW09QMaS2bm8oB
uZ2RkBdazeQWfqGUPhtWqZMFFboejGC0i9+cWapfaDqqFmE+W9+5DtmlHarwRJon2bj2R0wPkAho
b5xdJRlXBwrLgDEOX76QkT/Q1762TtY7N5TkOGGNqGiv7/FzAvCkH9n5tt5ALgmKw6TZ2KNkIE1U
ZcnPe0URvBE9gLK3xqqBTyd4TY5kLVLKhUXPke1xdNjgReeXzgLVSv3JrLYpGs+FOrrVYvBlo6A/
6B+kQ2+Ji5pGEJNbtCxdpua2i0l+qNG+tCWrnLRD+3qg7c+Lx5j0P11/iXHAz4bHSrzSjdeYS6bl
c94fcrX13fS5cgjWp0FXaTSXZMKtTpyM/uGh/T3tt/sI/b0CpnDMceObd8PXJ6lAEG1Ypc33fb7q
l1bkIzeaWKEA3XT1hTrdXTAjWwgd8YL+InUV3wwYLsLfeCI3+dODB8u4haQKYA7kO2kc+6pJADbL
5uNp8Ux+biEgJgZwXQvt2zREjjzb6jQ2UgavQQf4XLQu8dlRZjnk3ixd1RkpNvvcpBZJvX0idpAF
y0nc+1GIqKh+RERRjXruyymdOWafv5krzieQUpwoDHDtX9gO+tIAl4v4uJ48yI/hu8ME8XQQIVCs
4yGem0P+PE92r1wQRyo432eEtLL498eYjD+jZYxjUVih7pCSmLCuDIDRFC+mN6lMMtdFn8tugjpS
gI6rRbbFpyhDVbHNXabZcBkTUoM0cGXyNTKEdMQLLXpbg/c08S6BQK8+xF6BzecAgf0lE8eKByS3
FhY3b1MaymqOk3DCv2P421dIEVbXSxi4Tiu6bz2kRfe1P1WOvTKNWlc9VIt0AaxvdvnSYwnv2z2B
K7kVeb0sENwW06mllUpaUoOVZ0WDDTyusoC6e5KJwTYVN+gd5tL6RTcKHcpKocIK+28vaWk5cLpb
K9ZAtAh44Dt25QURy/KQOmmEesdAPt/SmbKT26eI5why9s73ft8d6b9txsZOW5a+UKMAItAIkevW
mZwat0S9GNM3eGPDspnEsxHVBx19TjRQl4P6CO/k4WCBFmcRT9YLppxISWzQ/M/uvdunGJPdNc+w
/cdgvEykXQh1qx9FttdOt92tpfvr645HYHcOjWJF0aF+fdnOX0TWJM/mjPMIfvOFmDaw+NCmrl+w
jyQBmuLXlm1v1bwpjX8NsGQjZCubrrkuFkEQ6DMtSBG/YDHwd3wxL8QIW4cnaiF85pvHp+UfA9je
S3jtzJvV6Fdf/AkOKNzH0JYGBHYKUUFtQLFgwf0CsBzTG9Zb04iyagbbH9wgAMp2Q0QFFkqECYJv
OPl9KXllfBpsOUi+El5fPzWf6wZvdQPW2WbnCc5MkosjDCxcIUMq/HBWPbxzIwuHevWnwl/Jjt/4
cosz2N7ey3hkWRgzhLDu+mz/bw6PyBaFcJHrgjIYxObqVMxRvOenzzZRBQTwrR8Ur3xisrZhab4t
ZY9IzaJ0ys8vPRVDqZVMOvYaBUP+UmLJaTI2Zva7Nq+rlUEIBLZ2xZIvttm6veDBzR4rYDPFhe4v
LQJeRjA7OQftHb3BBzOeui3ZNuR6XrGl8n6KFO7fq7k0capvfBVFUithiGTMhTknEyQrTj6y0l6E
TbVFq/1gVZtANnFXrypBIuOKI8Q/hwGBykMdEcdPfZAeyjOyxcBgkjqr9BIPEVvKt8tesP6lNxOI
1UMYf4rc5EG2f3V2SC2xax6PETUi+BC05BmtnAlPN4Ccy+IUzCrPIgtmLt1yfqXfABGbYyOC/Irl
Ka1NXowBf2FFlh2hSEtxN8WUU3TnhSJFe+TKtBoI1gRZayxr1I0axJfWMTFieKOy/fynDzfBIP6b
d6U2GwH3nAUC7WCDZ+gr+0VUYdgI6lmxdtBBLouD7IWNfc/MKkPo2WWMRkCIylM06p6Mm7t9rl/V
HJHgmPTxb25P+jKSje71+ppmCGFNnUtMSQhUMQeRdeeXjScmz0W/ac9a/9HIJMvtao2HdkUEz1pv
7cLYkDjDgzDJ8E3pvylwqIFsfDTRcUEDmavVXiwVTWzh9cmKRaYKllSvGDJIQP7eSgF1/dFH1SND
2T9T2MGq1VGYQRuRNX+jw3PX0WVRCbyQFUd5BjpxnmlZKSX+nv+F2um2VPELLVzj00L0svm/jX67
t/5VCYYgbxEgSgWH0si8FjZ6TpP+jFsPbxA1NjRHcHdAEBVnzouTTREMLZqmxze7tEb38honjK01
fgIEyD/FI8EvRtbiLxatkV6Akvwr1299z84CYnLTOkEFXkGXy+xspr78v996Ban7CyLZA3k2upjX
7NQVRzzpcPbGfkhGXYu+bvWhl8IDGyJl9+OjmQPYmOyED6hDbe4dP74tS0/kKk6ClwLsEAtVEHPy
ElXAS2FRNxrxViZJUGuml7UajleETtHCvxo24bbXzHvvfXXJsrOsZoa/VDf7dgqxshSu10lTHEMe
nhsBAEfdbR6OGfuxe4dm7vZI70yKBDJoTACCQRn/otrlzt8YtoAU5DZ3Hs/9P6M1hNlxAVmhreGB
T6UTxoFHtuM8Yq9P0YG8K4snjWPy3ZpcZbIA87csthTp4JkdkrUWFeucXzBcNtqtNafqfSOoBLFF
qJWKeKdCkBx+L/GSEqsXSu2p5af7MlOdCm2uHtNZPlrxbNnGmvZlJilOnGbh3Lnd1ccVdrHR/A2X
bE/l4j0JmP9dDaNKw0QI8Q75hQOJ8D/FvxfAkswVCLeSy73Noj/u5t9zsRFiibgaMOetpEW0KYMJ
1pkNn9gYwrDrmnuIORngGsvZwXQ0IbBygN+2cP3wKvn/JkgtTZQSHz7EFNZlyZ1ztaVKmrAmy5J8
/V00479Y7rIr4juXIHOegDR8bLIYoKqEwtezcyVf43/mPK7EBNxcNAsebdIFOJY1PFN4gTd5Qp7m
bBAF39tiUGWFcR4dE6AEhSybBiv89h19stl4oHuih8GHpjGfTlofdQlPijsF+QA1HUiYePKR23DX
y9dbyl2P5Okr4rhNC6Drpn84ol6eZ14EAeD2kVJCU1+HMGl8oy3CjJw9WphQAojX1iUmL2DuQTG7
W+wsWj5GcgtpGq9uMX30zuBtkDp+9MamArLrSs5q7v75WTx1hfdFCNsjn1vwCww319sa6lqC6Aq0
f8YqVoc5EqfqHWjSJzdWJeov3wF9PGdGbIimTpjlO9cbKOfltemaqGa60LYA4Wy7jDAX15xy7ufq
xOWU1YJG/H68JfOrgcWY98Ph6XteBtqhA5+RarUA63fO9+ot4e3KfI4QXGX/SMImkZQPa6xrM2sx
noqILv5NxTvlteN2ikm8a6Iu6PvKUDl29Rn1SYeEf3mNhIk1JAkG9Qvx/36w1SwjcG5MOToBOY3X
OYsOzfyZevu1xIzknKnvQD0wlT9i2SHVKPFrbafxQoLHwCDv6RTpMV7WJT6ue3Y4QjqDZYziajQE
g/K3/At7PV2jbmrK4ywYFq9Ho8Urq/ZgF4fsWXXmondncPVCIf3nIJxlgrCsezYbNCGyp2PT4Qyv
h2wdd9iOHwFBnzYVI9WxfSJzOC4LAEFr7nfF9vTFyIlZUZJ8EoLieh9rKx+wXtfBMNOOmQ/dtyli
ObztKq8IcbNNFkvyGmvP0Ue8QZ7FCdO6XMSVqXaV7v+UF3PyvvzBctfhslErb2Bi0yd2Z3pmyFMW
YW54qbaudxlxZ0lIkjo7SflxKAuUa3+D5QKP+xQJAFWBpKYS0ZxBhjoM1omhMEqW7VI2a3XM5tMz
vHTyjLSPbzg8gD1I22vhmuMkUDdvNhLaFL8j5oFrB1pma5aB+hL3aW/lHFqB+0pW/PMT+nTDZHml
h9+R+x+aW971FaOdK9riSjiLlRLO5jz/qusuCiDPmZiPhrYN+x2MSAhXUv8Vci5y4K3KsASIhiQQ
7L50ht3IH1h2iNngqEJ/+bjiBdGzHEbvF4W6/KC/LUmEWREgWgmB9dyasL7E6Qun7z4XjsmQs5z1
Cc7gZIiaNfGVdNci3xwaDfeYyLu26O6gKROCK900W9CTZ8GFMtmKjvXd784pgqe78IdhIEXP7V1Z
0UN9r8F6GN1RcmLCok7j74U18AVdOJapxrXdhITMJviZ7KU3kj7WI3vBzXd4kpMIYZy2vdOl8aS3
sYRnZlAVnjLdv+6zPLxM9sobGpKdkr56ojaaOVFYEJQoR2ltltVl0MAZmm83B68o3XT5IHfYxOBn
oXidd1omJSp6j9BWvv1wyh099VNo7/r/AfmNU+E1gK/YEFHP+yr7OlfFmGxZGzbLvBhNNR3zjCLB
Ha/iWAzHBNaTv1wBp/4PFlE0ooeKN66FJd7wBYwVUjAprT3rPCaRXu1e8JAJfXUNZgMH7uUJoJH9
sIFBWwFHWvm7pObyQcHS89gvgCkhjLte+B2hw4hjYgKGrn+U2xpxr+8Io2LMQ+ArP1c90r2xL2gv
3d4E5+rrgZjY6IBulEeetEX7DSQeo/Qs2asqucUVNOUQrxlBs4yX6GGztX1yVXXb1kONmsAHperf
7mecyA2O25iX7/6+r6jhgfoyf9phdN1JsXWUZ/qfhF9vMvx7qvdT4FSuVECEm122Zw9021Tk4ZjM
Y8nE/CS4x7FQqCusl2DZKfIuus+Ad0BtBunAkBEbL0oWnCHQ3AXKHtxj8Mzjq5dkdWcU84OV/RuK
srScgFPoXSGxPOMsNFST+FAWfkHdJKOpA6MFLDJPhe4lZF5qemKsRym5t6+57IPKZrcyrjXBFyQg
zkLN9S7rGNWWP12p+DE2ZaOlrdUtkdG1gU79rpSQoSGrcOw6y0vi1+EGzu3Hh3WfDqlHsyaUbE5J
ZOvLGTqELvioyQApGvX8aL0EsddZF2yHk1mgTSZW2dwoXxPJJR95mF16+GIMDbuLhGPKzRznnsMv
zpxvugxO+5jkd1tdB2E4eq52c/LdIbOOUkN6zSI8XCF6CXIZB6IQ3IYa8gXHFBjejG9KGprm58Ay
e4nrL3npk9xBsfDZJPNM5bPPMuYc32mySyqQa1d2XEuWDT7CNDCreylYn7ToXwLL6RsmDrPPfJAc
+K875gXMlCpl+973PKEm2RTzFYMpGSdBJt41Xe0hk7KnCLAE2vb+P4Nt1zm72VAuKSxz+pkeCubX
splEo0lYCV3mX8fyqvykgwd+i7k0MB907oKTqtxWDo5/qgsOvWntf856hG/N8b/S2KAsY0JtUDSj
f4KmHi4+3PwP8Hz/GGloqDMKK17+lCcBhod6LJeicXlZK3OnqDSFXuxQbzSd1xkqSy8yK9UnQNyL
tR+Xh6blc1UpCOW1GSAMqPWFSWAKhBEo+Ec6Ce6UdTGTiWjfOz6ArstSiy1V3otS0MUve+CRj/7G
HH+PUbzpLkVnG8qb8NLn5Mx+KlkSAw9V15qC1BGASPDYrJqLMBPuvoD3lH9x1JBECFhTllolDicA
DmZfferZ1gAyGKslb1ufS3z1hi7ReiSzK96FB0T4syDRWw/EsDdfZLy/H9cnH+crzRkGi6M2XN74
ny/mcnqaJOxdKOvGQeWj7KPjNQ0mkAeeh+7ktIqcqe8xzke6TUTHvNoBa/1r0c6/VBt2IGDZGTxU
Vi8kkqSQyZ+Wrb+VQsw72lzCHzNxfYTdeiY3Cst+OcYmSBDcc0VDYx+y2RY18XHLY7vTpZgVZ9vK
lMDAuoly7eb+MwSLlTmjxBE9oC7vCKOl111uxnOtyrzSygl2i25icC3fHclW0u3BdC4FDfMZv55v
2ZLDQ/D174qyykKJn3o6pPlw3t0ZMiAgK/uvvik6uq0Hr1xcFXURi5j8Dp7nAsoN7ILlUo6C5Lf5
F8Ff8nXAqzd38ScIPQxjs72SZJ2Dd4uXIQ1hvA/fI2dkgglgtzQF/NYiY5PrQbJCHImif2VE+bkv
iobinu217hqhvkG46ti9YN5Sz0qhbFrJhpd0afF4D+Zo5amH1Ig9xSpgEX8reUa0434GCcHuIh/z
ik7Evn2mD0r++IamSndkXySUX87nxLTSY423t+6XODmmXcxBIOR7eE25LJi67ppxg0kUKs0qP8sS
qSlw4IHU8vJQU/h+/NECQ8a8uSThN9G0CStYt0fsCONfi6cG/TO7gR1xzzEd62BT3XO1IZ7wd93h
yCdd4kUz2JDfImazr3HHPZ0u39xIPBJq7t0ZuYvx0rYj3BgU8/itHAkLSzwGMR9hbhpnMRULWp/2
AX/cuG3S7r/w++wvUoZidQAZ8PfJC6gtGQ7DI/q0kgGYk1rKk8tjKYXxoQoaclurfwhdkjcNgTGD
JQJwzQ/X6KFbPZP84DUAWHPxXZ2nF/qltnS7qkdSXQq1kHJrolxCEM/Xzcv9VA0SxFbyrMKch+Jy
WZcIHJpN8Iz2IeLTBBnB2Tf4O6RzlNPekxmPmq5krgp/XVa3F5azsmzFYq8XxYJFdasmn6+oLTme
UDDBJGrei/wK96AY82cPPSJUWj9fznKqT3JqaNIh4Ku1SqDAFb4uqZ8h3Sd6QYyxfwC0l9uF8Ck6
+QCfgWl3JE2Ky6Vjgm8rX7k5mRJ7xfjfk2R7XgJA+pv3g0QKADpaMSl6CqLr3K49cI5GFfJtdeGN
QGbstmr6BNMfWNAAmf5TakepRMKZ3x0VdjR9QBWhjPmGvBucb9U7m3IWhS87tlGxUw1o4Az0tQcc
qvrxq+ZjGQOX8bNBZb23/1i9DC+YTWiZmEppx8jRDyXxbNOh9Ie5VG63S09fZi0r4JRoARuAdn9A
835hh19spqZF55HS4PSpIZLApRT4J31uWWSwQJ2fvEMd5uuWM2OIKhZb3yjrGGAzkS6vtKxZXVHH
sSxJA3PmvQhRDZzJupkEACpJIw4IE6iqayD56Sr0qz5ZUuLtZr+bmBIyuwMlFXPt0xTzxNP3L5Tk
cjcWg/PRpaamWpXi/Dix5+8OXl6Dj5CLYci8pZFpqNqRhZ61c8rm+TxYhrV2KYF/VAkZmj0SceVy
pqhJgixIR6brBYT3BGtULxeiJQBWgn1MpdG64IQhu1tRBfGKacCcBg1fekb708vNaaTjyVjUqMbl
hCsob85ZBCbdq/j163q9Xln3It/j00oQ/z9mmxFlWd2EQGeLWBijb9/HGHARI7rQCZrSd9sRusNS
Fxpw5rINhu8D9K7DN7G7r0e5LobwR+bVGd5Ad7eUKF3G3Ee7iqknI4M6u2dNkoeK4NCFA9+SGv7i
O0m48RY9x2cVoWA48YeQgxOOjDX/Fx1yMdPOg2bxbnumjXq8ni5SGcr7JzbLH1h8VkBuDwC6Z8oX
KOzmgiJVYqOmkLmzQHeSR5XHz9YvylkMWaDX/jSN81Qh8ckkgK8p05y3YM1spnXaPBJjDU1DC9Ob
FDcVRYDXsAbfbzxF46HFmOMWN0M7OITc8RFe85RIoCakmjZYk9G0wxYlbG6SiZ+fGRHa/YOloHsX
EIwq26hYVI52SdpmPzo/2VCNj4BkOs+U3NSPj3cQoAd/yDccE6QwJtkMaeHTIKZVR6iyYqiUcv2b
by432skw2W8iot2FSPGY+TcuelZPIhe2j9Ll3V4ttR8t6AwrrBLlGQSdcFE1EeVinZvXK4ueuAXf
86ra0jST6CvzW+bVRwCjmuZbCPAHKGRl/oeNU/s8LUedS8sB+zh8KLF0n2RTXyHqOSkidz32A7JK
5O5i6QGbtIh96tx7lcVk3ZZa2ifOf4tUnqlTLmWeWaX65fiNDDg6/MCpzt2qhwyryiAHHSzNZqP3
RhiYmKg3Gyb6MOR+N9nBn3evY9dOVyRyPVuscUaoMPcy+kCP2VBUHU8oSiuclgNVuOOZzmyCQ6Lp
gFPPhujvEToVCY6higfohNe8FHgmQg3JOsqx0hUF5Hj2TMDooznQA1pS4UKO3pfXSawpyidfy7T4
/WRmX6hr8hNsljfrmTrzACDUMWXWJcdnyNB2G6tg7ZsEMK/6NauOLC1JMi3IWNBomNIEh9j88Gry
jwJp7K/CzEKTgGiqWGkTWdGYZBnqFo9Rx8JfeNNQRd4bI3tKbITd41a/946d0/62gqFbYWHm6rlw
5bzJuEmGzzXdlpeKa63PdRB7caCVNi5JPVh7juWvVqgR/B3szDO9mwYvovBjk2OU6+9bxqKJrzQU
oInl+JEYreuR2tQ0X5h57H3K95b7JWQzNfGvSOrDlXrei09m/4kBvCD8Xyftm8/PgcjqdzX29oER
Y7yBdhTP47SdDEzHjRgBj3hcbBNxFw7YZkD556aLdU/UR4hUpNbgJfuN5rqfzPQzpxyUIss4oQJa
nSNON2OJe4Stnp7HYNJm09iQwNzC0gxvrPp2csImEGJ7juk6xI9fePFbHPauEHVZszYDKrm8mVLh
UZrq00Eepkk5GzaATKNkJN+Q9i1mKm5LttclISuteu9fZHuAQ7fE32Q1yWRVhYW0PhHB4CiWkE7d
f9C+wVbwB7evC/mb3PYAHpP+Rwv2XOQWON8N+hINpFDTeqow5unpSnzohRxLE2etuteoJtVRwf4K
oNSTmeJ4BrUSHeVTz4HgqRhyxzAk2oLW/jacDW0v+pGaJ2zlUzy0b1csI5TZD69Jh7Mf4BS6jv2y
CMmhEMksSvucNlGk/sD2kFQWzNADesOU83Xohf7rrfgfr9fhDKLCO9lMh7+l1zSfkx26AA6WwPLo
1vm7EBE/x0vDVSbiFvtmoSJImwA34C2uI5fyTiOU4q/Nq/Tg/iXx6xuz1s9LY1X3dWVf+hR6mMUq
nMYhDAVccMApdJ91Pwsy9hGVcUdcaUvSleeYa1AVikFSg+gg1sCrtWx3m9U4lhCGJq/7QKiQoTBg
xdGjl0NmltCm6fvWkZvUX6idn018VXBVcfLcmrbhLYYZ1A4yAIv9pppMeEDDc+gl4UfsiJkJjs5r
lLCghuKdE2r4mve1UaL37eB0H9jMkNmGL6o26iaSLqHZ6rirTzSC9wV5r4pEm+dkhx/F32p8p6pC
HbFDgltZBUaBJhWADxC5QRfzOqX3u/Gm+YVaJmBgLE0/ryW306tyuM2yC+V7VP+RhrWbP0SbZ2eW
T/nUdnXmndU0fbnn+xTNAl/5IlIc+SBf3sAROTfEbpvZM+7U7ab4JhO2tcOUzBaj6LfCGQbK9ir+
pjo0LdQuo7lWxmS5zlWRo9L8rFTgVlIfkz83nwyf8vydPSCTId78Stl5mGvCQ5yKk5uOO8x97ptU
m1Bsrw2HVyopp1W1+QHwqMrFATruHT1rBXBDPf+08B2Zcsq6I17y1tmFak8AUNOxF/g3fDbekJF/
z9guXeM6jMoHi1cZ68edUWGlwrtfOVd/WOgtQvxYcOpIiR48zxutGDL18vyzISuVbuPVkCycsXjk
InLYZQbdyAuBE9O7K3L1/7/vnqRoBx5eWneoszldndKtjg6GSD/XINWxLlprFbueKvZVrGmYhRMk
Apl4F6eKqdSL3tHWhdlM3R2jC+dyI4RRolgXGfL3LJ6+YBcLBLdxb0rCdd8a+z+ZKL1rbVwGSp2C
2IG/w57KKBfRcwxhtCz6GbEa4OM2eT5UhHhDESLqL/ueYa/umEf/HMe5zwUeuO+VekpkPGtT2JXM
5RVmz9YpWJ6sHOjnHOlO80hthWtfTy3I1Mv5rU4+mEbfhYyOnUu+AEoxIxBaKpHspeWINv3t+Ezh
+fcDUR6tr2VYMAzdiVbwBLTj9JcWZv1uu50LgbRASqze5hZENLJ+LT4/eCbu7vu5ZkeuSrxL50/P
3pEqgSOnFTiRMDeBYn21eFotC+ZFzoUPG1xaX50ebUbxl9k0Ev0ePb0HhlOLbRM+vqQE7w3s/YIU
W54lG2WkDqgJF8x0TwKx0q12NWJSv461H/NjHh/uT7D5RX5i6zWYM1j23XFqUwblfgMV2rcHTpxa
TqbMlkYYnvCV4eMYHnTFE1CoKOp7cyyENOXd/FEFw+1ewNwRnMga+Bs2BGCD2Uw2F5mD4o3CKDUF
E5WY7KzKRlAX56+mcFETyGgWWiVMLR7UQd8l3etBQ0cwT1llq4L2gNVZrdMpzZJd5nBxHsoEtIgg
9SKtRLgPMuGq8SyassJ65bRvBRfz/BF4JbvE2WZNPIuWYPNckyhDh8Aj0QBEszL8mD4HpOJdFCS/
PgTqeeH20/eHqSgW2CiNJz+L2jTyQf+/2EHcnRLzhLU5ZmPJZzBVTZTWMRkr9oQyYg4yLY29NJLX
Bjxyw1aA65ooQA+If9syMt9wcVOoK+j2oBFE5gc+YV2Xn0M0X96OWWu2mLRPoKFX0gz9ZHvqUyaN
SIqnYgoXoB8mQovDS3WWrfS+e58y4yaLccjvpbVyvNBEAWwlMEUtMP3Y+ssMZD1RprDthX5l+0cA
ZXDwBRkOYAJ7skhmSBXEtE+suZnhy2E5/EYtgr1mYmOYllA5a8z4YHu0pVoZygGBykgNf8BmI7wZ
EX5OtfRTWgouQ9YRPR2CprdrwJvaEbxiiolSLMDZYV0QmXOKC/BNL89itub/LU2RvgrljRKJCZ3S
kifEt8peiV01xg27q9uT31yKQxBUghGIZ1OpIemoK3tjJeBWjwvyVP+8DCdpMckzg6bF6n2Ybt5+
Tf1nkCJgZKf5NMcb0lAI46G6LasDvUGic43pzv9qywC2v4Yl3txTNqinKU4f/N0fLGr/7Cwf1niU
Tg9Th8GbLBUlz2sOZT4gTUruuctT9A2UO+lG5pe4tAum9oi2iNk9A/x7s8lNpfZKmRaJky+zfNqM
++6dlZfSgSTUWoxV7vatkBfaLmEmGGmcRIZPcpooYdABbqP/N0g2oraGAerR1lFjJAOisDHHUWk1
AYhRmNUJU/Hrrer++85ouWTBeoVu3HxFFv7MZQ+u8wjRnzHIzJRjvjEUCc1fFXuY7E94eHeK+20z
D7humGJfHgFEozh6pf7rOjmZeVRHJO2r/ly4b3pbM2V6Amdp5a8zjMkX/K3dOWUbKIjx2k3b2usG
4ZsZISolUp0onsKH3JxXU+7l4IBCTT+WLWAy261qgl2z/rCpL8h7XPGkslVon/1/OjU/r/cya3EK
hoCnKSD3pD63wP/IL09vzHEjWyDo8aCaPYaIYFn+fjvYJg6kATCSo0SSSDjdcLI15+xAsmtv2r/y
jEv5gI+JXHDCbNTmza+KT5YO1PaBMOQOlwpYHKvCwyvBaycps/N0556lqmNcC/Hq7PmsLpxJwDxD
TclBBiYMie7eBszQKZF50x04xryDFFl6xHHyXz8XwXt7QBqYPw8mKOedYwIULlTE6cAzFOd5oyFK
y+OKGD8senZmyP4wBU67GLT1WJd9n487LyIzcsYJATW8xQnTFvrmTPF0rDlHDhqF1/iswDiMM/YB
yOZwwRWt1nhN22WoYRZQLMpnnQnMIVatDaVpdDMQrw9Y08wRroS+UwscoW8a8994Lpmgz5SOrINc
UpIh30ipJCUXUXx6gFoUmpI0hcy1zXSA2f7/5YzfEBnrOHnZMuDGV45vAl7Xy8z4eo+f4mUSDI24
i9bdZrlq4Mx0LvDkOh+hKQAmX93gPqxHH9hfeU1C4WAklCvCxJf5A5HFQukU9qWgkznhDXdiirY0
7503Zu4NMyN9TZDP2/KUixqFwHAIbGCyIpzpEArZQNRxrDjMxs+niN2/dXNU7INJMhCZUXOczdde
hQXSdC6kSUtjgDjOGGm8OvszW2MeCYLCAsXddcx7ERWrf2fIsHqlug2Si2dSUcz/EbxJVZUAMH1I
hQsb2aPrBiSLcgnZROegVUtN/H7LOSeRYB1grHFHc1XWrXNs6YX2w7PWDtAqaVxnlA5OX/KCSVRW
tUA2x47QYlfHQihnmIkjbFzfP9g4JHZgBI/s1KkCYKwCYkQ7fDJIPbYbScL0CWmanJsvUGEsHJg6
0REtGc+NSmj5UtxCszLPIBrsSSbEieKHjjmt7fjJs2S1hKvlxdrtPr9noC6hOFVOoTKVsXGszdav
HncAOfvY+yqkYLpIMf953QuxCADQxHGyl3k2FLZIknl5YTNMxCe1fJ618+3fxf1vDrwPgLWZGqgj
NtnafnHV/H2h6/PsbcdsK/iECABP/X8v87nFwzyWtPvKFJvw1FPWCF/ldMmTjLu5QkKJPfi3xG/A
oipyS0VX7P4kqu9IfIWIl7riLTq3xgN/kLhSAZkQICOt29ghSMTYH+7U5WjTz9BtjbLIqCLeVC53
4rQDdVvouIOZony1G14hFmoIIvk+Te6CJEamqXIPV5JYqvD7pCY6cfvRlHNX/oSTPEjN+Zv6k93p
LhIMw+0ZtG02ONkPsPAO21LJ1Xe9g8PpY2tEQW2e5jXOC4Al/Hmj3l2yEfbdu4WrmU17GtUFBCkv
iKcPy9JxMFefoxWrdUEv2nW/wDJsoBMK4zBoRY+Z2b7nlVC6mKQUseyFMgJ9YKMxmyW3lr6YP7A2
ZrDbmTTLFGme8BtCRR6hBHVpdL6r5q4vdmsex4hDvkDr9xEjUVjH7KzLbLdO7708cL9grCfRx5JF
vjrfF37RLz6A1V8q1Kqc/CVECye0VVFSum+zq37/2+0/tK7aaLRzx3E0Jmhlu7uptg/7PyM29zv9
ELlqpkwJVYlRCE9pwJvDWj8m+5mycrWptl4jH8lgtmEXrrgwmIgw7+FAVYCUnIWb0e41lTbZAhaz
2RridGPTrEb1dxCeesP48RHXMduHMZvyP/jIxPY0ZaYG4KXQO/vVFsWU013Jn3nSHiHlig6aSHmw
PD3VszyygfkRAgqN4jSg3MpmeR8MT4+YsYsqlEjbKO1ddj0vlU2jubVnD68rIak9doEJ60Q8kD53
pk+F2JblZqv5dDTPedEhTWI1u2qdebBmS+woqe7nB1VXSqHt9mgtsKcyjRSoXr2IWdIzoSl87CbD
DQIJHqwwskOJuegR8yftaEig+W7nIJXyR7KUNPQnjfrtkHevY46nFkIs+x5CBSs4i1JMGRwzlWbG
+dKFqZ55M1k3CumzYZT/k4O9wnEEOqwYB9FMYgGh5NoHtJG0qBrOrBOC5BUpyHGBWXM6jEL8uMhl
5SS7yqTE59IpVjGha5Jl1zz0+enPvsCkj35y2UuC6fq/KU3NnIspajZJBoGYZKinV01BqM4xeQGX
IswLU+cS4D9BEXMX9doZPlPLBXYB5UFQ8PwIOtnm95YGo313Pmd4qwj6VPVEAzj+GspQqfYwS1V9
RQqrGhXCo66LDlZ2X7v31nrwfxh3Vi64eGptpV/eBRMVbsWTyQZz4VSjRDrlWvc1dgfkIFDE2Nyr
wSKt1CDL5uyBLstQKt4eQ7YQ5mvbcBpRlfxbcKbVmNJTPR8GLJmou+FZo5QqFKLtFLfPm8oDUq4c
n2KSINlIN1V/WwDUkqpoFkxkJTzVq2wKmk0q5wqfXJrm77MiZ8/T1HZ2DHR9K1EFXP4IK8IQjbFw
KgzbQgzV+PW0eUIsu4LJWLIuFvuVLcZV9K1sbF4zKPFo164bUzQT3kJaHIOkQDsZqaJgHX63G3Du
nYMTsvEDSSoHt01f49o4Kc1M0bz1Bt+oRvelN4FIvoYlXZ8f43Cw3OFsEOIWuQXc7Q8eoYrmYZeD
afrsmVRF91mMIF9/Z1dWYRFldGAugbKrQ0Cv5ZDYtJvT3napVGLTvg7uMZK6CSspnfiCvHZARFQO
4yl0XJ48b9+ReaxPHSUT5CcSicwHPSQkkUuU0dU/D9NQUWcNHDcsYd1tM0QfisOj4q72NfIa0Q/X
jfUho713UlFFQQ55ZrEkxaN2+EMyNJDqWHodSucFz+5H4Y1/AhO0N4IitNa+BZl8wJTT4iajol5L
JVUeLTxLOhafBAh95qJ1n7/Ie4kUe2gsWgKTUloxd5+Pl6D9+8CGATqmKWG8CpqxebpAhpkjLTYi
B+U2bPpB8QjCPGpL/HbWUnGZUixsvSQu2VXxEP4jJbf/z1S3KtSysUqaV3ci5EBJTcJ3tilhLvI0
E9drW77w3mU4TOoItfEAq3s2NmKPvZplSjVzBYlXhWZAW7VMPJ2yHMcaSMb65ZhWK/tZUx83Xl2q
5y6rN/qbU+WqRIXRew9Q5A4JUcmL0O0BgcLhZF4zTaI1WDth1B8WtbvV7pSztzvtJYEABmk54ibs
/vhlgPZPmyBU9bxG/eQkVL/ua6FmONw50kA39li3qh5DnIacV0uPRXnnFq4GdlZQFDEZsnaXEcZG
XKoxl+qzRpS+WDqDMYkul0EUJVMZsV6GkLDaUOBkdi5NrQ7dnMUqNaP3juFAhALFHRD7OW7xDOjW
gPVLNj+XpmEgl/VjWdXLu7lepbLC4rv12dRH8svTGuzZrK5uBwOiRSZ8aKKCbRsjcvSLfzANF6j0
5Trkti9a6Zyw8B8RaZUkt5nvO0S9cfpiMLAgvreAJeXM1hIhAHdrp711/Jbzq38I0ZC+cg+5raNT
ygndFHYqh4L9BNja2ZxhcRNFeARyTwIdT8r9IlZ2FZ1CitKAbAOylne9khePWKget2vGBQIbiymF
p7nw84rJkfS09LFMER1mclrMoVCVhMfWtXuwXKMIJ65UxUKyK8hTb0taK0AewwUwrbjx/bKezSfI
YLtDERZTRC0cqpqeONbKMH1iluLPyrw2RQdsN/8O3VA2hAnAGiDqM1L4Zwu3fSQi500L+GsRtwGW
OZE23y5OSLtZdmOCn2sObfd4/fs7SPorcaos9HLRe/QwcCNbOjaMH/1LcQfThvkAgR6U9SPKaCHG
7N0l8TmjLxITI+XKE/Eb9RTLwQis6YJJrKIxZJ7hklCXc4IbwbJ/svV23FvrIVDawM/PMw0RaiOV
SEfW2Kzh+XuPRUt9cwIUpowxNGjW6MV6F2uEPok60J+vxy6fOTmXCXAAoaavC8aD7D64z5dS6Q6L
e/HdLnPc0xpy8QRiolxBKmorkpYWYebeCdQrc2S7s8AkUIv6fCIzLeEGjkqv8C10P6eC1531vn85
2qDiGMv0Tz3xoookJibpAHYVA83c7Qrjb/bIZqzt7BQkEqp2CGJoDYjosRp/xN/cG35RYVY0Rwex
/9jEYkW+r84IuVTA9IKwr+zeKMmQ4oq8ZnvekZ+9fJo3jgOiMt9nnjdxiKd3QOxuiTvTX2KEK+wP
QwhG8+Bj7e8ATgvM0ugfSuGXUDWTyM2157L4p18md4zX/XAw3tRLnanhNUHzQiHUPd+bH4/7VlGz
mgqkJx1f1rVKpyQDyiB7J0dqbSKzRjrteWgVkGj2xqrH9GcG5A2hWtfRhJD+WDRXysQ02Zics1TQ
+C8gRXla6jx78IZ+/+HarJMG5RK6ljHBd8AclV2a//ROdq6zqUwIYtQIq3M1IROpOXbHTi3Wtwgb
iny4m5aGY/bI7hipAkK6TPkmM+mTa3fC6HRzTgIu4LNv4Ky0SLocxWtFcT7AhqdstOyfMrSBVNB6
3UDcsQfdeZyNHg6/lYpHu4c2zzT3BESu7qoCdvCO2gyVZC5CcgtJQKtwaipWFYpvMLdtuHzTcIId
vQmLDxAuFshhHukdRcfcwUHCuYSI0wcpRJMx/nOHYtla0k9x4YDzRVpraxhW4XWuM/ixCBZy9jsV
LcTYVdV1qVTHjoU4AKae5IHMj39Gm9Yf8c986Ejm4hM21bt+38xFRvGzqJhBFomb7YWRKUfuAzsj
wSJTfGUelQmE91ka3RF/Xo3JwBXJh95S/9bAjkRusV4tFaWSlviGFkA3ypIM9ly5BtvvW5o7GU43
5Z6UyzCeBuhhQu+w7ETpxNex1VS8Ic9QPeUxvvLM6EU1UtDiuqptENNTb2hOfq+3rjYAsQMZjV9P
lwElMEvbFxNoamfCiuLTmuVdN8FsByLovErx69xELI0seQhitcA7feTKeEBN6cYVfZeORcGay9xD
ec1VLW5QmfE3K3nO3gD//Yp35+lj+bsmKRQ+7PXLNqLblUWr0Dw4t77gFaIfIp28NYGacEtXYjff
E+InEJXxNItZmKBYLZ9uqyNjboWNMA0U/k6rIEfFt41iQ9cRXYNYU39OroeuX5DWpsIpZH0bjOuR
zUTQRj2dbymPfxusDthy1ffDhRCmnr8UPz2EDeb6eHGSoCCZq8jAT3N0WCTLjKj/PKUvE9W4ugCW
JVXSZY7t9DaUbv3pTX5uz2Reg6txZWABFnr/9QXnG2XBf8AMJw+QzjFDVx1V0BMLdC3nq2XJeTSY
OaTItU/VMfscFNW+yM48YY7SpfzBkbgQIkl6pw5VPpwpSicaA80r5yR+k6klmL7L+5RkGvy0PJY7
Z/x2NHqEllT1DyJulG/Nk7U8iUBTxKXz8KOM/UamwVd9K83OZoP3ZC9FSDl089TvazZouCPBOjLM
BjfU5isJe7UMkokw4DL7q35yRdqGLrXmUShchCEHcszhTZBTG4YhwMA4bTYY/YyfeLsR11utjS7q
uhnKwCCiVsdP/DIWrRATuZoGUGdUuKt53ObseBnkTA1+bfVcHnpluDE3FuFoSvtvOqb1U9l1Y9jP
koKCHo8OmwsA1fwcDvopztw3IkLg4j/gangnN0YyWQnu1ua09w6jkDGci+2JLeMwfLkSrcwu1d+o
ABJg/jZ+3eajRW5Mgu1Zzhl53NKT49ygg5O8F/KMJeSjy6FKeP3fcTnAOnQox9MR6yzjf5uXb48Y
8crpnZ5X/MWg9YigSjQPS3JzudMJYU/Q2XVPILJR2uqNLsZeCc6AQ+DPdGiN8FSIUHqNixzBvPR+
MHkzH2y2lFBczdj3lTS/3Pv8gwqqThab8HfoWFlVCsyNIO5KmuJ2iaWK5bVGl91e9BWgscorMrVF
SIELWK8dvkvW0Rcn3z3xYVd9V2Bv+D412zPVTSSkmElydX3MvdSktExqerzCjF6noEuaFs9xv8Qz
5mdxbLTNy/Be3gNCxNTGqy500d+sQ5NRKDlqkjB3vUck3YGVkAWEEcOxKbztAxcfipJ9fTZPcVgC
DyFhDfjJdx3UsrZgvWPIpDCVwKbgXJ5fGC/zVbMECFUzYSxuTMRsIEvttfh/r/hNIki0IZlQSi2t
vIWyVjKRDE7bjsczfGd3b7noCAwYAMF1HmmushUCSFFSBZPAvwZKQkFMSWBfF1Zg3HRuwawsY9xw
BIpIGHrAyp+eflSafmwunrWvLcygUhntPqcbOnRyZJQIJ+RG0tkFp1BDPS5huX4XRnXSfXbk1CyH
5xkBPfEhbHZcOTrOwVI+x2tUwvRWyUwrJBp8N6AKp+3VZTf7hw53eGBdNZJw7jJnysrHpVlI4aP8
Tl7uxSlbW1XDeApHXWgpc4oRPO+Yj+HgdH9h6X5Q2WjVwuT1YYe+3SDAW5kEmUwfr1u7R/v0tr+D
G7NLOlF8TGlZXMsAbE3HAH2j2UIBSV+S4QibiRLZ+F8o84Rc/IQ8/7jczc99wKWpJJmy7aM2Vfhz
AH0Emw6iZ0XkuMgGJqEDl9ws6+vZDXBvqag9sytemkDxsRKEO3JtpXQFNqPeAlJzVuYvMFwp21Pa
KwTFR1snC8IUL77lRDkH0eySs06F7QawoQeB3BKd3Zvjn172Li3Yjz4k0Z3KCe1GyHqgBmMfkm+W
gc5i3Eugm8L0Pm1+oauSpLFPtT7RCn3oUKOBIOqrM09dcrPeKPLt1Tobu+X3jziiZHIkhFhmt+O2
qW/UdkpBH215I2BCVwrWT8Z1vNRcT2SVIvbDe6gfAi8TFsO0ISM+RnhPE9+vt/IrEISf/YgZg0vI
iX0spNikfV9qCeVP+ivTnEpmmjjosdgDMUDYcTZ+wHUF1xbnoxoez5iACULXzB8GPU/GfpzSMB/n
Rtxlzktar2XhKPpmCg2MbRN50Gi7wh8JlT+AfaOWddlfMXB8WZlEXM/rg55cZqI2hSRJhN3s+Lds
jvE5vpKxDqes15e+onUe1Tt+2xmMntyAZ8nZp77lUNnSLR/cE1Zc+g1zLgLlETDvqkyyRwNLYzK3
j1bV3s8DKvGwkTf2b/iQSZ58MvwetX3UjEa9rjRIdD3wyqYg9WwNpT7nIfQRxEIawPy7Rw1s16nS
d7VsJaNr+7M2QHDwleWXlzuEm3PC4yKz4/qbHupTbmQ2rdb28Ui/hDwCf9gYJdoRH+sBsV8zwQvp
sub7yPxr0rd3V2fFcqZuHIWd5U+Qup0b2QxPNwRXPhh3tRmGLK9YfD50AJigk/TQn4H9DMZb/LKH
Ps7iT6+rXWdmePUW5Dxqd8kWq45gi9DjKTuijn6DGAl8n9XtGsPPXS7fwzE1IcC6blYosZAscA9P
hJiLQX838S9IrnJRH/jAVrTmSryH5cZzc+trYgM2CK+UiCCRyJsVCI0OSFOHzu7+pQKF6lvq4Nzd
lkR7630S6vjTTasLzxis1IrEyIkYL5PcrSzeVVtlmSw71hmvTFCZuFbEMI70tYVS9aWwuuPC31Ev
w58+9L5WrDM5yDUjq1DJBxzf6DZlVyFnAk5PdM8boxw3A2NfBFUZhQNAPhg2/ZFlgIvyzGH+DRc3
2N+LzJ4GpZelrBJaeH1IYs6YE95XD2JtlrXfQ3AyzWIlwLh81XYas2od+60GXaEihD7JKKAVK9MH
W9CrOWIkTb6D6OQkQXaEA3bpz/HgkBlbUPrgm2u9SiLRDJXNdiOQMLuuNt772cwntmo24ELxT5OK
apVvRAc86PlGFvrDfD/RbLMdW/HC+NDlDUlTu9gyvpBnRgM6gvLz0e+uzZLpBV85pnMHmzkQOIWb
EmJ4T0hPDH4aUte5Nijn48ckZSRKMTB9E00x8pctBuF7hfP8pm5n3+JSQrPffSP6wx7s/CYnydTF
vwo3a6HRQ+JcYddmbH7/97R0oFZzpMm+B1V+2D1YC1ysm/fECEPEbQyLqzPgWlC8zqb394DIBcdn
3AvsZ5/8QZ0bCsALFlwmCSuEqNMKdqkoR8Ew9qzVO5TR9bzzqxUNIJUUvzQ+Rqg1j0iboEdS2VhE
hVDDiViZwE6hQJ8gEYJNGYt4L0lrASHNLiu2dr1ZKYChZVVtogt8phIyZg8D5Yb+s7Zwb6+3YW2A
59iVrjxk7S4VBoOwugTNpGTzzCuGMS534FNZ+wglzv5Pw+fuyB9G78rN6iR1RCzLJ+iO3XdWmSQ6
3/WgoOU4oSSzrZJH7r2jqfh4sh4OStIhSAjM780V+gEjuVHukZ9nO6ldS7dx+5o9BY1CnBN/2Dsb
sSPJZLp9LBDS4i2nXfjGzKVYv5QpNgd/+DRfC7tNRWE61MEy2lYMsXc5wYE9JeKssYatuzuRqnMs
++HgrRbPu3KCf0Zt6kiH/k/e6CDFA4FsZ/A/hNeO8ippbxgf3ICUxgZH7/a2GeLr5dLcY0AfHLY9
9y9VIzLl/cMj0wJ3huUvqtfor3XiImJreVo1hDk1SE239aqE6BWvBpmsEqWEkt+bQibrIXSDoYsa
vLI47Eo17iyf6oyV15S5RXC67q2Ul30i4yUkX9wqLvzZLWH7f8vCmiem9Loc/km+3cDpyM8Eh3xu
t8hNoo79wQpfBfroJ5L0rzb+qjyfy+cx1JfAIz/rOjmRsrUuICOpwrIfGHHWE0QfHoDLqkpk0oBe
I66tOP0wMcK0nz8Wu3J5AMi5hThcAynTz5A/2V8SNO4ZsutjglFilTItfPMwji2089steSPD5h1x
RKaEGej3CfE4gkmgdOs22+Sw9Dv8iSkuBv992zlAu4AxOP6Cg/5hHxg8TcS9oXoH2skkwP1HP8Tj
5QGlDjYqS6gvu7T/DUdlbjfd3a9+KyONFb/akGk9q4GCbMBC8/Y50G5DPeD622S0xWaf9xEfUAwR
UbAjpnto5ahrA5nryE6fPKRJq6cuzZ/asSm8R0Hc/J1XwiOs6BVrN7eY3/A6fl4SniRRaxK3+jXc
MaA9HYR/7YLrMf57a71mQMo90z4nwdF2sygM4UNcUQ3RltgXX/eq5YXJeK6K2B10vqqJUT2Ap/T/
e0i+HRbxfTADhdKBcid0siyRTFb9bc7R9Qs2w7OUFtnQVkd6alhERRsTnra8Np7/c49MBqHPlN7k
+UjUwoz/6RDmZwLB2Os7un6nlbGoxDvaJX7pdmoPPry7L9fbvguFS3izhSjgBidZrRMNKoaTlGok
/415EGWXxXYoZ1m6DP/kusdqoFblEwFtsUXjH5RZlDf7wb2Z6Qab23AW3X6+2zcIe+5bAPKwgRe7
+Sn3ADQ0Sy6ETEPKEb79Inp7spaJ565dKNpfKcJ+xGdnulncqTOXrFuvAffwsgIz5LeAf7L955WC
x1ntlELq6vxmEJW+fZoffUo9SDdn1wO0alWTMsZIKXg0UqFj/6FIjtiMH+GAx9i+gSmWI0mBts4m
fTy89a7+FX2EQETRc++YfTQemmSHJuJYt7LKQAprzZq0Iv0HTVpRg1MkQ8LkVnqFFuGP026B3CDE
kVilzF1TtAqDfws/r8yPRhlf2EV8IxnXhWPMPPDr/BEAH+NaPVzjzRz7rHdhdGBanfUWlTMs9kD0
aFrs7LfS395/WPKZ0G0hJlezon4DiT7am+p2DqfJMsXQD3g8HzIsTwBq+26dFcCEUEOXsHLixTLQ
M4iu1Ycb8Zz8Mo5bI/8E833y9l3XHGNw4CAUVdqetLpNAUSJyLJfF+nE55DpQYBXYpMdCgeFVzEu
BJP5TmG6soH6xBSj5d1nvd+1dzw1rxgy80G0PZJNdYWdUoOJ3siRjUpyMV6w5rOBydVwvKX7S5hQ
EuN2GHS0BeIZ/pqkd6BA4e+M1hAP0g32msWDCeidq0WEiKYGXgym/sJpDMi+4DS17WUf4MnaOoyh
fCS8w2aGZrw/f0FDwU6AtUu35qTqYUYbzgoI+wvsMktSgz0ZXGPEhnhdYPbeE7ycGlc8bAfKa6qC
vFQmPDMN/TkWM5QDYBaaFz5EQ0k7vtOL+v217YKbivyBZt4tOKmNVCHbvYOJ5Rgbg20AMXlpSXHw
bkQAvG+I833PahSjRUIumTzUxJObWUWrr0YZyA/jFSGbuI/CE4w4RVrGlzYmS0JzvU9CkFlvoVxk
WvGMhKwXW4uURGvm1FMJWd6GXP1Z0IBKi5U7xWaBurhtFPXShvNava7b/pH5jekU0tbKhIP98FAM
DCgf4qs9tkBh/ifLpmy/dls3/eLPj+xumLNRM8wvpr8Te8FZxecWjXvwKUon/bL9/KBsVbTj4cQ+
c8qRcHlPhmvhvGyRWxu4hJsYtbQE5laVwpbYrBZRMIHWNUC2dtAJUNDXdFwjWPDHKlosNH2AVqUk
vYCsxs0Wh7wiDCq6HCdtL9ptLACpS4KLW9z9JPN2JsLEVuC3Q5YYGYwMZDav6e9vzkTEcOj5efXf
hYEaS1e6QgLWuFUzWegaNMasStRBmVzdhAg9Ntjj4bG6n6cguaF4r07iNI1OiA3ffnvDlBJGoeDN
Pug0NBHF+jvzyfvcDyuWre3X9uJdebCyo2oMix0ACA3uJr+aGXCL7TlTHnpNCCGJrS+pmhUTu6H7
K4T+wB+Dj5dDDAMN91leR9kNVGWyHTXVcLhXz9ci/r32/FsKHYhLZSsebeZl5MgvtK9S0Qs/K65v
5KeC5lx1rzJvXMh2NSsKVib3/kskuR1UsUmKYw02BMJghYiQeot7eSXNGmLcAQ5VbgJEx44/fi07
M/0VTUikpWrO6RY593qvG0sVbxCB2NKfgouKUHywJCcVrybzQYIojVtXPGLGzHALNOdEfh2eMtFu
BXU90XjV04DyG6NneR5KGnYsFxIsBHayvx9faSM3E2kPfTAts5JN6qc/Itu3Z3u1Mp0fkIGebtdS
rEqaqcHIX96m2X5EZ+lYnDYtkgbpLDYGspi+pYKv6AgytrH+F3ehQIPawoWgvgaWi0yc+FLniZ4I
OI/PUubgkUk0aQlwJlpkr+1ldxoRQZiJSGDOFSmRKCVuJos1lDlxnOkHTNlE0FOQZCjawTz/R91l
UZIiaDkENmlfGeAdud1hZes2RDQ1vLmW/6vH1bTg3SBzVp2+YNoZKyD7LmWnEdUZ7ismHjEJwK50
qdkgOkhGBXeIMpq8iFo3Ouo3aG8qvKt5kv9ARaCb6scI+xWdNhIPfV08/ucPtUUlCAFKqIYKPNX2
tW5HkeA7NFytp/f5q+PFL+l/T2wnNRfeiOMr7fP/n7GWCqCACUwvcATdrvtulyPz8rx3AuzfZipH
K6PQk/A+Q+gwIhLGYUDUg2OngG75ZllPb0fdGxiR9JC0X2Rq30FN/9/GHAS24SiGF4qsVAxuZ3Ua
RpI4pihq8Cox0pY0rwz9R3ZblTAm0rfFezXeVoKUCOVlG7X3vKPIOucFt8NYf30wmAaFMfNFfVeQ
wLy9GY/cQ15LeHsMVzOVFUW3Rj4zjdSQ7FenANu3/4HCygLaGdGjJAlJ12jo6V2JINT1KdAN3mbC
eZdXOnBSzF1M00o5ebxGHoKfKvCQ4ViJyBSmbMjsQMTtGCBiYuvozSw7g7B+mJPolyvI6WSU+u4S
SgmKf9tG4bnLtRzfGTZp1yDUW6VpxX5FH4vjVwateLFqiVvqrgTY3F1R4hjYxyJUuRqZD5rYqM5I
k8YAqO0TVIoNYOOntmdceEoBF4wTfhaj1nCX7ndxWjOPAterzN25m68Re7HNlT0r/Z8IducgSTOT
mYxDUNMFZM/h6QNMPMug0UnX7XCuTDtqbUteP/2G2zLiILHMWQXlAz9nBBUFBwhca17UZCH/XOA5
kQ7Wj+ewAEhIuLDYOlN7KQzTZQJtCGpjmG/EOHBhKTiwgNzIdDAFQA+1iuoF2UKhaJyZhpCuzscf
yFkOXuIXyFs5x87D2YHMVyrUu21gmQqGXHGYy+rsX5kMoaXKVoRLkoySauwn6gg2O+GuB6Lhbak7
XFuWUjBesvSuNmuKTndVdWj3GlVvlZniHAFkgnOpMcyhDOSxii5uOHuSerJ5Smdb/7T4t5tyx0VF
f2Nrp/KOXz7cuk2UjSiM9UvCSBlJW9Ps0nQ9/7fpPl767qnBtTw7mQXcpI3VONmQLggth2t4p9YG
G+62km4cFye/wodCX2zIxSs5+sIpDRDVrWeGZTLUE6Fund8/sONku+ZfC+dnC565gfxgn7vZtyYq
VHopoKqbQKda7pC2R9qCep7kQrtEpBlJxFe7qXFQi5VcuQaS1be8LNjz7q5uVpqoPqDP81YOhF4g
7Mrrn8L7MsLqUbVPBto+PwbwbhBa8tGKTVqosrN44SHluVozhRvxrPpSjZA3zxf/Q7bATXzksrD3
W79zqzgQOofdV0CYuencGOePhPHUCqpanLlejv3Xw3z+QgqPIoOQKQ7M7VDbWPRHJbJndpKGYMjF
cGIgY/MrgtqHZsg6JC0alSv6MmJIIvkhBALKjhaMMwwTqeD45Wf2QMR9t3VxUAF7ZCYZtBjc4Q3M
lwg5I7ceD/lF7Bg0uiEBbaC1DQoPl07zKLmf7NAfi3nCOj/5pbIYSO2oDXROCw80/r9oPQIH39Mr
8CNMOnHEPhje8Pn/WqpeleByoLKnRlNWIKrfDWkvaK1gttl6awyFQNUZByWVDf0A7XJSHcGPWZQ5
agnFhVQKHWcBPKYYYqXt2it4kQecLTuGvdm7oBF4h9B/kVoTLYUSBoeVfQMYCb9PAQrg4G7c4DIO
paB9twlrFDdt5hXGRe0yA01S7iitwHWiEHchChPyzcD7f/fEWKjfQQKtoadrSVjKp4vOPSwZ1WFS
HV32ptr5epC4mgteB9rXRzYdployZi7oUhNSADQnBs9s3rq60sLy1a6kJNpGJISdeoFYftRjMGtu
JN1fEhBhwphhaQEgPmAEDijAm7YNQ4qGRXWDp0yTHLHa5aFELUt5cgx+pDj25Viqpz7gZSHsv3jA
PxsGsi1MTSA/lxmxvDf3Kj3xFOY3L0MJxOTbGVgnIqAhGoKZYkASsCDYy+FCYR5tumRWjBC9mWZg
8VJCKCMXRD84S7xlIFZzGVJSmdmk00KIaq/hsm6MIAOOM4vXHiv0YeohWQBgc/ctKD3TBCo99krY
GlIqTwDmq3gUjXwULY66RihCHNYkBG76PPUg6+7fpG3R3rbPf7MLDDdnhItHItDxtwBfoM3MUIfa
FiV7x3rLOcSUCjz/MJMAm0HIq5KuRjDWrCdFkFxRyoup1jOuc/NdhM/8C6eJ77SrdiJ20OCs6gQN
mklkpuIkesSzY1qeIShN2nyiySwPdxvNfxu1N8EAKNM0sFP0DQbLosAeZ9AofslBVZXszy4YGyld
h2nhkauZtQ7jWlyajGJxAI2tt2NAdxnmNCY0iB4xj0cRhZCMGS8/rDDVN4AQnbM1+9QYWEN7b8eU
JVnOusAIQO3YM11EyekBvjgjUWFOlMv+c5bp5/iyO4Xtm20HcFkw7Kk2ML4PzW0pTcF9O8PAmHfm
Kh9Zni5r/Jkab2c7HNB5KO3jtE7HLj3z48Mnyqf426v43uJ4aTiscRkYrdf3ntXZ9XjhqOXafq6u
DqewVv7cdhp5LEHSv56KbHsMTCA0q+lLHcbQOOCtV42IS9458EFaOuWNS3UHTRLSnzNYXJbjRay1
dq2HESIJ6zXNLT0rBVOJ8kFOMMg0Nuz7867jZnZY+Z2LCAsnBsF6YIzkcgQEjaXrANI/JRjZZytL
wSWenoaew3yc0dtYFpuo4T2eDRrwCga+SVMCkoWNJpZGf2Amq1yqg+MBtpS6lsvUtf0xaA/KcZnO
MBCGQxJkYTFg/Nu/lGc9LKBPCWh6Bj9NUq0bLwA9iCSC4ZaLG/xXoZmJKpRtr1DZEDh3+Tk1+wyz
ypIFqQ9vpMGZJ4XpPNhlssyqSG4pVdfqTIsrxq3CVhGBX4bCg+cNA661NfW5v4ZwuFUhoFAjleQ5
tZ8AMcSI13TRnCWsLr1kZvnli8IS+DWi15UG5v/ba/pDnRZPI6lVUGcLreRXzA976bWB7Wkm2LGh
KMgxAae4pH5yYr2/BvoGCHr73u4n9d0YG1KlhxiXPBxTItkHOu1ztpMMGgTySZVbvAQhoTAvWJvB
122Tstv5DB2+c2Tm/jEHT6v5UuATjFcYcYH/iC+70T89O+zA61qrQD+OmHwVg0waBiSvTvxd2Jb9
Bq/zWQyxalodHgDa0isEqzVjaNpjI6Y41WbUZ/emI1bdIJh6c4RLcm2AbiIroyTcNKQ6XomZ4zmm
J6JhDFZhsh0ZwHis8Qfjzm1GBOJQt3LN3fLlEQ2zVbTBWArK0Gl2y4ZbK02aSdu7JsASOwIauzEz
fFQ0KmGd4snflxCpFaCIrOWNEvjsU1MK95BCfNk7ZNqQH9l0zLbz0AYhOsl0O7nfqN12b5M46JWN
TSBRQgyHAXjjeE1M6pCtjjbwjxMP2VD86g8uj+i4FlKzpNfnkinse5aMTVHuWgHST4NUNUmZTDEE
smbLK0MViHc3vBMdtSnISadZ1z4X2LFKYHW08PIEvooz4giun4/kjMhfpk8nuD2A9cw8nSfM0Wo+
WJxRjJYmkKLR5f9ARO2puD28+Z5VjD+4arUpZGjtG8pfGc7K6Vv0micpxezw51XtraSPaeuE9KsZ
2vTz+EFVZzDYYCJt5pei8WL1Nejk9ggtaDXwvfpMXc25evw5OQxW8TJ+lMiVQXl3Dq4gR9ikRPrB
RQglZSPgNvyi9HH7V/MZNu4k+M0OsMUvt3Z0xbr2vQUtw36TE5Kv3aA6pm9iZ5pnUXzVIBvFnXCz
JlPnylbNVTDojrmIv6ctgJiDpkfRULb/92kwzUn7dwGNY8zIdVnuwuphtjqnfWDbGe444UcmWhBB
EcoHVBeyr0IwZMy6r0P2Zfg74yxR4DytcudbjMpcQHn4wEQfp0nTrVvJozqi8wHo5h5+UCi5yahE
klf65JiMWz1UcGbxTZj3/OaBeWWA5VUp+ox3MekIdZ97z8aCRJZUror0o/wsppgxR/W2gKa545xN
QzfZsow+WE9bo/QGjJVglo8dxVIbV6EIQVMOnSunKyTQ2aM6sN8PSWfPQ75dP7WR5Lo8GT0zaoPf
ru6qxSv8wBBAJ//1KPcZlsYL4nCFIa3qYfHTm5imFf1P88PXCdhqjb8d0ifFCcxMQUasByALeRlE
mdWstg3SE1ZOtZp40bQsmTfUYc0IbDGpo4QbZZJfjquhal4r5p8PCJcYeJjqETOl1sAEn+8qAkJS
VdULkrfhp5Uw23HJaKWFiCIeJgD2d+PyuHlGgjj14bOFJLinDxC7odYiog8YYwJ977A9UC1oHYSq
HXJqf8aQ2ZLXh/zZrGcH67atcbwYql2w6XIn0BqGPcDzP0SqyRfWSHgPZI1dm4kDXaK1BXe0HJLL
uW/Kyfe4ewoWbnRFSymUS5zSxkGDTN/mb8gcPbIDB0Pr0SgbAWvZFHZfVGSFYv5a3v040lz1UUA2
UVygmznedhogvC3YffQUTc+kMtfunv82jMI4XUCsM4oLcuwOI9zRC50fzXxPA55WoG173KsRNgtI
KbuFoX2Cyd66MZ7SEhZuSRUPCy8hoIQQriLPa/EeJ8KzHNvL7l1ZO7fnximQRrSp2RXMTJAA0RTE
ynGL/H7Glj5LJwBl7Y5KaGD8rGbRfEv0/PKbMKEI22ipWsoXUGbPXtEfnn3FyGea7yeEMJL1SSER
ljiGfl20Z4wJwR03vluCif9Rh3TgAu/V3Wvsbi+27sa4AgVD/XRdgOR2VWJQSn41Ju9p6kf7h2OD
tm1FsEptrRuBPzmhrnlOqX3QqTaNj65tcnPlvX7syAONCYSszfZY76SZlYfUn3Xhs5gCIbPS14c+
ZKOSfeHm2nyZWbOm/RSSpXSLvYeyWWKakZYH7KFVEPTbkCeRXUvLjq+SN75Wj/TmKIgsbIj6JSON
HWtD6gX1HAsT/a7y3cAMMbqlUkcn60+iAKQv1+luPeM8Vhl2YAFWSOn1W+qP7Hn0TS0chdN7zTqL
FnLUSygJ/oeRvyzOqg+6+UuO293YwtvRhBhEf3kX9kY3CrqRvRj2LLZ5QMnpggdvnmQbMxcooKl7
YMWddbhEkSOrSr4Ovd2uRVvGo01FjEeRiEXgMFGQuHrecifpqri1PA6UotfAS9jWo24Zp/0hXU2C
8JKDpJ0Sdt6FRR1G00Fd9uups1wamFzVg7i1goh2AkrK2QiYDNQOU7Sq8PsiSNpI9odEORcbw2sV
INIxGMY93VK6bgtrWTk07Pxrj3R1r8U3qz2p6iZ4O7tfAieJLM0JK1j62XP7/pJ0ZhFxaQcaeCgl
iIvcitOhqEYslTETHe+H1lUYtybKtfHKcQe4eJ7WD2qFLcn/6prRwT8nBDDuqzbNdKoamQDj/cJ/
1s1ZIVu7vpz+FCcFiUfFSJK6AkbPzvsqoP5daW9/RFZ5yVJltShIjnJVgGQYpfocFA58uSPzkOog
JARBCCxbe1lNX7gsefMEtfMDSC4xdAzP59GKBgthZtonFVRGHLMCTZfkkgeWFJn4fbqSntXfIy1P
ksBvs4Nsa3fOF8ZlTl6iYa83tpn4F0Sj9HIjfpTavbbBq5TOtkuqQhjY2pJgt/Avp14HJZ69fqaf
CiyF7TY4SJMVTs/UEIY8HAocnanQuCI9CPXGs/AGsJ0ZUSKe02VtIeNb7eQz29V38JR12PoIRVax
AtHzXrnyo84YAURHFqdraQCIEkgZAnEoq35r3r87ORu164fWd+T7V/pAjfcIRG6xoiGRePfuEPmt
XilWkcM1nyWwngwbc9Md+gUnfHQJiAWomF0Qx0cwW7NUOU2wHOKC0aFEBeMYojQDGLwUfIxKEUgv
5lttlsyekQJU/IrmHB8c+PxRMHMdCWzSI3Loo4YkTHc1G0xd+3tu4/oLpMYmvb+TenrVXACEjW1G
8DpibK3590dVv+LLAqEXanOc/ycDF1PLfhD96laIWo9SEWcbT6xLm13y/rr6zK/vYO5qoZvEv9cJ
Me0hdxSHIiiBow10uJS1BCQdaiSBQdmE19bxv2wDafhi1PebXvVuC/B+flkr9+s7jf0fdKifEnM/
VDxiFk5q5mJczlIu2OHfYoEuPFTIxrZXvU1xMqzsPMeE18NfRFxgl9PxW/AAPIasvOaGIvFQN6zh
Xn71eW/fwuTBToyGgRwZJpP8DGnofofEWyp6DpZ3C5X5FRBWzY0LoXCcdVVuk2+k8K+hXNP3Bdml
gvwSHM2JK7i0LjnaIYE8KFQJldjG6yxfhRDpsxRJxPec65FotS86q0HO5CsIeNIUKBrP1nKUFXGw
hF8SS9ARIvozIF4pwMUJvWPJMD+wZa8lva0J7mtvNstcsrCBXFXGU/zD2E48GLWUWmd5wb3938Ln
EZmFKJgz+IvcBuHdOcsEYyDjzQfKZrgtE+VV33PiAxAIRL2GGr18YUiD8bRsFrBOmgwpBNsAr65w
RsUKefH+LITpnzHGZ8KzIatjAcmDIwdVW/YfEywjZ7EVvFCgK3dCw71ayrcfJdLzn5MYMrNJlQ5r
oXZdLVKpji0iSUsVlAXCLH2PVxM0FqK5YnwTZbkEQ0Cz8wc+sWapYjYV/SMEs8ygCkVNAmQinjFJ
XT4Ovuut8e4PBepE5DrMbaGMIXMYWCroJ+3bJ2T5vIsDCeXiyNl4VsdOiWENvSmzvSEzGTvR03vf
38NMiWBjPA2ZdvcIZpORQ+mPF6/eudj65x1kvO1Xopm3lTdrMz2J0TUEtaAbiTIz7PCyEfc4WFtS
8oPJbGsTQUUrLSHQK/21zv81v/Pl6nPgzolKmgMr0xuxGppByuKmb4MP4vzk5HQrGsafgv4kGmoJ
r2TkSfc03bjDcT7PCOSxnCi4JXGM0LRGCAU4o8Hna6A7Ae+CfXO4Y0m9iXQeCE4H0KoQqQ5EKsW3
BMQn7AgCz987k1BIOQMJ6Vji0BbY3pMMzltA+MVDuYgT5Xt0Oc97CxEYxsPwY25zBWQwnu9nQs7k
zLs0VTMzjABzcTvhjcM3kwacHBVEeUeZtc3klhAyVdaYvysnY10oVTuTYwRp1UuWHTQ+21TSDp+V
KzpyIqcsjMmd0J2MFPXB+ksM9X5ssobC4MNcinTeNdm1EewVksw7UQU5d6Tr2+ACpwFA7C59P/LZ
/w06I58OUbAvNBhrc3HE0H+AgssrWvetDb2fJtlWR9v1CHghS/gpDGIkDibe2gLRJ+CgvAKYsZOy
CuEDKVwpdIDdIbzwuowUEHWaOfRvxdTk9iz3u0p0uFcraMU7kBOVAwqEgyLR5DGvpLuKcSQjYmuv
D5CuRcqoBah4wZRkD4eSbhW1fsY/c8FVm+ediXnu1FLqzLr5GZGDgOrgkUgY7dkE5wUACbjnoBma
8ur0w9sP9Z5qjRjJfEj9q9nnUZA1vZFrngO6ERJU8286jeUvZHxJ9ACGai2b7hozL/GI6vbJkKx3
C/UVNP3RTJ2135J0TeAFiFxFidyZYrXtXLYH/fnRqFHDvEXpHTIHJbY1BD/qj7BW/ge2E6xwIrEP
pVmfKg9yHZhUz22cl6o9IsS+uzOoYB0rTkzH6eu/juFNjx5Ahtnx3VsuMamM2J0Z0uduDfKxdiXf
FcLVqDU2NYfyQTq0RbQs4gMfP4MNiVhVl0PoxAuEwcPUBB1BDulLvWZwEV9bMyyrTXavrTcj8ndl
+dnLFrPI1uACN844qm81jWJHja8mnohTTaBFt5k+8d9gkKYOQNrlbZoUolhkwIX7Hoh7a7KaIVz/
Jb5xEofV/iYwOmxbKgee5k8nDDag51KmFmh+sufzqpIS7/BjgbzKG6bv2vOnBn0ZA/MMpOSLL5EC
Re30vgIFKg2izloIYSGu1JEEuP0titK3GHdeIrtYUbzDr8hBXr84ybKh7pZln4QTedqh+BraIo+4
INgM7gHl8gaPLJ1CTVDuF9TqWy1xyLnngTIkGBjwS5bhFSpHPBHBIVq3BpBZJZLBf5jsiZGdGMtK
falu7FJdV49BU2itYvchxeSu7oQ7MqF3juZPcS5hgbNiU9E9QUyVATDKjNjYMV5X8tjKabWVJ22k
/uksj65ppXZwnIPtUA6UyyOrcan8xZbAixj87JHlZuuIn78tMnKblstVe+UvzFxPijGMoB8Kv3ev
4B4j3tYPcdqlJwOmO/pirDHq/6iKBzyFvjzjNJuQWXj7Q4c/zric7fUqCGJwp7LuhlKrokpr/WJ8
yaxkwNVHvz9hE03Mrq/5chFSv+kmguDrHpUakta3N9gaRzS95Vyzrj39/8Y/QSr4ugyIBnuMwmXR
nviHFYm/hlNSN1UsWrUFJCsKh1lI0KzP3koivOXJfiuFYnttcX5KB47CVRjc6H0KROnft7b8kZ4B
woJZHRTyLyFY2T6Ktb7+ttR8X3ecUQmXMXy204AP3hFvM9FOKWc+/5YOXiJLNCdV5r/fW20w2OTS
xHBBG9IxwyukpDeZQiZ56Vz5hMTCiO2m/QLMTCmrI1+PMPmsbUF5wJHGKM1g8rVMFtOaG/6Ec4d/
WUY5b0iis9r30ETQb7Yrlq181ZZWXUOQz2Sq42tg1o7MnVJcslUScG9VJ8IqQHKg82X59P/AMaiH
hdkdr5awdve7y/PBgzwaCTvUhWEl3yeNaR9TheL32MhOnANZgwFZk07vpLl2EhfukiO848tWal9y
PLTyT55l9GZMk+3tJWvjIl2cxhNcjGd6vdmfyL+1/nsemFCOT9wstRJDYy74Rug2FM3iu+IIKxxu
IM2wEo2HqIOtN3luCqDWK1EGRV9DySDLrIWm0mWFHBDdS9KA0xyYylCHU5TS1bQvT5NcR4OPL91T
r+zYJ1cUiq4QRWnMjs0tmlnBtrgTSp3rpWIU8oyC8H7THYq3o7F4GwFQhI8HKP2GYzPiOApoG4U5
bQCwYYTMRWmaQkI4NgN2/DVA9XriI9vTbk8Tm6XFrO0vaWEDXFSIjFspGEvSwFaFQIyip41h5+/9
dyDzStVdqn+iYLTSnnXdGIWjhHtMb42th98xeCF+S2tvAt1dwiOyGY/+y98WoFQknbv9IAVrkFiR
Yp2uLBMqUYLnF6J8Edj61wRD8cq6SxYCpfQAdWIYx7AXtBPCpJPNLJ45IYkWL6uN+wahwTwUszgg
q9O32ywxensgClde+4Z6I40xt+AyRR1kiBhKy2rxO7Nk02qhSy5H+v9kSvnOa6/fU5UQEV/h/7/k
VPgPUAYHfTIwvlU3cfyT3fgZSERX9mXvqE/ktWFelWF/7d1nnFOMq5l8z3XuKZbbzBcW+7HyqgqR
P7Q40+mlVukWuPao7Vx1fZwrPchTc3sTQNcU0FaXhiu5hTGKfeLwwraTMRKphMr5zWCzyhBAjwoJ
rSfBhUjpqVNUzQUOV5DpMKQ6HCzRQePf8ms7dP/2xYqUujOSZxXXp+rBD3w7ZUcisLzADD7vlj7k
GaA5xIQgAF9NUmAsVVs4WxwU04hi4ObwWeCQz+OVahusgW9scSVEUAfk+2cuX19yB/MJF8nr0R7+
I7iOIaO2sRiC/0lycd75GKE7yoBng6p1kBZZ2U9boQb20COeZM6CzROi70MU5+Q+SHSfO2OLo0ge
noa03OKmUljvY9r1kc+MJKJDJruApIhoVzG67RYXuxiBhmL1j3J2OD1PXe5dnfoxyTtCOMFVmQ9l
VpO9yOU8PYkkq+4ffEsfOzOtYZo2E2KKqwVNaa3/8VhevBvHr5lUVI/ZMIHmkoBlHfWWygSeYWpO
9xD/OqxwrmS0Od74F9SLMAFCKr3a5L8GI1A1FDIK4fR4l3m6uLhjXtYTMNc2c5vu9Q0M7QBtkAMv
cr2ATb/xP/fxtSPdlfkeYq9gV/47TgysS6jzqxAv1TnV8bUZers6e9iPd7z+sjjRxgMT6AbjsqE4
iXyL7Bgy45U+ezhDz81Qwu4THC59P+Bcmv2BuM4+sQQqRp5T0n6BY46WfnIsfgHufXPReME4xnzn
MAMLF3N6+ZXqGt8dqkSLK3iaAoKkYTRhQ8Cf1XWtEbdaFbsaLX3kO3OoftsEdb/XcwVt7cwniaU3
kYs8nmbN06GPfMmRMIED9qvygpeEFZ0a0zdnO5/rvuX9b6RvmDhDK0DaTZ4Cs/wUTvAl+lD3BgEt
dZ59IDEVl7RPA885NbVP9Jucc2MF7FiCUelDNboWWtTLD2KbEdpg36HK60zHq0BpZG3l0e5vb/Hn
rkmxYlWQij+pL54s1M9szdDT6T41OuY8869djgzl+mQYO+wa8d1M6MnYvRotfbmyt6duPpVlUUjP
0Vigyn6aKR9TqD3zEXrC1/P4fA3dskRtLA57YfAX01NRFOhJ3NNuCXS3NrVyRZeOweGmvxdvOANv
csrNgZOkcdRWrVsFD3JTi8vWUtaynoCYZfzcMn/j8kavSIjrcwAyVcT4jWeefPHsG54MI5DHrin+
MwAioYFQ2r2CbA+KcdW4N7clctpBYkKkIzNQ/Vs0btLY48zJ5TAF9iY/gEUPtZpED1PuChesyFB/
l4nttsZX4MuD7rJ27BEl5YUNFX0tH1yf9kiZGx39wqwxj0lihu+ec+h/04DjG7fVG6o1oN88MX/C
1pb5L1LBRgsJoyPT5fCdgojRqJxIIPCkj4SxstHUMON3g2guDXQOMl8WBN34SFJZ6f7nHaov8zaZ
uXmOM/Jfo8ulkH9KPcY22HYwh9riXHGOEZleR+PrcAWNV4OENoTOcCNoNJr6YLkv09D1KOUUXe9K
Xb005uo5ZmmVGlRQ40WotjHnkIA7K9H/6LyadI7ur+gwtCzQwDB1ejl6CI9slBGhgMjG4Av/C5Ue
LUS7HuEVUjJRVkMkJ1H+3ukXZB7WyUQBAXBu9r+JF0CZYgjdlvNRHCkuQESzSnivX9bpSZDg1fgg
kbhHechc3huLxwTyyHqJd/l74yh9upiLDMqmXjgWx+KAaYah3YUQEuENSSDkpz3iNZw0obUHr/d+
1S5iCQNupboXWpJeckXKVfvBReJcRzYFDOR3T2Q+9a5botbjVkVtqtyzKtflQa10oGqTduGgtQEO
VnUnhGcZCo0Cto1AixMubjTI7Zv+xCQu662HkK0zhyyw8QdzKzW8ggMb7FonJejDZJf8vUCYNv3N
UD1Ia8ZyUxBf9VydfoeLs4xWYrZ0HPTLORdH0krd9PZHlqNGfjS37jLDbMZEjMBaot+AraaSSLk/
hn3UZ4fC5hE4liOjFYNBMeUoQddta0Ll5YU9SKqEugFlF1leqmYP11LRX2pfVQHN2AI1MV3vRMlV
o5Wj4zu+/8YUG6tKqA0tBfvE9+TVBaPDLIhphVkXL8EcDu0l2wmCLc1UdVM4xwHJ0gXPEI6Eh+Sa
6v+y0A+PbunHWcvJjQfWJGKHZy3ymgBE7a4y6i6i2DM51CSXJI40PicvP483oYQ59TPhpH/eR2J7
scLYPsmeVrc9Gg4dmEmNWRIUHhnnYoBl6gq/eh57tjuOTwXZvxmPbuH0e7G9J3tnSQ0D7lRxI4XL
ja8Y0+Y78yxC3nReeM7kl07ZOFGbsH57mCDWNzs59weDrYU8WvPwFQADwQfkFBhzPa7GR9uC9RPu
MG7vIHVurrZLaf6xuHU+1YQtuutyKPNX8pgO2c8bTHliLijRpuTF2OnVY+kLkxKpmSX3Hg2tLwq9
qe1MAUi5bIrUXhMwG0BUb93rH7Syj5BEqHEJvK7545mWe/axC12GhNXvktoBjFZug1TdJmPEEmMk
q//fuLXU5Am080WLUUIhUk6BcRuU41dCe9IvLqu2tE6PUE6Iw1/WdhNJPghvzvfaY0KCyntwfjjB
rsuU6cWr20mYzLuP8bVjAmzAhkPpGBRH5Dc4RFalmiu4bHgLjAxkW8Y2RRmpK/q2qsr1EBKxn8Je
S822FZ7JjSJvnCLVrljj8xw9z+EhrSAPDTCPCRJXtEfrpfscpK3VyBxto3znXZxIwdBN1vZGy5hJ
nedjz/lgpvc+1Uds0Hpv9YDb9avFhud8sSBbN2xdkEmkPz73VTO9CyXiR+51ReAaTrPYlig5DE8k
4nZdNwDRoX8HlHTq7xgUhZaJqEMSftZFHY6wGg3BdFl2EUsuG9gpr+sz39D86Oxj25anUDRmZ4DF
0EBQ6IRyiI1511i5SZlrn4ek8jEEpOgKcjLPCRx59GPF1dI7I/Be0aqbHaEewH9MAE6tjlJ7mK93
WcBiM1xbiaRjqBDCh0GidWQ6IaX6ahS2GhawYdrRB1izSgsz1itKEm3pAX+tTrv3jwvn7nGcgI9l
CIQSkZg1uB7lcSoQEqOoPknCNAC4KrMPUMLQOfgeoSCYqZ7BVuVcLN4dt+Rj/gGWrqZexpExCjOp
qE88GedOeQ4cMawF0+mi5QGMOCMDn12Bt/WBIfCBz11OH81eCGSD7RNKDfo2zY9aITbgOKwiBNCO
qU9GaIUb+l10woA8/j+rXjrhO6D90jUJoXaP0lRMoT3153mLcc4sWuPaIxGtUds3YEYx83sOdP2I
m/lHcw4vSk1sseMSxO8QfCjBNTDKRiTsck7U+EbA+/W5/apnf1Ptbv4qpTHlhWy5bYfpVFCXEM0/
w3G6AlGhzccR0CC1QORwkgAbOhI4f7G5JrAijWA1ZzpGBZfEv8YmlRjDI9UWRXuCPEGo/NPNr8qh
mxLhxJaDZioDKRKShvHumWj8Bj4LFsQ5PDF/Mw8QTprRwnx+/UTm8rTvCKqZ28+Ja1Rmj9I4negB
wnbN6zQx4x6qUlybjCnE2YTL/brnZiJzJeZIld0Ar7Nq3ypmYcS6Y3lqk1q8n31It+vQxCwdpNAg
M6aSKuf1KCWYcM8MEjFp0EBJGU7O8GgcatW2gidEMdz5PSIzAFjwPpSKBzYo19V98gedkkvjW6BT
ohAY8VTEFpv90uxWpqwMAZqIRrNpRRbPagg1/MEPQ86z3xIlq635Wtzp2RkkH7NNaeVYCEN8Oa2Z
yEtfYqPZfqFuhyz6AL6eSj9lThXt7dtMj8JYIXaCreJ85FmlcwBcJtGqP0iKDoQkG7eV9gd1ZRwp
yXRGCXdqI7au0SWYlal2hkxrCMNXf0axdGwLZIHmKE+FS3+4FsW7AAJcfHGaQAIvnDqbxVh22LMC
BsKKzf8z7AhpP8nkZB9PJ/SK4s3Qov5++JhAFNkwDzYV2RAnDz6IP7y59ngx2wJTx2BOSygRsECM
D7Q40GqRPt+IRIr4ytywygT0Fa8HDQ6zoVF/VOjq1jl0ElwLvS8QG1rQELAJU5OvVGL26tezJZy0
GaX6UCdUFokWjmqVNMe7cC8mL3CMVriHL21D8Amat+0T+C1ZIT/ftvjrMVZNlCSH64oA59xCwuPK
bhqZindx1Pw516ykI4lKNp5OPxbvf+PeOWMK+hYpH2jJSQzpY3lsZ+wccb7pqQbFsNlT4SO6pid7
8FsKYBrY5No3VILksULeO2xF5qPwc67XKGN+NRu8NMEk1Nb8RQL9O8MculyV2vlOcJUrcDJMrmBQ
CKtbN+m9+zPxZhGKuspngNFhmRXU3R6gNYQzHLimZyXV1xS90KRae3+Gz+4pSD5Kze4QT8oBcsvJ
o9Y9v88K7m2jNhGvgxdMLOutTjQSMRfr3n09fL2UQyUYFxBWgQ0cWCSo8/rZjCGTr8bORFLIaci8
K0fT2u2B1Xa70rr2JcQr+6eax4FkuJxlLtPnXoAWnExOUcdmfP2P9Lws0ozfd00BHDqR4LakqlwD
34+S4SO8NgayAZ7q4FW7/mnCbdfVSjF2NIk4q25r/eto2pqgw/uCSalgpF3+zD/wdfoZgJLWqTmq
UYg5VRdhYz7Q5PdJrBQD4QostidR0NIxhexpAgWZqqMf6qOX85m6k4fosqiXQcH1ijOv53Kje3zO
G8RqDaGD9xoaXxnlGjfiNjhQ7L2B3x1Z8ExKNkapnKdEmmuFcqSPu7u/YKI1mWEMqDjv4LHiUG2r
1vWcGMhXtWnRTxkk6xMQfSC2nuvo+mQu+MD0H9uPv/ifoVjmNk1lyH+8HRdlm4x+N526cnWnCITM
6dP+R7BMESEufK5dMtzBUX2fQO6gwImbBjtNWKwSGtA42EFDmCp4C13kbpymJiVr8CpCm/U6YVDW
UORsWrEwUo7TtY5sfAtKTuu4AXicY4dzpxnN0MEy1/nn5SKNzRXBAbDjlHLTW0tU8I3hvTWLoMlv
04Tcj2TDuMvgEKgDYTBDQugiHOqBS8RXPmYsf3GfIP3HFxT363L0da/WPDWGdgCtCgE7Lted4gnp
INfLbiIwzO9T4Qr2LngY8NHASDpdBf4XP2qDejx03MnIb1hXmCj3Hr5+3qQXH6NockgHHhdxuoOv
nozOptm6jS5jFVa3P0vOXH1TlkWhKZlQD0qrN6WbTlzqKBqroFnhSyRh6WG5Y4ybqeSUgfqPpzUR
Mq07KvigpQ3qojuYmteFoj6iCU9mLTfES9GJPDhY5j022LVHqRB9qJR7WTBrbZaKCSJgsSTprAQj
jo2EtVA1ZTzlhOshGfFgDbAJ3sBXHchDOn56IFz6BVbVKc46I8njlBI9Y3L10nCigDZRhHFs6vqQ
srieT92gnk888HMm1LaXaSgsaY55S3HITlzX6LXCcexSJ88ABiGAVDoRhgSBmzl9PnIB+3ZO6MCK
udktsJll3UaNmy151jQerbImRDfb47AQA4ypSlpbcOKwkvIUkJVWf/CObJZrdngn70UVT4DLPaCS
LhBP/v75cQBM4nMgdYXdDi734hAC6ugZCYkJORKa5gz2w5znCqcwP3iRvCtVSVlRCPymtvu+r/wE
JBe3yZ05LFXe+8MUV4mpQMKKyaw/ZTDa18iBtBsLm3bLX0jSinYmLZ9W1PWL/edcyq/tZ/8k7qYC
p6XAvcYyxxDIeKfvz9lEMm+2uP1QjWvdavMbEDsMZQNDXSJrUaurcvD3sXNIuVtHgDcZag/m3viV
p1ndNOxj0230YJhqC78JGZASVbbSz3sTGrrGnMoYtQVVNG5oKTlRpN2Jut5KOujguiB9bbZ4YxSc
3vi1HsTLbv1dnoBzhj/swVbb6+1neXE12nnhCz5aqVNJSqUkNPEAycVuN1cKxBMNTHjrqnjC8sQe
0pwtLwNextV9Tota6amyY5XrngCaenJypKoIFFwgZJYVk37GGvtvZtB5c9KhsY1ZwPrVsXeqZ8zA
guVnoXY3v6MP5E8JkpDXejnREiPCpnRuKtB8uzZcaODnUWAjOB62Bfp9+hLNiNx/VXHT3PsstI/K
eZssJnTK3ulqoXmdFCPmzjwYJcwJX5YKkFjQra+aaA+Pe01zFStlqkrC/xzcIJzBX9p8k1qcIis5
p7dln1YpZ+4sb6kUn1qKjJwfVmqHmUiZ/gsdFas9CLeDApV42we4c1TwrChtP0iiQwp/N4uyhVcQ
bh+pvZY+r9tZZR5QhEU4q9PSzCUT/N7GKBqIjAjl81P5KZu0eXITmuTy/wE/X69Ebx5PdBwFD2fu
EACa20TXdl8xY/Ik0XwkOn2UD4EIKRd9gaI9XqFGnGHa6WenLy74U5J3J2/qFPyaYyr5y063m6kb
e0bFHXJvbaotycqqQcq4KifDgBAxP2YWh6gb/wGJLRlP9sq4cJRYuTlOxbzAakcfVENPYrpZUbUY
Lkw9QAGZHpECw6Yfn6UkF79yoreFomiWqFnUhouJhzfHju7lSKy6r0Vn4cpCnows3XsKP9fvoypp
aMeSHP5B6WSj/R/7Tp37bNVbV8XXmT17Mt0bt8+Q6y1MjWY/WR5tx2UbWno7iUFEFDSq8fqNx7ih
ADtz/R/HcvJxvstOchsBCpQl5+2uBB/NeqwgB0Ia3tZM06xrkAIPy1jmzVy+U/EVWXaaNIAhPatI
WjUwbIvNdrcTYv+2VYzt/PqotJm5db2wAwJ8xbrUhLmfny17eUfTGDIffMd8BXsMeIggdlGSoStI
kuBBT0XLI7UKtoTZ9AEejq8e9/AmgYL2YLmnSOkrbhWev9TdUN/CQYC6z7oK5azCqjgHBeEOm6LM
bOa0NWcYAc839sOHRV5ACN7sltd9HYowh9S9S77Fszwk0D18aw60UGqgXxcvNd5Nf93c0scfNoRE
uuKLir3KYJ88RLagldi7OjVIVzhPmOIYadv1MbE5m4Lev7yKKLJM2HHoBHUiqO+BHnp32FQi+WgP
nsdirYFSE+0aPS0ajKFXj3A3/AWDlcYGZUjs8Ot2+med3NZL62g3An1oWa5Zmsml9jwaY3CWeIvS
8jyoR7qe2bdOGJQgqSaUF+7RRs+efBshVGTFjU5+HiwvxQ7xzaSRUuFzkhCH1FD0RIfePMg8A7ee
b/5TQtQ/iM72nsk3sEPSU+WtXMOFD/N2Wt6mY9Gqc4Dwx0vEHdZgKEQNaIrjh0QveVgzUycmpvW4
Wc7rbKZjJARfvIJJvGnzoXcKjRQ7uc7Vw/rWrnWxAl3bStA/5hxWhUeI0D8Iex4AT7uN/vqRto2l
6xwwB+zvPOhgrH0dlMEdwGtgPGfwvJjIWeL+oO8W8ktGekMPJgBzPpTUPC8cVBtTRNbR2Zt6Jpsu
BUPbd08/yU8+oLzP/WRw42iKhmMs+4s+Jox4fyuzU/d0zdjakvR873CPX/+wsRxZWh5kiswmqmKq
QwtbeagUCXAz71MfRNSn897OLNz0gAN67KrCd1b9/VFgMNFhkfvSb0FUhmOas0pq3idsHgx9AawC
uxUZNVyybatkED2YQIM9qRKV/59THQ7K5SCd2X9RAjYOA2aUBDniuZExpT9084PMUCijgsB6VKNl
xwwgGPJCVN6YB8GXZTaJ28sZeYjjryYarmjp7xJbs9XQKwLa0BHkOLe91CCDRugQSkUomCo0qc0U
8uZ0bD+RqP7wMwTQHAQK82Th/Pv6269KlqZHxOp/LHw2n89enn2id71mzQIb2o8GMXVDiTyrSsU6
pDzub8OG86I2my17ZDYMY5BGojP7c5+j6TWsUWe+QwYhbJ6lZX7g/s3GMxe0EW2e6QmYcO0+wq0L
ZkdLD0rU7EH0TxqVvUkMjIF+OZ33frweo6sSzLyT5ZTxTKINR/lY468l1LNd5ols2/j59ijYTCtX
vc89WA65VE17xh1Pxmg0xEAJZt+3inLtXDfPo7dBa8jnnZqRtRDBxoBWQsX3SlGQeGFkVc75HqQq
2R5WNIMLx8Kzuldjn2qk7tFFm3mJviH3txVe+j2PRDmuqkldmCxDSXXPLMX4t/gnn2N+01XHUuSd
lhYjzFj3M8m+VuRY5HAjJPt3ks1qbcbK3X5dcSsnqzLiYzv+W31+i3mLgp0ONNb74HLloy3OUNKw
m8GFdE4eSMu4jsmzqTq0pWLOLnwNbBZrLPi4f7VGs/PCg1O32pSfOe/99pMEsCxW0D0sexvdpVOo
DwNwbrlQhJJ3aVOZsNDNiPBEQtg2r1IJX7BHiHCbF9tMcVCzxnc60AWHHkqF2Slv8OlmpxmiNT/W
nw9UCCekODJ+f+z9OH49oO1spGqIrpshtn5ibVXnf4v1PVo29kN1VDqVxJguI870lOODO51urjjP
daabJuS430UUuqMuFzX1VYdJu8d+JnD7jbSPnQIToL4Y1Us3fLMm9TqVlHn5oww83BOPk4H39U81
dJtV5VEEnpBAlr9Djr6p/QLcOI75z/dEGlqQxw7TyECoW+NHTleN+Muj8hnR9qqWKB6CqyzMThlU
xi/6asU7EmA7gZBfqshij/r2KgNjFgFPzNbeGt9LllIAokxIOAIkdD9KuheJltaNPIhCeqDPcIc0
dHPD/koPTB53Yz9si7BhIt9uGy32JtXkWV3QucgKp8vHbQ7WaT31rQdMzpkIOytBQ9Wn/P+VhhT3
uy9MryXEKf88gVlDpJbAoFcrBzXMcH7957M6YrCIJmK6TeQzK2x1uSEWX14BseD4aAIqxp9A4J22
qPNg90n6y01tqPv4lgroIpCpKVPbx29TE6NedmHKB5L5vmkN1So/IGd6NGJbFzLfzS+03H1876YQ
Cj+PAJajPSMQLw7ptZFv/3GSDp0FN0CDY+0PkbiKpHATObzcmqKjFTju6YNpa5gIwscNsVwViW/D
PcsBNvoqCBjgpZo13wSupsyK6E512x7dD3sK5ENRLspX08VVmQv6vPFJYoBaWMnu3RpmACT5esIz
CbXbWZhggWa1kzMficRL0GOKD5a2LOT7I3M/9QwqNzoVPTuhr61wzMDn7DIz1djx9+CQmUrBw8Zy
oJhH+tX4iq14av//Pk4lCqr4O3f2DTq64PgJrTtYuqromDdY4QdBgS70VVcO+nu0zcMU2Vyai0hP
iCPy4Rs9IyZbWmf0KmY4qI3iExzPvFthgIVmvz/bIEWrG6oU/YfojKRBUhNErPCG9CKT5OhLhaUi
UblcC9FnLr597fFNCf1J+6V6ZROdn1BKuXAdtePr1/BbAJ/iSCvOPS8H+RHa+3OLGey25u5FXsmK
qPUqDdWzvL5AEanb2ob2dA+UNGhDFqnQN+5RaRkdaZzkUuaGxfgQqmhA6oX40gH9ByCuN4Brf2ZN
lzm2DaAQiGw4kxmyrBThobSgujkHcKVImhZv/gBujdz4UQGls0g5qrFbBMG5Hrfj/eAP60sCmSsx
AHSXEtIEwEIHRuUpf1UQ5QyamhmVip72CHZiHk9A1r04lg5EagPZEQnAmxCoMM9CgHKbLUf42aCt
H6SoIwa6NxY1kBV//LMX0Ug2g43iHKBA3zaEkIvDFnNGz/+faS0x24xm0eVI9qviLZMaxQrgDAY3
w8wT8psseH7wvsUPvRa9nqpuJGkIF4tcGK7A8dzSaUoIjC13ek09SCGAUcvjsuCYB7uVPahPAmeI
nLL4e+Wa+7Wvm9moFIyq42I0cu045yO9EnPV+Y/+lSFw0ylS/q7SVKSAA+1rHtQULaYEcyAzR+Kl
Tnz7RHj3kK6mwnc4rIC5zzzJ8VqPl12BD5/tJu9xQhfB12I6VW/viKxQXDf7juQt5LW6Vrygo2g9
mR/kXWZIwLR5LHzUHG0f2PBMBBKv8Dmbpv013F5cVVbPXF66hPgj+jmrWiv5YKJnNZRdODfS7WPA
jCMtomS+fiRGL5Qc2I4G2eOy30SJ+idAq8sW7sjs3fqDeMlfXoGopstEgAwlCgKUqYFRf0DDv94Z
dMnsxILBaAbE5xrU5/fEbZTBXDU30QQo4fWpLX4GTRpjb1uwxFCt4RW6sVSNUPKzquPWQhB1Gcsq
VFCNVcn/9XQqGydnY4+otJyFGcxOCI2y6dqjIgOihN+5IwEvtahab+/WFTR1d3BK7uTPycskFiom
848UGZVjyItx26OyI3rAbPbUtPKzdnL1KW1ztyikojYbhVbE6wabVZCMFraV2N1fIJvHAulizXrF
07/75SzFn/zXrJuWxsDgt2VpBFJ9Eay6j+zGpG2wAG39ouhkR8B0KcxWIIRJ7SdXW5I2p1FCEov/
ahGxDtFcF2pWA2NtLzIx9fvEXhckhq1nzbdVWXWna8ugknEWFSjRACaMXCI2MtAHZX4PIj+vSikV
a8Mkj7On5nUhAzShVDTWOBaUAlcgy/QVIj9Tz1b62cj8cKa3Ry5q5wToCBJqTdY0waXI8WbX98mn
cC2T6E/tH6vmVdlTDkwUmTC0EOwM3nqWbKbP0I6/tzHNATWY5s7mkSGB1qK5Ou+mDoVsZNbqxv5y
GZt5/WnMOiOUfs04rZ7XUP//84/4ZkzeiMRxItz+wD0hyYqqTYDYILH3Yk2Gwc09FCoI9hRqEZEc
cXYTSWf50ZiI1r2zPasut9cFx6UPW3YG3QYv/FNlnniTLT8uNJalU78jiZ60iKTG3H0/3xi+sMAA
4BSIKAZyooz+Rcb8gOSRbNTR2D63cgwnYXnGYCFCwM7A4M94KC3azg4D11hgxP6rgNEcS8TWJUuv
9jVY8mFE/d7thG4ete2CmsRfsoFDXZaglpEnjo0FUMBeW+rTQUF2huBJB8JHKnHtkTRn31Nw9XDF
uyB9Tly38IgNXicJXvyHq2UEu2U+1mcgQmpVI5k5Onnj4EGTKs2t7OcMVsn7h/xIDTsfavU2pg+4
Ffpy/sij7OS4kvGE79OH6H0SfihwtHzfzIb/2jRf6lpB/vzZB1tALvz/VFojTznA6mSYTPY+qztJ
aVzAy+aylWcC93j9Kyuf1f+i3aKN3/vai52YeR20Ef4LX0+kEXM5oHBe5WakpAzmCimX6GlJI4wt
sBC/FIO4Ww2RSNp1U/KmSl747R5NDDXNfK5vtO3JuFzx5n7L5YOpZ7Gd4nZjf6grP7LuOccLPD6q
z5/BXOSW2YaGYQjwlsspoF+q5gC1fWrzUcoM/FcB/USTZoaX+Ec9NnrLKZpKGW81CFqcu3XYbiwo
Y8mFm5Po4drXuCWeI6QPWkT4QKBoTj0IFgiKNAiNOGWSzBXyyp9i2SAPKhnIKyaakg5tk5elDZOK
RW23N3IwKxzv+gnsHPFgD6rwNW13CdbXmCG7zN9iXqGug1X0WyXpohtX5/iUUS659SUas/iP4Z1j
la0nLxW/V4ezTBW7cQAoplfVzN4PgfyDuRgrtLLaS4ccKt2nkbA5xPPlrlANgma8ITNHTaOQCICy
ZWvIzlVkcP/lrG2bpUxbaQkbrjFLa7s7/MQ4iGe4n40xYLPRRveRuqkFhk1EGBPYDqNFHK6Ixj0T
TBp6K9ZxOXRLIzVLXUBPbOmMnp9aRqj7+eTSE01oXf10i9AYdZEBwNra77l5GLT0wY1X8breMNJe
4nOlzBfXCVf/QwTqYyjtkOu9oQjrAs+aSK2jyE+j9d8sHuzKE2YHeR3r9e7RcMYUpifzXRRkFf9Y
lZu3N4DeEKACWP4HfL3kF732kjLRx1vDY6WpnRyXlZgI+rtR7WYsYAXUXHaOeTYCPPf2GtV0yKew
8IxPZaBMRjjmD9mUC0hGfXb+ODBdifYbea/0OHh5ytBjh9jEf0PnTmHmd8Dg0Rs/YwH1oyZ5hkwb
c5Ni4mMe/Wd2wZFryAj5s1hQyI/bm5oVLteozX4wnt4RZHRpaL29r3caXU0lnl135TQQbG6jbdiu
TkiI8GJILSBw2QIh3+ydAiN+xfYYz/6BKIysearUldlw+ODVZTtOO05lihPokzDMONC2BnnjgDs8
IWcTPVqw8AdzqavjtzLfsiUO/cHcMr+Vzo61jl7JWxXV/azCL0qkwIyc0svyp7PRhOedEoKt+/lA
YHtaQDlFKZCOhfW7N0KSU38yw7xGaHO5zfRYwPytqRbSXtPXGV7wBktACzku0bZ33NIuqyHudbzg
YlEEYlh6gaqVDKP/ln+0uOs9lP3MTIMvEAgdKO351Fakp9wyOuvMqvOVUj13cFtpd9fZiEEOzRF2
u3CZR4Elnf3hpXTtsEIDev3M4xJe2bCV7hMh+xcov82QoTOPTtGYmPaoVknBqzbgi1ubizE+AYWQ
XXTjnihUm4vavMtpPgweWH5Lja2wcayz5QJt3c64yNgOnGeFnOpiA2hbbuf2I0kWBvO5laHSLFZV
wVMzx+/Ob/u46wudi8YfBD1pdcuHhqu7ZbaYQZytsnVSHRJjIWaYgSKt6BNSxw6x2WBrKpa8HhMV
yt40D4rcgzjgJrhztarA643HyS/mxQEKmrshguGpek2Si/p52Le7FNZtInCRqzoNqjG82E5q4w13
cWlDJlwI9zebmYJ+rUaI+s2MvaWublSn4j6tOo+8be7QHv/1DgPq4b35+0JGH7HImoa1w2dkGVhk
nN1dSflumut8BkZC4ZVHeJMwLMwSoDBckFRZntixfo6dMVAcQGYgqdhvALhWTHj8TJMqbiqQRj4B
5agf2m1lYLHi5D5HC20k1Tqrsgd9kT3XAfDfwU2NyMWobcvo6X/3t93FUBhXTRHY9gSPKZNeoba2
+h8LKTsoRr0KPqQeSlYn1ZBGbqEeXKUw3Nd29WN7I6aAHWYr44isII/M/YbKLeoiq6IP51TrXnRy
yJ9eFajJo5G/RBG5a3U3XRJvqh8ajeeyuO082Ws36n2dUJbxWBEp41XJkbzAKTYPhpSTbCa4LCt1
cfXmRJgSuZlN7bDA9s4SAco68msaSpN+06cZhA7h/h5BlmtCNwHwXSm6bjq1M8gpp3HK7dn759Gw
u5MgCK5ANg3Qj4gJ1BqccuNH/tezjAQRRaJtv8PaM2bv5Csx/aG07rxjrjMWQkaYJ0xt84nSYc0W
Q+uO6XeP/o3hRJbh+EM13xKjwnAGjNDmRC8j5i9/g9CX1ve0Hk/1b6ybZXrRKzbnK3yW6Ci6l70F
fUaG6WNkc1wpEuXA0KfTzzl/J9Dadw0hSagqPBJjKDddQVf4FQU5eoGb+9seHqluDW8dtr/OWR4H
r/tqNbEkRx6e8wcyArc7w+b+nkwfn931GHeHs9YINKgXaPo/enHuft/hDl/bWlGblqsKkOis0vKy
u2XQHn4KGpx8CWWhpbTidlcXh7pNnzohL5TZmJ75fUcbHhwTX2mOBfiswmn3Te6jcQ+jxKKQf/8a
T96pU39OVKX+pq62D6C+buK5AhQzCKhozb00ZoGxYw+jtNL2my6Dd3jF3jPbLzpBsZIL+0fKxGMq
FnSAy/xpB92r/yggZ5gS4KsvzS5tUCRyUOqL7zwNMZy7yFAl7ndpOm9deXioQRlVLhz+AkHkiNr4
sGrdRvBkuVKi+WRSAUXnGTx0UKmxILzWHZkzpfdESYszaRD2e48A/95ii709GTDCDDI8pSEr5XPt
WIpGyPOkdhYdfQk4uWWzDcShOcVQPLXa6fw20tn5IOIb2X0VS0f56mAxN3Aq32mdKki8DbvwR7BN
UFFGH1AMw51yvHkgxI8QGsVgoifjjNPg3KRlhdBMghTUwFsKOsEh/c4loz7E7CerCMZEvt0vKfQA
UlvWuEPUZ4e3ti6u/yOzjS9IOAzllvOGBim6xqBRh2z/uurz9BgSz5fQj6uZw4ufUdcyPT7StJ7T
nNyXWe37UcbjSLOvWQ+QeqECjty0wa1V9L++Sjz/xixJ91SDMPtfERDBUjaj0hBonkxkM1us0PDF
Y9kylFPbTpRZLbmNWC7BIF4MzhnZGTvK2im+wcdhEwy12jxjKa0Js5Bm6Na3uqE3hl8JCRZo2wPx
4I3+psHhrVL64NX11Tbb4usd54pFyBJ+Gwv6uQYmonaRqaRY44L48VA/5za6YbonbI8r34OcvUN9
b8nNsI0Eri/ciWBbrQyYHwA8Mly9CoGBUp1F9ac3wSkn0De4kxn6YIK8szqvPfNEx6YilejeG2v2
+dcer7z8XBLaD/QRF62S3lly6q/sL71GfGLRA8VWLC9Ap1CkYjyq4uKFIKZcTsr3wqg0nn6IH2we
YVetOaJfPcZwBdvhZrsfjraCh+FhAMnRc9Q7XRVOCrbdoy1y3psGLV3Wm80XgtNYkq5oNLCN3Zhu
UJ4v/pfwlCNXw3JrNMaOIfveKCPqfRyqfKpdww6pxr8OooTp2rF8z2q2ZjjqeS7yaVKlq9G4iYOW
4FcLw6AGlO/X2m+xgHG2g8aVs43juuErmKobCKiyV7vs5+jQf6ZCCCFe4zOpV95yUjepB/U3wUK8
hwGbwtPvNOlu8FhUOhKIMMskUMYDh8Llt3gnOo8Yx9YKB/c25oa70jXumxjqZjyo5h/vO8TkoyH0
ePJ5flJGWib6Lk7ACcr12Qlwmnn/MoaGsyI1Mkup/O7OHAj6frZPrhuOlQwvySKd2TptAdwimjwL
S8PHgJIipS557LxkPfuMNwuqsGgvGJ5I+WUIel8Of7h05M/oNK2oClV/ErLBHF4r/CPlw3d0OhZW
xhY1oRj83gs15eRj4yJqH0uKiBckEnrIua+q65MlAfLW0bZLBDhi2dyhsBFC8kGnUdz/jDNzs0Ah
OBEx38OjplszmFJiQ1eORXFeJW12lg2nuIXqseJpya0WGoaeeW4AGUQgaRv39pT6q/ThuaIW3RD7
pEZ45fIhBQRLyAnBFoesyicHpyYnPfRVCcryXufy5W8T8y+nLm4QoaL3xlgyF99rfDHDZqTQhpOV
Gp3o9id4W8a1RN/k5wBMcHnLE40MqAa4FxuCaYZvattLwUWf5UoZ96K5BBbPqXmKtn3TWtlSH3Yk
/GpvdICPXqOCTHQP8sIs8t9aCkcS5ckLI5qhXOe0Kg0IDPdbxnNutca7MnaGcfdNUTfieHwZxcVW
04MHFoTtnH8GOktv0/l8pzF+LMd3HUwD0hgxO1y6lzOaYvLWRxW8BDqcb2jvxzobq0pnY4Lp1iBo
+ZluBHzZZaYW7ZOE5ND1/+2VoOyGf5FGVZv6BRbeKObt415RvO+5MOauiQz68y2R5CLMwxQtJ1Zt
GPxv9YcD9cIS4Cpo0aYSxNkwouuUiPOsBQtRQQkBHLxVNKNao+Js5EBUTT3N/Zq4xdCTGzQyzOZB
yVtKc1jd9t/HvRtjXFHPzZrdSSsrQsSAOaooUIa+ovh+Ln5Ia4i2r+gBwcvdjq3e8V8klFfYEg5F
WGshPyOBVYdb2Va0zjsRYaJYnj42z8NhIibynKmy1zesRc9AGUgQlZ5bjKRWrxeGzJIpvYJkMJcS
GUWLAqWZyEHKsUqqPTLoV3pnr/X6MgiPPL8nsjclIdUvUymHCEKzamQFDJBoMJdv2RSCP8s6bg93
sZxrxdyr86nt0JQ1kodyHHOw+gbpqdIXL3MYn1bHaqz6e+X0HozojHTCc3MVM2vocDwdxyKEzY3z
3oYVFLRDiXIVpqCrWnc15HUxisE4FvHsJCbNoBATRmL/aK22j/lT5HPze1LKqMdek5iD9caeS6sW
Pb3JNSzLKzgghODTFzTVtXZAfRpvqr98FzT8QpVfbESuOpVmREx2plJJt9woHicNdT8XB5SxQrjX
qCXHQuqz8tcgiSm1W08OQl5PvajMIGIYXST0qdkLJDgGryPoZSngPkBpdy3NkMwWNOKWM5ZQPFMq
GJ9v3fjKhO3sXyjMUytaA0dAKEWch+doNHDMfI/5CSQJG59YZYJCtGFa6XqBVZNqZQHHCs7PqXbu
eD08ilZiWAoGbw3PRMJBTY2Yt6nQYClx9S+hWLUl+icbP6Vz8e/sK2SyQ6oTTT1x8n0KbP47jQd5
8UDzP3bwQErB2c8+pl1WvF/kP/chhPv1UvFjuoNEvMablcOyJGsdvI+ZRFKBqeteSmhFSO2Fvt5s
i0SuDO4MIDspftBzMeN1zkxbglTh9UfHcGiWxqlI973is3c4ePgDpvOSra0Qk4WQNW+TuYMCMc1G
g2Y4oVkGBNRAblVr+znkskO3dgdBvCPDe4VSdMu8VaZ182Oca46w7gllCmhrOdLn2GWxdd1idAO3
qvXjVB3ln3c3CM+4iSWFmmZTtB2LmDAVpqv/okYk4ITJX0thyvfQ99F1mqLq50wk0z2f2n1ryVJY
ETrEorZg7cnQVYHMpBw0ydwCwOc/HtOweGJFpFDL5g1cqTHx4FZko+1ec4ZR75TY5RLDYBpQRz9O
+8/Pjvbg59EkYKOyZTIfk+dNb7yH5ZeQxxBeutL5OGF5Ujg8vNWjFVCZbVIJdVXABZSdkBAawbOc
6eRiOFcm0UoUGDEWGnwq3iFjRfceFqVG8x0uL7hfIU3uc8XU9njH/y1ekM0VjS0SP+wvLkWY+U7V
0bw403P1Sv9SFcYojNmDvLMM1GCjaRXawbxZtNLrIXB1577SMg15w50ZRymjOSDMw4SeQyxNAu+p
RJ4ONj049OGPqqkx9LlgOjdGOD4JOHkrR1PGtX4AXO6GLzhjnc2kPhhUkpZGbsnwIIntnHbYS6jX
mpJpZzLKKYG1dmeP0D0s99KfwMHJQu6G2wEWsdr+4iobelTHojtzgn6lAqgNhFCRjRqGr+s9SMGB
qnui5XUu4HnBj0STYoncfZ1/PdX7Xm/HlCjQ/O2dj7JhtJtRDG87OKPoMljC61n4wjnFCwpNym/O
iPOoT0OzQuVr8CKDgXbwpeSbPMJZ/yqrx/0ucO32KDkKBYeZaU0cDdDKio9HaCQQzJK6privxSlL
+vLe/+S5VpL/C81UZuY0jeoMmHReSInL2BUwsTqrDHokozUp1TCTGWXEYKmau54r4pQ4W16R+xWd
kNcSMilQPOy3iCaAXPRGfaVEDh85a0iQkHtwre++UiEjj0503pMsQ+JabSPt6CY41K9PcpVAlnjy
9bqWzC4et04ljw8zunDzcBbgHScN3Y9RaPFfI4i2YogKtBr8MYSNIrKfRcXjazi3rPQzLCd92mqw
20t1K0A5qWZkQHIMumnR3ZUO58zQJzcX30AjpQ8VZvN+OxE9z9Wzy0dtf6CefX2sX1eHtfwD691R
Xwy5AKrIj1nuw/QKn8N/ycXqBcIcyMndCsBXxs0X3tSR6JtmY3LGJrdyr4d6TUhuMdUOZRLszz0H
87bSyXe4vczEqpxnrnB0UChSJ8sZN8hUIQ7Ai5Kxt00J19YU2B2xN0TFfrwNl+oK48KetKc55Dvm
iG85LoNutUjQLEt16+OAYowB74eEDY+65HieutYD9y29o1cI6weDePeagfn0DQWcwZ+eci6a+eH7
F2DDhXQ1WNziNDlsVppM6C/h+rLBPoMJbe5B9fSTMR2OZr2KcimZdQKCiFyVc/0jXdA2gTWAmeZO
Dc2JsNRaqriMjvKKqLd88Y2KQMO/+bRXSPrfF4tsmm9MZU5IDQtNzHJyO2WmAJaKNq4rA4HGLaHi
LtgKVeZZzRe8FMmeB/MULuiWuG+MV+F/IjSPzTN6N3yGMlQhDPSIYylwgrZjFF+UCrYDQlWXpAA9
qbzbgRQMb2hgEb0Tea00nP2GliqX12mV+LudT0W3NdunkM0u9Iz6W+4zxrtdbQ7qrviPZWy/HxSK
QBWGll88O6+H5SjRrzUadUeh0afVFrga507Iq2u3l6myziLqZbSrNNKGQuOTtb7AuSmQ1tlXx6dF
aGFCARnIp+SFd1o4Wg2lDcJVMJZUDmrwS27dqrZZ9rIT+SDzMzyNZAk9/MwqBDF39u/E5apfH2ns
poTmMlWVGQ3VtAFfvQgfjZ+7qYLlJiCJFOrLoxnD25x6DaVdWuvIj/kJA+qdB4UboH1kp55UV/h7
isZ19H61R8xAKXkNCu7O17zVxjdE0RYj4pJAHFS7eOGhAn0nfL1a+wl8Pra1oOjMH0ylfJjhyfDk
PoFey1d03bGq4Amaf3a/hNpjcy3EfckfMNg17XooVQk1eMA8wKTUR6mA+qkRDA2J3METx67+Ztsi
OyayHBU/VTQeLfZ3vwLzfjVsBIOGd1W4I4zSOCfbXULC3cVoD0WRC25Nbp/CmqsVSk1m/NnOoZ46
QlqMTY14UWptPvZrF9NWEgmN7vpYvB6HvDT2qpwF2Ja8Yv6GFeG90FqCgT4vPSBjYqJybgOg4A5t
WQr4WlDbkzlqWCc/WBJt8Q/FGRCW8CE+z0IFbLZXHLDM4Cj3221mAOjF915r7FL51JPPK3ohZvLw
W3M9LDJ0gZTu+zx0p9ZfoEMGmFllVLxdPbO8K54LU1laBJq7OpCcFDAbjuYmbtTiMeku/oAnhEEj
+eBoZeNFHPawq9cOX3TnCD6JFmUZHD9j88KqgJihN8P7Nqrgyj0fZbTT9Tp4AFY7Pcjyk1ZOJl4o
a3kAboGwRG+Xaf3GAA4axJ15w5FWy2Xjs/UEOcaekzfnmBfAd6g/UwuFaqDx3z38OWbQQfdmfCik
oGchL0A4j456VIhuKYWIxuQpJiN4zDkMklE1tt+EsNqvFKyYaG18R1qNFNhfUkrbnMHhORdYxOjT
ncKnj8ByP2gCGftyLc3p7tXcg0iGMdKZfN+sEaVBfuPIwAItUxX/T1dQc79zJcAt/7ahpkesPuVG
r5a+xT91Zfp+s0HrQLxmzRDDWWzFR1e05LcIQIY5+VTjA2VRO1+cRG0xiRA7JFFJFxYZ+Y9uorb+
jR7mCke4+rMOkvPTgDjvoxvqKUosFcNm4srH+3Sctk7E/QWUS+M8PuBZFl8UmafUAfcoOd3/0B4V
xcDWq5qOlLPUt2g1xSFeYw6ZN71na0Pp1kjFmNr7t4JswSMltzIt45Zj/Ufxw3Jse5gH8IN+cTPN
1MI6A8uVPl/Fw1peqSed6qVYn8L2BLTPecG00SQpaL3fc+x7bFAK2tokTwJimckHNOsZaihqfbjk
ownBv7f7g2nTAUPzjYUi6oZoS7LWONbRSltGSTToGzlG28bEtkPytiVz7sLmBo3eVUgFVfM1r2iL
4BaxWvIqm5m5jWOGC0wj0nW9ATAe7wBfmIy/EGb/puBMOOrdO1Eql01qB2R0DFUjI+ZIY3lLLKQJ
jWrZfhEDCG806EMmXxnZFqZOEkpJFpzEDQBpkxizWZVu0NZvL+X2vzn766N9coqIk+jyIiMYAK5Z
u5eE9qX1zrhClrI8ohm+m8Hkl5hMxZ2ifDdn+r6+mjE+UFomkH/cfV/LbfodGkmyI9sbyQhaf4eM
eVG3aLuAhzHkyMl2fkoWOcuIWt5rhge2wFWsu9qKkYv1bsmUsIaEqlC8uAl5LKrfru/V8jBUcy4o
+9LnQ0/wTCgF5X5Rp1ANSGFp7U4paWJMMM+zSwrmCxsyUizxAPKhVluTBtendy8MULQVGNN9S9xk
bp0g7OPl+pkECDiA6sGn5DvS917if2Uc/e7WHiMXMoU05ZWOJH/gWbR2c+j5dukShE9rzJrITjm6
3+gcWQUTTqECoZacsKLWt/w2K4kjqcr9tlVoplXT+emLpvPq3MjOFQrMz8A3h7ntwNTX9Q0W60cp
I2yjlrLbHr+W+q61vjft02IY4aK53DrVjeqGXuKNPDKOu9Z3K0bhSh8DBaDY/QIJMEFFxZ7yCdMO
ZQcKXaj5i5ZTgkf9tNbsVs7GYOCABK3KJjp910awo+pj3J8g40196fKldCYvMBPwy59oJU/q/2nl
e6xBNyNUALDjGeNU/k8vZtp1bclhmPZHm523CatXNPnomGMOhEZKaKZIkM8btmRabgbqUwoashVM
komZqyOZfCItNahLcnMrYrJGx7G6Ufrzp0bBN9nnC59mVGvR2VJDhxqZNWHvRyv/s26rT0JuizFU
oke1mIp6UkfKRv/FouJRwBfBfrfIcp4JznQQkoqYP8yFlSlGVjaby8/Z6658VSFeRtHfQ35xzL4N
1rKPrKlSGH8wLsnOIJC/M6rF1pFCXtPfFWN2oNtvT+/cQXom+/BY19TEhmZ/FzihOY/VjI+Jv/hn
0aY0ho4etOt5sU0vNb1QZMsBOdIED8Ouz5AvkXIliYs6vz8qOf7u42FZscB46+nVs5m8UZdEKPmi
csu0BxFCo7Gc36/PdluhIb5bP4zZMd2GGdC2bldAMCUPvxHvMplPc5xkf73M4LcUJQEodDwB5W9o
6LdcObI6uzdFIGEpwz05Ib5aTbt4oucUuYN+F3KS1rKO65QmWV+LOPQ1s7JAextZLAyNmaazVVlQ
T213LVfb6OQZp5DqN64BQpZXx1a5ArSem5d9aLBvRsP5hlUe/MtHsApVkX8JqIohJGArDlIJaYXN
XPmpmESBZAvOJ5nMPRt6sAPS6/SqecGWw//z+YluKggihurQ3cKoUV6vjxqU2K20CN549jGRX1p9
Q8Yazr4/OzeJJBz67Z6Dv7ipid2TVNSlFSo9ULuulYgWFKlMcncGCrBTwqxfAl4aegBehKXP2K+v
9p3Xk/KAOf3ZDtwwEYcdb693Sp7BOEuJta6wO27B3bcE1pjvFhA4ynhzaqCtWgumj0XhkOJZx3LY
NSdNM8ZMnC2YTwUVML3aZ1MXeQ2BruxOA/xCWX+6ArcCW47kBcKCzTnHKzm7yqLlO+wjUZFxCqX4
WpItxh94g6rGDNF5ch/X8CtKHpvhGzXBZsSTv0Bcnu8jyp/ZjZZ1UFKGpk3Z6ZivNFzeYt1zWWin
vkKjMy/K33jOV323GVn5ml13r78eWHJHjRRWTPXu2AVv6bjsr2Gw3MWxx+zmQP3HL7d7E+z0PTPO
w9KccfOi8NVDFsGUzNpu/Luw+lGSSII97J64uQGfM6V4TjPqtvUryBKSG5RM/MKlFtQvr/FgX8Og
5EaKAUuiSVEJjmGizRTympD4I8oBCKteUrlcaWTDQp9b11N6GOYgp+YnBF0fB0YQjzEBEHbig2y2
ik/1ctmBJjy5NsvPWHpfJWWBjLdDHlWa2h8FeXwxojJVVL2TuLXeKI2biXB7jSO52tT7zY8hV6x3
d7/UTqGIkuTlnIprXW0tZ6xQVIkflilYe7A41UbBzZeIAyLBUyZ6hZJp23X9ctGDBZRhxrHJaON0
m2h49ou3ljCLyBAZ87FrWIeAk1/ahnLHTUeYFLOFL/qpkd6EROKvKCqcsRVhKdD2xzUYGMK/DiAu
MoIZzoRvnHpSp6XW7ZOZFXh9FZm5aIDBME7ZR6+RGKfjdXzbuYTblKSP6aD5BkxE3Mkfb0YNIcbM
kLI6/rvd4s5v3M3PkwG+ErOdnbkqh9G1M0CbaIc8PycqcaKmI2P28kuk2+y23hCiyPVxTOCdXihM
jwORRa0n6lAUDP42aFUGs23/re7onQIpVjxLPATHQYyefQIjdGTkjYbGM1i5awRThMmEvdPjErMC
AUNQS1BeShRu5vgZl7ctDLk5RSh4Ukh7Lt9hu3lUPbWvREdU86qeCePvopk2f5/JtW4CbdB7FJqt
KseXh5cvIo96Mg501zz8cy5UrvED+8QmL7eYgXEnSg9lgOfAKBqHuhVXyOCyCug4QIjI/M1dYC4g
8EcB5iJyzeHtpAqj3Uka8GzjRr4ODRzC0KaQDBvaEchBFxMLrBOUXYYA+za72iGUJ1qSfJ0/HsJU
0ua//aPD9ZwXX3BPQbuyg1/BIKquN7HFZvUbY952QfcHWZZmybmkvUt3Vz6pC2cB5RxghsjlwWZ4
0Zt8O0QW0Qi1HDHO5yLTF8XXOulOJWyPDxLvTrzWlTCnqi4YoI3/zuQOmLOaVM5VSv8WJ1hwn3Nz
X8SwI9ovVGDaSk4nhyDt/FKq5nmeoDntULK63P2t7Mmf6ZumI8wDc5HKeaog9kxK+rcm0x6AR0C9
qx7ZgOps4bR/OFaWv3dEC5JIsAtSh2OdHw9oX4DV5HXQMi/TPmDeBZGfei7WH7L5uN5OxIvnqR/w
u9bbUSuVsH4U0yqWoU10kfTlLvwlM5qDbG1yv5nYx4tdwsd0k+v9sS1SHyalqPr4Jf2TQhly1fSA
VX6zrLQSAC1IqLBUl8jMpLZ9eewern+0vF/I8hbS8Xi4Fu+Sr1umwc98qN6SMdelGP2BJwWkPnd5
VfkYTiwy4N3SIhndGzi1lYDCGQPLEaomjjKFRgqd3jUxkIRS4Ovtk9jC56sGk4IZ2ynsiiBE6quG
EcxJfJyKib2vr6uZGZ/jESmiZ1gDUn2z4pyXtoT/BwoEtDbc5wt1iMh+l7hxN+Iz4SCfUPTFbNJB
XbmDpmjTcdqg0wos3nSAOrBoPTFNEHnTH6+X2kcT7Q3M13OLG07SSvsOfFjysmveu6UveiNCzfU3
l8PMegDDvFg430oeStsBcpTIhY71r+a1I1wTkLzrv1Ei8doSpDnYkH6nSdqzUA1kMbhUVbQo3CPT
mVLI16lrdoKhA1zqsY84d/EE2KTz2YZWRk8oYI+FdRBpi14xldpll+gic7tb43wYrL3GYU5RPuQp
u97hWaeNx13hhZ0Rjse0RlGMociVZ+9UdVHwAd0bjDJ7oo1Vd+/QfhrHFB5LlPk/SNIrUK7nsylC
qqvcTTNkNtAERfvqujPIV+hVldyfFvWwyXpLUL9yw9PrqBwTgVbTtxF1/Cq15fa9fyON26d3iynu
EHVeR7oAzLgwqqNKWpcMpF8J8u86arQcWZdAAZkjYOzRbxKoerbxSYk3AECgRSue0eLxwgULDPl0
DLN1clSL9RGo3XI+O0tVluxNW5bfImeK73GprDyhA6BqDT2STF50dblm5MAq/mQi/BFGSgfB5+m7
iwMkVy+y+kLN+8ceRlM/ztRJ9BtBJrTE76Bskkofm57igO9EtsgRGeItc1eWNRcEROxVaEjhInBu
jjXV2kM001dstW+6owrLyiJFKSOZn+Eoc5RGBvESpd3J3HRGzwlY4gf+esn2s14qhbKyEZl7rM4Q
1roMT/57aynXEkSF8JcroBqqlFqYbSD29GilvRHRqcygZ5tiFZmVGI5VssOZUMGW24FeCVhXVoZ0
qBDZd8fH8FN6lzLrmzIWz8EFpxNPKfqt1XI2W7HWljBE3GpM+H5fbnmteerIElC8c5DRd1TYFhsO
9zb9KV7Hf/bAk8nEb7P/1IMeUSrye7iOYXqsXd/5kHr31pe3T2K/1OJfRk0SMW/kXRt5WlQjSgR4
KH+XQEreVlS8dpdzcEq0WAHueuzOcMRfTBkQK95McukDNGskwFtXktGCk27mFwTlAXhZu8CWSf24
9oWvHxbLYDiJKMvqpqhuhV8z+GOPIBTRbvAlKgoxl84LY/Jj1vBxOBvcGds904B2hNq4Pc3cv9iE
hJK0lykMNnF9mYNRH2KiAtjD7wcJ/ObceeCv4N/h5j6idWTm7Gb0UtjS3uf1yHN6pguZUVUuA617
crEHk4NgyUrZGdNCPBrqlBz8rKaWQsbnxPkl6OP8aWdP2XHKnDFbRoleDvsZSsts57kBf9M6i2mz
iQLyFilz17vTj7CpWR8K5DNZq0J49cjw2GbW5E9bdRtnK7CdM6MItRiWxW51RHrOzq7/Aj3OEKQX
8QGk/TOrh2o+Ub3FWc8fRZI1Zm5e1E02+/8LFeJKONS9QJP6WByL8dQX0I2iBH0YnhytipRXaWdX
ZtuizQieu2w4vEOVSv6xbT5X0YbFmQxOpaJM3qZ9R9ZjOV914iV8nUKFX7tKFKM+iuNXgvPYZEhU
R75FFe/m3kXj1+wF4o3Ios7eiPIwWqPhyaC16hlmZBu/Woiijf6Ll2lcE3j5Cd+3zqNKm8cg6Aeh
dMW7rHqgqtxDaWViSlxQfmhCrV5TqobJ4yROwEKPHdrqJSrh1221J8cB10ZymZRLqlt14XJpiTN5
AWXGMBjvNs8z3MmyTEwgCMq73QWY8BfuWBbgS/k6PheHexkJQ0Qi8ZN3qs0lJoiq+nlL7PK5zCKM
fVoCJoouuN8vj58s5frnY6lLifNNOXrtS9J6+EUJ5Vey/OaE72e5WEJvJ77vtgeYyONjp2g5oAEm
M8YO63kA6HGuSzu7cQBfdSY5qazHsGd0Lt9qt+GovY83pesrwlZEp6rvHZrF4aeeL8jNgA+lRB/Z
DXBeu0AoHDlrNzNwuEUEZ7pMqeIfcnoPwJxW7ajWQaXOkyNGFZv28PlJNWdDRSahZjVeXnDpU3Q7
JB5yhsYaX6lyU5rC/NneHMXp7LPcv5IFlAxOVVqeYrQ2/Xm8TYB4jXNg4HSDDaOkXWwe50LfMvoq
KP3R1zUxfxzrRCGFUDQn9/O2BaisrOjBepnxtZBbOawFNUePOd/FEqFkXaVT02YS/l/lhgyyjpn5
vdZ2f65iXESEiuesixOqaWnLKGARidKnU6sQCNmSc08un1xZugM9N+wM68UB9Wc61fdYXjq7sesy
veJL5gT03IqkS2U5DR+2CVKaEYT66ipe0RwHeD/tM3zSOe/tvrWRQGdEwthyTJaOsmFjRQLCv6Vk
rw9J/6nR5Sr53hIzpPnFaR/53KNc59NJUI1rQ4np2mNtSZEZUjI6Up0pt3WCYmoKalvMl+XGDwgQ
geCBEVH82b+U8d/7+YM7a6gx1IEQ/F+ivjTzCq3mB3vCVwEv5eb9G6BPJC4LBTvJBujOCl2HLyjl
7yyXDw299A27Tuvc3Zh0uU+94LSvtxg7nRNvniE9O7XERduzBS1KUsDHdWkf4ecIA+daL5QLvedz
4etPLkDwI21GVlXfFRGnAXi1Ch1XsaSzNNksBA02XFi4wxL3afkQL2ivW2Q0Tzgg4dw1AFxlH/vT
DL8rwDsYqeJOlL9F6X1UTnPkRwtrQAoJwzw65UqCTYzsiV32Hs41vckAvQfsTKCdDv+8RXAr2EVO
7djbRUrmIoCUCufqHEoNsQDQR99VbDZM9YDfyIz/okH+L3zmpjqYqJwxEWYG7LgOe7krjH/sKqWm
Wf3jEwwcje+ZOfUqqnw9F6ZsNS6kK87/oAcHQpd5VelwO8tWIrbN59QpCPkTK7b+WBBPkpnc+8G3
bTU6qItqiHLug+pV1M1hYkmSARQIAsxXioRXjGKmE2yCmiRO8Hwb+TOYjJDeATrRxORx4qH6zJ3I
0aX4iuZjFAmhW7/aERcoK5g5bH/2Y5sZsRkIkH5NRIp26GcRW9Awdi7VvTpq/qnvOwjejKstMql3
daTqlXodN/D2lrVIlzmiw6q3zxp1zHSstfw2Hu2ch1NyA7cqp7NoICaSqJUftjspnfPiOXAunFOI
hYjlDkmyxmzOlSS/Lt8Mcmqw0MZcQAiDbbJd1ZipNBdHYB/HXFUBS1mw0zo88sqcM2aXFnFp/h+T
WyK+0Tv93iCcaJB08Q+2frY5MGHGbPKH0Bl0Cbq91HsJEU9WwFPo3afXsvltpSn4BOeB5F66canu
u/fT3ebR74CeZV+SSuXelXt8rco0ND/mPlbPQTsYFdAJLLidX8uM4N8coJr5dCnDGI3i3tQLpAxb
5X4U8iCct6vc5sVSvlAIJVA4B5a6xKHZ2bfJoiYiratrm0VTzYMWWzAbl6BUykt69n7814AqQOQe
kwH+r9q5Ant4EPx+JD8mQ2FEPYWaB2EzRuERFLlo3cSiAURYhiO5uMg3WJQAVqi2kVMuawEYpjQj
nAF0+p+25OZ19AEladFWVF2fQmjB+HGqlVgloY1zD3oi7717SLvfqYFGxOrjP01aq10IVzpxdaEE
ZEljZyBHbo4/amjqEB0Jmtf7M7PlVfS/MqjEw5pivKPezIPHppWrcrTS+1JNYvLmf8Dog9wKG6Ft
f1gckaAxkyb1ilS0qgF9gdbw3ljutCUS6Z2NWEo6whIILSNyzHRKbyqw/bycwwYMe5GalU+1cGs1
mwAl8wmaur4CmxJYW53SJKFscP9/31bXOkl5llSmfI3BO39V+Gyuez0RyTOxiwNyOxhfH5Yy7Wvd
QnvO2Dg9pGTbeIl2K4TXLGT36fOedxKA4+U0PnCNjfFK0EV5eSH9qqU9stFJMj0aNVMnNDKyHh7n
I/OEkbRM71BhXn5mO9fldA/3FdPBP064J6EB+KpwLXpS+///vtL8fonHp8epDP8ybEOWQpD3qzIh
yjYu+UBHHq4F1jEq5ksSUK1O4cyhg1JqA2IUDTqy147Lwr2rtV4x8C1dSyyNbLjoNRsaf/78WPE0
9yKRo2cE7WPayd/n24zw896Cc2KJhD3ne8r8K16MJ8wSyJad6tvcow3XqsazMeJ0IsOdPPtDAAGl
6YCFplKhVMY0QIrCy4qw8uTDcu1ebFhxl/bBGTcLkQF28O4+cIm/1vxM27ByXtQu/l1g1L8iS1Fq
m4Y+QaSy157HwQzm6IzdgI4RnyIT6SnTo4BUu/kYHjU15dpbGNURyRRPe5zxDc2MmQc8Vn1HU+Qh
qYJvw6+0OHoNc5GYB1Vda9m24Xt3TOUbdawj1MPhroW1QcNBmhOXs0YC9AMlOozv/aMj9LAUuLmU
3WqEj7RMtsHBH1KNXvRGv4AcrP+aYhChcNCHihvZwtnP0/OwFtx0wHek8I4SuAEZCj1Z5M2NbGUU
yor1LUEVQ6G2B1K3dLNp3s7c9k6wWTOUsB0IM2322sxOwe3g0+n8QqItIejOYPOMHGts0HTaBlTD
lEoJHcO3dtZ3HtYKXevS2t/2F+TW9ZR95iYR9RMN4cjGju1y/VEfugxAbq+zj9kx0cngM4jbX1nv
TRb44xLHJ49hIrB4H30QtQyY/FMNGdJ/cPHzWVVCypWSoaHtiQDShee2xYyPmk6cOhCxaqLwdhwy
wequiwZ1BQQDJVUGg+IVIeSbiASEcl2IDBv5WcL3LY9gY8oZBVLqoAuQQiFEYwaf1gLqIOdB5W6t
Sg9vuX7LEWIyfFG6aUcdIsb7vKwu6yKdBmdPf+y/XSsUuZ1tIe4y8luYLGJWQe2eIkjUc3ytbOop
A4YDjVoqc+7L5NF1CeX9vA5rwXpicgvaFo2iYOV3GOMqSko4sQa7ITadXkg8g95qW0RNbDhyQ3Uf
5/xLZOGTT4UCQQh6vJdA159DVT+yV4m+mtIr3fwcgKaLEQ3H5CGeRuLhpxCSBROcu5A6BkBSxphB
R10nx2nXKq/vz+r0rCmhOKOfUpZUf71nS23y1mXRWd/3aXnIKJvHMk+Xjp3LxSWGxaCemLJhmHBl
2ObXJVBNaoVDJ2D3JrlD21w5EVMMeIIKLmHsFnXk0odPgbuaVTplJ982IbEQzaAcK0UX+ReXA1yE
0xwRtRamuqk8RoT2RqaN9fLmuuL64amxcfvTrMi6ARObKhmmFZhpYrB+51EJlev+WtXfZ32wuXge
KFOtLVarqSK4tgq/6CjVWxUdx3t3xc/Fb0szX4lUUE6td0TN397Bk/Pz91Z7O/7p+KMmRNq9V707
UF345WhXWvJ64zh1yLwynFesQZ4s0u78GiAFcYdX4fmrzMPmA5sfyrhEKdsTF3tWSj50LIIvmYyS
Zb4KhMdaIQoSlj0B9pvdwYr6rizWFg7Br+slNJye5ju+1pNX+7izeoZRMDt1hsAMztjCruAHs3S2
W6AXkWRjlEeCWDLuUELdFxCFMy1uiihLd7AhaYwki7gcZSJzZ9tkCcRWMQczilo0eI8dRRIQCWOM
XiUgBZdSoDzDt2gLs/4aZDcRUFY8JOmfnKgcrix6WKLFWmdeZBWfSvA0YJ7An1XcICiaRFksmU4A
TsZFo13fWsY4ksO9C0J5BmdHgE4XMb6bS6IesGvDquLA2qJ6oGT9Pbw7NiaMuhrxZJlHgTz2TgZd
F8FNHl6pFPGdTyPN1xir81DmgZIJq7t9v50on6MtsokoBEvWtnpMbVLTJlCUoCHc+ujL93cdQFrL
yfe58YKlce73DLGs1ErgGox3av/a48QQbm21jFtJjGjZUB8cQlnwM0uME+CsWiggcHhKuedLk5ra
34IBmgUg/jwBhY8HILHbw4nTypDPZnU9eYtXUFeK4pBrn19WLwvh6gldWsvwizzgK4qqXzJLutas
5nX8f6nUxqQYYrbzii572KLg4Dg3ePbV/w1OHIdfdPSlI3oQPFPsDsSYvzbGW/bteHllUSka5ck6
/bo1mYKknw8gwojNykon7et67F4nc2ZF6esDT7nO1aELPpqT0Eqhz3Xop3oHoIt/jA8xSD0uZyKI
SeCQATcNVHyU1UefDBYcluji0Kv0Z1OIFKYay9QW2Ph008pW5hcHYpvYgZNVWppH2KHnFcDx5ZOs
uA9TdAJJ3RpJwNTgLWO7+tkxeEGhtoHVDaJpZkw9WYZHaYEtd2PETctiMzHvNMy3K3vrB1uuEAap
ohRIlrpz6cNXfFbReOozMtYtfeOHWKNQoUZvoVFfC090bK0oqs91t4dLAzIPAwe0lnyv5AnOaxo0
a4VpnPzMAs9ROo936kffIEV2izBJUhIB7HD3H3w2u5Y3PC1Z8H+aLKRL0hMGsi0nMyyUp5tpZnZS
qj6JQn6EXVHHyAHhIQ4LO5ByVQy64RWIS9tOJV65Qmx4j7NivZMKCoLF+N/17rsBoYy5RQ2kTe8e
T4KBAcjBXiBr7vlgHVliT+Mm5LuPmwGmtisO/mEaQ0myve7W7NFCdJG8E49rRf1gyMHesBCcxanM
8bm8+b0BG+J+ELnS9ooASFpX5Bh30wqnx0e0FEyMqXV7CvNvtgn8P3GFrccy6RBHAjCdBt2Iooal
zGIqs+V+Q9PbEzmTtvKhOi8HOk2PhN+GpxJ4myERvyc2AUmwnvfKS8u6ED8KVumdS3Qb81wuJsjM
pSa73RzGXH9GULQZrRHEAwnvRWKAZtlC0Nh1qrzf9UQLF+Z27wQhDz/ahU3saNJjmouPUX1QookN
KcfpnyhLM6TZFf9zhJi6fxABDquc6gee37JNqsWS2wZpcKv1wmZIFXVSIpO8761r0516qgUgpYu6
osS7vGCHT3psTwJKYBCu3EYl2iJ8ZuvHJJ3KHvyjtFDE/yrcnxU/8w/ZwxBsNCx7EH3LgqCTRlXA
Wl93v+9YHsQNDFHNCzNOg7DdgJ72pndRJROWfVzPtu8V0lje+EyBmCSHdV0wAUbrjlgoOXhnkRIN
7I8K4bzVBsnyFeg7dJmr4KJnPHtgWEc/SZvC0wprpOI1+I55PALH7kXljUhscat3StT1w6A/ihxI
aeo3sUCTTasD6hVCI9GyQQugksqrT/DjfCo7mGEiUT42HDgqfZQrB9R9g/jtRh8cOI/h02AgdapW
KQeceLdW5uRtmkdeCaRpLy+is1bqieU4EzdCLDpJi9f44T9K9NpBUNhq/5j9bfMHrFnGjzWROzXf
gw8+Np1BgP71hX6NCeWAnXMGWW5DFpUlvbPpm+8nW03ky7NHpgNBRb+6/OPAc6TYUg2RS9qvkJb9
YH0K/Vx0+nSqcMTfEZrGcE1aKnMfoV2+zO3/5kMg163VMWbiCg0B/seS4vY0ue9BSvxq3PiOCfry
rn8n75eRzNoXl+CcwZnvf0hgxHpbWMxWKr8t+1gAdTFQToxUwz9+2mb2IDPCnGi6GhAdk8w+AwDK
Z2TBK55EdrMV0iN59AOGAl4n0a1+vWxksyx/4buBOR5NGmgumAVkqYnHi6NWFeXuxal4iMPjBk2O
IDBatf4Z0k4BrcGhxD5sNRK+DYWkFha65jialqB7c0ZD4hdhgPAjPyrfTXyXIyNcgzmZ/IMPMu0m
7eGt8yN84Y2botewiH+niMolg0rkwnP5qxnVCJzO22/EWXNphJrqdtWLvcB8+/WRthV3L7Hoks4t
0dnYB0tLNMbr0679DCRCRW2Kc7WK3AnFjSdLlnq/cirJekBZlXmwOgHfYw60mxufVkgylyfkUs8i
QgD9VB00sdxGQsHjZxnTPtgz5Nfvu65305XA0x0GtMCFtA6fQKxZzq9LzwydlQC1fQYerKW6wbxd
vubWhpEQJYdMSzPe/fwDxi+P8pOzuALXTU++2ztDIufYeSVTII7pK5a+4+KrXyfuXCGA4x4ndxSz
5eHv6eD9OjWNNC4s66K9hdFvN+4z90bP3zc0t0aZWhO7AfgrCilf4dVUUSen/auoCmOxa7dWdtBS
0RJ3zb2vtmAZ5oGV5WMhkjymqZjB3Gpn/2JvpvJwwonwDU1YZsPKB8JgiVpyHZQ/dEuPrbC4H6nr
djNw3wez0xZf+XNGifCmYVJ1spaOvW086KW+bDoK1ikokgM4/XbqNl8YiFs5BP1DXy//YZqI9fy/
Kt2pl1PFF0/Jjc8FfmiKdCTzU9NCQJbF4J0EmNfeboZzhI4AduAdvQhSXUG1ugTVj09pivy+rdO/
6ztXGXtxzC24PM9svzTaDXclkdbhQRC72abm4CGLiVzZmwZ//mOhkCnisQY36PLGlbmhd/f8shtZ
jZjr6DpMi/595qO8GaXvK2H4OeJVZvZuNV1UhKDje4Fyv5IShMkApu6gcx3ziRPaWtaHnuAxBotK
fPNR1QTdkZDI3qvQneg9JkQeN92Amtw+HWbB+kSfvRY4E3v2zZh5hF520gqAk7oudTaFdFeCDCIv
QsCS4kaeY1n40sFQ5QrD0/ay5WOn2ACZdY8WxBolGtxctvGRCLfJ6iK3dfLZ+cDfMM1BDBYn886L
jMSUYMlH6baL4mXYBDftVnl8Zn01oZJsaqA0SPU8HQDepuI8UdWWKR9K0rdb7dG+ml3CGtyobsz0
yjJaDU6nUMGnmqueIYKe6yJBCL/QYDYus8PpS2Wl7e/J9UDzsGbce3epZJFIXWhGfkItu9wS3pRk
0P4OB/LrhICEc+CxLtoEJvEKnkyT7CEubRflBQk8x4Df2aUmbWrUrSeRF5z2FqaEs8Uac3fv9Xny
PsjDQiLY8GbntAGgxaCULsGIDO/qgUdbO+7+nV9qZmiAKqrMPE7pU0MiIDdJMu+55oK6LV9NUXOv
57nv6IupxDLyuZUdcxzwjWBS3EHDUzP08xARe6j9wX8HVGfjWTn0xxbvXIqzB5Vq2uUynJZy6589
OHOXzAbu1lx3g5ZB5Kjwz1atN5YghsKoCMbPF5DTzHvrwuclsIA3xh9uDHLfJgEFZ1vl2ddHjOn4
mkwkCO9XibqEDS+nRKKf0AG9c2nvPtJfDfr2Pu2lsXBsx1Cza1eS4b3jrNrhMzkWu7Y5XCPrbE3q
4I0GDgiqOvRHgdhSX0HSQwTrWyJmb1GscQ61jf+RQn8ZYWT26gw6n8JE3/xwDxQK2xT/uoF/MVHT
zNIJJtazFh1+6+eRxC8+Tvc+b6fxZgqggh936Y+juCdkEkSOm/0ILmpSgvVjwgBEqWNEYgxbPttu
J1gs2uixTqkaZ69B8snPY6NW9Reak51IuHh8vMfcdpMjd9U+bgZrpWwMehsTT0y/4T8leTwT5g5n
7HMiFSLJLtoK27vUulIB4CcDatJXNm58/91NUDmDlklcSm2R4pmcDeUR5RMcWKF4Ydtq169pDs07
6jdm+7kbY7qUS8coWfABTGpR94m4yFf88+kNKA1xAKgCPEeOsfIgXGFLtrFIUfqpsNSn5tT/qfYr
/bo4J2n7B20mOOa+6JaCS4RD3h+OhnZI+eaZuHqhng83us91zrQVy4/0MddepAOYMaq1ttSoXe7p
0/KJBoirGjTZkXeMwIBWux5TYkdvtAd7mc8cmVxeqceIxPBsNa2SkDOY6H1tFvlKrU/SJ/yCLN9X
UFo6xYh71ETVblSvPF35ftbbbX7bkCJdzcNWdYBLfDwj1k+ZKq+5NPuXHoEUO5vmVLx9hLukYsD1
6RyNDE0vvdxF9//Fl7wZjr034xdj/qBJXyqJGpy9PLP7UPoLKpfhsTmtKyMZzLIoEvuP0rR9slv9
Q/j2cx49LpQkQwr8INqnQCsrU/5kXjlJJQAkndb6vLHsuqkXFVXNxnIWXmOwu10XusYy8kLp1cLG
eXgWJayR98Z9Hs3ndYO34oHvmklXbDPKrxNf7h8L2m1EW+72VN5w8yqINEYZ6QtaJnWdtWZEyKHV
sIOoUchUG5b33jWlbtModuv8p68jy+YLes/z+5M57kGuhwnPEJ0R22A8zPCevFt2449PDNLacmK0
28nKfL8q3SBJQyObv5Wtm9EclX/zQaZVxExoiR1r1f9x9iBIPvFhikzUPiX5v/ux/BYBrBkCVDBy
SwHiuiwdqXozv7JvAFnz6lB5N2H7bBn6ztKAWFCtmFuHISl8Hwr/sQfysxVYwp797rByIAbto+LK
UDx43MMj1UJU4KDwNzRoW5DjHCPJlIjUhSTQg7/NPE8vvg8D9gnK1AQfb15yGAlvq4ZvWVBiUoCY
1Fw5HFhIee2ZHTShQR/IogKydDXZXpo3LYlMSmLOsZS0ioPNDueAEkMCUpxf6J60WsJ4/ZLAtKAn
xeaZcftc4GBUXU2G2rq6nobeOmWF/qGMN0AYYjykJ9EL9FbZaGKdnTB03WqiK/FAG7jC9co5lANu
Bm7VLTL1zhv777RMDiqInXUDAUriSVAXbk0MxFCPBefgd3EpO9imsv1m3Zvo8L+hYVTOvO/FyWeB
jxwEPyI0Gsu7CfwBXLY3OifxQXJcVNCXxUkNtdWMcQ32wy6H6JiYaT0vi7dG4K1m2KiEGuA4dWte
l08h0X610RD6i1QnaE56WFhVCSEaLRpK289BejOz+tLNvUP9Z6HTN8WY2qi7zDS6Af41iOFSaaQi
Xzj3Mb5qR02Ez3Knvvx4z51J8vy9Sp5ZA1OL5X7aFvIqvPMX7Sp0qm45OOGvI9Cf20FCUAeRYSEy
ga2Mezj5bPMdSxgs+QX+vIbpDreliSrGWNu+JjGyWKqZ3HrL53UhOmrSSAZ1Cu2f69a6YPqVQ/bq
0tDwmldULqNNxU+wYG5ACjvIKMUotkxcNdwaWKwJL1H1nY1ciWYraX0pcPYGawQ8g/ZB+VsDdncx
kNsj6J2oe7dWoDu6WmKcNo2/OI+2KIwqKX55ItErE76dQvvCZJghcM3zo9Y/eQ/9/Rg3qNHVJfWv
YfIAEvmGRu7tEaC2rfTEmY+TsuRC2D/cprWUK8V0gND+hKStThLBAg4+UX4QEnQv7G8rbsVIXHZV
7Sj+4gP3oHdB6AVQeldPrhshpJqfeo4w4wP+7mVgd4dgtjIIat8YIkdnRkJe0ggEvkEZnXoyTn9x
bJijFNjTjMKHTKaHzkQlFyVzADWZJRTxHAu1SI48A2Dluf4jU2oRdEDs54cUQ/mZa4qZCkBY6lOl
wejDT4gE6HV6uNl5arUcKsz29znHTAovGe2+u6q0MqVCtOp4FiUK1Mi1yzj8PyhEYjZrji/+V6O9
TyeO9hbfvXJvZY20zWQHRFTxszEAIsGRsBrMTDvcDnXB0twHA32nKjrR1IvfTY3oAe/myolWTNH3
M2BlvuQ5+mVGTE5mNZAV6mRxq0vL0hUb6W5TbFxGpg19S6rTAqDFE86Lb1D2viYU5LpCY7tbJTUf
mDHwHG72VmidvfmOPuIb3RSsH06QwpAc8KTIbRbxaPYSbnMTIw5QUtnIY1rbTmHO0VOjpSZvA6EW
FqgxI5uixdavd+2sCkNZgNyzz7LlzX968tNFszbPWAGTX99ILR9fZiiqlDcqISsVefVY2pOnMekU
IbEiGw8+LgIvheg71YwVop4v7kY+DC8K4rlLhtUtimXq32QOgDeNG97PHfWLw6jzxvcg4zr/eGq8
A/fJCtLOKMpTO/NUWV55M3ZSKngh3ymrrpdg3Vv+pO71KK88FggT+uEYUzZVgjmhRbAaFA1rjYuS
ZOtUWwottwgfhVnbb+bGxcRxrAqjBQq2of4yhq8j0v0OfFVVVO7NTuHh/aHUmzErzY+PjeYWC9BR
rKRTYo2uKj7OSVArYQ2cYuW/5xOYPIPd1FDXP/m1EezXS41FgS9C6BtWWCmfqSPZ9P3p7vaSGofF
S98/Yj7MhTgY3FT+7BZm8vJfNdT5c35Ga3xJmWOjfbyUilTO/qSLZVmdgwkryo1btoHJujuP+H9Q
NidAyS/4Zt3yhSuX7Ait7q3y0mkBrYxdD/xsF95t0vgV2PfZ1+Ico6Y5DOexG0FxNMWkcf5gBbJs
pOucF/agSD5kuJlfU0CacVnf2fcswp0AbQuSxNqI8PsV9hfYYz+1TIhG7DM2WtSm9W/4+L3P3H3Q
enC3tSMZ9DDGXtZTrJFU2YW+DZ8w0BrztNVdmZ9lsemMy5wZedMhXN8DVClWkvo5LJzvu1Gpete+
no71GpFFhkWwisZ4U/CmDLgNWX0p4srp80aKya0KzDsD8tP90YxZwYfzzzICkDzfavLULPmgIoib
KO63j65280XsSSkESpPeR/v1iaZfIRFfjHrR7BThduJiPOOaPrNXixrpaodhqL4uePR85fuQ7d8T
6bLAgxnpPUDXoJ8o0KGqNgdL/6LjX04xXE69P5FvxhkRmXkf67tf5pna8epT1cO5QBs1X0ElV1oo
/RUXjHHRoDFZ3yKF2B/yn6tQ2zxhEcL+FZFeT6hzTzSYO9pZqhFJM2jL0PcBGDZMMHHCY6k5nZ9M
W1zJhSb4DHjakJKVokWzG+KFha3Ye/D80Nqeg7viT1lGjSCBS6QnEyEZ1/4j0957iqlimTnxUdeZ
u65Ksazvl0JETqy+LQNRMxceICW+haSC49O+JnKlPLCow/iH0HsUqjygATE5d2zpKHKNhVsmxCjS
ETdNz/2qtIlLEPi/F7QThQegtQgoszXLTNXs7EAAO8qjdQllrWn1KRoJIMmiHHo4wKcjwGum77j1
uhSABZgjV5NQ3r+9PIwBwK1UvbCce3dVqIsMwthV+AJqYBHUMl5nUg6OrT/d4qu8SY13L/gzAQWZ
tfkFqszAfbd4P8+rWTzoIMc/0Mwhxsyt+tE4w8HI4Jcn4rCBfSqeoz0h4nOnKyB76oTm310r7gyS
QpN502hbqDRAF4VJUkhTsz45UMncjdDNhPemZ8HxR8LewEHfVaW1ehCEqoKWvxXaL7hLqjcE8X9q
IWmF2gXgFsdc6BYYtROgpTKTB+LYvHyHJi0BKmix5gVpvBSkOK/NRG24BEhbiN52h6cFCOtyN7I6
Jrc7WYmD7LgkNI5GYouWZmh/pVDKA4FN+i1VBTbBCOXYU8+lQjUVCbSIA+otJ/wEPYOHJexmu/LQ
inisRF7rxBF/DAA3HmLSpY+9FfyROO82sI5EkkeIo8T6PaN2rn1QC05sj+g+9cyaj7Owu2U86A1Q
tcfJ7FxxQLAttgPytzI1XwlduOfIENmlCsi8Os2OwWmFyGqDdH9W1sSZMeTzZ4ZVFLlIaeyMOAb+
PjbQ4N6WOFpjW+htCOvvLmUpCjlBklfh6YqqtOxEgcXB6anTjT1MwPg+d93ulVbhUo9SgrxI9TCp
/RYdq6uWp2opNN+QYjWAXpNjMkmTovVVF/nhjih0EkGEz0v1GBxUSOGcNobIF+7oL/hnJVHMltna
O/PO9npuU+xDri/RH1TDevZVizpz73HQJEt1tXyewR9WNXxvPKfzXIocpK5gIyjTc7BJko5k1v0b
0k+s8UWK5kh8GU4aixfh3/UH3NMBFDIdCL421YyQ78J/tjF5mCS7QvP+CuFua8ODg8hPOzJ9WQQz
/sgyi2pCXOMlRXCpN/cYIqamH7xaozBW+PMtOJbIWlMKHdepFKRjfA3qNG/f7NucD3Xagb2aa4PI
fn+tCxkpZszGhg0h8Yo3FRA6S5kb2ZMxzIu+Jny78WUo4O5RcEhWoi4/YlJ9HsrcmoH70JrrRRcP
9IwAXkRFeQpaBYxZ+4W/UFISkkGrRNhGcafb6lhn+rXKslLYBvhD7TgxLbdxcwRSG/Nxu3ukJ/Ki
KPo+kbbHlvZSwD46IGguiNvcgQGUJqHFsyedK9EcRq/LqstdKFKHXpEHzPqVjsdgWyOP3b4iiQl0
If8OIDCL9P1CKZD/6VDd6ugCVDtAK15khDEa0wapx4HHUkIJr7FRaDnymXduOn+jPYn5J35kXSZx
DutnFQ0PfQKj746mPQGutMXH1EwOLPBiX3MQghg5S8hGOqzTiLEXHJQdUYDYnihBHJRTpO+3EHT6
YCDNcG/114bwRdy3AdL6ZTQCL/RZHfwRhI1uaUKeBOBd20jGWO5ke99fZ8bHqACFBKE3s1kliLwn
kwq0j2HRhZZzEd3ytYnoqRTeYfwuA/wjMHk2s5H4+ilwQ4cjYbO/ftcjN1eBewxpktxGgYquAR7e
mPigv3ndTkOSHAOQyTHoUAOSYVpx7JhimYgmF5zeRoZ8FkAtfOhmzWge4hNawao13sE4zwQJZNsZ
PmtMnPL/huqeQWHT3BggFI22qCwWNTqh+W7ytC8/qS8BX958NmOj6lD09Z/JOWbLZ2DqDbUOEvfi
Rz1k0rT4Hbnp8l5bdgn1YWcwYYmZLIQlC20mo8WYxPvEDLZyq3iuImUAkjFF1LNP4Qwj7KuwAcEL
/JzFV6nGbUVVpAKVRf6zuSmzhJq6cdZNUSVJDF8/JrDl4V6QuQ+qWDCsKIlaes/svYSqgo/jA5VS
JkLc0IlK7Ez2vFjYtYTqvmmxWcUmaJOlfmHHdp1rtMYWHnPExSN1P8zpJtgwKcJqDlab8fHjCmcT
UnxAo+gw7YQoZHWPAtKRsLsPAYLtPSLffdXx1GK8DaM5HO/Lzv0w4tgqjEsnrFoybiBC6aAz12R6
TnSokusVBRt6lGDBF43Y+NvsWx9rjoV3VNTUD29PjfAyg8TRuM08FNG2VQxjJa3RZ6wezBRLyuuV
BkcHRl5iYulu0B3ubZ6ky4ThXge2ufSW1Ror3ZDNc50KWRb4HZtu14SxtzrOp5PELz1czg+KuS+T
PuffsZq25GvLvhKqEwJEfQ16zmCQSilV3ttLlrRVeZ90Az7QQCmgC0yFfalcHhGKdGW43oqv0La5
MvPT2ThyqZhBgm4fAUqbwyt20rlJb0VstsJ0nFLF5dEOS0o0iVakcOX0RLHgRLgMDWYs9rOTEAwp
BKnGsMgmKBed8WwRwgBjTwf+aCmd+E8HqfjKuNjUOWSSs1l/ZXbUX5xrNo5MSHjfxWJGw9gMTxrJ
pMSxgia2SbDyABfhbSBF173fPMrkITe26ECTA+9G6MCp5EGziuis6DJix79TYbZttj1JLhpwa5uG
Tidaz9zkUjmr/0cllacR8v2i+uCp/HS6cIfM/2k/7V1k58g/tVOjk8AAam3UkN78B8tzNVrqH2Hj
c93bbw4sQRIoPHMHM+giI7JgK2UER+UgxNo71IrbQiG/4BIl3q+siqe0EuCiE/cICaMReAh42kzS
RGdto9N8TKnirzfJNt6ssLkaAQ0S64UxOHKEFx8MT/krX+TEOFNWMDgPBZ3WdINjW9ajHbdAwG4+
7l+sqjgZxZ6EtemMovndxFIk+DxgtThUzQ9fh2peNn0FUd3Z2OSv7OUTh0FtSrcmI4LvPwG8QvgE
7YIFSJJ/7D+VrrOXP7xc53uuPse/veAeYtdlgb47r6f3R8jGKj6CupwZnnlFd6pk93I9MSYLpgqF
G+ME5HiEqYGUWM9oQRrHjoenZeB6FbMfqzNdzIGbvqz9ZBeWd5bc6LclpHePvA0TWDsRB9L4lH2O
kkIEzBuC+zhdHOoNWhmE4aEK1WR+pTaDFsS79N97k6L6mYHbfA4M9Nmuoml25Q0A35bf/tfWQ2fZ
XsjHxs8pIRkDYMmManejwgMS0oo4vmcvIckxDsSXsQvZd3XCy6HyGbzMJpcoBK4yDI3/iPQ3Uxv6
cylH58Ss4YTum654tzifmrYQ8i1zU2SN8JwrHGnWRtaJufcv1BYrwNQeyhBNfFr8GkXCLAOUc6Ru
qB7Dbl70Yub3Tv7int1VSAu4ydWZSIomCI7YrWxZjh4RYpcrw0VCazHOsJpO/0Z9tLxs0/uEee4u
Vu3f0GGO6OObYhQ9gP/1lSvO+SgfP2l1J3ZY+iZVP3pSK9nPAQFztZfffmmPEL+R49OZA+VFxBpT
yDzb6zsz4JXdFvu6DDjBLbbRiXkyy71N9mKZApgnmeNonFQIfDza9TPkyEbI8nBgkVB5m2MalkgL
p8ufAZMgTU4ZusBHLraedMuieqWJqrtbPvI/0BmIebHSfzYkTPHwEGMAQuB1g8BR4y+mw6dynYyA
FbTuxqLQ1iD018nkDk5ufpPQRNH0jXsYvVrlt+incqinro3LN3TV2YkOQ9j1MlBGY+q1eXAB4AiQ
VlQmIXJloolNTE2u9w3NDAAkGucvM6EzMCTLywSKvW7xrvZdhVlmzjZwph5jCYnKiUfuCL22B8Xe
G+QrvLuxq0bVPPRawg1rkuTgV+GDrxA1RFD2JEK/wCBm7OXu+l6jLNh1owaEc0cXGsnRwRS3eBW1
phja7QExJvqHUfMBWqwd5HBlrpo+HXqX04za0JNkLxuQXd2yxL4J1TsJ3NQHTdRJyVs3VYgexlwg
4BO3+LDYkpdRYcgHLqXCo8PltLnOba6StpoJFkncLNwQ+xTLJJ1M40X+4zDMmiLKFJuYwrHDzcex
01ajxnvkCoHjq1sC9LYcW/in3QlWY8sk6oZvTEfVLD2Hi1KWz4QTyDOHPUagDMk41/i8ZLqkAhkQ
/6GWkNQDqX75jOEPQaNoiGrMGz+JSPJc1+HpHKwuN9HJ9vIwssXFjVSj5mQuXqgKbOnyzo9TUMMm
ATJ6tU2HK5cl4eDZXdXDuqEFww2mSR3gGtwhws3LBR4qGnQ8O5bBFbDZT/ZcouaCbXWz2lnBVy2W
Idth4RIUstWbskigDGNoV8enNRmt5WEY04LdVtcTz4Aq6NlNvetnHi+mFx4oBLDjYvIAdnV6zQRG
6yZHVTAByBytvFwmy/oiIQo0Y5A+uv8RU3SV6uwH1+EWUwhvCTpcuNyVvj8nRWA6jhHsDeIbS5hb
5NwI9D2gqcB2XGNyySq57jB4dUa9szBWs6+mkdtNXppHGq5IGNA43ot22OkcxJsy9RvD7YwTKkW+
iS7359IU+2IvvK/kjDJDa41oR01c3wt1GzR283kwZu4ApySTyyFdKjQqvBznQ3Dv5u/f6UJUv61a
6tZG+0lfF6yI3Xkl1VtkUiK1O7UFvXlToA6yi1gisbJau+D8hJVrNXMiHwDxjJw6Eh42/sHewfNn
namT2KilhjUjk41YkVNgFawV/+1fFn7yZXvEo0C68HxU6Wg2AceA6tLVLZo1xVNEYBw4utbaP3lC
Q5GEiiqI9IUW7dDjdp+leQ0Mit8O0Hq1AYo+GBO73hDCLIb3gSMcEDrF4fSal0wrGRqYroNsV7jU
qqikIJoxXPYcXSorSL+Aep0waLC5mhEvnyGqOjt9mj/BT2zodFZyQYB3ddev5AeYHek+i5U9Rx2/
AQxmZOVOAVsSm7nXQSWRAId3THIEOskD95Cr6i4myfn3/i4skCwIkYRKCQxu28AZWPxjqTRwOIzE
r8DbzxSVbf31haypstPYnl0qEy+z96mfUpWqLz9P4yR6521pQtBj9l+mr1cgye69ud9VGGh9TKfB
kQ0+jdMQfSGsACl7A4FPLat1wo//SovoAWSySsRRKqeG1dQK0baAjpK0a2okfPbNuH5AMirJQUSL
ScVK/bOztO3e1TZBAvGC0mPbk5YDKzHYFVOwzl7O9yjWUbYxb0ZoXSl+8TkLnKFult4J7P4rCfi2
fPzANh35IUYN/vSKxtw6Pv6c01TOgU0T3I/92zWdFSJEAxmGczrp0W3VZ8EkRtz9o5Vb7nEmYdd7
mnfeA9DqVWmPu1+CEY0/pySXSkV3B0o/YofZabgSY57X7L7bfxfwdksUPbBf8AeVswSsJ4rSmdi+
nqNSm+5CuzB9em+PKgRFy/53001v88VY/hiCFRfNEZtygZi695C5jvrMTBAEy3JekUljqDGdNywT
8NQG/ltvBKrNzXxKNpqyzJ55IWMiqEeHDH0AL00Yj6/85NAa3oGsM9JgG+dP2wlpqnQOkimYpNYG
F1T2fh1zIMpqM6IE2k2xGSkDOs8jo+OROgqUyBu1Zedj3QpYKlGDKTvUPu6uawpqXqPXhNJKmPe4
UvwyWebJDq7fTlfsyOv2eshmmD2QoVKNx2hU+Jhc9U2UWzkQU4ncuMGzPsQ/taljdtk+MeCOCD/L
o3h0j19CA1DzJ3dtWR5sy+9GCOHudD2b7eqX+IwNT/UaaTupLJ/Wce5EcQ1n0/DQMmP60Zw7R72D
aDg/cmIjiF5P+BS/QsE7N36vbHZRT870JW5br3hgW4xA+IrSDHBlgSUZD/Ci4XPeml8tMwTmOAJs
FneqBFi34wCcoGviwMFRlXFGsvwwFEbjhIFgCtD0uTRms0PfJTrn8FoDnkPUxO3+Oq/4kjO9ROiS
GgOHY6OnwnsUDxoHjPjJzwdfxrTCu9eiuyuoBKLfqeZ4O5m8JsPkkGJjJmzAa5QVK5yTNGLUU5MF
82EQ9OX0WSRHDt/XteVb1ZMvIvLoZgW6j2TJtiojnnMKE52ZmoKlXZr/gxZkXRqSl1PeK+uYhn2F
q/f98UhOtlRk8mrCq53/6Rg4E4IP4SC4qXysRiYDx6CFE24xGcAfz9ML3MBkngCKDl7qG0nR1fpp
WM2PNDrjmLnu/mjJMj5yKR3FyAVpdWdL1ZD0iP1vFCmpUrFUC+TrosNz/AKECd73ZBGKVVskgQdv
ku+/Inoub6HeKsDhBMUfpStNybPnmp+wQoslhLGTJmImGC4RY0Fs2r1Ao0CoCU+aZ2iddSh7+9y4
BPkQx7mVsMym3crjfov0nCq0sp1/ALye3xkqxLBthTEqUFd/ZDCPr5dzKM12qBc8QIk7lQDCcZvA
NIWtLl+ftsV2BQxL+qE9vcGojX/J0b4/Vg7ILnd3tyueGJ0Axk3IK4CmbLeXBRETvA6NPOKJyohX
OHYsgJS12/tBLy0C6wo1CMZrv3Oryk9zOq0PnLT1QcS3uJnkle3D1eC6UBuUlbT/M888JGjeye7o
qgTkt1uJ/Wl2mruO9yNyQQCC7vT+SXeSzP5vbKPnjtPDZE/x0RomuE15ZIOeYv91JK2QALNLmsyV
d3t+StA/REMmmLot0uHpyniOvXDaxhHoq3KeQd+BEofSZwDVehrjAMP5/F/EunC+62h5oDk/LozC
pz9eeNV0lmzlKg/B3+WjeQadSeDGoZ981bekAjeTkbCd+PJprrszE6VTVO8luVjQ/EA+UamRRcSZ
tgoZLOzdOGh2sHtf9Cgh7Dp4ttquePEUIBnwPi5DF2sR9R/YgDfphC0xWH4YlNFN/1wkbnEtZ2Md
r2zM4vHsm5zC10eh11plw8X9lYjY0f3/lTKUa0EhtbbJcsK8VjxCycgSuZE8QaBzBbMecRRdIUVK
TtUdPD/qRTN8SbCqAE7iYi4yScWnRCbEfuaalJmgQ17LiRFKNK6V3/OywX6XnLQ/KzAZl4+9lEHw
abLuXvp/o5owqOyaepQhVsHFi/1lSUST1+itWKjom4ZQVNQROj4RlEqlLF6Yf+vmINuPthUvkx2/
9azx6Jz1FwbCUqiskmtPP9E11KdBikATS3UPLVZwoD3/x+W2PZuqVo1Lt3ORc9elYJFN5hWQpdXv
vtlH19owU7coT8jdV8wXNCSZPD3ebUpkknK4rR60hJ5skYe8gmu4T+50pOWyXsxb3uio2bstMz0l
AV+/Boz1v9F5P2h0C4mUGwnrWXqxF1YLTDyM0g9+14jwJWcoQV1DQdxJ6H/81qZF1xBKTX1Y2zIM
b8qqr6uqAXrAXs+8zyP3GtkuxC2w+FF/8jRJ8ajFsQ1kvdot+VPjpGB8/mzVTInudAv5F2IaBZ0D
4NFGVvlxTScyxk2C8kumzoWWF0mtMogiqnmjhPqeHTXAtiu4rZKWF1x78SD3fFTjIO4l9Zggsbcw
uSFsIeQ9AtysVAR/TeJjNh8sx94yjkScrOV350PABFdXFSp7R7PYZTmEE7PfB1d/FaZFzskOqLb+
L/NHEkz7s0zM2qYtNbGIi9hhffsDjyPbO8Tq7Q/DASMg2J+Jd0tQSDZY5k/Of301YTrxX+J4PUBp
a2gQqNjeRCCQDwtFwIPuMFnBf0hoGD4Hr2SpMTrZrjtAFFHTuRm9LV1BTOJd9Go9dBCINSA09S9B
GMbWuUy6yOClaYpRbSBjC5ECvQQY1W6PCfPj64NwrxEppsupH4VQRHwihSsD8YyZZ6LVFWrEY9oX
OZ1ZNkWlbuEOGoa7kHrgdXTK22Er4Zg4JuOA6jY9yo2zgCQT+Xm2hvBB8LcZB56kO/9MN335drmM
MPYW0Xw8/Vetlhdt14/G/2HaOnzCP5jUjEeay9ANV9D8bkHOIjY90Z7PWq9bMdaFnFt0MFeO4xCu
XkpJWF9y00xwq8Oh96P0jTNuJ1RAf85ActYflP1nCNqt6ttAGkKIZqm2GpDp02/oX3CRNb9LaGKr
Hnkt6pwDwDfbBXUrEl7sIOPwyQx6hc10Q/FJaYwifTLZPg3syWXCFiitB8b810H0w9Xgm7Vd8q6x
nCF0kA/jRGxC34dM7qqlvgu/hfRlT2uUDTk5+jQHjClhW47c8YbarG7zN3V2PSEGmSDKhkz232gk
6nDmwWpXLEbsnRrcDm3eQXNN4NDT9O1VK/czmpsM0zBaJdY0m/sqfAfGOnq7kEsOMVpPEojXYNzJ
qFf8xMcZ96AjqPv9f4yfb3NtyyWwJr0K6HPmhB9QWBthHrUcwWGWzB/McV0FAo2o4aJ4GFjJnCsO
9+Baomq98ccLagzeMMQdni5rJ4XxsHvAkJUhcMP6uo93DTSxw/0UVKsachkKwG+OW9Lei7XEftBs
i22UOCSX4ikvf8bybRf/t49Vj2J4jsFF7RBGGI85IpU0DNGnHrLtDRjGzUXZXB7p6hz6EMMVOiTh
W385IDbg7Btcb9gBmfPpOa4SpxvECIPrlx1q87rvsv0nmcFzozT2b8d4J9eEsxwhdJ2dYuDAzOMO
ZQGOBGZbyxaOlnVmSKCBErOWinCeUVIdrnt2zYYzFXBSppV6PC/T9JDRVyO54HGNiaQp7OrpJYjr
UdyhnIyArxTEh5/eO/3Khg/1Lp1YzADRBKPYEdE9dsjQ4OKZQ6UYOo54+1m7mhQTAW5YykYcXlpe
HO0MtTyUdQtPXj6jBsrb+Q7bV10FTzgxVCaBQTXjcX5ll18Hr+Ss63FlijYPZhTmU1JeJQOunqI2
rcwAADVf4IQ34LnSHJxc8f6qaFxIqYxmkGUo1pyztBJXyucf09abgoFR29uWQBhkkNI21/bITqtY
XJMlubqeN46GMdj0p6TrguW14OVLumn77J7TzqDEa+q/zASGxi0RTSt78yFjnM0JbpwGgMPJ6HPF
EBlVQG8xQwsDHLpmBzXo39g0V0p5Sw3V6qS2Vr+jdEjwCHoeFNN/HBD7KE4FcNC8nYxwOscFI2IW
Zae7EeAuX+6EykDsgmvBfEVfRa9qpZj0dqi8scXT+PO2qSjBKvgth6rQGsK6Okq7UbzVh3Ldlqvb
WVRG+lVu0EpZImY+QpFdK6v7pizchayMkdUW5Dsl+IqEwhC3TkS25WvkywhqOlUjxPy1HNyCgTYO
oEMw+aslTIrLXHuB4xDCc/4sbkhERI/MlhqQE3RYulTD/whiLE/F7dYxBDMAok6iCeqJW7arxT6K
h+cNPn+LqB7leclbVT9ft35ybpCAHtEDcWHHX/QRhmiUswNTptrUY0AcKUjuRM597pgxrxAVuVKt
v2ySNH9NSe1y3oCMbqvx/o61o2/RvhJcWPMlDk7HDpHxzUI3dyH2fAc4eQPypdFQFwVRf/sfdKQi
U1GAs6Lt8xg1LYZjz67nhT7aSRc2dVqaSppiO7fnzs7JmXFALhOHzWffjSu1n7u7QYwes7fgAUK2
Fpuo/XNRqgjgIKObtLi2WmMOHjjO2Lgh8OyNnv3Alq7fnzod8GRw1kwjwm/BuFJZazpRi2n+fpvB
je3mCSOIp6ataM2G2Xzifal3TRgUfZR7lMVf1M76+z/4E5tnIBDLeyCcPiFRKZ5XS9B62gmlsUjU
BT4GoYVEnq30NRLMp7q58jA7X+4SVOBRVWw/UioR3yl7u6FKwHYiClFiqlbwZuIeoVxpOVOcxZeK
OvKY8cqFbBu5psanrUi/TxGwIm2U5nJ1CQirAVhjRbErP+4clswRfp5oe7mKfMHoMvdFMuI0YfQ2
6gGrvUVITtSB9aT+lVt3CAxixt+oQrUOwxWR1xk2BcDRR/0JPlNscTRbR2wHnXcHZC1IeKnpeyFk
Nf9VT8PqowmOIIQWBDgXflX/G1+jKl35UHOlHckInxRbfG4NfII9V4fi1uHtrqIxaXrZlrfIlWnI
fjjMZsjJuXpQRLWLPyMkLIeV0Muf7jD5WI0bIcJATptf4B7cLAU66YYVUvRt02y8gSsPMWVrAOu2
pVb2R7PD39yxr3UQmDEAGLsZUEqg6Hp6pDL/lFT+tPxrrvWVVSkVftb0Q2g5ZgvxSghWJc0Hq1DG
VpUVXGFMJDGluEj0UxGHXR2fBtme7c7sTK3hq2bgmMjYaWdKDavwKD5Z4KWwag8OrWVjYuoeZvjk
qUyzeSC72TvRKAV/5MZWddhbZUKcCE3RlXgolmCA/3c6UNUUr+5pvQo7DTIWyCnJiTY+gmp0G2Bn
N7bBY1zylnWNOKM2tVyuVVqtvEnATKR9PijIdgpmrNBi082Igm7B7zZtYTk3bh5mefRHgyB/GvWU
gaYjIrLoxsepw+7aiFxFOW3QqzaWBnsxAw7fywsbGh+gHBML3pOR45sdalMp+ToBPoquAS2EeEB6
aghoxwaIJO7dOeHVrlGg3ZVWPar4ZZAXXVYzlAvFGgWpHh1sHBOBK8opnJbMsEF57uKO/SJUbye+
t0mKnlaaQmAmlH75nqgBttnnxgjh9DTjqu0HLC/SUKNFVj3GD/dokR93A0Qr+WsgIpbKEJfUzDzj
H0De3kmRb6m9WSoWD/hsxtWTGHN89EFvmIefzlSHuS4/gGhahV8VnkY+ckkAR3WKhKkK9YccbJWF
qWji9CNryRIOjb6WodyAnhWrdnPgzZR+o+nAu/ZXvnpZW1++OAdog1PgcClKN5AtC2fBakS6oGiw
D/wihoJLhXeLbLz5TQo2tJtzCeyyzv9n5EecFWvRMjrAw1QcqQmGkyLt0QSS2n0U4QHkGKeYdMXh
aNmm/gebcxiU8XQO1D9CKU/qwuB2+/7wZq7WVszxvGJeqAUYeX2cRrBh6IU5s/MTD3heOmhjBoPv
MBEquP+kpi6hOpUgaKnlW8AY4j9kdBQN8iggSHbILFLVQHkovjRCdDwBf8no7eh7isMD1LWpezKs
ygMxijOOL/9FxSfjg6Kcm2yFTEWKDaf/2YiAqZboaldLe3K9OiAzNXrUpIxeeheJc0teDVzyyato
RH1tDGn2qiZu5/xgedTTdsOetkjsvJ86txDQVuP8+MDGt6zU8h0kFAYN9Z6FDVW3ylXWTpwrdt0w
nw5m/l6wkZ6A+xZuqyG2LvJJn3FuC8314Ux4RNnC6AjOGNd4CBD1Bfde6GwV6UsQeSifk35spsx2
k6+erof1MpLz/ewXKvBSM4jHWUYL9qVHBTA3mQha0hvSCe7j/mOVh/ODT2o25TIPJPvDT458jUhB
RED4ScVuy/hYF1NvunTTLxM6t2qfpRI0kGRiIp0UoHq+kRE+TZfFOqKB/KodG/w+pcCswPojvB9b
Oc8w18APIyO9hn5dlYckd/YQOCO+1AAK0jRjnfz+O3iba3DNo9eM45MMqXYc2TXycMLIrrtm1gkX
r+fAncatG7OfDb51r6mJ0nug2sVzhfM2Va7G8BURb/84kUy2z41OqCgIny1x7adluk4HVe7hdo+8
hddWWKPkQLq7uZ31OzV6hHs1s7VGKjArG79nhJUPY97oQaiE4DYuv63laAsKSL3eeo7dRDwQOSMX
xKANLfMxOJ89S6EnvyYjwTuwlj46tjls5U/coyGJkjsqC5bjn5E96nlQclw6/VDwR1keOs6fKmc9
ucgGfLBvAb24kkuJZkxNuC8d7k9me0kSnIpR0QMUG2giCTdDAIKglKEG4Oed5Lb0Ee6v41Nd7V4m
HKQfQULxLP33ESMfsVhFPOwXUDx0B9PaaMFn3SbjInQxfv6NuhBZw35w4GEaPjmCLpCSV9cjG3vt
zrVZUQi7WhHWZkU00mLgVJFcXvBwO1HavoVnUp/l2H7HM3vfbQ6p27+MFWJQEEIw0c+HrS8LHONH
q2H0Rp0sA3lcyuOTKtfD/IFP1TWZ6u8LNbd8mttGEVXybqBmZmx0wCFPHbNB4+tjoTFxc08Vgtze
W5Su1Lj7UnAWVZkNz5bE4UAV37erDH/h6NjliQ/nAyKoQz14QwDm8JhYYRV8PrS1lzvCoNBQGXeg
Z2Z1GuvmIFm9CUP2WsQlEIus3qUAsRJfQnhpspURXbVR75TjO1WI1nqW9+HF7ITRbVV4iPONLwTM
o1FVSn8M6aAbwDQ71uXnLG699k3ABUvcp47D/fBCdDWSEVKolL2LNZqLtpSzc4OqrOHX80rTw794
+z4MkM3xAyQ99vLF6EdlwgDPRt8RVVTDgyhsDfHL8wAErfWD1sR9nq2cGb0+T8SVAVpLkyhyVjSt
2uPcWNqVsQulZK8VN8NNZxDSxRsMaq6T/tMI7dki5SFHfX78WfBuLbsIWVqk9c9e9wlfSKUEaXpm
xSvISS+k1mHzJe5j7kJGAH9Fltt4fDzuIUqZ8TxUsGelqUhrhdyQXUV4Hhn3SyJPo6GFftfEnJRT
kHfTvVZNI34nC1Y+yhq9M5BvqgWvUI952foM3MjSPxhnl60qg6n2VGL6DxLLV/b+BeDYebvjN2g5
YDHpmRkriFyUEJoAV2cy/cy8TAm9Ppd3ip6Yk2LrVK3W1ZBSRYBr3ybodZ6bekbqzgCtYlfWSX3v
qqUDxO89toxCh9kqdmkDbzDot8OAQkd/MxtixDIM3UQuqB47ATRr5mra4ob+Ft7l3SyFxiaBN5lM
gjQy0vRqXqZ/nr+VpRzZ5+hlSj6Qb94fNS6sRX8+845RdQC9WitC6vOHzdLo7Vzkcwl5DdbIakdZ
mVtdxkr8jhcXGVlwk5wh2apvDEmd2q2alBFHDWTUctWbdfFgEt/xNYQn8Mzz4fWxdpZe4okozO9E
X1iQbxipCKPpWH6y8juTMOZXPJicrcftwZR8Uxliu9JN0ub9e6tTQ8sRh1uWFXg4LdT+lNnIfh75
Qu8qsPOA9OpDlEkTVbv4MY3Bzv7+GpltRM4PV8HwI3frxXF+mv8mjR8TY3QhcGgweckd72HS98u+
wwcFhAHikxv7BiAA7qfW/g9evPZlIXiabUE5DOt/cVnudzlQmwmIijBHOPOqnWZnHRqOYlixiFAB
5HHrC6uMreJYG3wFCLcG6o4hDr/q5qeOXHW6mDsUA/8E9Em4uqEIiYQyMXzFctNrBCZ8cwm3/HvR
wDn677w3ZZH/O5GJ+XEsagJOr/x1qzSBHVYi8NjEpKvso5lfzYMuM/gRrOzsj6BlNhIlH1IHCwa+
unTHvsZ45M8g9t3G0nJnnFEa6fl4R+k9V7iY0EXzudZVx94wWOUwV0MK/gcyldoo1uXRhs5yWwYA
ZcsxZoYkTkLXbA11BkFJAIuiR1d/hIxs+5TCSxfwJcoSY/dq3K9nShxCJ8KQFuBgTJJWoH7ggOyo
eKaXoQDnOdZw+4JHh0VrfpbXHzXt/UYCTjU530SLuDDSJE24+UgXJz2vLZj+E/L6T08nNuYb7p7P
qZ9KMoT03HmL06VzTApLFlJOHtUeNckbQ0urmr5TR1RbwjfqLll0MT9eqHY5u5aabtxgOG0xIkLr
Zht1c29HSkcPpGmwJV0y3bV4/7yu23xfuIieeEYzFb0vcF8be2Gj5S95VhItcyDx/C/X5z8OOgz/
XRSo6aOMaUJ3jdWzpqoo571iNHvELmV0SWHOIpbPW/cWlC2/EFU9D0ijAmsfYMiKgjEW0nbbhI0E
inZ8Qf8VB6NCUd8HuZ7iSDJ5M3MXLdJP5sJamlLmInzm6fnlb4a/tKaUttCCnFhg/WO7httnRsvf
lPc8fHVLeGtaqFRSiRsKmoU62rIVY+TnfZaFfgFEG206ke2eNHcXdkNBA1w/89yskAQWQQPEflyO
OQti3Lf+EsNU6Y/vuyPwGlPF33K5hcctYeLoa74xtfvSyT8LXafv836Te9tHBYFWX9BLFcJsGXIj
Y9REK487ndvxEXlZspRfztd1eJ5243O+Hzl2997H6J7xzYu1GaP0Av2jZ1yhs9WdhQMkAiFyxLZZ
C5sQt1BWfgekp86lj/aVQfqypLwfElUOa9/ZblKrPUDv1OsipGtLIOnVuJd4Pug1QuSJ3QGfDpcZ
bPHYXyRnWEOkKpNOfDddRfQVHECkou/f+Ihlpoxbq6gfIhQyGgdwKOvvT9hCQjKvwJabJM9CAWtB
Kekz71pHWIiqRjSyFJ1ptQVS7mNKom93TRcQ/Te394F/HGVw2t92z49KZCR8GQ2adKJelvSqhGfL
8T3ji27xtZi0ORpPBKooWBPU8y4IZlHPYEQuFiA8a05wMfpC8XuLyvjnpQp3VhIZwW51KW1lO+c5
0JHjvXHOgwYqzN/koyJGnxNzQNhD4B/cBYEj4IgzoGKVNnVezL9gDSgvVCRz7gCdfTcP5ib72Hk3
qBw4uT8SqP8XxajHJ/TGcqQUPFAfyq+KIvpAOAVW0Ge+usBhTQVlQc+dRYE1hLDXIfkBxtjMraAR
j2weD8SC2yohO/uB2MzwKuONqlmTl7O39g1ltUvcxewZJmKCqv2KUDW8C7SW0Zn41tnMlvCoAZT+
489JOSWSCExukUVIhtspPy0yT23L+nkrqKffCFQqHWQy3PBicfZUQgbunQzqUnMAuhj63BrtO90U
FpxfWa4h1Zcpi1P+IL2ERunLCJg214R3FL13v82N7zXGBunpy02I5ZShXNGuXHV/6Qh8wmqu4aow
JJ3tiF69rgIE0l2YlLKnhIxrJFCYuGtzXm3ZddtQ8PGySK9N/0vO/x+b5BQxhixSsH7pejq36CiW
asCZ5lT/meD/MxJky+I6nKP1ZwNDT28NkA5HiUQHR3TnG+UIhpVACd6Rgqv+t6VCoQEHw5Wg6AeQ
sGjzB53YZ07JPqCmY1vPEp64Qr/215dEOAECDSsPT56cMJcnvi+Uj+vL9X5w0Rd8ilT2lrRiXQpk
jc7Ur17Ok8t/VcKpZKThGISmpSLpnmITiq6sTUgh3QavqwRv8U6XA/BlbB06DunL2rZ0d9BcuH/5
W4DCxjPq53z28DIm6w1PbAZIBrKXud3pGTkE3sZeTdokCBiSHis2w0rO9KVOK92SaFrvWnDPWUdw
c5ZXjYcU10Fv1P2wXPa7OItsJnYIZHIE/r3t0YSlFlrtgy8tDSM70DNXKjJHifbUDUJwpQFN0pHM
gJ/LYix0wmOHj4MPBhs/b4zN8jmlJDGNZ+hFh6dbUvxuZfudJdc23+2t2YBbvGMkqSYq+GPBGLJ7
cRZknrpIWp0RrSNF7npD8svUBFy6ZhwzCcHiK1/kT3G83P1+lm9PEHd6mA4nn1FunqAqpAy+07+8
UJXfxubVGIYPYeyEbGiDS+YLKS08nVg+w8Dccp/Svc4t9Gw9oxDETbAwqCmuXl1GnlPVz23WmF/C
5NwEo0XsfX7yFe1JdSEl7uq77KZ2sqp4kmdtnkMQlITD2OF0Bdp2We1Z55f1nHuGzltCEJ48NVSr
iL8ilws+Vsooa6Mc7iAUmBbfMxax0/QQ4crvzHx1fzN+lWDxp6zojbvTYrs5cHmjFTGg91WSc760
WfsBSHBD9CFGQ3IIuSNGL5wXk+ALuz96hIkH0PiG7pv18Q/WiniCee9CtZPb0crQ3phxzy2jYjhI
5Nizh13etiPIf/8DELnBC4zg3LXnTgnZ4Ji+PdXiKzNAAMC8aBeWByp+XW4OFJanBYfQ6eSUKkpa
1oabfMizie4RJqL/qoAsQw4uhT0XHNgsVgHzT7663Ox4hN3e3Ie/NMZ6PpnzIyve3JSMl5mKV8yT
h/1/+TZvNhuSWDI4+xbGtzau/5UhczbNCViJAIcsWwInHkESEBLB4luN2IDnBmyCDYLUSyCytS10
vCenNc8QddaiiN6mZUXEEjWE8aMnBz2aWEKXmYnH81jUnvanFLbK1WY1fPw0DPvEE6cbqiV9pXhV
sfpQU64KHFE2f7bGq00JKa1uNj+XdmhpHtPekuIXXmDIxV9sdp0Iiho8+YG9H28riLJsQj0IkQkC
vrAzFUU8FjJqvbgJG8wwWdFW8FFBeP4XDlRtjrcFZ3JlHQGs6aRcyGPFFC31gzhOhnF7UthBYLWP
m2wawdJpuDkFV4PZGAPxB0J2/8uJLRgshtDOhqlzsS0F1/3dqzIdjtcj+had71d99/ip1t+fg9Mq
xsamATu9ry93x08aZb/m/JyrwAeHdDBGY1VcAkJ4X3Tn9rnGYw30F6uPuEn7goLEQCIUhjmP8O9P
y12k8UyeO3Fgg3628j2bHZ459IMvRf4ouJozmU8RCrk+32ouuR5XPAmdZbxw1Fshjx/klhY+1OAy
kdtYAaBYqHXtbXoabHemx+1C9SyB3qy1IOswTh6nst50hHFaMwVqqP0z4QSPpS1EiqgWJAeEiS1q
qUqHUD2vGYhZF9dsztylmpO4hhfNlWqOV04CR1+U7NmPks2Hr++iP7XuBzrNBVPaPalt7blxsxX3
Ay4PjRur9DvUgqxY2rHfSdDoEdIBWZ2yIqr5JqB1js3lzoIg1k241P8cDAICyGHaQlLx328Bbbz5
AoN37pxuRpNAoHfY1JTUy0otvs80jPQjM3FbQdEipI55ULQOddZh1vtKCbouw77RN4jaPOGCrPBn
azqyCt9uoF1tIsZBpbDEXdJ5l0cNmnm6FuKeEIG+FDhSgPy2GWO+Lg9GHd41z/LsXBN4PulECm3A
+pQ3dB9Mem3gtv9N6nTaIXJnd4RAw+7n6PWMZ6aGv9Fr52TAOn6c56HmwE1rk3U/tKP76L132D46
qHIdB0V5qAYKQLoHZg4xy/v4A1xqy28LZQb0fFFw2Kd4nltATEk5wDaxJorKvYAR63RfFf0DKKUd
Y0s/7p9Dy/fj3qpT/bZHZ9fb4kuebU6Xv0vCnP4d1qYCjLOJsywLpIQ7uAggGI5R2Rc0mf/mrlCn
0t8vDV988z7fFrP2RceVs3xBmkeaZWKTywYKGR43W1p0XqpvVRiJdJ3Hp1FERVWJTJ/i1YN2Zctk
bVYkxmGMiXKYSdPgj/az0cTmDA0P3K/JWEoKzn3hNmUC6OEqv7StnTx73ct6p1QMv0P1OeuJetnn
5CevmEUABg7dGMr6WZcEsMZYKRdrcmooCCFrlAHOOy52FqRpZlWYl0gX0bOqob+2hmtFtV6AdngT
1A3SUkLwus6cLXvv16zYy0ApWE928/svmmLFx98gAKWWG8zf+cTBed5J+WOvbvw/1vaKN2IdQCno
gEuJvcdGmptopxQgqYT3bgAOu7eoIjZ8QB8y/mEjw4BW9VGf2wclsY9vk4sJdXn4bU2nMoXtvdO9
G0s4Y3J+p5hne+kF1Hj6YtZ04fxx9N1Zp4ZeWJhBVXcmPEyZvbCBzmyZkbz6wosxZGJHOzXKmSPs
7O4keb/jFFtFOYsipZkKZpW+rMt6yN/RoCXkTAKh9mlQiiwBoYzmsHvZT/gUyE2vAwMm3co9EbvZ
Wtbd8/DmFnAdFEAVSD6wCX1mWCo6EfxKESjUZeog2dH5D2PRW6GN7REL+Aah4qpLs8qy2Num+sW3
YBV2YVPLLOzBv85XXSHzOq+sx3au8wjXUwQjrR1J3OkVc08k/3/uBcW4Q+vJJhb3c4sy+7+dFmH1
Ar44aWihM+G9xDE1y1saJinTh3hprrspc2WGCM68NQU5T9DMH17LKoSSkWfHBjM+uXb7DeTbxjP9
xXUOCsy9n9H12RlOHVq7Hq//N9QsMX7pkiUHyPqJ6FZdIIpfxYnDBBGfrVRUeA5Q5V7Z9OD/UuUz
47vAJgmcdiZSIM2W4HMwrdEi0cI2EP770iAnRoEqXvN3jsbOskKy/q5kXdb18af0JP7NVVWRUHh3
91h4wKEH9c/QK6mYaNG+uoSBRZZ4n64p/6PVzYxC0xR+rkSLgtkfiFMXui5W7oX9x6CS/Ei1Cqsz
gmApm5Dy/pxIheoFELcR/arYcGLj3bn7J5cCFpjTdVVoqwgwhWd1+60bD08dJBnX3T0EMuZjczUt
Pd/oJtZDJVgALmlhYEoCSbz3kg7kMQyprfBIaM6hVhJ6XyZ7JsyB/S9x0PFTqsD0zv6sBr0hFpTL
vRQI8uoRyx0FXtR84xok76YsJvV7S9JTbbioQPBJgF+CURWnViq3AQ0wTWo2IHlnfuAAliSGPvfc
Krg4D3U2t2RfRYVWS026PO2UzztYeXBZ+YGh9Xt915BIegHg43st3xU1+rp/rMXK2qkrgnReyeWa
f/jE2aH/7ATASc+R2E/acmVoVPD2UCGpuSuSuZP3Sug4TRNvkHWCi+ddAGPGWfFISlFjge/YR7sW
uLaS650K5m6N7izNlo/Nm2FXBFIfL0p6y5/5mRKED2rAyFkbZHnZRSoaeaKcJOOp0IQBHDSYgZLc
A4kiZfQUQPhUCzJjApCgpwsvTJ/J0081plKzS0tyQzZYfK1pmGCtFG0xcfw6qaiViT8Z/+vUGNZn
UC0tW9pbp68avZrxdeIggS00HBQo6mndA1UA/P5ajd5LOY2PA5KAH8YQBocnYDNZm308gFfGkeDt
T7LTIdk65VXfOj+3NsJdeDTgpzgeOMtwAF8skVM44m/7b2hy08fOQuYUFU/qGPohhFfJa/IC9byR
k7EHgeu5K8KOfp2NQWTQNo2ojrBzXwgtb5lvAwVvH+lpomn3s3YSMMRBTgBVXHKS+v3ljbB40Ph9
wAsT0j/Ahxw9ONR7pbCSXSmyptOX3pRccr5XPk/M8q05TUC4pbX9g87mrx4EzNslPxbwJY0tF1I+
xsTDNSn0eRq01WHAX77YLM8trul8l+UrRZZDzPbA944XH049H/bpXSJu23NGkOhbzCLCutquIAHd
Y9X24ZAs/GmLLgiIKvNKnYDsZghKgqFbFLWXVecfUKGZI2zPQsf4kHTGNL2mgobFfBZypwHLLLh6
SeSmznc8Az0V9WUrWcL7aeU8U3nE8ZZLHUhNv2qDyZA+co16SFiGaS6X3Bd9EzGlyct+usAjKgk8
F7sd4Nh4yRsX0GITqaoo/6NZeXKH9RjKawssc57+MmmfIqrSD/KJXLzsmS7PF+3tJDl4Efa0xY/B
HFaN80dmgHZLraMiS1NY+KKuguhKEYX5Da2dTijxEABWZrcHMWRM38g5cBAC0SlfvVu1t+5vDSPJ
EeY5kEUzCUopEERgnGa6ihn2Dswq0pGJYcqmfTThueacjPJsIxIvVG5ONZmrY72kIJjkajtI2WNp
Ji5Vt0VZqHvOHzVNO4pKEGn26xMSo2kQwip/aq2S4GMl75fs69nwq9iC6uX/OBmWttRzo+t5rzr2
hLrWXA/OppORT+SurIGaqghHLENqF0cx3sGedlV+3Yydswpt2BvPXLxTDH91o06mxQcn0U7w2Csz
0kXY6E4EyVsbUGyHfpCKWRQxB8CjzjgHruQiIt0D5sRCdQ554EnsCHYZX+9YBoBcssBd7YFzglzO
z8vidUrlLN8D09ygBFRcTk2bdkPEcUjwX7vLD3GP9Q6mSvOOKOXLVEPuqU42nsB5sG5G68leRTL1
fPM7Q8LTzgKmfhFIPdUN58ulY3OznBAg0mz4QnFy5yEX7asJwIn+F+FhzYv+HH/srRFAd1iAIpq9
53t9SFyMsRa/6JPk3GqZDgHnSIiMx5asZvBKBKgj0BnGrhwPXfwhWL/M6yDQxflrRaa8hDiCUmJQ
T1SVm8lU8dky6MKabmz1Yr8/R6QybGOD9rvG//z/thQ2hTZ0LLESjYFcz9hYwnwnN7yFUrsubZEA
q+O7lR+B+1zv6ShRUaq4Td4G5yfpUmS19p29+Ppqt92mGtnfCvGu+z/xN+O0GPODYwd0IKJrGV2V
IX1x/x7fyGBVjzWISjYDcIHoQoZvuNJT2Mcxsyzr8wBIPPXgvLo9Ow0GHOzMzTPUJyPX7+EG2lb6
yDGYwPpG1DGLvZ2T57gTR6ElBfVk/OJN4bsKiBZtu3lbso/aBtGErXl7CU3/TDp1XZQ4Tmzr7++l
SYXgeIWg8Y31ArmIOsy64QGXtmL4ck+SbZVr1QK9ca89TW+XZjf16lZVx7Up38AkZOQTGSXtI3RG
doGrH2q2CJa45uROoJxlJ01harZzXgC2zcEcbT1QReIFUuJr4wW7+9BwqiQRMjtnzaPeABF39doZ
5mEXswayMsiVsBhIyUP0RGdy2qVCMP7G9IjT4YYpyk4jAySsQ7njoKhIEhC/n/xKVKs9LiLRsyU1
1BCraVaWoDYf706sTZYSZ8vWKFuG4A6cjf92fsBPA9zUAdeOJkq4Kw0R/jgerh/FHQPDjvOvxQC7
+i2yUoZ7osZ0+NRpaPbELca+AFuCHvr+bbXoAxh7c6pgPuQTRNKN4TRX3Pxb5FooAqU+zjxZMBM/
hqeu4RZhvq6k8AmpBh4eCMZ+rhH9H2eqYkofXNTyoSPX6wLOUbYKJ4ZOyEOZCn8Jp1K/kxw9+/MY
aopbYygc2cDHxwoHCKEddLFv0W1m2VaYc0jEL385opAyVwHdRaSREmRLFcw/oSnPkx/pD94xv9cF
cstE+GMs/30aueMhpa5vADGqB4DIQSvANwnEBf2gdOHLTKdj1JWH3/6ewYLPhBfIb+1UUdFH9YMK
p2mBbQmQWylx0qZEIRvk6ydG5RICNO4Ex7306tGUloFYWXwAnM2BwNOs8xHy2odGolHqXQYlBVmq
03lVk2NVuEfWjeWL2/Xo4T4f1dK9gV9a/S7o0LMUFgbPRlytFNsQcql7q8TMMnxaPpriZpxP+zt5
nBmho+dghA35ZVBCHC4Yy0ceX1A7YMQ06fZsK9CdaNIR35x5H1FOm9V/G+63iekrEQOGDs5peWfK
zv5QAzbjyKqa0SxAYaUK/dWAo7H2Rz8OqnQurQdNQUUNOivjQnbAKVD+cpuUsj8V/O6uW5G9Z/sT
jrEXTCAAXgPBuiSq9Qidy/fXLZT6cK7hNaBwaB5dnTss0id5BCA5eyRpe8ZPFjYzgdbmFNSMDVI7
Tnjv8FhQT8+bTzVk8NzfYj6ImP/D90kzmTS1jlXzjE1dle7HkEBddkUnkJ5N38XDIcwhUz4J+NEV
B1dYBPSh6TaG7d62OK2S17BXRt24oj7+GBPFBv7mXh1kP5r45Q8CSYd4JmnnYtPrapZE7Pqvh9TP
P6suLig7+0H8Jipf3n7lpCyqng2Qfef834ezq8u8mCplY0URTft026azYY4n8s5OI2fiq3Dg6F05
fowwBR6wuSo7ScmpexehgDehWpRypqHaNeB5tzKApXqzum3vUUwZulSpFVzsXuDMaKKs90+OPcJb
nK0bpG8U1OClhP8oUNsQGIIBIImGC/dawa9rtx9gzmsjijTs7QYIDikQ/YrGosz0w0ZzSmjP8Jk5
G4QbBXv7MaAkSwNnAv6fvtJ8c4mEB1BvP3iTHKYqtuUUZxSGXZOZUAkIIxBziJbbexp+gstMsYO5
km09OZ7BGCVMeKukMeWSnV0ltsIQmUsw2Ub3qNPRfhOU0sMrWC02u3L8QqtwgnAYjZZFWJb/EwYh
9P56ojSEyzWKM9k0rOhwoUIAW35ZuiNrxnCi/ACD13ZI0T48JSEDGWkFST//mcovn6m6lRBfbwJ2
cRntJMU01k0uqF5ywUaljG92biePBVRSmfsHO5vuomCx/kDkSGUcfhsH/XlkQyj54IaX79XBtO/b
pExHLMxbCjCNqqIjqB7j/t/d2hHScXbANByatGs/SqKcef9O0QXjqDI8F0nPn++YQlFDOE69mQl5
2SsP9zcxALpdjdcTEtB6RW4PN0f4rSMd9VeL88f3x+29m1posNKPBZugsCd16kPUMNGq1nhMYekk
6Bv6FyNkRChb+/N+xCT+gepHE90fXFjCV6flqN3Q033NK0u1wEqc174sxtM21qIbnzWcA2IAXzFS
HvmFUYg7KZeaHj47nqUGD/iL0M0WydwYyy5+i7x1bfKc1kOTJMBEeWBe6ndWwfXwx66RYxG/xYA5
OES94hW1FzkYCL8hq3opRtHpja3dSgXBQQEJqaoItI7l0MP9TMk8f0zNDJP1WzED1D/uFxQya9sE
iuLrLT82aRRuTuKBoY/ZOwEXov9cNAIxL5csHkIhDSkyShQu9d0NQ0qH4jCLlI59HrAfyNS3a/QS
qfpIIIO6Nr7LLhgrztalgejuQuLY6HYgRPOevnrgxMZwFa+QxuO2IJh/ymgiEb0zTZwuVJszaU+K
UwxWIu8tsY3XDWsnMTgaqfSyJBPWDFfbwdUHXjOCjxaG7TpYK60nh07RlloO3m8tPStiCByyxZhB
utJQ3HseRWzAoJqInr6RWu0jFjaBcoIjvwwGqxvaM9duMHXA1OUgAJlghrDCrR6V1LvCevgqlAJI
+pmXnd59puf38z3KDaQ/sS0rkHtHF1nTdeaXXKdXHjUwFfmjWAGjtNHJDqIfPm7Cb3+nPVKKI2lE
4CdUPv4Al83myLolF5493bhQj7XJYp5AQk3MjJw7C4zJaivNFrySv+2elKjDTBlFcuXWmly38K1s
tchHT2OzMsddkzRHbk6trwMohHa/Bh4KMrK+TETZA7NZmBSbmr0Mll4L0PGE7a8bpDgqZg+SUBWn
TPYuNf7imIFsVYngdkwlNz1H9mFSyD6KxbAjPnyZiDUfBQIpteYZdJqfupxRs7OTRP3DG2GRLmq3
rC4JdWldqWbSte/leBCxsFhjM6ASQy/m40KeELymDUZZwjZu5/K7vPstErFU9ay84QRQV6KQl+R4
qpuV1cJyET+ZanKSDyt3YdcXKm8bIScbKoDT5PhLLsaVxdDVWlWR+n/UypaqP1qO2U/ZhWMwZ7jg
AwvtHacPTMs7HPar2QG46f1MKwnnYw1P940RaoK8im0UW+AgaJhjyC34J/8R03NqlfvtkkMjIa7z
uTG2RMZeiY930Gc4iYEbQKw7506q115WlCYsX1g7pT9B+JqNVkGI9mZB9WyU/UheXlz4xwsM28U1
IC8TngXYJW2YKr/s2XKVChHJR96VCxcQonawANQh+Y6tSNgs8fKEDDX8jpidjIyGbecO9imkLPla
iF6ympuPIaki2yhSgLoGR0kJJ4IpoXbFhgiLHyI92ySoh/kxhEGHdTwcatEZV6b9E5wvH3kQ2xRH
mX2MihVzmMEDaY/aIsI97gcCZ6j63rghaOUP8PcKPFh6W8YJE2rw66tWeH4InMYCpsq6P4X7F0cl
R6r+DuAkInm+pfs8U0foT8xgLXkBqBi3PxwWqx3jQKOI8cUuL9FBMRl5Y1atw4U6Texy5skVpmQb
RXxuFMxowUpz0Slp0e49fOJykdl5amStjM0AXOfsC7AziFLAigl+bg9G6POIYKDmP5Lg1G6PEEtr
k5xEMwTrOoUP4a4b4ORWjGF8Z0aqGhMqNJczwaUbm04tOU/CVVFkrADJVzJz5ILBWQMvjOp36++b
Bdr1WPuLSw0Rk3lld9BEnwru+CuPUlzJKW6i8xq/UFIHdY3v1tkKqta8cmYK19+aRyMPv2Q3Z/S2
asgWMA5+9LcG+7s4BVHVIavp4QDNEj7yJ2FoxG2snYbhX39oniycqCLqSCOtjbhnkDNAsgjZ8JQ/
m1ok5IqlgnJyb6dCt7La436TsVf+LbxjEyJGlNaH6W7/vi8r6FcNaCioRQ9e10+g/NbKfwhAicpo
RIOh9BNCxBm+lRrh1Y1ys/WWs1hThXMuefcmBKtPRum94CFoZoox5ChMt/rYK+R/upEArL5YuJI0
15aK9tkUZ67CkLrIaR4xgRp9clLhTq9r3VQZw9L/fH5jIaNrLTDjxv+TpWaGj61DeajLUgroSaqA
Hm8QaRmUPFMBYqnWOlw0Y93m5GMmzIagrDhtmL8xnUvCnnWhXy+tDoH0lRwv1yCQkfR6EKaqlggm
aFbBoXsUP3NhR/DJyuLshaAgLWKCbaYR50KIntoDpFKsj/WE8Kj1wyMTI6fqD1lMZKT7RFBvdlFX
G9ZzoYPewr2/D7rhCw1Q+abtW0tRzu7jJt1vkgYNbq/5xJU8R3oyOemGd7eR0ke7qA9RZi7xkIkU
Hhw5vorjkvMLb+XPAHP7rhCmFFj5eibd+frNA0gs5aEi9B56nyyIhvGNzcu4GUa3IdolZQYFXyjz
5IV2u6VrmAjo/kKpjwBEvgi0tnvtzGOnNl407HOZIRQ6iRicqZkfjcUGSVqEShrpPTuaKmxcqNFS
Gf7APnHXOgfAcU4KEpqPihakagQJ5UowRJscevYqNOWNFT6TlDXYoNIdjBX1Mog68pOtc3E6PMJS
Om3ulsPfkB/1+rGzLQTKoNNzV3tGp7NlcOjn4nQveyIEnmJfM0GnGCMTE+WGeRSO2KGQwH92w1Lp
+12zVZ7NuX9T9/wu6rghrw+HkyUli7WTwMzG8cKgYwRvMVKVrc37wSHRVw4PVLt1P2+3VaN+3W3U
m6Ofnc2vPvqi6uhgJQ83DcoelsmFlg/36uiQ8Z9/Iuos32/UQubSLzOhSdJZDxNFtuOhXMH2lacy
jmMbS0EpVGIQmVgzwkYml9vQ/+IQ0RcWeV222LrPdavJAi5uuRlNr3OcqsSxca7hTJaYE6PDHvI0
8GvKYKg95GWuEdIPSFCrl0NHPnBrpLqCNmrwHLTYKkEEbqdW6U5EH+i0ezXZp0DptuG3hpZUrXck
D9jUFWqvUMWjEW4y38iPU8nBr5NAVv2ukxibGyL12lNCkq/ULRaJsTy8aOd1r4RZny6fgJKOHbsR
/VWK7wPlbaoRjXIjm6O+0Wqa3N/CWWpA4Eb8Iyhsl9qy1jy5si8ar+RNqY60Ko7QRL52t8LEDRog
AJAUD7U1rQ/jBuBsxi0L0VdymbMMOlFVK+qGm8jtcv8ufoOBcMkx0Z+3wFTqfGgkKKjfVxSybWt7
rDGISmfFfF/yZkbP/X9nlAqOTRbVYCi/3sCtuIANSH/l6htaf3B8P8LhcfiSze5iTegqWYhDPRva
xvzarCAd6jqYkA+uTx5gm+wxcmXkNNZAX0VW0sSFy2n5jT18zCIxuDQDo+usPQC42B5FRjOEVg/N
H08Cg0vZq9uqRkfGMaX8mjwIcKc3pilwUeCvrHr13wLQoyEYbn+oywRbF55xkH8SMy/8w9rrkCRQ
JFFG6heSJwAIHQRqk2XkX2t98f0h9PUbhN+vCJCDgvLuk/2TtPRtXHZbm5qX93KDLapvIErtweTr
xJqO48cXQu4j1dIxrZzXv9o6SC21NWO5THObyjlGGAK58XsJUnQ8aBoDbONKRDYMQ3QIEgdXCsrW
1JIiNvuEyXufUZ077/8Cr5PSi//wanUmmcwyeGj5nOp0we7ke7HJKDMSVAg92QgcmFOR1bbIFmNA
8vyjengQTKIQHFwRoE8hVgUGTf/PjeEbspMGjs7hsMj3UEC8peEE3H4VJ/0R+dxrIFqfRwb9rxB7
DS08tRixG0WHSXqF2MMTVdNVa1wJYe9DvlTtj61eWEcqXEm3/S+G4BTN71T2X+6p8mLJnufzwDHU
j9RWiXqoBsFfK50itewgxMPGONRxT6Jsi6mlsbjvR0XEOTiMJtbp+fM+XR3h8PYUe8CLoV/GYKI+
c/8Ca36v2DaShFEYgFOuqUOD4Z903MmnjyKbCFYUFhsvJsV2e2NL69BfxjiOuKWrqkSyQmz9S6U7
kaEKzofsWpqN21toIoK21MuZfzJ8hkJQJJPFVGE6YFsiil3QV/nAmnsT8VKuV3YnGz+OOc2gBVpn
1D4LvRhfbONWnTkgH7YQJq8lZWOrb/ckopijSomto8/0Ki2PW0seSvxwW/YiwQJIAf18bcGSXXEt
f5aAi3XfoloLRRArBMbBhmy2H3Pc72YYxzL1QVeua1FpBlX8RXNPsqC0NTy3TQTzyF3rSnxxYCEs
wx4kkSyrLKHR/PZR+qLIyG/AJzso3iTbmbLObmjXUDRPNQJxjnBv/AoCmbTdhA7JcQ8ohF7AxSUo
1/uGKWG33kPUXWNWQ0bnsBczJ9HkabzKJg78rhlhaHQOpLuFKFArxIAcCz6bIEy2vb5QxvBXOE0O
UVvXqstZJ/Fd3MYmeDkMSPva05dUXwd2lhQU3u4rDNGqsPfdQ6xK6mskTPp84KSSDKh8yjONKGWM
0LYa3swCjrUm5duGhXEcumoUFdFD0EkRzJqxgyXCpgq+KERYDklSFuxEKnGm6BQzaW1Df+uNXnct
06sxpl4PKumwq0cnjqniDlMBITzi3ikBvzqJWc+l3336Evash7IBf1iJuaq0GWLbFlaP68l5akQR
Fyp4kKC166Z02LHJJki9s5x0L2Qe+ZhTHmN3E+/P+oANjZeZb3DAshZow8Nm+hKCk4cOiTYzxVGD
PdbGcDes+e+gPeaVbHNpNxBwe/yc+oQoBskYYPJY/bjT36dDiRSW2zm1MkpjhWsgCnSf3ysbudfW
hEDurrc+3DQG6W9kgs3rQe5n6LWWng7mR4bCOB2TMmI8k//qNDAOAYIuoK6ANa/9CBC3HuuClIr5
LlTx24HrH1PWSC1U6Ukm+q2vUpQITIlcQMvOderb3v+ujA5cSQXmixwYS54rUAPNRMjpJw6krQbX
s59O+fOBhMeEgL617t5xdTbL7Hhh82LhaBHO++RNBt0yIkRhp/W84TOAyF2miOxLxeEr3po1JH7L
7u50CEyyPyrIaWXEv+Sp0eTfFWUq2dkbwPBCKtviXUvuWM12MUg9rhD7VXHOr2uJwCIVQWKVRgTe
VOCuZ4nBiAwA4nAeI10trks9HiauiX275An0ngLNnFsX9fPxeJzZ891uilNl4OICSEBlSFaxLjgl
Xbmeok7RaEEGqIk9edkXYRbQHyetPqgMqX7+/4DkEVZ5BbM/4qbD36uTujO08lKuD53416YP4Hat
vYiwNpEzNlX8ryfwjkecx8om486sI47vBAAuwVHGgu4u4OCuFOwSgXQqlqk33GQX60ZghHS2NXbO
4c6vKQwOY+fwrFRk3sv0DGrQWnWgLtNP1xlYNCdme5U3acO76qhfiE0Ygc21JmGAngtZ//F4YODd
DysJ/XVcbdjSgxY+6qS7Qc5VIC0iSzCGqbUlseC9zVwDuLiiRApUJAlrHvxhMzAluYz9hOmK/Fwx
+K21QzUeUGdpEGmXk99ohJCd48YuNZxAmwYXAjUFUr/0TB5+8c1mnk5pqLQ+ZM0R8uaB+HpRt9UE
sumYilvnCxSJHwlJe2+aUUjOAlCG83ODspYLyn44TjvHw6Os0nTk5qlOEZUtd5mBx7X8AGi/aKjB
6NRCb2xIyA/Dm+dX+rkP1TCDb3wxpYI8xC0L+LVhihW7YKEW7KQdQmyh4hS6pljv1tWueAA3xWft
MXv0QEF8UC/q/MohNkT6N2zvzcAvlqZJSTvpEaEImXIGUGaZ4monant4AWNSWmCDgjHfXfPKMOe2
gwaEXK/Cmx0E0zrPBuC4VJrCf1Wka1+yfSt0Dt148kO4WwMQs0HGSX9ix4YOcFoJ/PSB/68/X6V0
Mqh2G5lkn+C21G62Qnjforu38QahpInV+uXBfp4HIWZBMtIkl6He39phABSQGVc8WK7NJJoi8USq
MEaDUPlQBM7An9bRllSGocIAaNKhuAoScXHWMOAoCkT+bym0/9dr+Htb+7GZ1jpMOqgH9R7Y1qyQ
Ex+k+o37JEskV9ZGB91GZJw2wL91DBR4EV54bchcLvEbsiPmQHCC244HfUEizH9odBd6CquUpoIN
pLRIHAeUjU/zJAY6zqxoModDV8Xv9LTWM6qkW2uOTpKFl2MIvG5Y3aUqAhpAEmUD7L1XnXxr9Rmu
a++mMZMw2mJe5c4GNt3xXq8J2Hx+yzRHHvBZjyAh13NQTM8aQKhHrgJIl5CeTl5pfVXmItXqv4om
lPm1Xrc0+aeXSWgEhjAFlGQiXCkdhr+akmVfmnvM/e/PNcsMYO6h8k3oVpXk+FHR1SPrn9Vw9s8g
D1t6Yrnl/lhggSpwWKp22zYHa6r2sXjpb2aE/sUV/m6+arlnVm+pxSqRs0PurI2eh+fkDj4e8IAP
XwXUN5eEJslfvr064tLj6A9g5pOxfDCKXd2UkCwHb0y35EIq5D/MOeBgRGPbDZWjTic04KWo67OT
bp7AXPDBzpU+rdyILVNUGrwdnv6p/JYjY62py1USsQEP0NvjFqsDe7OZTae0oF3Lzl8ji/ZfaRA7
7qdb4/hL/YNKU0iIqNleOmFCu64tEdmtB5h4Miwem1XDXvQtwhCdoRmAQ+fyHgAZbmz4P70IyF9X
lnWZD2DBH7QMYj5dbe5yJ6kb9bfFxRzWllrkjVIIYhJnui/GIM5jRkzp7A1xiDLrmHqKdIbdRWqe
kJT8UtuKcyCQU907EA7bcta18Hnwoo1K5CoaQu552viE8S5hOYN6ptS3jHGZHhMDPcHIdlPH2Smn
uKyT11QQRTfCkXXGvJvFHjlh3XSOK8wJk+mv8wxTIpP5ypjTwLfY2C7pZjnPWGZm1jmeyIrM00NZ
tiq1NUfnc1TpHkNPY2D6f+EjpfhJ2s8gat/7EbQUe3EfycmxU7yfrOo0cfsxa5HpUDO1eSe6TQpZ
k+aaQW3bTLg02/GiQZSeQXBpSBcMJys3l1qXCx00l+6eTsxnuLm3ZwFvh2fPQw4Ah32XEyCYcAns
S/ohbcsr8G9e8a9+kTnz6PUdihaURPSy20WQU0lyJK4xd6fHiRelyOiDg3reaC/Om5LmsYbY2uZ8
3wwKf342t2jZXrnW8v7a7tMdndEMWo7YrVtxSK5V8cNhoAOvG/XdoK7y/rBTJwA7o7DIJvJM6A8H
NOaWD8m1PYSbdHq5UU//t6Vh74ejD4SwL/tp+mW4UIHzYmZkVO6QO2dcL1zu9WcqGQwwVM8DOZAv
UXGw3SfXnwyQ2H6WV3uJw9dzzHJ8KiprEfdemD+06H45FOvw622V37ZUFkZa8p4bT5vKjsPpTxsO
ll0/Nb/bAPbNpUQIKrxssPM2IKPiCxz8tKB6a3vYRJnZLqAzWxH/01nWeAf/MPcYgZcVO6FIqCGC
agfYiWjD3jstkznkH+Gbyw8YJQ3zZQz+CFS6rlj9jrmY/Wf2POutSLiefDVJdyiKY1QaKkcNO/I3
KHvWNcV1lc8CnSb+9TofOqUdRjyYRMZVIk2P3rMwNfjpuMDUnlwKQ9SnWbC7kBdj/e6hXzpc3Uh3
shXk2u2rPbL6MoBF1neAOJuKbsXDYza4xGhNaT9FbBbd9O1x3u/Cm6RYNbo8PW+i61V5hl+eHW13
T84V1zHl5sOFv/QoQSkixXuZLLPGg/fbNmJ6Es8bmJBkuJkahWR/uoTGn1C85Fa6+ci5A2g25iv3
LytVVpalAWQnDhKF3/FJ1wRJfRRnVCPUlwNzQLho7dVyBIXlH+FHTBwhp15PiqtQGZ06poWPNOcM
5ohcz9lYUM1N7uqJMNog9YTipa8aM+R5BXhlHqdl1b1CmxznuXjfM1WmUkMfPJxQQSskFUklFbjJ
qOzx2XycfWYdHUXkDhWXxFetCQ9G6Zi4civy1pWRhijnTuQOuqXffwF0cJu2GQKTCxlqK2dxuzsM
NckF1cYJO6uAy4UJ0nS2/HkZSt1BGQUkGT9qNEJMiTYAh55JzPvrHgrabRNYkQjKigYyySdr0eLp
tFPH59R+gbLrtdLN7a90Qj3BiTxxnOwcv7ZeczLFFOS2pf98eWruP0BpkWNfJArbO8EvtGKok+MK
9bbX6RWzhNQvKMgSP8ofUH/qRZjeq8Mk8RejuPcBlhz1DoW3VECqWVRgclUpdmlmcBC9ONEMBDWc
u8t2XyGUNeu2/Z4xiD2yzy0fiOC6UACEo4RZOUuXMW4BvQjau24Jj5PpOO1mDJ48E2Usnnjsp9CI
rTcOA43RXadDXnlWZpjDl5/pBe/hLY/GV4c8BurrGtBm7/HiPJOvqX4wqyP7FCaQMNcaJ1SNiss2
gHlaRu4zDDskeSaCbDL+Stonp1XN/uuLQWUfqG66OvegwYkS2tDKj9V28+S9G0FIX6iv30t4sLp4
3MSne+QJhEWcYbTmv8uUdp3NVEXRBXFlkTqBlfa5NxI/NwfTSRxGYxbBFRFw/69QaZhWg8kdHuj0
2M/2za9/5tllN50aSZfj9RM88PaUGFxeGDPVjqa4kwd0t6iyCZoj9nl4Ne2DgLOW+onE//Wmz3Ju
z8M3eXen0megnQlGe/6bQkfIlI8q5et+sSlv7Wh3m28dVVsqoMTClPFDSs26Kp+WvUtzvqlgTEsW
KoWzYttdVK7e+NBvCNCK4SPceTv3FCJcfufpBDGFC7syfhkD6a9Wl4WXYcOVhP+nnmbRkAHE+M7u
W9O0Q8f1PuvkTG3MRMx3271evK3km2SDhveYEuzV59/T4IZ9SQBpTIlHWRdGwlDW9RzPkfZlTE0a
AePBMkSPOsNDMrt5iUQtJ5QbWCV8KXjHufh9ts7SCnvKKqwFrCqxmwePz47N18JCNX+xf4o4B2m4
f0uBOH6PUV1Xg1HdWZCLh9BDIuGFzycRo6t8qlxdHNfojnCVu7s4Z0E0yW8cnihsVO1Zotgq4JYx
mSdFau+tPucivfh4U1IORAn0YuGeAH38y8mWK4zmQJ5SZekgPDtbydKpRhlK1010xwBNUnZqJFXd
DRQmoPB80ng1myoW6ppK1vBubmwtwjvvftiYOYydJD6qEJNpfoT4q1NHNegRS5OM9h+WS9RNoeDz
+Vm35QxpYKJbdOI6uA3rsKSQknhW2LpQzQVmzlDMAwv9frtDzeza9Vk8ZDymcCuaZr1ZgS2yNCJQ
QDxyCmksSq6rDmU4JUIi5tjpwZx2z7kzaumt5EOby/ypOmHMPd17IoymRpNdHNbKaefEzDeB/Ago
485+80/V8gJgNP3KMhkDwFgf4c8INGZ/eZkjRbshibXuf9wXMuZvKpfNTDL2WslRyub2Opj08qXe
IEcxnjHA3qvWJsaOqfWv7fAwY9tkiV8+sfcASuVZJvAuMXbd5m4X7N+HqnTjmW0A7xMa70jIkrYO
y4ibZbOFbRHa1tmmeAhPESaI33QyouLNS7EgKRgqJaYOnnmcPuFwJjxHIR7dnxLm4HNro/Y6a8Ki
RiFFnGaHFKgLGFPf6nnAMEsyFMywapkP3CjTTCRMNVpPAT4M2Tv+ELnkMWTaKJqLunSuPPfF71fJ
y/KTRXGdGdrg5go0Urp+oMlrrJJoljW5PPZgiXs3H9sA4iP14CryJJQ1JpF1ExDQK/dl7v6fGPD7
QJRTK5VbP250Vw7O06SOpqxZsJTXkSyrZt+Axu+G+HHKpsaGVVJPbiUqvoO9wzQKnvmf4+qYdSAO
jnyZPQ+VkUK58m6wfFFBRtiIu01GFXPYOjg4HxQe4kZENpA9c+cRpntfWpr3tHI+pH7Xfsa/CtTW
FX7FU/mgcl/2+uqljwCGiYKEQ6dl1tw4iDtEe0LqPkbsuKRkqlHC312dKWEfeQyx4nid6trOBpIF
8DvqArl/XFH19viq+pB+hJMABVGmbhwP4JHgEs3ztL1g/8OyeVAnENUufeh1CLY3CyCDrZ7xafGU
1KlJ2vRFWP2sOSf5gj7znGs/oWY/kjMhO0qmIXciqbHuR9P50pXKC1O4UDGG+omQmVOwkiLGv4Ot
GSs96TrC6fU5RV4pDZdMOygGlnZllTJrhxy4wOkxkRiSDQ/hNedW2rGGZl3mdR3aZGL0HK1diCya
z4Ex3rWYoeC17JpHXfzE0TwlgbuEh5andolszfYugsrWj+nor+KX1SxGwRaxunSJYCDDxHJA7wTg
VqQY8teUcm9gG/ofOCqwFrSTwolv+6m46jcEN6fxKI7wppqSp+pEtK5UdJGNF7pCvBRoReBxRUD2
UXVXf9gqHGGABFZpgmgL8S0RkFEMldpvxGghjADpBISolfuX7ZoboDGmcrYryNYWW8JYJmFirfBu
zwpAjOKesbtJERvIPPaQIGC5DIjj959wLRASEbm/aE5S8hhUjO05oIjyGVR8XnskA67aEHkb/ICC
DgOWAof6fwsNxcy/xMcQ/V0MUfWZg24Zt4wLi/xhq1KddhlJhmey/B/OeT9qtVA0uSYwU5K6+GvB
3nWaEuDEPi73YvQiKVPKAwY0RdrGrnJ8dh42yP1tZjWOJCSbbPFq0cQYn3Cr9ARnTtH7FauPdqUm
wgjs0ucmYvOG1nT7XSklzvfPGK3IrY15AFH/OZpHTMFyusKvZzlvoIqD65TpFt0n/l8QqQtm35t2
HTf+5ov0ptEilCsxOOW4KST3hSYmX5PFgrpecT8do8n8J/x+aJq/sRKCKJ9nMuNTKxoXy+aT2y86
btJxx9U+2lsGs5s+s9pctYjz2XDjSRMulqGHRiWnhxsk7o6r7PEi3Di/RFykDpg0oyNHLMJ0nkLD
etaii0dv8VD0peQ8gFPCtGtdNv+Y161PrtNwk/Dc8iCgGV9Tyqnkn2LhGiEu+mYw3Lq3nDZNazog
SjFxYG73795sJoaleLLCprg5ia4MWD/Rct2iKVBG0N66pkfoJXon9shiK8zahtUhxXqJl6d9/Bcm
MxE7Q8UWQ0m1aZE984scxRXttwPdI7jSk8Xaprne56CIKMWJF3XtWubDPNdV1Tvlfp4+ifeRrc5Z
LFMYdLBpZbS88cve5Id/RHCDd/RocJ9hApKARU1E3g2uWwpvlhSh89k+S5aeTORUUnfoRQ7QPU1d
EMynh25nEgBj6d5vZ5gjWGpQzYuUs5VDHQIy7RjOFcnWsVf4zUK5mvTf4hTe3vJucAACIiLSb1YI
2QxOTwe92/ZBcVnNnRGSC+Uu87n7qr4NAQZ3+8bnZsi9PmfBKlJp2E68KJ5oDqkJ+dSe7tOP6nIU
qFYsrZnL+lmahygRS3ugmFKMGTnFs1EmtvNHm++4DZzG/+vh8ChFC8Wt931gbg027cRgfyRO11QL
XmHZAusJH2f5nNEKje9euRSgwP3Jixvd4xZPB2ZtD4TUVBO8ON6HFsW3r8MjlZZify8B0ZhZqjhI
tMinFWM7NSecV3w3P5ywMQVBk7yz7l8suQdeuDJpOk4ocy49hhxIwgoOUxBBxjp5fAS5xV99uiUG
QoESCAAj3PX+1rFhwQj5M3NyznVZq2DOcb+K0N7hzQBartNjAyASvEhQGvwSHKBO5vpCaiLBqs/V
cu0wnGc13cypXAreXk528TyPF25OkViE/GjFFhDu+bKdUgrODxA4RMjoGUwTJr6veLNVL7Dvsp5e
6/cM3WJVoDFUqE0P/3SLhd0AYPwITY5W5izydQNXxS5GL2T3F8Rh+DjbeRLl4XUcG2Zdsu9j4tyl
cMDss0OxmvYfGK2msqZID2YGWgat9NR0XRmo/DoktkywCXWZWO9s7LPH+vimXXBP/aJMdjNPOI83
ieyTnGrdWPY+IsaEYO+QqsTV6SezAXBX5RMv7mzjUDcfKrWtXV8DBwDGAZE2r+EV1wLcCYwL1n4v
sY+hLSrTOSI/4Rfy08NVXlQEEXw9LsQAm2anucvL5rwfkPst5XKmtHDQWvNRvkGj3nQRTusmGNVU
bag9sPzzZUF6FWgEXoOGD6xuXh7hLKXv9trrxlK868o7l6fi3iND4lRnOQKdLgQuVCigHTS2MXpP
S/x/VDpXLwExlbLwovLyG7QyOWkEdO2sovNXLVJsiRHgu4E98b7DzCyyejNV27WJo1fAJdeAQgm1
Cd3nQKP6+u7kJ03fcsYQuQ34FFvF6lA0n0EoJuucFDDdzbugaI9yfrhrWHm3o9b5Vq+x0nEzxym4
oRoHkEdApTHBiMd8/pw0y7EQMorSzyKgw1CKBywJusxObSRxbebEiZwXaBxDoAL5L3wykPtb54rv
nx8A+YYsKfmm5ur48q+GFlJ7EWlo7KUdRz0w8yPNAYe5wOC0cDTi327bntXQJP4f4aB6cHF35iLX
rFB7klFJIJwU7jLKgOXZ+axp0I0HeMV7L6G6Vb3XzHYhRmUo5fM8SqnV599rDSIEIVvWgcuHdecQ
Izwp7pw6NWDp2FWpsilbtb7TwCOSMfXQQ9G3DKxlUn5Mp68jXtMppzGUUVIfte/GHr83T2/UPVrs
/x2qCnJASVVt6BD9e+3GBS68D9LSrnyN7oPy9KHuEE1UA8k0RLylp3aefFDc+o758d9ZmQp01047
jDXaaelyHnRi5kR5+BF8/bwgeXzrfZcIq+a5wIrhEDmkg64YWuv16g9LLpkT4FMmqxI8iZp4ThZZ
9gTyeUcTtZgdYoEAEk3g2BUzhgdQPh7uBEzvZpO3HR5AIumB9wwHJ0gMDJ+ENar0C7PtjwDAG+yw
oB4lH+955rLRzeKE9AY2LJdFy0h4wR4hLTY+I5hhaAa3bny3KnsEvAYBT9z8mLaYEnUnuvh5Tac2
Nd8NP7owOkHAGcaHQ1Df9qwJw8jSyo17rnU/dMMf3a1XDjiqVBUFcu/cyhxOiQJwRIOzl5n7I0fS
H5APdWsS0X403hw+hVnsq2q7ZQkwv1wID74Kuy7D80pJRXNidNx5kPj11+IzGpF1lm6VhuZk6uV/
bTtvSijECXPCfDoK3VHirVm1bgc3lC2JuZ1iwOye4UbDuOUT+3fnuWdquet0gkwptzkSj0lf5jia
HkNiHLxKKF6Tgu5thkN6fPFY9H99oBGOrJbLVXxwPWJzhHgLyvHGtXaP02TGemi9zPxEyTdpbFx4
GuUXWStDZIsuCwktoaZlr3klAKgkGFz9eU0za+uSdaU+GjseQNfsD0dd2RSGZKpvi0fRNbE+fjhu
QI0qrMKdUEHDZ5P4TrxtrE/ZFOrftaPZcbZThsflIqFmN4vHIhBBSV51UWjOiJ9GlGmhXtYZ41hw
B9e+5/fsg2laUU7VTMW8KGRQDoTacY9onhbAyDkhcJrZixlspYtRSomhCFRLwXvB2IjLViPkjARD
WgnLLx/13i3HMtZZsbcgdBtpoZtHoVJLKmn84qYAawQKYvXO+0GTjkUkbzd/I4MaFTMzNk+jgMSJ
pnLJF8vMAPMwa1Wo+T2n3tFCZHkWXmIcYhGYDQ1+2ikMpLKH8OsBpbA25CzoDXtMJVG8ouhHOshb
DoIM5sE1fKvNgx1GZ+O6pEbFN7Ng6mCvkbyudjXA7VOKHl6QCeaN1S+TjWXizLjfTZq7up0NVew8
nlp0YHT9GfXPhIXrLgHIHlvoe1agEPl/fVyI+7AL/YtJDWWLKP2ajqXXNFBHrnJofp131DGqX8Ol
VpkQmrUpSnK49cfiu+Sujh7dMTSxVAtgAxuvuW6QgiYkhyZrJx6MJjeES6GH/qauCL8JxZVwJrmy
H+iO+Q9gF+hx2rnctUcB1MTCDtspHREiozssSlh5mfAzW0bOwnBnPc0+jvow25ovrGSg4NWDTjFa
Mg7X+29m8WTjG6uiMSk4hvvpt9mRqgxw9ANmwKS7uxra6L2PHyAHgrM5wotzIVHRCH0zQPV9MgYM
kt6VtPrOXqqPaM+WXKr9vTpXr4lQpLRmFoY5PiOQv62+rGIWZ8XCIMNpEPRE6dBNVd1j3vuL/DCY
TcUJJAzCwlaX/qgz6/I5n5craG3YtmY0dRHOQ9+2I+qBjwlkAKNdAMEifU/Y/mCyXztsb9SRU/m+
pO2pSZBylvlmU4oX/UXP/YfyC/n78Z2IbtBXwl3THMNGLPGwHFBngH8Q/FBI9PAEdb4McbidyjRs
PAw0QMapk8EdSt+TQRMzL9RrUBjpOYM2qQIUoyizLWs7bEY8AN5jdwH/1d5WIx/gP7ld+cmIxZAa
6o0MeU7xYMp6cFzxgNV+0Iyxr4vIQF8MtonR4vNDvhxMCoObtjWPwmFkvQ7zvk957lrKY6NQisBy
XOQB8dEklJsux9x2JCaPsU3tqGDyUzlWd3q1ZBbkd4M5pyViNFaxeaqMAtH3vFplUPRUtQgyW6Cv
CL6WpXSpbzRi4oPDOsZ6PTd1ySWi2rKvHJEAw3w0LeZbg+AtoBEG5nb12HvRsJrINrRfZKhuEub1
J8XC3IzBS5O59tLWrjg9qDtGSb0GUiLrLi+vFM3WvLE8bYGTOHdPp1kCP4trLnH4XjHkEGhfizmF
ED2udvBmPerfQVqdlFk5aPdBjts5Bu1f8kP1k2N7H3Y9abeoKDB96jDguoG89uH/MbYADyAnsacl
THRq/QhBX3Vp1Js0RqZ21uO4q4JGnqrSlNc1e57yUfwAuVzylTPCVPWGm6JRh5p7aJt7N4GAY5Mf
AQM2f6vagNbQf9TyCga7TrJiKul2Jq5Vl7k6gkBMqezezJQ0XzCiW8+STAv4tTuiWwvBJgG+a+gH
fnAuD1Eozj0cVKBaJe7FIb4S4pG0i10D/xzleUzNIpGSLiI6d9vRvKZyxAXLe9ESHIx6lq5Mb3It
DroUK3VRGJMhgcvlEdzNznHHXrOsGroazUwV4Uujv/tIStVJQi02aEEwr4PootaebNjQwbNFL18n
PjM3HLN5CuHpBkrcMH8lQYvSfaDBK4MCva7MD+Bj6sehIQfPQDraDCyIkM2dZGPMVO38KSmdssnd
TbGUv8vthfrkc1vg4ccvvah1S29yuqCVkvgiTmgx6CJFlKCxEMffOJ1r+oihMunbIAnsEVpeQ3jK
U+G0xjY8PGQsL3kk+mR7z+kArML1NEH4YRW89IrYZVnkzfQi1U9gSFGjr7mlJKsh0q8l5nE6WFyo
8+O6efgWnJvoI1dBR+uw0wlgDnWBkiAXql1oCcwm/7B9udl8qUywQSj7AyvbzgOM3Yzlm7IH3Zug
K6iNs9d+PGQa68xwbPP6ovODC0B491zEItS15TY5Vg7f6kh0sSges1bNp45NcTBpFhNSyPME0N44
OalfFKaJMpSCmKkaPo00qMM56fN3v7l3YmENeS9puqkVKMxlZNYlwlH5SMtDKKyo/xtu+ErkBHIy
PDC/KAaxfjsVHrtGPiHg+170OULA4smpmDDnXsASg/GJf7JEiVKyjgCEw3AsMIMytzD25xsZ6d69
/qGQwUcxPj4VD5EDOSa8JLM+FtQApziHp9csuJVoJH9OJDH3sR6U7Wf5dqDZ6tcbAsWldQy7y/6b
BhUjwr7P8gz0rNY3+Dya0DuBe0ieTwLrf8paEqQMdDfnbfQhGnDnVIQsxQPp+zX7RNmb352LrDHZ
O9v3voAMwl3O06xhu2LdzKwXnzv7tjyT6juAM+2stAVXb9vTD1BKgnqAYb6yX3jqSMBO3QWuLDrv
XuKeblLyMt7bRqohyfmSMvFJVcYV+YXA8E6B0jI/eo0WDjiLi6/13fKm01V/aFhXNHO9jrx39ew2
RazKmsTzI/HRTTawjRo5pgA+saDbwMRiiyXy9JSHxZSqFX+oBNTWq+8G4taVmYAdDTKoQhJLySuc
IZM4MeHCC196OWVNNXicWE/VY2C3l97lq8BeI5M1wwk2ujrb/HMHlkz4nCjCpBgVSS5Wsnr1NSQA
IuiV2gv7At2xdOZm0vO57PuNzJhXvyvjedE53HyQqK86CYh0j3QQNAmTDzNqMe7kw4LQBysbz9XQ
QoAxFdtFxnH+UrXw89srYDfSvytE9NuFU03WDic3jj3O6ncwrrAm/JzqBydUbsK/8bLgheHBCXQs
uzwSjM26rljUZ83LJEiGi2UWyucr2gkJ0PCu+pJzCtbBZf685ghV7ceSx+cnfjChydu5BvWGqT31
gtiOVKBXDua6LIiDEghoetBO2QNc5E88HF+r9vD93P4SO4/kxPRPWgir3nazDhZXcfFT0Cn1NZUr
ByBckt+3AVxeSawx1/mEju65+DzAayxYGv5MB6Be1RRo+WXDg5xoc4mn38jDYF15sT78WBNpv9Zq
c4HVoxTa1UKNVe/No0DBMu/yrPjzMY8Gf/yfIm8npip3blwlDE1uh1sqY9+gfvuAmJRvxIuzk0M8
MsytSiQAEAoOpfjojGhI0L9JB3/4+TCITw9lgjiYyweZ5omJAZyubvzg5fID4adCLjz7YY+ow4Kd
SHxUCAPawgGWqyqpjDLwuQrQz9kSN6uSOhX80IGXVGgflGo8/PUW30qoDa4b6ZbPRNsVzolCT/Zz
6kldyBJxULOu7tJHTD3EMUtrPdtuwJMt7wljpAGIRa4T+bCzjwnq6oyHYaLqSB7d49laJE7vx0iv
uxe1kC1AEDiw5oFewvzDqKuDU3FLYg0+Dy+veIkDE2qzjxaXymu+pSVo3TLmX2FlcYTZ1/Ubgz/y
aLpXTNEG8RKBygHd7DHFRQEFYiKzz8x7tOztswko68JxvMS47/0AN2r5UAJwcOALssKR0VMq8cHU
mBNV+4Y9PVKadgB+etcdUOM3i7VJq4oo+iAHREDIBB8Z8hhe1zBe2t6WB3vXHT+NUqG7YIHa4/TQ
N/+jIxut4eEJfI5tUtVR2Ra1krwuoGzWFDUSsZyFCLo4VakEtbdu4Z2Em5jHeBdr7g1kTrkDe1bG
Ff9+EFFZBw1PjqyVD5+ahJTuSUdHkPZNpetiCeupOqF+YXZIKpkCgj4RshBBRK9fYJXtcKSnWpgv
FBrQyJxyNLeemaBZYm1HDpYWgwjGQTfJ14i2RoAfaW9C+84b90MtqrB5qYxYkNydlgO5BhRpT9d2
8w+2F0gXx63HuAGt4pmwmWvCOpGyASHCCyouQ8Irr+oe2o52v3lFUAVK7BjIaKQJvgJItijP436L
NJoxTwf5aNFttQw5epIun7OlmjaYYReQ6kJAm3t4Ylu1PlUuztZCtSs7/uXsWC5gdQwUCM92gFxe
HPH26hy112P3vYs+ocWpwV0WGc4tG6zCnU6G3CYD1CF1BMJqU5n7TbO0NTB03URNX062mcEvQbsK
DPXr0l8RKZNyC8is9fRMQzMNXxnWRP9WbpsNdoPhd8bc78mtCl0/6gad9nn4RSVkJhOm9jK0RI9Q
w5QbJ9pOUrsm0CeTP5g3td70zLcccwKpl44a94Q+gdxHcJ3z5t8D92eKiCHHexxcyGw4SL7NxEb1
WGaVWzzLhVR/mn7Hbhu0e3nCetd3tNu4ggL7Mlm+8vqazjqvZAwgiNBSbse6bsLio669BmtMs6hZ
9+Qb/G7GfinZfC57a37bHnStgCCF2fz1Km4Ua3Orprph5jvYpvuuT22mFBI3RJFBmZW957YZSqfr
naSlcz5oJRRW4jEm+HrOn4NAABE+h6SdTYEWcM9WHfrwklKJpuIXyL6ErhCrmKG/QZDkxdd0MK1M
Gqyw1rZSapDqrUa8ob8F4FBB+sDKJS9IJ6ecEz4PRnovWbBefyzrqzRFI6GR9Ohgobx+098M1wZV
rPqpi6AAy3rOdfR1UZyoo4ktIzT1DERKN0U48Wghn1jRbY3lLt4jVFrWozk/2zMCzD/KLXa1RZTy
PMiwnU6p+//c6THZGthsT6TE0nmYkX3arvvvuWg/tXQRL/EVCdGSObU/1aQPTlFlIDCTTTEEcABX
B8f7AzmUeEC47Z53F+Rihkor73LT6sOoOu8ON/r24IH9lekboGStqEaQSKXPjrnyUzDnXwhIAE1l
RzTh4vkgws4bhU/lRxeh+8rTAHXL7Chq65rZCGceygyiW8cUmasU6RttwaBrFpXKzsZsxfactKkR
MJ8hhh8+KtwOHyuOSMfL107gDVhlcfpnPa+6xTUzxe3/nekwFKNsswBvH7ZYWYpqBmkCRc/xtA3d
qigFHi6naVLhZJJgxu5ORl9OVaqYOeD0QWMAABJNoHItryApiVo93aNfYHn5In4Belgy7pRZ/97A
n1b3S1nRRJ0nQ4Cu0gsT1IXYkNcbe926x3xkHtRf/81F/pCdzgT4jvmqXg2Jg/4L0y7yYQWQ9AQJ
/ix7aNJ5GLl6nVV58xsI+PixE5rN7uJ90rdNiIkyr38FULVy8t0a3g8zu1ef0dLc5HYvRMH+uYJ6
27Gl0jiYs9qsi5p4w22oAXjPkkPQC5J5O8lsKiPOr51L2D4ylazfWYjl6VsBjKljEYJtCHNnUY2f
xzFKEApRNgm3yg200LGL1Ssyh9r+Lw8TyrjwaopuMnWQk8O2z1Zjmvoz76p3hQwacPBTKX6yh21S
kuceYSXJgapXuFZ09Yg6O42tu5RRCdIv6ytFyUEpEepQCV4zDhbjHeL5tnx6LlqUKIaiG+QDNSEN
GmbDsOG+ptFWLWZRmDgCrEO21wP/iblvhOGSX7lLQSgeacVi8xnEaJSw9NrF+s52WLpDk/f7GQoP
TKIn0+kP9hek7mw98/SAQXyVBvx0ll4JNK6c4Q/evMJMyJacfo3tBxKKFp7Ikyk0r57VsRkC5fpN
w7dmxTLHTkC+KWcF87ITlwaYJMy984AkBhyN6v+VmGbb4Zpy9nXF/wxCkFNwsHVJR6iGh938w19S
VtPjO3/Oir8m1yoWeUmYZYsrnrVVOeUAWWjfSmcPLuFDkBWJYJ4pXxgYAfVRwYqsGmQe42sn6r4y
cgZabYuKnNQCyY41khDQYwBOcaVSK0ImJGQBEPXC3PXmC+O35Q/R66X5xhBZZjCAjP9CPzWyLW3f
bDxhk7Wh89HDxQdNTC/Tt/D917bEbFjtPNLkdb2vt4MoewoFljUEgVKhsbaq6bXFFf97foq8s98O
sx02mRT9peq+f1aBHF6PgyfJTBAIE/YiP6bJ6xg9S6GqPgyI0c6cIn1LUMm+0AtY4kWdzG8VJyVe
7Fr1P9NLePmEOpXOiDA/4w2CvQ+20Yt9AqzKL64RAAbAU0TdKkOT56JxzbvW62zCJi3FUjdl2f9h
1A5hwGiNFCHbn2C5T8sXRBbeRr4hSMAZf0k40LZwFQyZ5s0misplTowvLaltLfzakw7bi+Qph1hd
QUcAH1IAlryBOgg58Im1HkTABiOaKOQhClhZPn6d057a3r3qfdPNl7kUd0iKFTEgmPwyS4u/EqEe
FX50n822W5Ohcc5DvTk=
`protect end_protected
