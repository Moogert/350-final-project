-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TQGyWYLmJBL/ipsxoDTFPC+YAJIlnxxENRyyrYV8vHhD+yNOwYMiAitu9JrIPDCq6pGIHpwjHRC7
ZSauu0lExBRn5v8W9HFdLvNF+BGhhXz4yP28q6HWgDTuHgHz0kiGR8yp0ve1bgtGFihNIoYw7JW1
wbil+P4qmcz4L3RDwMRrLTuabsqLPbA1xrXRQYJmRbV2M1MvKcbQ3iEeY5VRFPZGDnQ4Xur/XX9M
DTD+ifdsj2cs9rJufwDsei0NFPZEpaAxXEbdeeMR+dNshm/gHadsSLkbNfEsMxK3iIXXocf8DAxG
Fcsvmwrg0neYrN1VQT6Y5SFeTlbQ1RxpoGHDfQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
hPuY0dZJi2tk7G29t0G9fCzQVzrQwWT0uxWvDXwFBlaJQ+Fs6vW9u9sGo7lH5r6nt44vfmqnPBa9
NUKpR0euP2k5mGa2pOOXJPABF5L8Lz+zcq/LwZ+vMBelWTfAkYGoxVUwEw+crYeWGctTnONGi5h2
ARzcDiCZSDsgBxUGFJdKkpT3L/FLe3m5Bdlm4ffSMadEHiiRHTUkKFpDcNbb7PUAScy/gYShbOA6
dtpwznpzsx8NOTl2+Uwt4DE25G2zzpwTfmUiILurWyXogeKu5dttqPzq/1frUsMC7Wd3RfsVdWNW
n3HTHYaxAfP02pEZ7K/gNwfI1ONtvmAtD5Bi88EU6vslSwlJ3Z2YRKBanwE2VPpjYBKMpoA/uIxq
c7Ifjrf2rLCBosiWXOPKb294dHtbWoEOK/RNwaGvf53u5ZL1YIhVSpFHfOb+Ys4SxscKzRlOP1cP
BaYRH+5TjBOhRDxVElUsjNNiERjaCu9xIe+Xf0ZshhkHU6dq7z+RRxx2oRYEgOHGlm+DLcxNuaHf
/I2JO8rmiLb5GGw3KdclRyEOODOGjMW9c+JUe0MgC8o8aPOP3XPsVUyj1oEO0pHw6JMkJaagOxCf
f5fVYtEQ4xk+p3fLwFg6LQgPHJ/or2jbya2BmMQev3p8veIRDrf5JgIAd7kv7acEekv/odmY+asb
TjWACJq4qbnRxp9dOKUCxL8qkp3vJ6DY15SvM1P3gMIo+vnOnbTwyrVpNsz3Dt+PFs62DniQDqw6
Z1CEH88khxqWq6PE5l3c/tAdXhk6wZx6CZra9s8WRWP6RmOq5/HGCGEKeIzHWaXKG0n6U1huVy0v
Tc2c2nViZBbD9yEJ4qPO/g/eLja+bnaFyYm7gJrupZ3aLJ0RkGPs3UuqRtKQUx7QOwuALK9g47ca
ahSIyRGZOlyIo2LSPPXCgMU0DruDm/3bsiAphQDiKDQvQN0Zi1F8qiHanSP+eeMK97zuSHDgKgu6
HN+/wVHcgYUvjIjBZLo1fsbw2rFNUIbLICFFeLS7L3Npnhq+QP7VnNjPuWs24YkaYWLt7KVm/Pf6
U6X2pYU2jhWdQjnqNCVOCus9W7a4Ym3YvTURoWcQtIQWfGz46J/Pn4cfYPZS7OmqU42YwcLz9Kyl
eKrsiuj8Q74tJ4/jh4+jMOUPDs8aNdqvyh/0INsXEpAxG9GGkWI6ji23ikaCjAMkqxR7tQwoUljb
WjDXQPQlj872D+ZKXkADf2PmilogD18XQm4/Gu4DoNpHndKYiyndmL8N/nqo1jFrfEUQMSaweIsn
dBQJFc6OXhXjyyLba2LMiRIlNuymoq5M61QhfumKWj58KCfc/5lwlyHVTQpkZwBgJXWvZZ8IGi6E
B7+lPFXWUhoRkjlogpGQmHRatV664p323CCJ7p7h6Qg+YWgVM/0I0u3uaujiQIffs2KgnGU3wFe6
TVgw/gPFHO0Iee6PJVb9SOB61XrtuySlliUgx05j5IWJInDjtwWiZjqk2xrnyeEF6yRaneGGAr6I
fBSme8ELW1slcc6LEbigvLag3W6Zg0ZaN6fAYFpmS0iEbub0wOLOEnrNG/gvALdFIa6NPMyKBnEV
rB/8+5s+morTNTXoS+/lTR72IOAi0PixJKWYbefsUVXrQ20Bu9tcd6Vqc0j8C7Pl2OwwM7EuKhm8
OeSbaBd2UQv/wKuv5SPqoIMOvfcous/jKM0osQ08WpsjDJGWWAX3G9fbHwOmC7SZ+xFXcn3Lf18M
Jii5yNFTdPOkRFyJpoOObU3SbSIeUQ6h0LORRYos9rUQbbkQ1STOXvfdSQKKi3R6OMJEr2ihKznp
iZjMv0NIeYy+t4wA1EXGYXejG+lGl2Hr8r8DHPMXjBgC7R4xA5k8yE9zPq6TULm0p7Ok4xbJbtnK
vNslHDbguOj7Xe0qGWyWzNku2EsmQbSiZFm1my2EpR1HOe9UYgo0hKNvdJpy3z37IZS4Sz/PGU5z
UYfCu5Cg/1OaZEU/oaKfp5tClvIDS7iPNya3ImhK3X1kEV8wcpDgZTE2YcKILP0xssdTXd3coMFC
m6zlFuj124p8dLx/ecA0xdDd6EISHp+rniQbr2jx0zwCy6UEaHwmA7ET0bL0e0ZcSWl1WtySwVh4
EhxaYBW4L59eUKPze4q43EzJOCU2oSHa4rcUY3N7zJ/aQyWX1gImfLMaHnP6Ss5irWiquK883LgW
YgmrHhHrMMZ8A6Gt/dFDKzzmq4ps6VX4yFNn/8a5073pXI0ekAGGOaf7IKKV4Mm3IWxPLr30PJeL
iwzEQCMpbpuG7EuIx6gSArFbMgbwamEr74iQgXMtuARTTCz8x1fb6SRYfJF7PXfpLKds7lNdf4RH
91oeX55fH/3OQeXTs+MIgULyX+yuJbyvFBqPuHyUcz42V9Owo2JEL2EINZrdS06iT7pJ2NJZ+Idm
ubP1MDcjFPik3gkv26PkAjHhFuvVLjij/61FczyyY68Qx5Dra2HAv7jab7wwqQNZBMKwJgZct1En
yRRSrsIFImrWzMhCxyrLxKtFdAsHZy1a55gbmzF0+7c+1zd8OmyMiY2yb/LJon6VizMEZgWkZp9N
xyBXdwLf2nttBie5Z/PUNtH2lwuDThE4mU1skGjEK0ldRMTi5ywOZ/9ofyFqw7uHLT9u+sih1Xrr
/aBkq70s328z+uj9nnDauzKClxwq4l3gBwXjRIvi57d37QAiJgzdbVG4V5MuSJQYnmGeqS8+OQ5i
amcizS8u4JzPIzThmA9NM/Lrwvr6nB08flIZLrcgzMnYCY6fyIvqG7gQ8vDHYZfriIdM+alam4ym
WmTmmbv5rbDkaYOq68jTvDi5nnEZPyJce9QCW5xV3aRrd1Y4+odiWLyocy1KjlH5b5Jl7NZK6H9q
VVsealtukvbCScO/46mG9S0+hnFrmnESyuH85aTa8TFf1L3hJwZRJL3jogzaF6REdllypuaolX6O
K43pRIwNez37kl1qiLL8MUUFVCSef1bh55AOIdzXfi6E5PIBYomD9VZtGlYCXVlimS4jxb7ClYeL
5TszwUFpwoDa5TtB9hsxtqCrqlWaOAuGO4A0UkAttxoasu8g7S0xu8PqwkA60rNsGbNRAzyZwiPc
+J6D+SXrm6uji+wtXKb1FimeXxV+otsW7EOf90TGY25NK3PBKVgsQ0DcgDw5iiVx+CqCRdM4Y4Yf
bg/AM6SvbZ78Y/sVPb/RRUrCQr8RN6Tb3sszYJf+6CpZOCiSuhlFWMKIjl19hfjj6P7OTDIF1l6W
MNKhW7wThYE2w/voV+GdZJ+R8jrw3B367p4Pku87sQxCRHsliIm4PfHW0XrwuohA7eapViPV3FMQ
zOPCHtUDCFGonNHNpJMLsHhDubCSzgT1W3x2jrle3Fw8zFtibw68S8ZH5aACvZpfO+yVyakeTk9o
yZ6uCNpNTSo8zsHsYzRmk9mcrI+XVIQ4WxKmGSA/x0zl9Bm9jIUMVDtWsgwEqmGn8J3IBXDjylc0
WulCuM3jT+dIfTNnUQTjsRqMGUlYs9lTwuEDuTzfvzajweu25SAvFMQJAevLt6AtOqof6bCEh9z5
LZPFJl+N+sxHpJnEw2E23vGFc1NqS7qyKIzKgs56GsDpbnVSfenGxjwYDky+5E/XKb1cF4DNB844
nWUK2+P5r2WV/e5f4Qj9oVyRFu3mw3NZfPQJ7tTdQIjdTPjy2V/VKY9lo/RxhC8o++O61tBmhBae
fbbaSf5mQ2t5y72eMNtuz9qvUm1LDKYpboOcb5Xak2iC/IbUiX1ILieIxwNkIR3fQJEV0UsJZVK2
C7JMyillWgOPBfcIULZdZR2zSS2+8Qf8mMHZ+lBTMZ0u2dn0cvopCwS/e5sat8ENL3n4l5XSpJLf
SHDDx4P9UNxrfm2zSl7N2UWn+QoMYVNnTG7fsA9OekXj8ufCDcWIAc7wBtbA2M6r6NB1nAYTDDYu
b8+Rq5fLs8joA5Seq3l7j615tZnD68MLxC3C8X6h98iN0ODFZlbB5rUAxgrRh2qccCGYS10UbUsW
OepR1235b2DumB3nCv3tZhJaphvpirxaoWho/uttOs8Ldq8C62bjZDHjw5SujyCPAgFiDa8C4TdK
9fdIwh5p07npBpPuM39q/vpMPqmebvDWdx5excQOvRR0BCOtpp/sOTfV8FzOx4fJuT4MdHeygcxJ
NDYEJ5frnJ5t/B1YRfhOQQH9J0m8d2L/8tlmoL8uTZ6RfpXUdIdjOYmMA5bvYxGyikhP12CObdoU
XT7vVbCMzc6Sm2svdqr8HcordkZaKML6olMx8y7MWmqltM0of9OANegjWEDBRGZ0dYlvgcz7cjTU
wiJmi9z+YpKeYL9uhZOkshXVW2XsrPlp2MdGRu9EwJXvk12jBEquPy35p57Nyyrl0dfTc4UPDkrw
VEcKR5PFfM5Qmz/GVfUvbdn3PcsjH6U+Y5A0ReFhxsBJW3Krke94r57Tq2YeWUJ1ArHOhfEvrZGl
N3U2TqoYiiwdMcit648dhbnS9Ha3SQIF8lyJ642x5feHtcqVAGGGxS/vzuW+PINH1XMSdL3MNGmR
m+FucjPYnhuWi5kQwxbcztgU7MIyBPiu5MA5TnYYmHKuI9jy7b1pHUq5vdSZmXt7SNPHv0R1Y/Ff
UQlBNZXx7qrEG6FHKafY4smO7/04U4+UMFERb80xG7wes+pGF55cbkaJKQ79MjEr3daqbJgb33Su
ZcPp14wbnjbT4P5DGPN+FJh1Hz/0zLxAByZGJ3wRltSqYj/XOc4Dm7erdGnR9FeqZO0kes8NIsm2
Ud2ZE+XQYlYymYuzvrDIo0UvUj6CZWIh5pU6brmYLre0qxcFFgVF23IQklFUmZIP3kttPtWhHWvV
X97qQqlCrPPcgZD8FfsqGlx3k1Yldck6fQpoKbR9mQqWC9LE9wWRaJrkEJbYy75GgmtRor+h5CSv
i5MgPGOX2Hqbmj1iOfoG3FMmdQPVn0TW3yeArnm/zOFkUpJG1TcBt/H4As/il7764a840YOnNHtm
FrGvInY52iyz6QgDiYDZRaAhkM5gsw8iEb22bck1DQUGsqZzF24sXOD0+AyEb8yTWidfdPd4AgkF
/UYQVk/cLGS8a+RFlFSyUspIrqkEizsPL1RBn1GnCzcRXTh99UI7KeaeD4G5MFcDgdj+uNG0tp+F
3zsZuhzgmHu0RWtqtm72MuklH996zXesQlKiHSO6/AOWBjanr13SwNuqi1/izYMaiFXYpeID5v8F
u+VbSGjhs4/y4BBhBp8vgoQxg4+c+EoloF8LgR2aZn5QtEXQRza6FJeOkZhPls2rUcx0cYd42UYY
zcS+R6FCt1O7TbJyixrB6MZi09hBRBGbqso8QDZT/DKVuubroEa0vozPjndiTt5vKHYclpczcWcX
jVZM8RYMOIQdTJY0odS/Fc2XBnq0ZOc6sD1MN3OOAfTMCTh9NO+Erk5RpJc2n5SRScP+jLhpf5pk
LL5Cm8voQnP6YL5Sk5LBDk6ZK8PoBhgvOGWRqaYWKI/5phW41/2ZOXx4+PHeH84XRWk2YGM76zWv
entIOu2CJvM9akyTxGjytVUrw7J51LmquUy2vwB3cCdVF1dVvw9J8STZE3Uj9gWcl7IaKhj92Ctb
hS3pbHOZw0SMw3jkwJsqwaEfKAmD2EPqWF0AbXuLedvU2rk1w3oDoHHFriwHYbzTIVmSNkBIYF0P
0YeGxOvKQX2v7JjLpNjyiFsluFv5Jyp5+zLbYMwFjMaShjA2t2lxYBNUNLRTt0UIfi/djsiyWmjB
nRyFfe62CEE9hkSmHPRHNmZexK7FjfBa9Z6wienZaEJIEbOBLEQRh6a2JpHN3CjoCDyzRg5BPGkN
EQ1PU1M6ZrBDfhkOXw51M69WjgQQfGdxg+dVMLTbXbGmeuZlLIS71t9wOEfV75kgbndXlJdoyL1E
zV7SN6sOGN8TWLzLVDZax/jdrRqg9KCCrapX6MMMgw/TWccJ4iHJDYj4U0CLRA9QWrB2mhdUTvfz
wQ2kHXDbgYWERuV0CtbfbyVic07jr9wZ70+Rxjmrz7mfGminXaf6mPg4TvN8cOYRsooLTKxfFOjX
k8p38sHBKEuBYfccCX6KxnIxedZZnMFgBjxJF7D0Zi4z1ZtMGneBwtBePgC5nXDtRF4rOGSe9Pzx
T0oWa8qfPFpucRUB5jrCNkz7/6n9eYcc09cFosF9/OXDyxlRy/2G3Ow8FtWLdbSymj6GVhkTepI3
6YNaugphYADGIm7IIsGpfS57/EXf1cV6GMbgRMJgMHXLVsw7NAx/kzFyIyeTNTFMIZeE1J+UyVIk
u0q+XmPP9xg7Qx6oydodilxTSFQE3HEUMxmQf9lHpThPGQvkhturuxB1+S6Uy1A9FDMk901vKO8+
imGFxommUhhWG/kprJDLNXCbWIJdBB5Hw4QkOuADiBlHTaiBnrFtDiG6l+uwiwN2W5eFp+v8PQRa
emXuGln7JLIoYblClExQlfoy+sjA/lFuY9G98Ptbfu9GfSuGHuR5MhF2K3I3eIr6kmHSr4s4gXU2
3Ua+6eC64G7/3+sIzciM/Dte51rUN3spHqaoIXqa/JeCqHcxm2wlpaQiOGxmPA8xhxBRv9e5tPcB
s/dEDdwnouOMdSJ4UKCf3tcqUqqnmbhusR1XGrNurYJooInWaXGOe71z+c8dwnJRTfcEf5pLARqI
fbAHuAdNe9bXOLjRMuPSSNmCzTGGCKkKXIwLoiKaxscZgyI5ABO/MsvXRE0xkIHM7rpO9JTPVbiz
Yb5DF5lceGdV4FbUm59HiLn9o3hLCKt1I2XzZcuLB5TBjc16zRggpjtg8VmfA3uB6kcIUikEsY6c
QfiSHaVTaOF0lS27cAJB6enChDDSqKF/xQ5UOEM++A62TfAaV+FmFqsQ/BMFuswxCnxyKocFBJou
+UXtnF+p7hp6jKM1DQM5GJb1pCfnVDNexsFhGGfT77p1Ms4fG0Yw1cR9INKjN4KguyHY+LFd7SAy
7l47BgqAqh2wbZ9+RONBZJORjcwIp6uZdr9secNr6AKJYK4KnuvXO+D6nWWsJWHPjJXumoOUx3q6
ROAFNO4BD8p0BL9+oN3gIYoAuEPyg5RVUM+MuaauGes0BFFcUcuq60WV9Eb7jxQ17MSePGC6kI1i
n8PzX1KN1wd80NY9PPevj6khOIXkZ9x3RGIhsZ9nL0nQZ1+o1RzEjMv6XpkdSVukaAOBFseG8wY4
mcsjpkKFcCHF8KpxeovEWRsasIaQXccfd12eIB5XwJEiXJwkHY0ZHqOBf1XAxInCnLMaFtbGpaNk
4SYZQbdwBAyYN0a42fYW068jtRPpachHt/4lpXk+2psJIpWazzxLykUXhY+oh2duNWSZR47RuwU2
SFStzma4brXrvXDPUL6gcLr5kDezdMybroqyRPPpC4VlJs5ktBO8sI3Cn2USWqPAVQCZ0W48gsv+
UGiGwwB8as8QIOWPSVnJWzWuQtL80IhPkPN6ftVLfG5wqfc4Nv3JCAyNX/6zSMgvouTzVU5dXngQ
2syzjnYGEMFO8yhv/6ThLAwaAFEKikvrAtnE6qWt60VFvs9Egg+lLe81el1KPLGKWa5ywJDARc0u
MEVKgVg9lAI0GYDRseezpxhqXcV3I7RCZD/AGUR4g0b2SKBd1jIZqlZT7K04a16Xh4I19CW4LDgO
uWtYwLjb5oCBf/lVMpPsATO3WCnYFkEEbGN8sd57EaShhG5RfXbqCozScx0OucNXL+v3i8XOFsEL
WAGwQWyphL2bZ8Wta1ayNzL8r9HLJSpAy0CbSeWA/XVLvDFqXOjX7By9LIdiR10dnQJUlnwRV7in
VOEJDUhmy4pKoYZvgbmz6w5bnft7GOVO0QxkGDYDTSq01S1jxKZu7hBu8gWyVnX0oLSH8H/O+Hbu
ioOOIMiULeCXl+Emamd87bcWyC7T63R2znlIpV6H8l9Q/L4ARRFZKpOq3cQBRo/YDo98vZQHUqtd
PVJ0agY6tvJmX52uS0AkN1hl0sMRUKDz5nAbbxge5MmWz3u4uwmh+VNO0YG5GRfVq7zRSXxynlbq
iWCMpYBcAx+xS+vhXeGN4ATnftw9bfEc76h7ChUidvkceVSUAQ8Xvd2YKY4kIaIXpfbzpe/qn/UU
4/O2bBhR2TxNzSUp5FJiZfsa2ISAp01Ymmx1xrwqRJzE3RlnDIN080HxUJNWn7JPR8NK2yOUYrOO
/0ZUmJV3VHPH3z4hc0A1ovi/63/PXz+QBhdj5Vc3KG65mfCm3hNUiuKgIbvXwRqgEEVElh7xOjHN
NMPWzpxL+H177ChtojO5mCBFHuHt7vLMcaeTIdDuvg9W968NOhMD/7cTlrFsJLaSOUlNir+GqhdI
Eh892Eaon7N9aWrJS7KCf8FSIA16DJxqDdImiAJOuxfbqmVNam4ATem0qASZGeSpG6jeErag4rH5
9D0dZzcXsPJ4XHRwwNBRAnY39AsqKix4onOUsxaEvXLzvpRCU47OVgl6+C0Nu0Vl2bX/B48AvOBq
n4M0QM7M0gHla8aF2Zubf0SQ1GrVujm6/W7b3MU3paIczn+aqYlis/RP4WYJlGJQvkYsIGjrylE5
2CgdEa313cfDARbxJfEYkZtlSK0fAHJumRe8Xf2IoCzW/R4VSTOPBOsk6ZE41VgvT/uDQsKvNpXG
K0o/QFw5Jj9dFa4DNA4kHtzhJCIUSs49KhN3ztDxC46lkjkZW2Ko3Kqp1acEf75DB/ayzgd5/oFg
xyYOInW5bsaAxWjEtfsUvYRCzn4+9ErhD78fITsR66FVypEEZdCpKU6jMVcXZsbW5pFqgmsPDtZu
e/l5RzWkfEDTqCMVfkUZ7u9+bX2vxEbVzRuwes26bYLJptwuJOyPcJRpusxSibENV3gVxHYqZGI4
81eFdR0i6OUym9sPl4bUG7V3fkFSwk7+NiiddljFgqJndAoFxaq84i0gpjBevownL/hbKAYWGyiu
g2Lj6/uK2zdbaE9ujXtT64mY2DdQovTg92J3M3BcxAEWt5QxZmT6AePiJzSSntYmX6J5jFOlGBPV
aTJLOe/cX7ElyEhuyKRijQGyKxpPptL+lFFPJOR+bqRqSKtOMWLnk7YbOLNvqPATO+/qyNQi9QsT
haLpyEm7Mbzfg2XeC+5QDGqjoCMOQPoMXZnD+w5LCd8b2Z4z+TumKBmmtHoW6UHy8VPzISYlbivK
BZdMEyAu6vQ8medSAM75LnINJaqGBo5ndx4oYj3LPICixy0tP4pdTC4iC0lqRwzJeQ7GCUHdcFrN
qyGZxso4G3n7OD/3xHCrfraxsDJ5VdmxOr87gx+SnXLBFro9vDu0dAg3yHyZGlSqkykIjQgvSVsV
iDBDUQj+wJ2YXk6Wz/6v/FxYS7R9VqA/zpIBvqd9xoBol1wobtmQTFWfe+XBLEsg3rR2WTVpFBJl
fza+wOB1cdvdObvEEZCMq0jNERIG1hET4h55s0oApuuDNc+I6yunBbKOfOVeZ/d9L002jK5nnQBx
45e+jIYDiCYOuai9b7KypRIyQ57/b1J8bFXnk8QU36OGVU7VZSRwbWx5ov6NhlxMKReZO0gNHI/T
MO6dU+Pe5s1mWeyFi5uW+pN2iSJIuPQt3EDa1UX5rNk4bOHcDPq+qQgo30512johW1Kk7mi4pxBW
MztCCliSX1vFy0Qcl8YdN32U4LXQryM8pwxtgSYWzCSDSOR10xSwPYH8I5M4VNlpjqjf/4RKV+Ga
UumGK7i4jXAjgHqwxBs0W7W6pII9LSR4cXuf7/M5ldoDTo741qEkeitKEVTpd6EvNAfvbIZ2tBZx
8P3VjyOm6tWhwTg0sIGAlp6dW8jQ2nzkJ/IOyBupIRiFvOOFbZETDi5tMkzZfN8F1V8dXRRH7OLk
DhJUaU/H8jTMJKkP+YRg/4Kovd6s9VlUz5cFHNdXTyPMO7rywXLGOL08lCU0ZvcAqoskgO9fndPo
t9iM2j7My7UXjSlNm4lOvageEpXPGSXC5ZAzCeBh/jnLxCd4fx8YuDpq+ZIFxnt9oNc2oRi5Acdm
Ad5aq3ml1lfRlucglBZ/Mb3A9J/mfWvKj+9f87CqlRkArgz8jVPFAYeX2wA0w7DNXrAyMn1JvcXZ
jBmQEgRacALKXD1YghT1L2l7l2rVFUTSkoDwsU0MKEEw57P8ja3Lq12b78RgyTh59OYgDQ8OMNjR
CHHFuHcHDAEtB1zSx7fcDVM0khkX4FL5Er3ovnhevHwXRAUst+0otQJND+ja7Mxf3cGenroceJuN
cXgKYex6ttnHXUtZcBrrpDybV8nXAWqdnZTFIKK6TaypEs89loVVJaN9VUvPsafNQc+ahniSRsvo
80eaogXtwug+O6IjDzMugH0VOGDmtlX/m9NzeftkaFgWGbG/THAkceeRyOtOQEeqHF+TgY3HHXWl
j47wVn8slC+vSiLzUx/DGTMLwe8rB4NoAAwZqJDWnfh0HzRESnFNB4UUvnN1g0zxl+Y7w+WMyg6K
Pv2sRIj0jPGG/CxECztmWXsuSPJt7TXC0a8IDzVLfbUarTw0z96ZkcIN3Vw3THS8JqFvbasntmrh
26PYbAennFFVk5VuLA887piNYNJytSxLa/dAoYANf0FoKFcd27LNma9XRDn209eSH82xAJkbf4/N
Xos1Umk0p04HecXJVvf3zMETHKsFpaclrfkW1ejjpoMdL73Eu39ZAovT23etSFxKU9hdoBx7YO41
s2LNbUkhO2XblQe8AYZPgZ/zzEcMI7rblkybtqbnpLlbn6AJNWzhbXTHk/cbKhiheDaijIDODv8d
qnCD6mwDNSDUHA6TKNNfgUsf1ZwRDbR2HpPWyLB0tj63KQR7ycnpC21DnAyFG8ReCCi1rGphxeiI
4cnw71zVzbJ4TmRYx/al7GONmQMRXqMSim1BJ81Z85EWxGmgKURo71dC8dLbbdfP+WGKs6+ObH7c
D41DeYpMAgmkdzQFEMhfOnm48F7RBRsr35YkCjXinwk2ZrGUADphYteAImPYProHjudNYV2ySpiG
X3pvGS62Eb6basGPmX1qCJB95vaVBFUkGO66aztynYbuMljlrY0D3jkZuo1jDD7NhNJF/WigA+Xo
PoAIRaj0XNJvdU/IrCKajznZPy1SggUqIQ3FvSDyvatMhEnu+uOQ8aqj9sHOhT2af27qyHNjS9Si
dXgHJIMu8QQB4bCVHGrmYpXBq0xYuLRm3ZOvN7tj5IikR/ukdpZgOQwoQQ5AcUhX6l33ZMyJmKzG
SmhzJUiybj6Ynzbu/Tx2hPVKgKRKRIWDsnZy3AUFlZZBfYV7UpIBTvQTdeaprSb5o7gAEscNi4tA
KVBbPqeDyfQU0VVwD0jC9FhKXS52e7O444VGA/CBZTiNJ6OZ8OaU0a+6K1aVCmNTMoz1l7/rv7z4
y8S9qCAUCJQ9Dc+Lq/qzUB3vF/Sl7LUHLfc4oPKukZ3cueA7w5x2zjPCJnaNpyYrhJhpHzuVkAA1
AybDu8h6Rn0nKcW0Vv5I4QGCyv+lR5VPFTOpQeeMuynUo5gCmfKUwLZI22XmNtewKj9TVhXPRX5G
o3TFIFjthxcuBnaHtVIDorRcCvQYROu2DEtBgH71iVPf54TxEW4TKVyq4+axABtUY768nScCltWc
2DWA5rzLG/9EnC5M+FRKKTMirb05XfLn64FAF0XMvkVPXY79rOdohCwadAHAKifnmlVCUB3CZO7Z
efGikCT9hHNvseWlU+tkB+az385aJQksGokqXbnCi3apOYlqSIffE9XBwS4S6U4Mw4ujsZYvAVf9
ZqSWY8NxPUNh6kyjsxv3/Hy36WY1iPKSKs1fjpjFigZtOPE0flR4pqNc0oWl2gFFz5CA+ruI2h25
mVOoL3i7tjxgb89yKXn0w+uyAq0VL1Av2+U+jO+z3TtQw9YUl3UDxBgWi+UWBmLd6SEOL1DDl7YE
YCkeXmrso4IQIXBjzHarls4sOrlnM6zGV0C6/b7HKLinwB0jde/Cof/J2/yivgqNPVFkwwNN2Q7J
BdXrsq9gfep4xX80J/eGO4v2i/KGINed1/Shfke5RhzerwYKlIC66qsW/rgzBZHUGc3zMbatBjzA
f9K/gW0SJqxmxszh3zqjM0xyh2dBDAiun4GLKE+p9ToLcefjt7Lqva5h9JsdPmjqmUvt/vxrZxeQ
nEHFwQvEFSQ5uDeyMhbtCzhH1ZoEx5BttaFQWlmFgIFhYy0XQ66fcJLChfSTb3gaXHPPCEG3s694
ma7oQktkDp34iZ9ruDTbO4yenaaa02mf2uqEpgV/Gg3/tgmDJ203RPnpl/ykbwUsrg6v9W1+SgYx
H4RHgn8qq5VZrFDP8QEe0021lHGR0dqwSPG9peYg3CF0UbJX6aoMVOIPu0YUZ3hj0pDy1PaLQaXH
enREVS5iVJL9Mj6jcrkdgLqe/Br4b9HWcmi/ivtV2xdyam+S1nlZU2BQVg1LeQVYtBi6/2CTsuxp
Seqq21yfnDrASFHqJoApkA39jOPrX64DldGfvKxJN5mvOPZuFm0poH1lPj9jDMqqNMJbb+usVMXG
OTO+U1gCyQ8M1myIpSvm45gfwlA0IYaS4WBIoigjEp9eyN3lr7+renI1k/6CsWd2fdt4TDZE+d95
n4SE4+VGZaHHKcNPuZAkOs2oA1FeIezMQARc2YGSGCffi2NOA2bPB9xiH582EnuxLAgMNyhMHpzn
QiAyvaDglovPktSYwz9S6NtdFKZzh7bjVg7B8Fzb3aK/XPsbMnV3NAN7h90OQ7BRuOlRkbs7Wql0
dzjLyjTaDwDcpbvPs9DWbhyoVIGib5giqyRILV9M7g01O9jcy2ojS1UtLxXTsYiymj46oWWsqHz5
doDtTnOFaK4r1mrV0sVm2+FwdtjwSYz1L8D2yz9lOhZfA0h/vcfgFi1g4088mDktZCCA3bHHjbwl
USPTUqhztSIWPEIykWUCSan/sF7oD+y3RxDbOl1fc4ZIsSA5vw0DHnTjEOTgM0/IQfAQ4LXWZPYg
1T4YI4J45YRZzmlak+MvFUpxR5PSDnE/Tcu+vgkTlQk+HUz+nehotmFLxBI7+xTfgf9gD0uji6pq
aU4fM26YBSzcEs3r0O/YldWyw2q1O6W1ANMu50RodBw/9NJzPW+wDtZNDWDjo1uruilNXUMIc7xj
K2YGfEvchjTOugm970u5zUtB80B5mdSTwdAP05Gkbj9GzgPWvcTzhmOc6YZdbSorXCDWNC071RzC
jiVnFouZsAv3dxwX34NK8M+Bc3IQMNjvMhCKnyN6fi4o6tC8x6zj96lxhqWQhfJEPvfi8UepdQTh
c45O0p69jnt6GqNGTpWXb291cUFsEmXFyQMmllQkciw6BJRvAyDtVzlD032njVOxcq94yrOk8H1M
be0l7b3Q9uDjsvSHXpo4j2SIlhRykomXfeOCh2jH7LzK6mv0oRImd441LJQXq7Ob/pN3d2mx17FO
/UZUZUh17mS3dFse9uxeO2Xq2Fq7Ky627tFGGl9XOFKCN3rI5Ywox5PtISi71X3Re2+/EjVnMNCd
2M0TYP7U3pRpblF+Tl4J4C6MqFNG4kUuo7JObRIZTYojmLje72Lme+S2ymQV7P4hEXDdCPSdnzmS
QknKZPKaqG8fQwpJnkVQaNW7Zh/yB2bYP28rOWZ3lfYvruNWsj94bcd4DrxyUUtrwocK5EqUHzMs
MSOkaROhI9l2mD7ml0/13FkEgal247z9w+fFavsXXhdScQkLFKkd94tKECmY+eqFi4PG2YkhdQ8n
ZOE1aSU+2J3Wpcbs4WDsBSj5fxoXuJ/Y8VtoOqjFLhJcDkZhy/Yw7mKb9QCY2qk/8b0tvLkgpjh9
64OysWqGiEgg0DRYte6vNkVDZans6wZAZzpFk0eXxblV+S9RE0/FQ+dPt2wSEXOUIZ9VjgS16uqh
Ef9h9BvK8eqBrsm63L0FLNxcgAA3JUDerL/Kx7Y5XMpoJN+ECCoX4eEeMUNO3YBC7iANEmHrLPLp
jXlkQ16KE4tI0UtnUnL2ga/UBMcz9ZDYmU37ZWp3G3u0hMQImBmQAaKd5Si3zg39TqEVXDU0K6jm
nb5YmbaIqnVViLiWKnB5gHZ9200ax7zcMFCMZC64X9i+vRz7cAnDYSQc+SAnkgUaLy4O5ACeQAc1
4ilBwxu9
`protect end_protected
