-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EqPhrtK3KyDOEqAwcKVUwtJAuCHdXvoEClOUQz1Frn5HCPkTaAlaeQThQyJ/CQKUyFbalXiUqkq+
+ae5hnouxtSf6/NLqGL3LQXSq8Ki3c4g6X746yR+pbLyJA5BU4EYEtP2/+XNU10qF2ukZ2aS4u3o
MQP7Q1kE4fKtlewIlI8ZDrheroEb0+6USu5b6G1supi0aEx/YsWHjMND+6PrNYIYoOoJAtVH837T
Bt+fTdivNj5hsuWEYm3ERv8Pa5TOxGBSv9QpmYKmKvOJEi0h6UpyBEiRG5MnRZV2imcxZDYIPIYw
UaFpyvePBW6nHYBQNG0hlGXG4TYPAt9M00xT5Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2976)
`protect data_block
RlI3VeNMSbpW+WnEs3pO7PpF1F/cfB2NVJBSFOiYSTKVxw2nDlFTZHbDvt1BGxkWrmzKqvcs6DfQ
qYKk0PXtn1QwNbKe0spMMaioQPIpuWQBfoyuuL061CsXYc2FVcqMWAzv8ZmPBpe1d1fRk97g4vq2
TgLSRXi3DnPDE1LsXr99ZpQiE+iqvl+pq/vTNy2KqCTJjUQpSBlYK3fVBPqcU2zlz+cdYqb9vkwu
cnStn0MmTrvU7N+iWN8adX+jYcH1VBG4EPxDk7hNlREDqoZYNmvFyo0TTbv0LcZw7IzflGiTHJBB
xo6NrRGttupakfQ/CqEtdlVjE6PDkANh3b1JmiX3D9Zw91yhpwl8H+t6rq+2Sc9AkapZ6DnLCp54
KeC6N/ltq/UgbIMPjP8rwr+k+UDy2huaUoTo/9C9UgN6IFqkfwm8d2UFmad3ewe6caNgXCFaAg4l
SrIQ/as+hoqdN20BlhvpXEUOGHRmLR1y/XpT4HW25nLrdEPRCCkJXOmwpXRjUswifVrSZlVc1w0F
7h7XbUux3R14r31KvngvPfJF2LZfWH1o17Hm1NF+DqonwzYvbzJxhU5IWZzydOWdkWWqC/wFpfMh
0fDvDL49cg5YSgGJBh4CwK1xnhzOO5JYy8UyKYHwWng9w9Jsm5hExTTMdb2Gsv8FGMcSrYXjpkwc
Cv0b5A7baUxEO1OvU3kQMDcCQUl569o0qsNBW2KgTHaUK+nVqxCR0Oue2TRX+TiTIj0mSfd4Qge2
VDWP9iuK2cUBuJDScG/D/nZGyQpFF/cflMpuNKisGfmpoURVa27X0EzV7k+51HtDf1IR7QhE4y+O
jXGdx78tsCr8apvXtCIKRmuwkHLrm25JZ8QvCq46FdJxjPenVupB5Oos8SGsZeZV+StxXYZ1Oi3v
PV9K/Yt2uQo/GlfqfV58N404mhyiMUGwgPZPUNRc/JzhRoG4pIuyI3H4WEtgWBspQ7jeXN+rusf3
MCB4aZ9U/+At32c0KlPzWXleYd35kPkDr5OAvhk/7wLtxZEp5rnmolbf9/fkfFq/6QtBzsvbNtsL
wUSdLHRIy6tkhO/o7F1SuQi/LkfzVtNLYD7YoAr+NBY7JNSJfZEUkniH1IHk4EvW678xLcfvHFaC
V8Ulx4qPz7z9px4NTofmMc77RU1f4J8/PfGjGvyOiTZqvwhodkH/QMQ/aUUeBJTQPB+qt6jszbNb
3itTqSwBsn58o6c4EXyVSUJ7WEGw1JasSkz3cT6sxk21sASkP/DMEyJuAHOpWEYz3dIU4eDnIIYH
GRoermTJDbjPhHAlNsBuxkMMAjPLSHSYmR2MkSuR1HrxcNtrO7+tViMuQ6Ue04FxSvbi1K69H9e+
ucjbnHK1/rZXVa97pnZfLNW9rurYZE6deOzVvnd7unWaeKFqH/XHgk3iZ8HzGcjn4ge/mQ9Bkb/T
QC1GH1f5kSIJMQH7uqY+pBMKfbKksrntkYjfmB33DnQh4+2ox9P3S73nM9K5CbZUGeTaKBVG8MLc
hpOStYqToUj0p/jP0/GLLKT52AB2lmfdSXlrxxLeShUCUkGqXKKow5IkdZbrPjUO5gfzabcF9D2m
zKhsUvhWdmehI/ml+5WH0IO9ZQU2gCPbU3i42HBJkuLv0/JKHTb7cwlp+NQU9rGnrVTcrPo5NPw8
sab/Ed6Atpg60zKWcCAkBegWAtl/+r7vhYnMP6dINeGN1qbge3+wKJf0BhWHMMDCYY0JFG9H9Kjm
+8Sl7+W+OTZ1oe4SXIHENemoSuTKPOqsbccdol1GxqHlA8awS5iEolhqh383TIGOWOGdav797aqZ
AEj1CdsirJbSqsKRpjnTL72kAv0r54bq0wMSveqRZwBGQlOCLwPEu3Capsz88qPjYSX20bG5OAVO
dGbslPOB6ntv4RYA7x9VRI3TY2tdfj1diBtXJcnoWZrf/IlJ825QPf57UchrMLdwSxCL2SmZn/5Q
SI8yoO05Esd9G/04ONsP51teimW7hV8Aejwo1pidEss57BdFPOS/4lcSCGJgfwtASyYWBJCgoJQe
dX+X4OZ0E8lb/wW9Bsa+upIjoshNJHUCl3GE0juK4/Nrr3Qp2yEp2ZolLYpE7nmix2XsEsjXVkBz
LJqBP9X8QM00kQf+sMF5y6QlqeS+BtRAeB3wJ5NJKS+KXvSyvUwfVphkw453tTbDqXPNGlzyLopA
OZdb+MPJ2rGeMz2BYebC+8NDUKPqm5A3kvoaJcAWLf+0W7z0adRntDBQ4xZAUpyNQB6maew5A0BM
/mLJS3PF0ZOkrBLq9u5mmr22nUiHR1m4KjvDha0NWvnVxF5EPz75O7cgdfwrGY9SdqMjdHD+OOL5
ErOtWdORwKct5YqGQB1mGpMd7j3ILtA1gp0dT9COqXqWBGwX+Faz5b8uNH8IF+9PLD8v1hh0EPRO
yNhPehj4qP8SQqD/a1rYVSmP7buATUCRQkZIHj84kDHqyG9BWgl/7C5MpDjRemTqN73kSzFco68A
FJogNoLxU0atSO7Kep73GV1afnWsVPOkTnHewDOMISCt8yPKKnzxY8m9SverePJqA/AwckFRZg44
G7NtH8rzYw3cQrldaV4j2FNfMHSORagOYhnmlkSX1tuN0IKxtjEBHSOLYWuBBwBVm+u7NFy5IEr9
DfNQwCVAKIS6WD/dlnB43CSbEUHHncYTMskvg7Lfr4sbtpQpR3TWXVoVdBWDryWFc87L5FPedMv1
cS0pZImBpr8JpRT+WcelIpdaNNMk8L5AI7VU339qbFmiu/Js91bBkyvB3loMliuqFufs+WUUyOb6
QGVyzAb/8XIGJEuuAgt10G2GviVAqClHBf+xO0gFJfRUIOBilvDTSI8NluTehOiVYqMhsmG0VqEu
xvjUA8AANpxUXjuTRHe+N87kU+a/JtkuwV37G3zwgq1+o8WBH1gj77LifIemI+6eJO3HpGhl2LYo
LLbF+j8h6/eIyIFPx5XzcclW3j07WAiLTbuZqkL0cm+pAvlS9ZOrIOUmO/vAHUlWet5jop80lcW6
BC6JExPqZt7hOKvZh+VaztEQDaltqcPnGLrzlhYyizeDMCmg6eLKepr/e9qXcxUoKfsn9PtJe3CQ
RcBfvKaUEfNj5mHH1vYIV1+dnB3j+2JXmfm6O2QKl1adYOe69UIdufbZhgiXxUfK3m9MGHm20Pt3
6HLc09gDzNy+xb1bbw/vunNGo2q7+HS+CGA6WsJwSs/1JtQuf3YlUxGCvVBEGfHoRMkSJimDucM9
symGYk4xP3u9ifndhhyYhD/7YqVZRwan0duZY63+xkl2HuunFlZHGHvNIuJNsclIOwOWVvYfVMjY
yrsQV/dc8Uvyw31F2Y315bV1Xmi5kRzatP/G7vAAyJe7MS66y54ZFquFijOr7c2lIPOccsydl8Lt
yGWCV3tAix7yIoj9Z2rZ24hXxNLhnY2tfX1KKlEuZCOPX/QesDhCWcfwkvh/kPMSjve7YfMKt2eJ
9BEBECmgJs+j+EcwX0T55mgfDETLIE7IeD/ia1B4ni4r2KkNP7u+SZaTWLpTSXApejuQt173Wnzk
HAvWB03HlycjphV3SQ2iD7zY+IjYuAyCqLYsshAJ3FSNTTvOAdlaGEH0PCVLbZ9BxcDz9TCFjvFz
MeT7sTH+dAmYLgMULEz6+Mv5B8XIWAnJbk/aSz037xMCHHqyp4BWriLgHRXTUU3l6xJ/G7BircQs
sV/7rWMG5Cva9DBruFtOtgLiEAU1U/LZ2N01fV7dhC04V3QS31Q+Jo5A+Q0jNOL8iRR8cDyPCiuT
rvkiA+oTkC+bRqonZQRJwwybpupgneM9WDJTvjIVYzCEaFSM3U+IL6wMzulBw2PYGIB6UEuIvJWV
m11g1v9WyH/tJuRtLUX4fXEsHcS+60RN9HwJFJhP4vsJqDUVPEPSC2Mk38jjrj3h+Wp02VrNKqho
QlbuaRU/N60JPMPc
`protect end_protected
