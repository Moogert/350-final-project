-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IS0A4c40ZRKw3y+qQfNbHmDsbm7mU2n/Ys09OGOb3WqRd3g49bAbTeWCu/UPknxTFCvPc6NkDyrO
jPZkwQxdIwe080OhTYaIlSUo3ZWMORuYvygR0S8TWzPo83kV2PP/wwLuAkt+8ugvYCESUofyZka2
B8Mf2VZClgjMBGI4Tg9Ki1WYMBmWYqAhFwjrsWM1ZmnZTZD14B+pEGOTcA9uDz14jqB2NufY7zoZ
vHEz897F4XQ4NernP8YIFrAd0Vtb68N8X+QbEV/SsvekEhX7+mvcMezzl12vdVG4R7efVsw9Nr7q
b5+VDAyb+FKKwFFARDBcIJi1M9zKIYWe1Y4lfA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
37Ltmi8j7D9RfnFOjKZiB9GTUyKLHWWpxnAylPwGbJCg5Fz10tI0vhAKp1+EewTCdXag5iKaeVz5
3l2lRkC6SYbgCQGa/xjNuN7wZTPrMWRgHscUMO6mHOeDseCDoLKXTDrlia2KM8TIxSww5jFROVpL
Fl3UG9gUMnd5LOZ6PlhRPEUKDu4675vc5Ri6FeER8Oy0x6DwgfLklD4f019tB1vNBTijaIOo2myx
x5tFU1BTq3uID+vCQGeifuQW2xZp5IAUm3948HJ/gfrtGolDCPxMd6zNMebs6MxfOXOvfwX040lS
xRSYFv/DwzuqhJsxpiggmPTcSuZIH7BLRzFl4UF1iFo1yPWIQo6i5K5Old181opNexjeFtr5/NXS
gvK5nAk5HczsjXOmCncScm0USqn/T11bJCkxXHI3quzBEesNVWoGVLHbkNhizvxtXe8ayivqnIQE
rxgWeA9r/mt3caznZ+xOFxavySSsOPnzgLarAkeHrMimzcYGL5js86cMFv5X2gke8HpYZj/nN9xW
5NrR4m+7lMPdCUnj6Hl8rnHnC+CgmKSvKVMIx1z2MSz49CzcEdAfrL7RILAskcio7bvkGEKD5Tuo
+46UMNO0xM6OVbCLozFSYOKIHlV9fRNx2q5NJR5ISMsfDCjiWk4ilvJMWtOyvOCmgGlk8T21WuIO
uaYV6ViOM33naWFPDu/OGQNlMbWw7xpnD5Hnyq6x+f/t5WTX2ZJPvi3902DGlZZIO6FdyWqz9raT
yKUtm4Absqkcu7MdzkCPnUS+XPw27Ns5GGM8Xyu0gXcoZUyzgs9dASRZBzrZ7kDTCXpxJunHq3wH
5xLQPDv7APquAIwnWAGB4/pkEkHuZ8XrofApZYJ9q0S04tA9x8S2A0fQJSpsbqsT2WPXD2tS5yn0
+itgUyN63Bw0a+RY92L6EuB9u8HwKwGeopWdnDAEYQQ8Yr6a669+o/6w08sxnlmGMMwsqwQzIGgB
dnEWNn8RY40teE/QuLE0yvPSxFaZVYSJsBCDrUk+/1rfwTP0v8rahtTQgCyteP+ezQVYEh9+S6CG
lMYraPEkbDQT+34/J+FujSmJNZ/9BzfxkoEU4TWaE8BoHXP+iytMcZSeCuDshuZCdSGUDt21pBsV
ZX1HIkC6C4j3/aLjdatkOxChNSQrjQ6JeOHbPKNXMpgS+4wI18Vvvs3Cr1YExYdAc4MEwttZvG/9
xvf77iAIKzvCMEYoWrehO/hnQhEQXKuurCPf8XIGEgyQoRIMyfpfAJqw5SB8FbN3YvJEDoWGuShD
nu1ClwgcqmCqTeh19uh0GD2vv75924nwsTJbqTwjFRlBD2Du5EO0F/qyv5c4jctm2idoiRsFmWXM
odTsVSfcaXlYkcFlyraQSSvFthpuo/4fK+4gXCcNWYFEXX0AiO7XkkkwY735Ptc+8PHMzwgDROwr
/om8gIvVCr6P67rpS5nIuBvcAzWQjI7HB2xrhQePIN6V/tD5Tm/ZUgei3FGdwyizYSrxUSTyT6R1
Mhf1+QFgG5Ro9Ri4+4P6RhkdBY1SShO5w4AIi5SYmB+Sf1cVhax6bFwvxMYthjKKJmclp8IlBCbW
fFec6F9akX7Agj2nZyBvr3mAZ6vaaf1g2490nYyiEsW2IHbbCcXB0p7yfAbNH70zs3pSo1s7OvaZ
+BK4UpSZUwC9MuQrjAWOmzof+0jcPUXwpCoGz46/U9PmOezvrKw2rg5i93mxmawjDMx0aXsQ9k15
j1UCTgM6KKQNjyN7xhKMnuCCYL91hvih3dd1BUwU1gCkgp5FPFjswzsYi6sZlRwNyLzfgu+ZmCJS
3hmvXncbg9hGL9lOZJhyF6/+Zt+f4MEG6OwOC245X6O2g0LgkUICTfCIt8GxJVWRWHw3b5CKW7Bm
Eej33wXmpHiR99m+WSxbB7nGsbnfLIMQUalHvtDDGo5S3R0THkhBUwOospuTFeaKj2X8t+48+WYg
IAqfsXvI+9eWRbDEJjBSFndF/W5EPbvlh4NJkkv6XwNpB+veOw4nWjsC8f0Z+vXjpA91d34C4pCO
ZWZzQWTz6UkPcCt1NS7BQZp7md+NDFjjOpD9UsXmuaRjpIyZrQXbAbX3BKbgU4sJNJ+DJZfCfXPu
aAxM9cLRki2u1pBTfp/QFXPuq+7c/YQpOqTMoi/bbmsMh7LZJohn67i3snD+K3YISykegVBAjSaa
1LWO/GESL9AenboA6wh79x/LcFCS56jQLj5p3v4cvjFX1Y11PbfzIhDNfr+G35VAqHusH7okls3K
XUIz79Ghw0Z80ies4cdlozcXreDEEEFB1CdtRnQJDW3iu5yg7duY7j77AlD3lCd5wZ/oV5VQLLc5
hCn/EmLW9nZXDUuVD/DPuaQ/DYonfoUBQG18HMFy314Oj/mDcwsLLfqCT25mBaS6u5d12biRh7M1
r7aM2cRGcSVfNbwucx5kHt6RrPMan2725X9NC6/U9l0UwYh5fw8Z/HXnVqpugMD5Ye4+7oiAuULD
xRVPAcYEOaObzy01RFSa0TEI6wEKs0C1oQYk/XlEReXAJdLCkwXWK/ps3OQxSqyDmukwfAL6sD+x
d4aiIn2M7r2BSec9benzTT2MbM+62nd8sm/PD7oSkwIf9ot4BBlG+79512h5BfBUV53uWoBXGNYa
RXG71UMA1c+0zCcSy3YG5CzbGGy/AmT3nUYr+e8sXxj8kcUC0gn9EuVs9Dn90aYDf9Q0kjQVmKJM
kBW1M8nOoxfhfsis5mlsMBUuVkAjmQTA8G1rLz5eocA1Vut0o4gUXCLail1ZpWPFYK2Izhc/pqUy
C5YnvnK6GXhhHIF/OocwalZ1qK/dp1w5cA4NDQW1VR/4KSkMfPF3VGRfwoYPBYvDcPXBbB7bQrfv
ccG8R6S04g/jwAMjZsd644uLFEwkhdA4VPt0SOO6rkH5rArfdxuaC36F20CYtm1N5ZMcryYvvfrw
lKI2uTF+Ncg/l9vnYSd3XO4PUjdPvzRYPuGQeOQ1gcsyQMwm6qDccG2wSCnv7rhJWVj8ABbz7jpb
lIkTOox72YpR9LvdHu1Gi/SQl7sN04Leq00AYqeamAoGvl31fGWhgnK2HszOK51EmewVZOyc6R65
j0Kyxa5xrvBGveuWGc9xG8RuKrQ7u4fsNQr4xFbnW7Gg90DLoGkexpvOGUd9OGbCRVhwp4wJeAjA
6qFfqVMVZAyRaymYPGe9wNw4NiP1tK0NGSvZugHV9ER56sDsxQDP7iQQJo7vL1nYOW/GD1ez5Bxb
i2g1gN2Al3/J6JoxQvqaHJfnby3rONRLotGbRWFjaDQEUEc3Ko10cY7NIqa2OuAtlr14ogsnJP44
uZKJecRb98keRpq4nMwT4xApRhybwoOTOX0//BAgPTGx0NN80Kv/nluMbHxl35zowdBiF5lsFqX8
dfiEfWeHZEGr1aKC0yaIOUT9Yhm15tl77MpkwVnMdNmhk8Ku0EFPv6Cwt1AhOC9ZqEQ3dWNwZz1j
bVViUU6UkpY6iW81M5EWCgRjcPfYVInJEyefNBA76TxkfkNn8O6gAs0lYB1IEiB+goo0vyJ0O0Rm
JH38H0acIY2TZqzZjDGTlFrNMOl+i6yXAUvksN16VO7CRryCV40cQ71dAaBX8HvWWHJErcyPKDk9
H2acqhW8C1xUFW4Bi3iSQSsmLQ567+bqdnHyCQj4XSd5aJL/sk6v89JO8BJwRcKTUsoRyEQbwmKW
cIYOME7V2XQq56H2qJsVQhRs72LXD19a2w9TyVgTWgE5WP2ojyyYoTUkDTjpkt73dKP2raRvLY1W
zEeRvy0I4RF7m940U/PXN9OadQnNWHuysF1x74kW4ERrpTlx5wXivHUzWh6ci/uTsqYSLCT0ch2v
d2LF5UWpJwKTo1nrr4t/PbnsMlhdrXDHyyG6qVaT6GYJGpcu2eWvLlo3/JGgaOiFfGAgU2YnZZZ2
sixNJk9vyiXKe9tticKR2RyK8mhPUvGLI+/e6v0SObVQZjFyBF6wE26C3h+ldQWRxeRTd0iMV3Sd
rv1C3IDeeqv6f8+9buFTeJyMtoM+eBV+Z90BIn4k9FI0gRJU2ZONLFWADjqB2oxS4XFAX+QWmRw9
TW54qZqnNb7btnvefOVoJczmFZ0n3j0Xg9bzAgaViiDpe80iZWZJg3eoSdtAGLTLbttDHs6MeZUH
4HyCYdoIa4AfLpDAlHvAzpAwLg9BWYdLaS/mxRpEOL0GQlFmx5wVZgt71zddkpsQPyoLfGh0KtDh
kdmXWVP9LAmhqqz46/3uEJsu0Af00bVO9NXi7Ifz/Tm0b02FiuWft8zkBtNVpKIvNsz4DG78oruH
wF9XkHYpUffcL0TpoxL8ApGVk9eqSZBHv3Ay0PS0Dwe8vkCXlMK/fn7JNnr3AhgiCTXuYG7qwwIC
0TJmsY298d0U2jXzjCQqUE/AssSfKJOFFCr5mpBfys26v0MyLgMAM7lQtK47xblr6ornz5Brbsnn
5p+s6loGVSvy3q197C+bax/bg7eCUdfB50zdAOdTg2so50KBnLfrILObynoLxFZMBJAnXZZWfbRB
6Q+JFw/qLf4VNX3YiaBSg8030Nm/39O0mQRxmTVLH2taiTLrbtvZWseWle5Grwgnix5IrrViNLtB
AyVMhZ6DUvHGY8NqKZyoWnutQziUhb6pitv87ZhUltMELZktETHQInryjOzkiAq8MLsyeanzMdnQ
bOLfRwHdWXW5E4vCbnAJHo7wFHhOrk+cnRzXwyPLOQ/qQdk1gnyU2d/tBi1JReKt3rNHf5HDmmpI
or3IH+jucy7XtSXPc+5+myA1fp5A2SYRQsM82uYR+4N0Lk4XXcxX1KsXWppmpXvIC4m2NL1luG4y
fYvcxaFv67uuMOK1v339vm9fUsqTGeVXGJjzOsH9X/PHpoHRV05tTtmK99HxqJoCP8meoIpIYj1r
IgtERkNoQH0sEWesJx2INuEWmsl3uTHoTLJsiVc7IheiNMy2JR+/yIIBmxlIk/teNGEFfFX3M2VQ
8hVo0eYp1uQZylO+NWGRZP1853ogDAHFgYeMP9vU+1eQZCpuxfGB49BIqrFQTpvsYwOZYAmXIyWS
EiacSrPSikpUxZ1Rn5sq3RyeZeLcWOceRdu2qRSjKeefSFN9XDHfPZrphoNrg+mNtmjzkEw5Rb3F
sOrivgNXNY2nEVflC6rjMVkvQ/nVGhrhBzIwtQ7YrFbW+bYFwGFiKnlJ0Nk8RFhg5CLdSzS+Aoil
c6IpqYQnmtKvXYoXFyIC5oZqsRVNOw2IJ+APxs1B5BDSfsjjKN6zJaKBOW+3GjncVpW0etvnltjx
DINqyVnudfVunck7ed92a40jGi5wl5er3Ud5MN437IO6UkyAcjPsviMglkwzHSyX7GCMjlMKIQfO
lDkSPTR3JfJYIXmM8uckW4PC1/57aPj1P5ttkOEQSrz2NLa1+Hx9Jjwvhpcy0GQEQvEynShSxF2S
zaPHvdmZGpPWSdCP9N0AmXNdUrdoFkeSRXbR1QDV2DzCLqskZJaKjz278piA6YRzrQgRwBR/6CHJ
l/0FF0T+cYhy7LsSH2g9H0itmEAX6cfiXkEEzWzqjJQw8ErgjFPbdiXXfU/2wEojneUkVbLEA8Bl
gPMQG7jW1YAZx8XCi9Hb9SPj8NupIVya6omBuuFwt3/HVVS0SuuCTFMkK2cN8K/iuVfquoIOBvTg
9lO/ZF2wUieXJF8vyO5yvlKZBYlPkvz3S3TFw+gNBql3OxKLiYQGCrut3RqdgFA03PW084NgOBOT
DFWo5K9UaG2EwYMXJrePjMD3pG4rk0SduZzVl9LW3yA0YrkwDc0uxDjuJT/mzsnlEhLhXevQG6Ph
yZWUY2bZNLhg/BpQU+D1gTUgqlBCnfxlC6+tkQ9u+ZD11ob1V0GhA91ixedA+PmwUA1P3R3bn8Gl
tWz0iAFHbhyHPUQFZM55erTvsowYhTaijPluZpTRsp/aflYyiXNVtLBAD74B3Pjq8N2s7cTLiXHx
hhtmOsYUPh3XbgZOQ1HPb2zz2lgCNDa5rxbB2Cpp/2eQYh+GlYUydmDVdzVNft+V2X8zgN2DeP3O
/aNUbUJvtTuj+diztENNuveNNxpUebJaWvS7eFx/oJ7GxTfLUoGm7FklTBSbZxzow0mHzke7Y3rL
l+zFP1tOp44k9SUMV7At5Iaqg79hYfWiKaPMqhp/GsiYCbjqSp7Qv6b1ArP26OyeTRf/HCeSxQQP
77aubt0iIODof0L7PS8Pb55HU4T2IakyhRYcLWpajlSy0tJRBILUrhfHyXfc5iHfKJ160vomQzqX
pAEgdWuwlQ4EXIMOdYkdDcI/q8PKiZbx+Oa8AgISEw3c89QRTnorieOsLNiBae80JymngjHgILe3
fQPo/QpfaeEsqKG0M8mooBjTiu9BsOi3upY+Vdh1o3BCFwVL1J0TdjcC9vUodByn9TQP707GtGSY
NNgGXO8H9K7EWzxOKbZBAkXr4i5Lrf8dUDvrJo03dZ6OQwtwGmNTuDX2vja/sPuFg3MsbFG5Ij2J
aQDPv7qgWW5A0Pv3wuMlFUXBfHpTL5fHeyajUT22RK+XM/IfQ3WZdfbeydU8nfwZrbe25ScE3xrK
u091ZeOtGj78nDZJ+GWKTbR/exS4GG51uqUk0eCY8pGSE9SLnc/eFy069r7wEH+hdEJEVexob2nI
Ippe2XrXLeLFJ+cwY1QSvoyQ3g5Y+M1e/8Z2weB8YvfW0jmKaYcvgaC4d1JZJEpKQT1SNaU1JQa1
DsRnfHFfNh3Ec4zsB3Wdp3WcrVcQB9DKq/h67vMFWLbrHZm8aNSefx+QfyOYk1PuheDMaahJayoQ
SjKbNFvKOgblfv5IRXiWF9s8bGX9QKiLfVwO5WZK7l3pVe/qIoC7xffZYJuMZIJlZeiWEv5UpObR
aefb1nMCXKx9lzPNY2pIrUCXZrkBas/KKPoPEtAV+vfvWZN6KdxmePs+Jv/YDoQ6sc7SzJgH4BlV
Z5ep8yVEgSusPKhsMuDrsT+K8YfJrKZjWnNL0I4Uf+Ak+3b5zsSI9NM3GAbYLENQKhQWcJXt2Trx
uJvli86UfRIhVxtbjI3x0GbTaYDIodWKEUae2sNRxxN7Z8wINFmVS2Z1Eiw6dWmF0ifznL9PBhJ5
GfquBxn/rfyV9H6keExkuVWD9jGcZJx63ArO2wA92utmrWiRoB2OyUYvOB9dbsGtYIsr+KloanFB
gVZreXgE6/AlBMgLTqqcXLdihwX8nZaRpCbUCafj4lXUYDW2CMnIAisG09UEC3grP/t3L2HYZKr6
fC8fwM2pIgLMvViFACrF8IgmgjvrMXiK3hJ7/uQck4WlAqtx9B8xWb+UaV8qBKWJhBQWkBryk/PL
6mVSJgKwjEX2UCLft2GgYlpngXFMgJIeXzNej7wmQY4PlBAUou5wWyKmNWwZv9nZimFrv2xGvECc
qPUhfrl+OiHAipRRcTBxn9QCo1pq92W41C6niywhXLu+Apn1zrvGK49wPMx4ZpuHz0qav0+HmrV0
LGkf6yPBsvWG/4aMG9QnXGBtlwSzhRt4kug6cNaJDcZrfZnd36wSFOdbH8kK44uPN1LMe8+0QGxf
hs1MdbvMBcn9OvmtUwRku37zGR2nrnEF/lBqrEuWYjZT31GJV1X30hTFVBlKjFKlsq83fvqrorFK
wRBc0pacO5mx9TF6pQB+5uMdACZ9gk9k4W4iP7FcuOKDfa9THUU8ahEkWrt96IZCkS0Lu0QaYj5b
Tk8TGip0WjcJ8DZ2GGvxo05gqbVwg2BXNQ6NKJWY0i69K4cHti1K5vSzvXkYO9Ckrh4sJ9mHbfNl
hdXHBGOJJZG+q/YxPp86juChrNDes3z8gNlt8aTyIJKK0e2bk1Y2lExVUb6PD7Lw2mi9gN9NVzxX
I+bs5kLyQWYNjJXuMog7DpOLzp21TL7V76QYP0MovFKhTfGzMeHouC7PtpIfrC5Zr6AihMyPIQhQ
lSbUpiDWCWiswwAb4BrBiUYhdIefX4o8UkKAPCAucYattYixvnSfaU4qMVYuN+0V66m9/qwnav9z
UbHzxmL9foZ9k5ISO97i3OBUw0mylhdAV0A4OHY8CiLXOFwm8AHFfwPJKQmNHBh9tABAfKiTjLOA
sw9lef/Twr53En4vbxXKgBjbFwlce4oWy+P56XMmQ0xMWvfu2MGQU7txqJ55Yo/EZrTf/FXKe1tK
YbB9j9tLI9P+piax0lX67SaEVj2CI8awrZjwq91zHTpUb5dwYwymsb/96xeUVDWfyVTct3EGLhhR
RLV2LfcZ/vatv6LhDr2e2b0YCHXxYIhAg0/awgJ4YPfEQFbxLafUvm0F/+87/EI2Nlll1LJnYSP4
a2oUGq/b2xaBu+vKHCSG81EGu8Q0WYHiQNzPxriMlx9OZFdZqSf0/dv3yVVlJKW+VBvwTrvk2Tnp
MQGG3hPj2snuReKPiJ8UI5g68/l+Gmkt3NWTYnf31oRF3idgkrX+RECRgFB69fDsIhw4bHr/Gb62
P/XiKteaEB3RuobUyln57qX99ms6GwU7PCoHBTvjB0i38M4DoJgrfWk4D7pgdXC0tLEFU8lfvt4N
IGuLB1kKaMQwbuRtr3BtHq5m9RHViRLUcRugbuOofmJxT71lx1FN3M2zUbModFTXHphLGD+6BeU2
8EujMafxQiGQH6/D6kKrvZ2hWH9yDFKkR1xiGftILYkH1W4bSpcnWr/h9bfUIw5TKMPEEZZvbRI9
1khYwHoVQCqyPBRiGaSQXhCndVKy4EA8c2kgmmi68GhNyYy0r7OD7wVty+7/UrsIXwuZ3zxk3ZsS
TnHPXkusacbCUivy5HI8l7PtqdAKJvMzHTaBycY/Bodl2f+GtDoUa4ehhgN8P4QUffk3fnvCfgce
//QpwtwmLnYnyTssNvgC1UFCvmcsHicRpsArvlz7vsIXkztGYAxjePovLByVimuynkDdnYV4qQt3
SAof0s1oxO7hLv6IPG43DcEg8UJfDx+cFDQB9s7vKUe63aO+JBgMhuC7VeVBrXH12BqH2ItNrhZg
m6y8iPk9HaKTjRSXWYMvStexgrgWl3z0VYxdJTyZDD9/Oni2h2XD8HjUI11qkAYNWr3GI6DrTwja
ZMMWewKKWIysX8lD9+BfOPBAbyB1xvLiI8S+VNBznIzokBcHlVM4ymEfbhkRft2ofyRsoCOb/HL8
01HggsifhiuYQVM49APkZTlQH6e6d7Ms5i8oIOvapoVrGnNEGtuDyssJ4C8oSanxTFAXBzd21/0x
RRFmxu5UOs31/T1J/oiXmbaK9HRQi9mBNVAO0G5TerLR7AdylGeyN/lQPNOiXgzEfIGPFe0dDwrG
DCHM20QoITpFRlUelOg8iEufmXXZHqdPQ5gbPnovCjyjV2jeyuuOeQ8IQk5dEkWN3MYEYYTvM8po
AWK3AK/v+B8S5Ec2I4ymx4Ro22t1OnkoVPa7D+gXNokEv5W/s4dd77ipSfTqLruQp1TPIVeBVCJS
MO5Bo3LwGppjrR4j4XO+QRg+jM6HVJAl5Dob9sDzsa+8VyHikfdMxnmxhbCAleDx/hbENvcm06vN
k0gLCOFFevyGLhLemZT9zuKBF/PNAUEeKiHojHOOeNJFOa+FN05pNTu4ccv7EhZywesJ1onJMi+c
H79Yj2dXgySzx/Kk+0OibZRZxFdHG9V0lG3auJMWmnpi2TV0eT9qj6uHHFGzRwGz4KyQ5YO09Iwi
zNJvjRFf2EYAITEkgZXHGCeGnxBEcop82qWpDCTQAXbXIKzZveORFDq8hHEdQdFUqhV6zl52IVcI
4HcwzKihBouAmqkYvhkQVTmmKObDFBLAhx0n4Bq9JYPMLareCMhFjPkAPbgWdeMmo7LGBTn+MUEg
7LltDkmFH1CNW6L78XJYqTjra0JlWbXQ7CcA8seMaedn2SY00QtGAalYJnbS5PxuFMlbdyJlAWpT
Wk9rllIwiyuTPwoh78SA3QBJOeW4HVpSOkvIeipFpLajYmRdPaxrQm1l5xvDcVQY4gJZ6GnLyatZ
SlciojXN2npTJLxxinS1j2eCyiX2KxCjpR4nCi6xfTYBBQLixt6vKK8hpDzlowxiTcO6re7vhc9X
uwcKYBSPBXHzuzTHL+3Yo1P8Nup9CIMZXwdE+70bQDjMXKRobAZ5q3O6azQp5ZcqnakIM5trVzY0
g7+ctW3f5TVNXSCqDh58YSHB6UNhiqzhL8ImAGt5I4gIs2AOHDomu2fz/8bvbUk52oX6lh4ID7UT
DgKmriqm/kE7qfuhVsB3EHj/dmWbqgxPVpFSImge3RpYkAqAvdlpX9kUyDqzPhDcO/oz/aBOCEi/
lZaeof2O4TkXHmQ8ZKiE71D5Bgz24hyupNRRRJKjSs/VefuWtg8DgCe1DqMddQ3VIDXitKhqkBjw
Pz8HypGzHIsQzcD5abn1IhbgIokqfeNuy8kz+v2NSQ2b72Ux+RpWV2Jlk5SQj0hqT/1PVMUuGleZ
Ayf2OP35BnfykCyvJ+UtKUL50SM+tqBhBxDKxOlUb+fEO1/+pFUVPJuYb8awwfe9BdwqmSWGhPcg
jraVSgVzlhQZTvVQkmlhBbquv8t4xgAlcfZemZjqf9FhqIRU7m9qV62n2CWUPai/1YSIJgaoqT2q
1xisBkLEuV062KbIAzxhI2eZRdVMFa2uEdGzl3fXJfmdp9adLGf/FaZzVApaBG94aC4KwT6oAQOb
abxQHuQUI63zyBEBQf9PHnvnEFMtvSF4Mw2suCtVYhuCk0FCp8LCflE46iXC4aV0X2u1YU+63r2i
t32ebUPUzBQ814Fi6ejXopM8z1MqquBp3GP40kZGvsirbtx4fU1mJ7zIxwEtNV/QnNplsurLvqi3
D/VFBQmnis3d/G4mS2n4OCSi/RnLL0sTubrw2GlebqVFdNDe/Tb5Z7gDeRWky2TJqoBSnJkeqmJe
c6VnDkGY8s7onbVSziA1SISft9e3QDXFhaplE4rZftWHmYrin5eCMzIkwwKYmk034xi91p4jGG56
hI7FlV2ru9RfAINxf2ERu6LstwnpSVgHmRkWyPs8kLnDfaQV9p1OnlITIiE9yTFVWfTunrJ2USmT
jJMzxzuydA5rYL1copzTC1Sy8/mkD2kLkFDNckUH1xgJ6ygYr+DcwEXyUIKo0/fb+d5ovqjJIl3D
3tkfmuF+2iS2GvfYo3IeRQiGwIN+ZIUFtoZNdd3p5aQtzh5F8YXvAVzyO74ZV1ZNzX1vKm6BbdcM
V0UFoLKEZmxM6hihlrmEKCPSbvu4csJKrUxrc5LqT6+9Z2kJ6X3c7SK0azfa74JZsqFtFEUytHc+
fkhFvsLmpfMSMmDTj+vtxIbJjyEMPYTurVNCYWsdKlK6ykb9kxc+00ALebFEXbgEONP7UTwQxu7v
cxeDvbiAPxL/qiguYqefm5BLeQ+63QK4JTH8EFmtc/J72oa0bkAy0nQHduMz1lYk92vAuzKAoKyD
dtI4aeaff4VT13q1V2/Ym4AUoyZAt08sjSMUHnuvBePfUVSsIa0zLrKxeqxHQVzuYg6gKIqGbZ6W
ZYqqw+wlMvB0bkoyrgHUpQ7oH/tfAD5S6+FaI3tlbaVCQ0BKWQsjGjUAP1JexfvGDAxMYVDHAP3g
mcXOPRdgZXeTc1npt9K/kYnO0N7kpfxbuPXB67nQQ28CxDvJM7y2qli+m16BrSNPzLpZh2hCCxFu
yY8VlcMz9Z1FabAk3B4lKE3SqYXnKrphFnhcGPvqAb+cX1nPaqrprMZSCrJ18K2Jo54grUzAgGb+
nhtiu0N+2vDvoEXsH1EzOneTILhvmobxI7IRCjLLkmOzK3w/3LuEwO0J6rq3
`protect end_protected
