-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fUDZ6HEmHGrOg2QLZjpmznhu4WAVcRkP1/I9eqROiHDFHR+DkDH/Ds5i0oi0X3aFgiT0H4MHtPXt
0V3GQ61jr4zLPsxmgjNinD6+J/tcrSUUZOHnKWM4NaMkAv46hmBAQQS9FT95ZdK0tHPIkj7BM+gm
T/oLO1Q+N3QIUdxtFn6OkNHkZJlV+pJHtcMFcgiArg9yIGBCdFCM6ZNpji8Y4s/OD7kjPhqgi0Rv
3Y3+oTFnB3/MC8dvP1kBkA7HQfGostFyTKqIUs98Ysislg9Xjcd71z6IhYdaRyqX0R+naVzZmVJL
+KUObImN2uYBja5eox/SryKHuf3//yH7ZxahNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3008)
`protect data_block
lvfQVzgKt1w8Q3iuN7fuAWXKIKWhjILbbGDA66cOEDNXqA96WKsJsYGDZvCzaM4gTwJcYL3eM9aB
kP4+xbr98fRk1VZ0CDyaDnerQDOYq47jCxNdQVYkEacJy6GXcy79xci2SRDWgUrU5RgyaqqpM1B6
FXV2f5LjnrnFEWyCP703keeiTQ3DHtqIuphHjXRTV5Z7UodICrLvuKMDCHVr/Db7bQfqlhTln+x6
luWJR6pAZEjlrpRydq0bI6jPVMD4kbUh3Mxx1P6FxqcXWOVf43jaddxrvsYST+GUXtLKk+sx56Wy
o5lE6copGR7FCMTXYtxC2/Y4or5XcRjOINAvYRiKsihEv8rjkkzaI1W1V8gaGu0yiakyoemxMb0a
rjqNgS5/Y1pGv6F5Iijs1nIlDUnT2ZnkbL5zXdS/09LEpf7DJekNnrKjWAmWXuwH7sR7qBpPZGCx
yRhpqVwdtw5dLxL1xeJru38+3K1MSEF815nuYGUuV541ezCnTUcAUGm9Z2RyORTITyc+d7orKGZo
zZsFrW8ZpP7uEV1P/hhQmqEAKrc+xuzDeAE1NwmN+xXC/EXHUEaqB6MZ9y5EyZrxz4VI8A5atC2g
YJLIF95vDEhwY2TFfFqH1PJN4J2E0t4Hg2IAVNhX2kYLVvZmFQmrjmSV9TIMPT9tH/DU+SZxdW/N
4XSNPAFWDKAByeD9k2/c9kAkPGs3btNIj68E3+nk0yyABoFAHMuMGF1HSRbsPfH7ZyJgnh+jvL/w
gPzf7xO6HPumGKgF7kwJ030j5nmboEXDhuinD3bTT6t1FB7LIsAdSdark7tpPqdLByp3gXu27thM
b/lrL1Oo0z29lE+MUyBbCyiU3Z4usu80fwW6MinrZ4+Xrt4wx/q1/1tDaYugZlHAq/C4IeLvxvG6
lrlqpgx9ivwdhYwPS/OzYjSitHcT9J8k0Tqf31+CAnjV7LQNWVVovyOwvnCZCRg8rqtMPKzH9VPB
ElQyODZUgWog7VYlAx15ktgigNNJJ2xd8Bi1GJcWQ9wM0Gs5XuMMJj7JB407T06xLKgbAxX3It2g
fufyJcXF9B8u1f7dwPvj1O80o5OfNeZv+Qqj0+GZADSAH24O3g5vdGqDiUPlXYT7dV+E1fmLrjEx
luZLNRwtJB9Iqc9Vrz5MK4YwH7b1AcDUxKOh7+xgrMe9snz/JzqBJEoUWsLJealh4vEgVTX44IkB
o7lPEtL8Ls83qnrWy/f2q4Qu2F+vTC0Ga/8npi2WcWiaQHu1hqeyyMFFQ+u/PomDQ8K6Wm+ANko5
RoFKKUPCuNLegK4ZL4txSe/1jxJTITWkXMzo1b1dJGd42n/0X33++FvWgVczkMyCj2MesUxrKZGy
fF3nWjt1VtZh9G6ZVP7/Zl2RT5F/mmlw+23EUB7B2TglrH1kSoKEZk4Jj64IHYWqitZxqaI/tDZC
DGp6J5YJRz3UXdxlPqCi2ZotUEmT094ECRfs+kmVC+VI97326v1u2eM8Y+oRbb815c+QFn+yAY6c
6YrDLFnsSwHh2QUbvei8OO6MWvsnRvDQw6/FE9T1z1aGAdPTKaZp6K+QEwaPZC9e5vKxZHYamfKd
PJbwNB/9CbkSNT+zO06DvTKckM99+BLD/oXeeuBIfgHt9yBBcoQaqllJCgnYrFIhUsnVTbLJ8zd4
tQCEjL73nJ97mqjwwTsZtZNt/ajibS8osBFxPz7r0z66PZia4hRBduTAFMxCF4StJqTYWSYilNnG
0EiJG0K4TZ9ip8x6Mxx7gsWnGNPoFp5MBh8VQfeIvTOCKgLdc5wtXlvsJzENGaG93YKmKZrCdT49
bEAP7drnONZjSnbdKU389vTgJ56kDMg1noHi/fLeW5e3Ah1i5nLdjzzx8C1b4ppGtRlagy/P5VA9
1lYZr/eZGtWmHuEHlKwtrX6oSdCRmSdor/rPSkMeR3/dZLLehG5odCUPBIbZX60NH2CGMMNpGcy+
7MlkU/zXDdHNhTeXtl7uE1sFaSmuxTwxpvBzTYSld5YbXo82qSRjyxVD/jGIWR+wb99RCkDLOYCg
AU1GmTE7NIZy2oPK8JIPS4Z2g1whT9g+OKndvb76UE5qaIE+FwU+tbTsCHqnzmc/h9sOKBOGytFv
abu6FV4WKWF+voscjtsUtHYvvAmtxq1FKwADj+43FOu4Re9+2NAu+DHYCsekklvOKPgub/+25cUL
dwQ4lP5P4QbkWXJ06KUKZjcMW0ODRt8gNURVF3YrPv0eMHZscihPXgIfoiwHSIABBb1gCi+tKoNV
RCqsjeUxpkZg+raDQfJ/IJjFF2h/IhbfIjCw164ihXd3PL2wYFUVIgtZtF9rgRTYq2SSOjQZv/pc
Y8Z3SDBqpDdL7btwErgUDOkwY06icHZoSUJU3YN6kzu/le4fNxLcXnspEn1KHXiDB5zr/gK0IZuT
qmG/71OVbkZHS3zI4bK1gtJhv8+Pje9+AlcaRH+qg1KYILz4Y659OlSLCd18+/Ko4zH2dgWAurjD
HaRXenHrZBp4LH3UgmTWP9hTcVbzc1wBc/pNuRlBgyskcPjS8Qp9RWJqMNKn3oVj9SpICytTpWG7
0v2zt7Zjwe7AxT3ONXZsjNSJmEJEtMZja3R396hXe4W9k1uG2jtrURrSP2VVLFKz+AzIhLfNVnuN
n2A4qy8GiiV/nTTMrzCyTyHEf/Ss1HyYYDxHWTctjzc7norvXnJxFMYW+batcpT4xBTAd4+mYstC
QiV8qhQodiiJ2ldJcxHa5ZutbZQRhEAmFh1WH78DlQNb8l2Ej9KMpZGJ/XhsUdf80dvHjVVoPfQN
cq0z8dhJ3XX7rqPTIjvHvEssnqTVQZSfBbQ+AXqt54zh9lkLVmSmbeQxuDA0dpAEnRQGnw2eiHQ6
48fj7/0OxY361K0zjyAtSoIe2cAr/MN0L5F5xkPpgRMOcitdyTTc0afImNt4pPAb2y/V/K9WwWcE
XycIbV2t+2ewjOKbKE79GRzxBQ6yn84K/283cLUEA/3FgEhh2aGxNhfTIcA8fFCuqNL4CivzMlby
CZ2hsoxxqaH6VpWiX1ArmxWgTDcVgJzL0R1EAkuIeeKP004LdqmOIAl/i4XL22kpKJO3AvdXFHBw
YpvQvCdLbatBhfEtT5Kio3suT7Sw8aSYD/IQNvAcujAwRWFgvj3a+BRnTnFpGYCgGkrjaWBV3Cqc
ZYpFe9Krnx/FlTUm9SlzTzdYYVuqzDYKDc34rCruhXjyFVbqnzbU4rrmoLMyaq+GCE700bJyVElc
oCX7a7k8s73BoMMsAb0T+S4pKhtYF1jVm/Eybx/r0tb2E6i1YA7LJ78Rm8l/pEuCHlFdFLgIotq5
lW9kkoFdoIwus+z0WpO9pCvtBJRHetOTtpydZzUMR47W/thjFIKArULXh7umioPr3CANU3ka0Xhz
yWlIwiafeBnzylQhibsFv9ubI4bCA4ihds5RMueWa2cxQpQl5st6wDP3WDH07HApTDlaxe4BxpYb
zCtKTxAQknrvwYXpQzx0/X93mGw8fSYfC1Ske32Hm44VPZxc8UG+m2eHI9RmAmNiWwZEoZ96LYzz
wUNgJYAtvQpqpCXsSi5e8LMRM0x5R5zoNUNAkwTZLdqCr+ZAhl37QEAsaokuJ2Y/pW3KX+y11k4p
gAVAvzmhCjcVV4fR27BT/s/TeJYXkrtT1Mh7paqGwN86Ve4poZetTnfMjWCsamwHi5ey8Kzbwojg
tZBdXw9uXhpuUL505VR/D62ZoUsA2rQ8w+KZYaufFhYqwsDryR4gTqtroOnxrlx55PnYWSzeZDU8
aIpSpoI05ghNHMJIRgbBPpt9/CqOwH7ZZw6uZIwLIOUCGwN46qO1uPDJlI2sx4/HauofdL9l9pyb
Vnq272XYqpUsavzDu7c6P1zmF0adBM6i1gCGGH48ru5Psj/iFE6VSftwPbDQh+CtEq6I9qEX0RwB
02H4aNfad7bX6yOoOJvwf1J5YW4SQSI5Q1UgTW9VHPTYOfjSiiA70ct/4g4=
`protect end_protected
