-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vt7KCCT62NBj8u+hiw/kWADKRPmUkQYb5L25XvOkTpoGtmk0wlXEGUTqTtD3OQ894uEXQyc9MFi3
6sU41NDMOJ2AdrNxA1+aXxDr3/JDUKghInYk6vWta1R2vSlvjvgoNtJ+PVNSvc8epVw056CvnEJr
0EQw8BcpBpq5k+ftkYnaxgCclgJ5ZHDGJ67Wwtz9SefIeiT6UhToeET7tEExllAmsu8+1AlEQ7JN
1UTT+XwHdnWer7BIhHo/68xWLmN7ZJftNfYZHO2FXcNnenNDRVZSi/4YGgi8qrgAOObA2h49jUeu
n0PBKp6klL3hu6XOFnnbuOolw2y2YAveF4s5lA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
SOY9sT04XM4AqofDgdGUBgO+hvpcPfor+1T0aQwJA1plpD2n5w5gceAscKu4A29XBvzUtQDWxOPh
XQ5BMSxTBu8pL7+/LqwX1AMk/Li/xzqrzDqumNxT+l3xDuJzeG8sF5rsJ8iSn2SUca2HOO3cHAvk
YNg+th7qxj+Pa2Z2/DOYgVT3PhrxJ2WmWOV8cQb1ARBOhwnG8fB8m/B7xbyoJBm7EMilJL64/cy4
6uimJttXnM5nDJQcoPxrMwUeMZGzxJY6ip5drpXQsa+HETpjeeL4MLXQQUxCBrK18jy9PL8eoQ6D
r2ybsXrbGpCKDMz9cNGX6xokQW27hIqOxH82bIvALwWPxV90c7lfZV9Y3+MFYhBdMQ2FfplcIv+L
Dur0Wntaxfp9/527i0NobN+h0+epKsBoHWOf7tzfh4TwH29zx4pHUvamzCHtTDo8fuje77o/4+IO
eL5JkljcUE4wAzvmxcD1A6DfoPYeiGIZIHVEDCGBsj0axPwuuC6KXuiIQ3BgttzAFPd2GHtuYX1L
I3URmYS88Xb0lZUohu0DL1do+/Je6byS2WgFnkFB1l/JBQBwyUtFh8q6zeIRdJPKwRjFYLTto0nl
neU8KhcGeoHfosikhywitkWuye0Dvg7H0ZnXolz/SXVSN6kgR+4pjoRJt1voSN0ZbTBz4vXf9SnR
keoHNmyKg3OHSyS1W3o1EhasqNP2EP++PGdqSux1gyBj+HWuceifoSX8aTn7fVadp1VpEf4K27di
s5cDSEN8UbinV9DG0iNoO/7MqyvcsVBTrxmoPbF+Sd0vMCVy4y/ZIPs8o5aaLPAeOPnChEQ3NKWz
YXayOrPQsg+JVl/JD49a/yLs6K5VonQpLb4xOAiGVxt0z8X2a74VCX7CCCZRJQ4Wmm727nLulp49
Z2NjwntSjcJrVoAtH7kVYEPi1JGcsC8tnMoJQLLV+snIzq2/dsoEaH2xSBlBY+ZcliDRDp0d6BBa
0EUiWCtxD/4fEz4ZIpz9R2Rx5ZQhcZOyW1qXtSYemUQHgUNkQQZ02QuGpLyFrpNFOocXafFadxlE
WLtEWJx1gJqljKXoGh7lif+Tob33gskIOlDC0mAzMRfQCwBMVxO0V+Et19Re/nmLVYxPKP6MpgRX
0Gv2CBgLGbBVxTs3NsHVefre0kghk8al5KD5lnqgzuJHiv9KObg+krmqv1EJtxGvtQmcwumMjzJv
gLyKz4GQ3zvmcFF09D9GFzzpJZH/rxUH7bVljLifUQ67pBP5FPrm/VgeywWmfBjihbeI3lAicv+H
fk2+JyS6A+vb4CVYv7sZr3u+YELZ/VpSR7rgm9GcJHTPI5K5zEQHsZ3XJKDOy3YZPH9qhHNhS2R7
05zq36qiMGrUvCRPbcdcCiLBTEaLcbTmmh2Xy6cG5zdCOED+dTSxnd/TxymdmBRC8rtivuQvSL7h
pEMI+vuvXNuzSEb5ij2c8ttqVE5eZg2xTXKfs/ftSQtvGtoApkihsTnEoelVysjEMgdK96LVz2gk
5r41SsBkwdJsSjlt62KBs9vOiEi8mn5ty/gaH9kluUCkW8QH5z+asGC2QFyUgPagkk+mLHTYGIVZ
byEFf+mbpwLAMEBDc0xA9hYIdnYLAuyxMfwSOl6+T8LrgABmoqvERa0DqK+rxJFzNMhb7/lhI4N+
d3R49wtdM9AFoqmppt93Mu2EC6YUDALeUpfBMltfMTL4hAOSjpN2Bi8slQRIsHi3eNXTMv13l7Qm
kC0HjSMgtxfTypuocyXyVHXOqOXFhTYSMLu4sCEqahko1LQ9mv0f9YmCvWHPueVJft1yDYbF1Dli
wPZrBIozDeg9OloCi4QZvl2QDzxsCmDZUoS/SlXZvuU17Q+GxgL6qeQ4PYqErjjyx65QAHIV3lId
w9vkm71YUOrjF/6u9oQeQ2B0rCUpimAnSBnOJsTHfiU7zUwFLnUTDKNOil2PKaZRxHZ1ljZ9ZzGy
bjPH4vZYAc4aYeGCmsvq6u25PwD+R7Gmseiim6kNNRcFhDF/vyUV0sc1gYehqaHMFMiS1GJqWGVv
um0CpzLKCYwyo/YrVNvFmVG5xQ+VcKxN32S7EMX44TsznTb9dec364dGeCogVBb4DIA+K2bfDeEv
lsKb5BB8X+ExaI+EvhR7qpso9xKPxW8flD7RldqI8kw3KDUphDfBXSlCk4+PoLWQQ6+yAeNjoZs7
23cx+0DkXSGenQfcEbRzWb3j9Fs57813VagYKz6byWBMCmi7aWlSce0s8lrOYsbWi6w01MYrPUHB
Asy9Pg+Ka7iFXMN2mYNduMxPQYJBSpjH5RtY0uqCL8y6gwKY58k2MubvdTz73vwJiDOeCY7cBJLW
Im4j0owyjxlZ2U5OIllZ5AO+/exlsc+r9sIKOtCQbYT6BbJQ8EVNZ9NVoIxQCR15tQ5gIkPXayoj
sg/GEvimGnYSuIIhgDaiww4bshG9dXLZAYm3FzoDIot3XcdS0r2ms2Nsd1hiMUrDO7Jr2hiqkBj/
pFFasRGe1Aqy2BKHwA7Qx2CtzGVO8RnEXkpN3JZeJW2KXndJTNECLVG88zcwX84Fur9dL8J0GwxR
43a3rZWO59LYeazDFFEhtFN4hj4HP4WsOxeYFpOzBs7Gb78wyvmqaB5fc45AJoJjgxspafZn0OHO
8176FFlGgrExsTW46GG6L5sapgK7KYeiYZ47uvnjCbIBiPViunfU2NrwI6w+t6O7s4dbF0xeLcEs
nwCG8XxNmPtj7Gb2DnjKqPGlFU4xJzf+NVxmNs7mY51SnZ7Uhe9goyuR2JYygMq/v3/h9ZsYUpus
LZn/lMW0hHFrGVI+JvvMXtPFtQuw5eet6cifzXzsXAX7m6JHICvl1Ehmg7l/i44oEaZxh2S6zTvm
5Ve0WTiaYU113/eWuY7pkCT3lhBetah4sOwRK9ZGPRxCeMnoPwS4buNdQnD4XpLTB25S77wHsY64
5kDltqREwFLlfysDcvVRz6RZrMAGPaLzH2d5Nfpv2m3wkxF2yHbpzn9itowU5rgkegIuSLDCs7Q0
zW12z8tJdhqjPg/Vq84b6ow4WX70vn52xSe7w18YRjZtJ42/TWG+cxj3w6qkY0B/LsdUDxUbBNU0
K+9aXAwGXrMpzD7HpZn+hYxqr85Fig9sPr1FssyDFcnIhwslb3D7WSwBBiw7pqhohyTd7mUnaqqN
N1vwHxYXX3dMWKUOYusDZbStdqb+CDVrBcNcgTUUMGAU5rLdV3jtsTl7RNDyqgr0TsUNdc/tc3He
L/7+WVKJFzK6yJM2UfGLNfpyOF+gvjZArP7afpcNgVwaCprbJFkRzGKs5U0wIKUs81Ni6lI9WP0B
BhnDuihTTOQONgS/WQwP4l0kfTRsrbRgUCTNvkS0J2XSbCGJhiphqQmOHZJrDCovK8Sx2MXCe4Nc
RA3sEcSh+pdX+/XbD3MaRmBYkEfY9HeRFT9XjCsBTn82XDFwObxL5SKqL+/SVNxiYqmO8jazcgnE
AKbfB5DBzyBI/8UdfCDS49Ge3YzyGklB+l57/5Cq7WhIPBOnIwE8zpwdHHkrHw9CuzeoSyMsqZlW
kmRxjdcwZEcUhse6wBcaqJu+qLQRCRrzyB+6fj4aCofK+IaGXg+tBMn6pjd+grUxUshlMJ228Ysh
GweSMd6U2K3IzNltEtV2K0qxJobo7GgWXRvmLdUwVRPwuxfJDFKAFKRiRXnnHY3eK0lA6tb1y7ig
n4hV6eEhQZYWtWJnR0+jRdLZulkrYVmggp2r9G8CcGKUPUVSwme+rgex2tIilX5JZ26R7Twkv/cg
1vtPdnkYpAfCuAzCljrPeBKbv/n32GkHSAH/R7N4Qn8dOoWtzEBJiht583EZXKtAdf94fKhxvsQf
FOzSiXwrCx7a4j9RLTxj/fx5mah66HBb22jjSGkpllCia7hTXkl4T2cFs2Lu71t6Y20NRQI75oKO
VSOcstT9ihWBCOgMMnU7FtszPIX+npqI2v03/RCkTrSgNx07z95e8RT2IU8/ahUSeYkvEe41xmsj
7q1+1gL9+1xQ2nXooxGZfc3Oqj/7dcRgl5XFpy4R/eQI36IqdyKx5PU2QHDqW/jKippUr9NrheH+
m9PBOoJxr0Lu14XqH5mjO1kVG4QCe5bSZrKyw2DIrlGtuggQXWZnkJXs4E5XVWKJiaqj2zn67A1V
OAE2ftd+K73CKOMP75uywwQI72cVrRRsq9eNrZv+YM2l7ctXrtSWaOhW7nitSwZOOfkzq3DLdyBE
wKR6lEEZAPqEpTSz1nG34acIo556wKrVG6jGDJq4IaM1RHj+U5n8/st74Gjs3Fxu/0QLM8gBXbpl
19suKQT8k1Tn9XVZCpoSnswdwIurZ1g23mvnRo1P7P/GQpfUU8+mYhJytRIFl7tksQVniWFhg7aO
6NABS5RlDxbwnymRWMoU92wxW4oJwJNIGfqGGCl38N+aFSWfhzV9BrlZTXXzZI/S9oUK403hvAf4
l9fRfb6Iuoi0e8krlz5feb3zPCB3JuDcgNLRDx4lh2QUaHqjVxIYyVrqOVnfu75zbsveCW31AVb2
EP1KtRDka7xSV9DrM4oaJGymzKcCIZBrLgnzB4vK5v6m1Z40JQM76h7WoY0b1sm9NBOWBU1ztsQW
D9ZVLH+l0X71CC5kskrPbgkoGL7gX0YlWnnwCa9lXfUGhwnnMWanT+jdsDZw3kfPTmEVyPVeCGY4
S4gd+DP4+4NRiWWLjzQ8meNAhIatqUARFiFk7dT/5HAzdZ6yzT+HZZJL02VUcEWJfrf1FjCbHx2O
vQ585RAC86lFjjaAeE+wTpQ4P2FLQNdVfO0GUa69WLsGGdPLP+SHqUsRbaradawil1nnHZxUDvKk
sjsRL79UzKeYq/MkgOHYvjFCqQ2XDgToYks3X+FGW9W3k07+Q8uAKj+3btsftnQPDMJHXvtSAYAJ
0+hbiSFalXqcg8U478A+dyztVkmHLd4Bi5B3hW31zchO1GgB/64J//3EDjLk4Uj7oFCx/q/cYoGd
j7YUtJVxxGXHRB+nxsBaKgUM1BzfV5EnsfmV/VeusRI+xqmRO107HmSf1t14L2E77KRYY77Ezhwy
oZc1sonRsM9IjkdoccS3sX2/lqwAZR6fbpjO53mB6DQYTn7Bi1g81Z0kfB+FODGpXdKkCb9wFaVm
18FstF3fnChPqoJiM86ONcTuBOH/DUYqZae6CzJsbqMSGivdrBwiWBARPkSlxuGxmZr7V2zV77D7
VqnMjXZ8/wZ3jM5degEHYU+DH3654PzAboZvj5jGiwfIhxm4GnIw1dwSmrzcCM9225PmIK2Op9qL
LU84/k+qKiFs2u8D8aMOGbB0p1yXmmd5ca/GUe8ZLdrsLFJZJcpNNjzpmdDQC2Gu/0rGtDlIDvfz
u1TqBTegFHCupdSLB8nvZ+yeaycpbNJSfK4ehle3yYWPw8h4MvcwxSdgpZ082i2DycB+GuHTXtnX
OTdFdw4ypPNQ8p/hpOyjVYaeexvFl6t6dZM6qn+Pqank3M0oGY/1jCww0Kckx9f1XiIizsi7L7SW
4hwueVTgRdxqIlnWTeMjj0LolN5qBJQVr0Y0LGdeJgKVnBuxH56hRy92Onp+ecTbv5KuqG9aFi/Y
4llOHt65E0oBpzJ8rluAtCQAlhKTOBFlsHzW5m4cGyLHfJrfm5ZR5BwPIqwQdq1HgK3dKxhD+Ujq
vBPuzt0BM8MHoKpeR3NSSLqtRQru+qaoXKf9bY2FyLSboK2lqpfV/5d029snAGSeqXKqn3IEHs3W
mn3xolBuNZ1K6rFHa+wm2p+g9d6F7dVtdI00zYMotUFXF/oc0tke0+Js4vMsK41+s4EqaQlQ3x03
aEYa14qy9+xDivgoNCk4rFYz6tPKwjD2GbSyRiCjHG88k6FB0PySEy2lnE1ITcdzb2VudCFcoRBF
nf0e5ivO25nloUEhfndFFxiD7SWY6arQgiJXd97DwFXjGP28T8dePX4Ed8O315gU4pfNS48XXBn1
TWuB0YR+2qR5V3u+KPt+O89YMZfmxk4b1GI1daewY60ogZTSeSlGGpP1R+vpJDjGygqd1Ptz1aqB
TftpT9Ifbhs3NHLgXrWs057VgOS30WwQQGqRfhU3HFWK5DXzi0ReI5ONyy6KM7O8+3c+/bbxrMRb
Ocl1Sv6JVZ0KfAVKVyIqpRFJ1fjvaELoasFcedO6PbETuM2a/xyK2Qoyh0LAw7TP3k7jTC4rzJ1X
7Y2QgPl6l/B2A86FYk8e1GoWBcyZJj4f6ewvq1svd+ShkybwnRnoieQztkO+npNgPdZRnWo8+DdH
8rsUwOcMgvmIE16CPeBXlayLAhO1kPKNukam59X+xHSBGfc2Q0oFLYGzfs5qP2yTrFD7eHGoFx3b
kpR4PJC9hwv33chcbcVygh2gO/mWGm5H3NAnBEh5yg1CXC88YmtgjF+5bPXd5bS5UIfB+gVP+ItJ
PAXsX3KCKhczOrGYuuYX70wAAN9xyck0VvERvWcHkIjgRFMYDxSZdOtG7hSise4oWdrS+2Eaaz69
2lVOKeLHgLHpvlT+vmxZPePoY98LVZdhr9utvUVUQ4Eudgd7bZV4StweYpJMGMVu26M7TKBoYikW
KngvBTQToL3AMb7AsgNE9DYA2/QOOgMf+lAXw7vpGBAdl/tIxH1iu9LVt5+SyZv1weiMNbxBOGU4
OEica8sbcfhjB2mlONSRM12eBabDEnqhxaJmj/Wsxif50Y2zGrYL+m1RpxBRnZop5uOdwQRRWJHn
nl5ETIAd0NFW8nkglMnmHuRLBmh6jwh5aDJSMUZ3qe/7mha2yLlSqoGRg892lTEinD0ipBoR/ZSh
X0i8PySM0gw3e8I7OloThEMPkf0t6SP1HzHDJbl5da67SSp7QoYP28RgugXVq54eeiloz4JqwxMk
PiZH123NUx7IiBTOksVC05rrAseaoWfODY3DRPKBPH+dTz4YrhaL69bRfZmgbXTWap1uBLvjOP0t
Ufi4MwnFGu72bIq5KQRAEnzHPKi5EG/yUspvf0Si5x9kAP1SZZ1Zbj+ILzjov4kmFDcE/hhvBFW1
f3Qcc5/xM9hWyHYlbDA7Tvg0K0zOFvnolbh+gMmFO/0hlFewZV/UPgVOTo7DBC5OFhyNYKNweute
XhWxdvBbVDpRd76ZBfVFnRn+R1erjFARAh+lQ3MJLpTX3ocmj4TcHI/Zu/WEXYzcIAab7Kn1OD0l
VYmT+VvZp7r7Qjgy8sjUG8aXTCrXV+fYxKAkXyPyl6RhEC91ypBKlgYThi2Q8HxTmDbdTHR+gyvf
/p2v5bmPWy6zw9CQceOVpgokDkyctNXewod+8BtoOWhsjT9IjTM82POXzHv/x2v4qPXZmjsfUKbd
5V07HyP9KvwmUf7F2oG/3rv9wjvSukTaEzESRd0i2+Nsd569SMWQbm+r0g8NiMKKgnGMv9R2tqPs
4hvzclKQ1N53oKZXo1rt8meZY1SS3CsFxD9s7EG1z0MlAWAMhdTMEK+NF/v9/oTlNM9xYvRBBM1b
uMehWUI+7J9mtDsEVP711I6WyOYwEhyH+4NXUqrXCWFUeyxdwQLppnAGGSQHSQy3OKZ98lpQhyhi
AeTYjHuwWYQgPuBzd1YxdIKF4zvXc4nK1hPnD2CoB2PWuu4+PpP6MIPvFUd+B11TJZoPZzVdXlbf
J07eIYNCFHeIzMmYAB7mWYh8p8BtLaZVVfQH504yPzteAXm3LN7WvkuyFSe+U4ruPuoxbXJimLQN
yjKVhA1f/iIQ52mGR7jmRjH+eXlmUwnRJCqws8hWCGb9sR8AOAyqvsULiwbX97hHBo4uaq31wv3R
6KUx2Zt8gAodPDHV5u2PlJJj431CIepP7gORcWkr7jWm69lgFC66CGhBuw4+ccTgf4OCe+AxtEOZ
ztT2BkRfTJ08H9iF+QAusuYTeGYmEWdqM+N3Yt1KGSt17USFj5GNSw/4m6/b6/BVZnasNhEw/iye
ujFruvnH1hkW5hf6ZN0Sr8CihERPYp1Emlj3i6pAFcuvOrzNe7jpvcIWwEmmCp5pMHpXYxoPchO/
8Luf7n3gTqok1Pla3PTcYVHMbfW9FsecObjn01I6PlomUV5E/AEuxaH8bg5xuJO1taOTCWkZ7k0j
08uS+h4zgjhnbQMJfKXpT1lHRel3xpbcm09js13m0QBR3+Z13fvvl3knPwRAhgHxKKiFzhucEssc
VaBe6N8GIe7GEBFzxO+o89Yct7cCLa4GQ3d8XlQHX16ebTAU7pEzOOHOrj+3yK829iMwIylwC5zm
0jJihIXudL30BT2SxT3DZoB8AwobMcfy6OkWtbQJxn4JAMYzzT9AoV1/8No5+DU+HV+yXbxPeK6s
FFQmvkl8HTRJFHDgw4UvORNTg4SiRKFKexQwu5vRX/u5b+44bwRAyOEP1QWA3eOwQDSLBx0O4E2Q
wv+Xd5UI74rM3Se7zzU97bNffmvkIJ7iiMeNbz8Bn1+kp7gxmS6HN9JRzk70Q7yqboE16NmdqHMt
b5tnys+BWuEymRCSiBbO1jZXiRAD0nvkuUI2GbpnRP1nv3a+C9PwaQNW6/B1ztuIDmjxRdp4qrFI
KlN+EDl4keHrfy40T/o+4c6dQKlqmpMMHBXnABGgvzoC5XjmVZSwRLtHzIXlyShXKkpxZyCDMfTW
LTZcwLL34fhXrDSeY+CrU1t7qx/yQb16Yt2NYjBdrAMNNiWHasb54620DzG1jgwQipamgPRnJiyi
Ku+dLfeGb+clm/aeRtk1SQ3Bq62wxkXDcfj/oJxfeTovPi3qeIN/skdMIOMu1pi91Hz/qP7fiytP
ujNThGW67FU7qLIp0/n3QImCKTNiPEgtN9eV+n20Eu1/v2m5RWOt9asERu8jOqw03BL2Fjd/kcyf
mJFTjB9VSTNw1o+WkpfjLR6gjxpRv+7ldqgUCuhZnrGzTGZDuwquIFVBQywq6u4b4rJE0lv96pxf
Dfxx95i3+ndhJlIiQ0M6LEbMSC5fwXifK9NsIHOghbNHnCmVtd0zVkD8fDAC59UxKLLKnwxRjpWb
0HnBZoYvq792nHblQj17mJBiZmbGF+ZtbH3R1Q9+Lp6PcctV9bas5IYWgLw6XyBUkgpElfMu+DHR
dXLXs9vLoIkV56vmmiO/CbitVfMcSBHODwRnRV0r8+Sz3IJhYkHLXnYY7Ns2gycG/HMnM86F5m/R
kCBKcIkk4rQ2M0nkxU1w7IOEt6324ackpsbuoJCadGNc9YNykXRvwU/VonSlgtjGsKPvD2qm5r0x
eiHK/nKZMPyDBwS1d9HvmmvMqkruQ2BDe4imXd5o7aUcqIZZ0MKJ4eaRkdkT2dgi00qJLNP2b94b
YCSHTdKk/eSf0+6T5dPlqpWpPudHPAna57hTsnpNfReLOe/yTCA0DcOSzU5LjKuz/rI1cXK2T+NT
/+viZWK1jqPJQpozsyjqZ+f4mrf4OCuRuFdc4LueG7yhj2E8d4mz4RFYBzCpwh6Clle+H7ltM2Ee
RYqn2B/M+ujC/bE9y3sG7joOrAEdlAilYlqXo1njonWosNMv69ZeAi5+YV69cZLBLlyqz96YS7iz
4G/FiaJkk+XnM3pJ6acxg85sbzSfIR47zdzSpT67UQaBivt6D06QbQfdOACWe4ZHSj2E4BCpO6t3
AwAkfaWoh6EGac6v/Zg3pngcqF8oteVAabMR4kCb/G3bBiY5jt5AhFlkoeC4Qr9Yhh3kYIL21Ky5
bd7HjugR+D+gVP95Mn6Z3rEZ9vj6mjxrd2Wh+GoqFluj/h2gVr3r3eht5BKlwBs08WdnoCachDgR
hVgLqRgU9yVBQIuou05dOXRV2khXBkfoG5i/GsqCofoHa8Id2zLj0Sccao8vjCNF7NwSq79w/ZOK
0x7POkGYCOI/RfzKm8lccldZsmCoXPJ/reAy1Z1Wz+nZfqHZPyuSFiz4Wtr35SYhJ/eU2tWf0LCM
VAOv9OsNapeU5wfoprSaSFBuIIbTV9shpZRr4tJECHvFT78G/puxK/1LRG5RaiFAxyl5s6heniMz
RMKKeRJ/TH41fY5Tk0HSH4Ib7prb9SNTlQoW7XflUREm6gY/N3coaZ1RiFIvm1cFDwkB/U3MGD9U
NGQOU8pdpEwpT1N5ewPvRl2XLI0PYcC20LafJvP7HcPJ9ND0JUV7lWD3jUfp+ksqROkCOCV1M26x
vDKXgUNMhySrO7/7lj8qa6c63r+AJJpy+X45+iSrUqp8TC/60PmnCfH7zYKtjj1RwBarhtvaB7sI
bLlfZjpcaaQxyF2gnaE+f5Lrsd2y1xAefLZrSyEJl1rXs9aTpM944l42Q9KsTSuF4Ishk3sgRsdc
2KBIlswInnN+VkwnqNn4zUWJbrHobHs0kwYy5xvcHVUDExvBf77ZE+k8XXRVj9GnK3lob8/Og1bx
Cr1iTVrd9XONh2hKDCPSno1tTw06rX7EKgoI1jpaozSHcNPnlwdvv+RbI1r2WB/8SksjgSF0PFdM
nGNqPASfsVOjPMcI3I2KsxwhkYZexx2rS6J8hQ6NiXV+uPb1yjaE9/Fd2X/nrLb5T7jDVNji6Kv0
4/vutJc0846BqWcQhCxa6wux+2M3CByWvFVwiv/g9S0TeGNCrft+ytbU8x0AuS41+jgqW1SXebGq
MygNWkFhkgIeblzsqX4NfxFkxQ0n5gDQtWmzcbGyVhNdF1Oveo7FB54WTc2bH2n0nIUqFJmzb43N
fTd4Rylox/f2TkpHt2JsJgEwXrdDXrc4CYGDK3MXppf7xhtn4PL31z/G5CTbXAnufcV8B1CKwz9D
93QWR8QEa93i/F0EOzenl42DJA4xxXlahWDNgKmCMh9GvO4DOJDTYufYPqcKygxHSn7w+6d6+dct
sdQFiNtqoCvlEjq2hRP+oM3wsLouUOq6womkxJ2M+aJ6cVhJZidHNi45YxSQvIzA1h5Kgw+ojtSZ
PdiTQf6ykJeKqWVT4eU459swVVMWNq1cfXSjMf6mbU37JNzC9jkGHJBxHEurZWpZbUmvtDA4DDni
o2t9uwWfVsNyz5rn2oamD0ZGTDTsnzMZyBQogprynvI1wSKIY+4Q2NaHAA3ob2Ls7LEOzAz1Hrfe
CZ+VE9ZYQioM99/RFfLxYvJb7Es6AvDVTNT5EU8i8kBrVfueLdoOmINKyZm5d0qZjqwXuTLNTzZQ
US6RdzaEgieqhEX5EwoBc2AjgKTXdYE+AJZqp4K4M8kOCMAkrYdISBiM/FAvUiSOqa6+zL9adgC3
rS3yMGdZnYho/Ynu7f4BaoW5XZM1UYevY5Hpj+riZGmDxv7rvnC3PkEuyprmkTgkxKz+OgGwNxdG
mu1BhUvklOKDcsHq4oboGAA0OlTASgtRc+PvdYkHf8p49OeUoO1PeelV4rIqCIt8DC2MDFDEepnq
dLvQJXdKIQ+qDKs3ldliMlFOyZ/qhtuh7TyafsRGEviB1sF+TsLBqkQzIycK9q4SmbXW5Mtbt9iK
BCNc9p6e8y4ZTax7Lrx0ya0219Cj74Dpoy4aWDa0CmYvBz8eoEwEaK8ZbWK0RLO4UxxFVskCmL8B
snla4gLAeCrVUsWpIweCTdP2KYKZWouuzJ8EpPrYDWTOJxhdhTddTfZa91jntgafx9dtFU/6Cr+S
oTh4TMJ2QOSsEkBqUPXcIjkuivXBDD/1dtv9G1/8vkQg1u8MP21DgVuymC4zjX3r4oUeHKXylNl6
XN4w9EWIME0nDer4BAoWus5K7ZTcDqFd2b5DUjibqCOfxqMoLDdKbz6zY03YMWmYcS8JJYwW4Lnt
VsXheRc119DVYC6z0C1K7/NSd8rzA153ZUxvg878Eb8he1zl0qtxuuv/jPjljkdayuDaLKcNA30F
YP5hctUBTVE73O3ATEfmCFlN7qZyM6ZNHTQSIQoSOF6sML4IOC9Xis9nAWrlMMPkeu1W27u0Z77G
bdv5/J//K3O7JPKDx40gXOI4wg9pwBCkMkReYvmxCRQbApy4kK0uqjugC5uWiZv2fXmwHtfpyoSC
CHqe2C0vQd4EzAnHIkIYp1QI3tngQTOo8voe9pmxFAUl8utNHh8U6JAZmRHuX7GUOaIMJYuSDcbF
SnLj7huA0epkwW1Yx7d/ZyqiiKaVjCZbJX3Q8tA7C7C9Ofpn51YVpSnS/sjI+9UBl8BLo8eu09ul
00MTuRcCFJYy1ANp9RQKKizsvHZIW3oJuwlF9D8GXAx1/LV7XU/d0yyuqhNbW1gpdMALqPijLtPy
UZHm+nJ5p/ks1A5CPDW7+F+PiwFgPe5Nxlx98AXL581rwb1hjnp+LgK9KRcQyFQ//YKvL9CxB4/1
Mr1Jc+Yrae9JCA9wVI/zmRzrddkMdU6ZMj0jyeLv9lYf4FK61zae8w+45eoeDeoDuq94zQXd9yC9
MRB6g+IEfaSSk8Xtmm6SpTJyNLSk0FW6WJOEd6gM/yh1jBM7zaHHe3mRKFHNygNIInvaY5ivKAFj
oMppn17q9Z/ENfhD9uDLscy99OcGyH3G+fZBCioY7sKw1FqL3UIv1lbrTER/OCrwoAxWGiQBeDec
90eTOP3kibSb+cowH3Klm/tqepMQnZhY39Ef2YzMtJ0W+znE7tR2TVCp6p63NHMG5cDT5TsQYr3U
1w7deXi/4IF1lH4aXvcVNwCyOVhAQ48oFs7UC+ko3h2bkXWCru0kxA0tXPkkqS/JcYUJKavaT7AP
IAL7zPvcoPQJRwM6+djgYkIdAreKj2UU4d09tbjacqk+INyPIMxCm3UPOSPUIZS8QDWf2BncrIVe
tti8aittkaXBI2NzPhrfsR/P971fEoOc979dgej6oqgQMkqTqaNnHglyIlJoBFUI5PQfV1WF3sIi
Kr66lKxarBMaowsrFg3zR/IZpy3rQhs1L+08V/plzmaJokydit9IdPUrb3eYeNJTzPpn3jzKp4Bk
gnbD1HKbBA/4BkWTJMbOMgoaDbOqqE5K8QuLJ1nFsbtEhnvk8KoJu5FGv8PftIUdxwfyfkKVgzhz
H4rgxz/I+T2fHyu/EPDG+ceKuHhyzI4DLzaIjEa7VC8yfUPc2p5MAKHE0W8FSTBTbPun08x5d2F9
ft3/EbZkQqEXxbZdIZXKi9JA37A/MmagM8OKvCgDVhdWjnaO9tqfceOLpg5MbrYY97PzbtH2rOKJ
ZBokr5GAONbBctCfakzs1oWnKLTgA6xXtDhFS4Oz9Zy5c4cvMHPOl3bMuEd6tPAM0KJKY7RbycW/
fGConKikoSjqPGJJ2vUs0CRABryCqEwlDjQiw9q9gdZ4UFoCkX42vahRjMkxm4dwCxzJJ+Po6e2M
kbriFEZmEq01RBTPsM/mTzj1xV80pDrVWqpXLjYbLijx5uTa9V5ph2kI60deWy5KG4r6lTds8jCe
sGecjIpnTPF6qk7vvQLrTo/rVnH042Q1nLkfwRLjdUABOJa56QFOHTinvdQu/Tx6BvhSN0xLRhYj
mMGDEnXc+XibP5LQ0lb7weea5BX92v/VL9x3wfyvGT07+cFtiVydks0jlNJ0rswoudciQHBchky8
k4bMjv5P3WdGCYxdGW4yArL/gYTIIjOzYyvIKLSYbcm88ZL+EGkTQGszZTWUO6IGev/I/F8zZjyZ
hMcjnaXKdFcNpGIktkWaI9ZZX9qoQDc8XKbVYICWtJOjdOkgZXKsvaXQ2sFVJO+tqiu3/V2GLubr
NkcB4eucmCy76a2PheUT+oyy3IHHmx/xsZHTdLnw9YcMkHqAGlBqN4jmQJ5OsUTsWuQweZ2Wuc1o
Y2HJEosOykVjyaEx6EMzXrd0All8ZO6LS+NI0anX7yniPvygfJNLb33XXG5s7G9o3FjTt9cQU0o9
VQnD34ByMKv7QOnp9QML9QOT59c9/rH7J85iK6JJFdHkGe6mbvnxfoD2L1uABkwXULLAgnDtGHU+
MJB3UpjO326u0q9RWhO+L76BtSKsY1IhDsl2EN0T1nLoUacCanBxE5SrkZ4IEXWPxO+Fa055cjrD
csONFwFoXkX4X2t0zSWa9UP9I8xuJ+xgQJixUkUB91ee0mgZ/OgeYlOLt9mx9FIWDkOSgUXHJrS5
q5RGzzOt2jlujpJjJVCLR+MV/k9oCryA0wr3WuDayBj8FFTreDQduz8makLc64NDXRqD5+K9bV1y
usUnxseHiPQGtu6vIKLCFOdfWvyjf4qTlZPXAuTdQ1jR13pc/k2qwE0EEfRbl2iQ2fAevZoG8zBq
W+kB4Sti2CZlx+Twl+Cu1N9gx44/8pfpt6BEMGpG3zClUGr4QMzHsPVbnbF3JqW2FEulw+y5Vn+6
BLYFUev14Z7Q7uDVY4MbVOfGcKgpPTC+DZ3YE6uKVSFmKqko7IxlKsNUzGK92bQXZm5c+m3oTDYF
fyQMC/zsTVjpmO1gDy8cmWIjXwlLKPNiB1/YgdCorWdyAX1+SDEr6vRqDq1wNaUtILpXZLlOll5p
XSsxZP7kXyHo0OdINkZnntucLYExziTdL/mE/IuFFPbc72gN9BV4EGcGE485MWfRFmKOvWHlo2Wg
UKpdbS2Pa+e5DDbJZ8Tnt9dKILid6J61THQ/PfHTZEPsuVVG5bW+9ExYRw4PH1l3BTVq6f3XNA/S
CxX5IegZioHoBGvqKUgSyCj/5JK9adJb3kB4raSJc5XxoBJovnT+P4G9nI2/l+IRh3Y6liBY++59
X/1VwQTpvEwo0OA+EYZOkMF4CWlKnS7bn57B0PpnUBKUZkPCZvr6YRbsJqrNzvpNsI6DZJFq1BQy
2TfR+BPT2qAwdTsC/VsMKx58I9sdbpoxSgPMGhvxztXqcFlHjL83LdzQCuja3ypEgYIS6UeZZsTQ
PXzFnCzfbPp5PtSJBU9cYSL1HtsipeCHp7xJBGy50UsKBNhVqWemKB2VJW1EO9ywNSLm+QDRliQc
MalkC5mrcUd0L5IALO6x4uEhOz0mTJWKQW6GKV63noUqvJ9jU5RAIWuwgzLZDMWOdByekFZLViWB
YSKufIrYOVQuXSDuzVjSeePhKy1MNzPBRs8lE+JLn+poyX4lCa9zhDqjGPuf+TmFTA+P1GE+14NP
tH6wmb/EXsFJ8YSQOJ3P4Igryrz9IORH3uOY+xrrQl6R5MM7UsNWe8ety/Kyu22b8sIGMyfbKJhO
zwP6A4aV+EBgJrvygqJyZWyS+YI4zheMb3Tm7pcy4CJiJ9ZGrwzE/qdbP5TKkd+7/frPcC9nU4Mk
qcRiXuSG6o9HuEa0Iafvz6q4iZjCkdwjLt4BYpaXh/9EXrVfSGo0K65XaZnOqvwboAUtjD1ssYMs
HnAsDpcpKxC7Vx/uHOpL6gkXcYjOJq6ko9brxvbpRh9zwVmgAF+WgVrxRw9PVqnshzxnmQ7tIslF
peCvRdljxOf04Np4kfNt1UW4pRmIhTI8HQYqCQAYqx4nLTpL98stoK2x9fDBUFOW5GVeUNFcxLaO
cem2ZuDW0emUAHzVj3yMyg89FaF2Ay01uYsURhvs99+57lsd+oIXcTewCXQ9VvLQuwZ4lGOmq5kA
42Xyf8Gx24FArL1U/5A8kRsstxSkF0vda4yuyxDiJnY5ijHD7kn65e4JBl64T7EDE99SuWq/TrmC
i3YY1Nhf2a7sKc0TMl0oBi+k55DgonYKgKAMjCiO0fTtmPn9lSd0zf5YxB/p3JxHMX4XTtVpSzQw
E1n0kQVwMeriSwXEJSiyfeenAsbLoIXcjjw13s+HKtgNzcRBB3wvEum+LJ680iQL/jpGj7ZKIml1
wQElgptsGWecOAwlOyJAnZV4k/3I59kKyOm/u+qL81as1UeNl0P2z5312EeA6SlQtUU3EvO0hsHT
DPwD7giE97JlmKn+qm2T7mhlMb4tHrTsut1iPBBNXYWMkoMOhTS0GrqfuH3J3mMjh6RK+QhgVNel
eCvOB5DkjQLxJ2SQxwekYjkZGE/JZEEmKfYDA5Uf4NyYq7Nz3mXwbYtUkhCpcG2zHnYatAFfiVcb
iQOyFtKk6LjDr/Xj424ukXKZmy+nW0Y3DyRzTxJgrvq8qbjTkk9SxWv6CRWpcwdxziGynTb/xBlL
dcTpOt4cC8TGlsMCM/zM9UdNI0XXXUbtN/qlUx8ACQQElRhjHQS6OpNFZLbintfFJC/uGKhH9iIX
WuPXU52sbkvoFr4rAhzX1yW6rzcxbV1/s472VDtIe+j8VQTalvu1gZ+GGoVqT2Vzj/UGPr6E+NvS
uUNs9DdLSpVWwT4mAF6uCiPLT59Of84u4wLhQIbSxnRrJzAwZf/Rsj+6i+dAC9hnRJCbgsfpXrcD
TmYUIyVYPfWOZCGD0mRffpCVNBDQDg+Il5Ksur9apdQBbXVTLnAqoX7DCiB/2cKaTGRDZb+7tHML
ToHzI691hQzTDPvpYTbzttY4IHN4A2N81/72oqGbGwJNioFA/wo7TFwHJBGNE+sV7PLahDE7qkPc
UM/MukCwHBEqA5QOCRjRTIpx4wBvWzu6YWPL/yrpOMcSVaRlcOycz4q4z93+aTQujW0X+nPbUsO7
Et0khdwFs3dJkL2GtnV2PfxygKkCsTcw23r/4LfWcCeUFVgLkla9Yt/ARv0EhfHgYud4nxkDt36a
KZEj15xkrigw79VBt0W/YMGvzcza772zSzR3hqWn7z0UKWfSFDswY2aXYl65s7wrOdAYrDe5z/q5
M6Ipl3PGa0KcJzYiIF7ryHiHCylX9mvVLOCWChoXXoKXlT2xGU2dAZnZ+cfaC1v/Rdmv8oqtkd1a
sOVZDmVXZ39UW/MC7jzkrf3L3fa98mMA1C5tRiE5vLihJPD+sMV257r/jZuiHtiJjEylLzbCrfzx
+N+ipCWApF5G2oJOCLL/N4yYZVJzgWQXIPclx5zEbPTNEb8vzO6Xb70KkJ5XDwGeGvZWhf9+UrZ5
XvI+/EdfxF/SnHmW52AJt94cSZ9e8xVc84/DHCwxT5QsNqZjhoVQmnzvhXYeY1dBFPpQ8HY4auEx
vJ7iJuRzIMO1Tw5vyVV4jmI6OKaiDr/68muBGNFNFe0yClA6bdI6313SuFYM+NIBFMwfHSQFZc6K
6JGBgE7luKVVFcZNvQaQEXLtX+Zv+Zf3UQs3gC6+yH7a+qcUtoi0e0/qs+665ZRP2BJgiGYjvzcB
nof8x7xikj+cfEm0+lCEW11RLi0AcpN2l/u2gbrxb1Aw3CwcpBRgs7k+BlZHlAt2Q4WN1o1lYx6L
2Nbu3YJzWbSkLQzb2n/I3FcLhk7bt+gw1bK3i4SiiKWRjOz4rjk9Y2dWIBwUqA1elJz1xBrv4K4O
/U5FNIGg+cqdrD2P2ie4uQLu9ntN/DU4O7Z3204NB+oCPjGmuEdNZlFomh2ZBE43m55nGyL24H++
rXQDslu6t5hTxAzd7HqBkng9GB2KR9xeWJ7pcKyHODG8qyqd5PEPn7lTG8ktaahux0rQ+akmAlmM
UDhIw5mw0+nK4yZIO/kwCFPtws9Awa4ydlYxVjmhFrJiwD434C2ZGy5UfoMBmGlgjVm+0VXxDXdA
YnNK2tH2XoYouiTb3ZrBs7H0WxtrDsDHtNVcUVJO0FSu/zdfHWhL2ySGp4Hu9wZrhyXVKt2iFpn8
T/XB1L23fqiWGBQw2w41+m32Bw/p83KKimxdtZ89QxRgqAgii8ngL/UEBEK7MlRoQdnjjGf4w5s3
vBPKWLggKq0hZOzNXDnMGpexq1F8XN+bt9hISZASBjp9OUyW8CfJVDkpO4ccM4ZPHprSv1yZzOhU
+1maJzGYDnV9x9F3IywJg72UDqbG8jR8BLnsJ8hoFkS52NggS4sA/iqRuj7AnmkE0b8awjXuVEQZ
xls/sYkXplektqFnbEbJhOvbbt23YFOm1iuVu1wj7igdp4B8x81A2SasNmjPF5Mzd5AvOyOs4mEN
SDX+Ny4vaLHJT10vm76O5e47Cw9bazzvhqpfxDm8OxIWFsETi31nl+DyLWzGJl8bKtSl8MjMEN0Y
ENgYqLJZnThGe44fzuATD2kgVjpr1Sbnxr8bi4N2Wf4TNQfjfkFJ/VY+a0MMLJSNmKvr3Nk3CqCI
vKUNn6WYLMiCGZCjpb3VehahJS+foewc1qHUIYEhg0Mf7flwdW9kBdAC8Pj53sXhTQLDwW39U2/P
CGYVhdsD8oeKbNQPS2QncvDm5fweiajwkZ5kywwyAOFfnSndTBjE0HXrPq0lYK4F5kQnHvAgrYsB
ZBTWP/qThCehWynK95xV7Sa0Oq0m/UEeCkDxDNLxJRl1y88d9e6U50kq8YKyQmMREUPPqrPxMCrT
LO1rvhj/hc/Rtk2WMcQKFAG98sfLHtcaGTDtT3lcf7dQmjFCtbh7E6HHIe4fBF0iaa5SH3eV/fgK
e9F2BvaWt9IbEoly/U8TmqSQuSLQzrj8+ieFjMW/2TGqfiXRITPnkxznD3lIq/xisyXKUk9xTxDp
v9Zsi2ZAgBPP0STASuedV6+gJfNHKEULEc66FKcqiBIWdy7Z53sBD/Z05Jh/m2FDsWhpvrpi4Cps
nIUlutCNwzSo3c/gjmA8s36p1keHslLtH0u5kWG4Or/GqdiZECjCIsVoyhvIFPYvqk2bvVJGcptB
BqFGFa2LfdpD1n2UyK6w8EOATPExhHzSs/UZgvYTV46kY8w/G2Yw4d9Vzlj+6gzynPqnrArSslgF
nSWfBagvBsQFhQP5d2BmnzdMZ33MWXpuWc58FhbCWNgSWyVYQeOvAsWorMzRFvKQXQxbgrNBycN9
6HPza63A0HAkSUwGszWFD73D5vXGFZPy2XoGCVlwxuW7pF0xqQahPH+AX1i4XfkoNPebQQlO9qWe
r2N49+AIYoEMCKs35+8H/iYE/kTHnohiWxHU2ex/NWBR6cYR/E5cChLwA3BSIiLOpTmQBcJmDFKk
m/o9V7yjUVA5+zVkOTIduBCEFxfzdhTaXTYUqX0FEo2kaJvdL1LDgPD75Yuro8KDqvZWL4XNldPE
l9tDxQfgAVse8M2VO6kYw7HhFF+EV3q/+zXKtd5UMt2KpTDsSxyNhRKDGyJQi1m4FvtEQfsvvlZj
ymWNhCTqdYghu9fRG7rK2FFtmiq4Iw3UPTubzRQdqteMbcG1wYjY2gthB8Jc5bDYLsSxzIMwNz4d
9Lizt5Uww0e7btw8Jee1Zwrq6QEqqhrovdU0b+uAfswK/KR2z3nneT6wpNYAJ9QV69EUDgsTAQST
xsWww4s09xONT5GO1IrZ5Slfke24ceO0zZKtgWmbJJSBZZr5BMJnsTkz1c9qOSf0PdMMSaUpcLMw
I7Eec8el3qJJ4IOoqYaOvxzd1SwWvOysh5uz8MDeC6cNqSq3TVP3lK1bmv9zwjVlLTUy9E1IX/D2
rZlDW1PfFmI5vGiF0+jyuMNpJT5PB2BCUbSWS1BXV0h7QEIkYpz+N5pgUDjk9P4LRad728yX4JPq
NwGTQQ0pjXNWdghxUFHhxcbmPMGm+9m+m/2HL9XrD0VbJD1/b/wZAZ8YYOzBYca+TcjJ5fY1EVsN
Qm+X4OfJsCqyS74G4qLjzPAHN61zMcxuj6i49bkBTftSrrhyR54hWPYnKm7H4GjVAPXTi10exvGJ
DzMyMLQv+WR0EjaFxVZUbt2kUHk61LMxsGHqBJ9TJW5X5IKOsHTeF13PwzJ+c14BnLWjQ7osMGPV
8lTKVTyZmyOrDnfpw8DmANJNphlCfvERcunQLN+Cso1uaRhFYyDhr9Sgg6KiGupvSqGJJ9Tg6NkH
eQJfU50Kl2/c7cid4i0aqhHPySsvsFvwyhQullTkIybdpvdBRXHhNWisexf+KCOfSH+HHuMi2LAl
3JVDNDDVsuqkGJiapQgWRBF+E38hU/zF8jPtp5CAMVy5gY4Gw5LrO4vKka9VqZahK/CrKVkSU5M+
xDor9SxF4StBSDXkkUI3UD/ATMUrhC/dFslHjET/OJFgGEfMizt5ZufFfpUaqWWCoBrsr9vxnZ5k
DVJTpBi9OYXBbkJA6ndlhHKfBM5bQVzTsmytQcTT4ivKPn71yJ7LP5QVzHSec1Vue3HEPB7F9rke
3DZS3Ladg9ZLQg8D1gyWRNcBVWmgseIKIvA7XcHD5hjlpQW0dUoOBRtFogdYm1iqtD406giTkla9
gExZ46AeYkiBrFl8hGAweo0ola2viD4X6nYU+JRcRObehU2ITav2PaXH4ElevxnEmhdhIbB+hzUO
CHFQQdkFJ2rVm7cDWWO7BjyQYT0j5dlmTX1Ecqufs4Heie4t4luq0RFFh7b+/ewsGACgGJG3Yk9W
+4c7vLHEi3iqvbY4BIpj+ZFcjIFUh20lyOky8c7cAmfWT1dtOm1EH9CfQkghzGx7yA3nVhOPAjpM
Srd5y1mRjVGGyKHZyTLsV5I9kjwi98pR5LF/NEdIfCtp3veHQdYEhtY5p8ws7Z3+R0xYk/imdSXE
uuiDkiCAWQ9uUtT1YVWnIxwQhKxuS/X01aI0dEA6VOeIknjXZHPSNudEmSCJ2em4lU7zkozsRxQ6
msikP5c4DUYFoXPSUyfYMlMnJEzmm9XvIc43vQof5Kw98Nnc+2dJfqomK+JqftN58HImncljP/Ke
r8U/70EmAklITp2f9lbCNabh49Eq3OJ6IsYtaXKoan32Abg2e5AvLYtKDzNJ7r0u7smrLXist3z5
3f4UKbnPgbnplGCTC6adObHhS7Hmq60urVXMeUN+t4+xBuNWfwenIrW+9qMyYdwuWO1sCtHiOLSk
Dt3jtZenUaEgaD7RKczeChEVofXeffaHO8imXS1Z7OdCJLqKTIZXDkkvPOkX0znlskgsPb1ekKxn
1FXss+gPqjNXS0vnbWolDPnms02f87NZHr1mZ/v1LU3sVIbNBfqAXg7KrZ0wUX+cGxpQyxzVuXDA
2WhIkyCaT2cf+9VJHhWPZ0gwSeqfZCsp3aYCIdWMtukfVh5fys8Dtcl/Pf2kwnMBfQdzCiVs01th
UwzUsus6AtJr4xfq83al+sov0pNDg71hArkuaAfIoTeCycKTnHcymegqtHtOIgDfuUBYlDjkt+d2
oWe4QUfNClmawsQjeYPaxDL8qTxraCJPYxtvOk+Jy+OxNGu4QO6b3lm5zajUEBN0Y2j6fb5cKgIi
3zjZNXgiRakYcb4INOhyfJd24QjkE4XkdVRgkrVf7EvRFdLUj2/RDC7T3uKPTEXaWrZXkkO9pDtk
uppFOO6mEg8yYX7YY1mEm8SNnLrmonrmxTtqnjtajaVqH635J6nKTgpUZUlUEYc5xpGja3guDlDB
fC5ISfo+JlgeNIyZM+S4v8znI5KH0h71esMrBQC8x15X1x8Ng6tTiB8bYMk+najKuLG8tzTb0MoP
Nbb9VzPEYp2oGDgJeMsT57W2tfA0q+EcBzFSJl9Vb6RbRdGe802/sY4jnNiYRmjjVgDBYSU3+4x1
7Pjviji/VPy5aBBwQYoNAq+1gw52qw1O+tpl34p36xZIFum5/ydVmvUBO8BBaHjBuyRJOA9WWeqo
7xnn7S0SlvYMU6j8O6DaN3fiIr6+Pchu0UR4+VCvuRQ6/00kt/qbJb/atbzTqXmwenuHbAMisT8D
eRE73+f6G1dI7GhnTq5TuiDr6yBZUVuoxdxdB2DkqWw31tjUpjD5/pkgqzOLK8lguz1BMuIHX9xg
8/sNiBO6ADiQ4tUgrhwi6COPmI42WCEO5vp809O4tBiwvzHQrbLmx7bXhJl9ZKFV3sz8xwKKy+He
9Md76WsrtmniKcENZKBREYzn/vl6O/soAnVo0uSWw04aH057aHvsuum0ZUA6JGYej1lWu03vuHOR
kK9XPpkPx03y1EzkMFKUj2S2je+uEBKIcssFu1LFqMWBcEshnOUT4gJYn0Twa+aP19FOacyyA8Sv
KF8Sz9U3D5F3sGyrs7EXA1c9VhTw50ke96A/2z92Sf2t97TnNUFY7kSW5F2J38bwI/8DmnBZ4Imq
ndT0SF13wwxMsh1XOHjP/Fig7I5aK6OHCVoUgV69XnRSbiu5JFXG+awwglm7L27eKtgb4C+2d09r
5T17q+mSrwEuekOhJAYLxCKVTGQ41V6xr0v1+GbGwBOPyXkGo7CzFg7X0YgWDn6U9sHAqmLydCDq
CeJqsiT2HGA9s8PBYzMAm3FQ4k+Ucur0bWBdGORQ76nd+YDMjM85yR2iP72PjkpJ9TAsQfVwZzF/
LKLXPUnBeGAzB7ObwSEJTudnaOcEFo7Y01MF9sKcjvKcKU4mwaZa2MD0QgJWE04YzlswTQWPDR/I
PdXZqISUcBkitp6RoHu8XpK4cBVjsCAnCY54P07sGc5tCc8k3U5tLrZORBfgc0YX5ObKB4lYS8uY
Q6b5B2seYGaGBohnKjxEBOd3dHxdVKIotBUK/MZAo3AxY/aDKpo1mcO8M5eM/vWdiZQmQd3ooMsA
xRyvQHgaH+NkgHplnQKQATvPXNz+SoD+kbEnfS+rKXBpV677q+WNdee7nZa4YBwC1brEZnYbVcj7
2oeQQXonYD5AiU3wNcmtHz+sjNPpnQCoDTjQMESlfsvJ9MukgNZZ3fz7jDEksOcFnYVzaDzCCYbg
hXeiUUMy7wStCnAlYttF1cKdOkPShY2XY4jLb7CIk6Nvpc/VtkZj27PAcarXjDmsbz9cqevcO1zu
1Pvej1Jj0Y4cCPnRDjTrytnLEev9DmzJfo1VhIz6NYa+n/CAgcZ061xeZOh9lHUQ9Lh/6mfwVigI
A7H8Vm7maPec1xo+I5EwF+sanm9opgSO2cNB70qxpedHFzIPLr8R97SYT5rZt10UpHtQGtTqht7p
hhf+lmYYxbJN7CXIl1l2YbsBzqjjtiHs6cB1uoYT9m34dRREOqdEcwRYxJ4DWerAUeZETySbt6SM
W8ZFfQztG4ikJE7ZndVmPVJb+BYdycFAmxWXFNJkqr26J9Dw+fXs6A0m4oTDpw5JiN306gO2OOgk
rFlArsIpSm1pVVxAfXlXcdKRkEHJcoMBRcT44Xakwg2wyILCyoDw2zN56ScVADXW7joHTmDM+Whi
laMR1aeB7ouQrb7Ipzihkv7o+AEE+nWqUxJMswTR8m8+g1ZMekLr+W3IXkIBqCzZX+L71edDK30L
C2Fs1ncquiocLzZmdVRfhsRZlJYBekOJlWYYFykyE5GBfsCHh91WaixeMLQGUckgZaIYvYogcF+c
amNKY4ZzMxqELCFTsR89nsXE1Xj4bq5d2EqeJOvP0njA1iU8IowEb/pcm3+ek+zOdd1ceDbqciSr
c04UICZsOQTtocXfiHdGqtgfrzv+kZ8k35bAFwiU5BFS1rP9oIiU7q4o8DxSnlC1C8jky8MFZsLa
17vQy6/1tgz8VONw5k/mxVcTJU3ZJRtZ+YJ2H6WKNUDyyURx0lJRABiP8IqDCZVZlDj7il8rZ3BV
YFoUZdncxaCKB/QLPY6C5fSwCqSGxZDYTxYaYrmj14xzCmu7bo8puKmw1S+Vw8e6qQaFeEBrTvOg
Oxcup5aUHC6k1kEBIvoizRMuQkbG2W91xTqPOeAVTc7Ggnhn9Z5k2h3RTcYJVGmE9r7uxMrPh3Uw
CkYVSnYDJIqnMxOt+Ncz5UF4eH20tLoDAlk4OZX426tAO61aiYPnVOpK7fsIDWnvK3mOi2m0QMVA
Y/mjM42RIihWX70VEWFcPOLNm3fZ0gLZFh/m/FrcCWxuMWaGcVslCFKwltR7NdMKMXs3jTItYs4b
fCDILt4HNmIU3odwDrUg1OgkMhCecqi7KieSC4hUrrVLNlO7wTw0ItBOEcpWQ1EspM6B+fhB3NmS
9hZ3EBUHJF2BpNHxeye6PQ7oyqa+/YlYH7PLagMXvlezh4D0/C2TkaupgTowoCVjC9SCKfgtuTYq
L6vQXIQp27F4kUIU76tg67AdEOpdjE7WfGSBf3TapoSxTNu1flkx2x/2/6tYMGey/1OgaZuogvEr
aWJLYsdT0D2eB0GvOXECoffO9CMYiYhMjOQhZLYrvOELv7Vsgqy5n5e8EX1o/YSFYvHAOwfcsAOx
z2btiBim5lehIdkldWyH9cFdHyf0/RGVALXNSCfWEP6TId+ZCas8ZLdiCvxv5jNL46h39TFOR+5m
k+Pq3Dw/G+pSQxsG7Z9mb0ZcR0qqpjOTuNtCVbzO0emro9fP2MhijptzcnKpE5TqHX4sHBH5sMmC
NQRVxUcQgxHRwuA04xvb0nJ05iVmM+W5NuDRI3mhghmnQW17nbuKwSqwQA1tGGyT3yFvHsAlmhss
gQOZ3BRYFUERDWVeL5e8n1Xv2u3u+38+gjb4IEj8Jn0Ja0cJ7wda7cf+5EFzULw6fh40r4F9etzd
X3mfwubTJ9hS7hkjjxBYyiJn3vrP7UwZu9/swT/6KpBzSswNNFyglF5PsOsua6Zgb1+7tSSyvN0v
9IcjYjwxU64ggavGF2lmGdHEGk+iYuPXIlrnmUy6EycMoQkOvlinRvyCGRWCVPmapXoCA3gXrj1t
t3u5H6HcvPYqin5xUS9xRLZ8hLPny/yZ+4sMnvK2GzO1L1kJlBAEfVtV8QDYf+EaYWZ4p3Zcl3UF
aPDbLU2MRUitcarMtEkpmCKXhZ9jxxujiqUncCtrT81pqCXxPwbFYm9/Q+OEOVBhm9MHCwSOYw28
OqWC6KtcnB0U9Bt+YiLKxwQKO8sG23wNQU4l5EyhUGDvq3DAZV2qT0BUzlod7j+usOwFFM6Ym3ot
yIpIpDEfn8yp/NooiTEGt7Pzd8EakIgXXGB6QsI8qO6cEogv/okIToTk+R9j24pRh+KJWs3RrltB
pTb5j1CicCPeCmeVsnuqLAE46376xIuk32RhjRKkZi2Su2vSrvO+5Ht14Ba+l2rTwtzWiSEkCOzU
Kso4Py1I8fRHNpEuu+iY6ArczMS3TYSVMzoOJHHlrZA4UbZXii4mbrudoVeZZOKguMaVwtQpRirB
pgddvmlS4wGMtHriPqUp0mh6vXtuiijjBe8roLBFmh2McZBPuoz8FO/om0UDAVtVkoJm8fBlGilj
/X4RAoI0hIfTKr3jBlazrUs7h/I4RxTe8+qxSkigwbGH9ujLQsBnSbbNaUFIuT01sY96NDhh1hyk
GnLhiEE6MDr9sa6T73Hd9cY15wWyWEYwveLnR7f0y2c54q89YDRH9sNPQCA9gWyNPDImLJRVwgSX
oKZQljO5tdM1Wkku46BI8qt6Cpq3nWVqkF+YxDjDK1rRKfn2ALs4IC/3o7pcuDwsVgzdgDlvhoFW
XMP3J6lg5fn4CR2F3/uXTQIPC7EzSiEdTwIzakppR00vGhJmMskBy2OMRWsLN3K1b50cQyYMUu33
BSYSRiVfdLHft4Yivd+2Md9I+viwjw7ZSR7sSBFTtDGRHS+XsO7bAwxcStWr+8Ozmt6uqqnMC8G7
X0wk/UP1CE5Hjkby+iKLlWvvI5WUkmwuR7SbZkf/IUp2sKm+T0OKpy19TVvNR7nbZxryv2DLP9Tl
ByqtLp8Yn2jl5+xFFtOCF/ybXJ0DiofMp7YYyLEuakj9Ir0Svwf+Se4UM8sGD8eEU8QxJeCDZAa0
6hB7IYpliVI/Z4dS47XyAuVeIyxhINMH8s8J2ytyPVH46KbElWG32dAlSa5sVo3yiuPiOXmhex0O
lXq0SC/9sJNJZge9ahG6KXKMjV096BW4MFvwDreFY2JNO0GXaIBaqBvtEPtrCrI6/7QEViD76IEY
cA5snbjPaAoPDY1tC+ehC2p1E1YvURWGfHjIxX7DxzoIe9hMLgbzv0R9qhB55LrOX/Co3XZlG5jO
yalXyORzEZqpuYRv9/epVqUXd1hTC/MF7BZOZLNQBxtgQ7B1UWt5BZTONQDWY+I1NTj7P6+kKacp
3p6a0CRD1zDfRTNV4gOvxx3GbTlZrFPoubkGcOCJzjzLbVdqBL+euysikPXtTSiqcAOdU7xUj07D
Q68nVUcMMHeKQlOIZgt64qyk3Lj/9oW+9Lv7gqVMmLKtQA5lQIYlYBqOxiGVtP9h7IIFwrA3X5S1
TZhoUbSX0Z1siascL3w9LdH1vBMQBH0RU7+sQH9yAgRcMBSYahEY0w2siteI+FCMwZJsYtvs0Y1y
icv3MF1AxQaXXMtdaWZrk+36QzntkDXecdkDlz5ywNeFBnFCMmZjkosrrUhBWqDES0BQ4d61ferO
7t4z3Brax5RIFJZATMIySmOjdsShvALnNgyWu/W7N92awkq/SCPFaIN4jRPpsgalbjrMXVmF/IOQ
J3bmEhb82QHYrHcSY0ruvebQgSHTr13XL4anzUrAoKBlVcb7+xNOArHzsYWkhpfDSbmrpeDpcUkL
gqQLGN2x7YBLgm4HD+bvDQVoZYkHcRDEytU7DCw5d23sgcWZnGd+cQXpOC0ZugJKVQqq1jjAZYAS
ES9xrfPX+UgVnTmvkgp1tCbdnwUMzTOTvC2zczyJh3b9HYbIy/qxEnEdw8/qQUSZMOXdR+h3To1V
GI8VkrWHza8GW/MKaEbTXaBxwi0s861ZhdV1urQq6GAwUz+0euxheQ/vDFpiRi8gnjq5NTHERb4t
meO9sD0pO53UhMqOfjMoh4TDIcp7rFSPq0v8TtW4nd6g++RcMnYzxcvakS7lsL3PsM+mnuCD3X13
7mcg/Lk2u/LWyqdDcnNbHebZOdKc9ak5SF/P+ipEEDRaBjZ7DILo5tXLIBPJbeWhHWuxyJv7KaKV
z7nqOKytRiEQUFJ26IWnm8cBa+9adf3l7kHDCEttzA9QOw7IdD2Rux6JmGnyHwxn9uqH3CoJStBO
HxIN5LyucNy3IgHEn9h9Alx329a62E0YqztaXIY3Ep70PGuW0BY7MsDtCF5ql7/j3OH47VA5363j
8lLYzwnIkOOmpb34K0A9Z+JnUgaW2vPJjm5KNC5AlqUK0OyoCk13WLpqlYMk7sCL6UGo6xNeC/Zx
rZTgAvMyDTYhex0XDApdgX9hASr3+LMshmrOrAXuujj8gXFqYZmKe5agwfUAKLJtvolZNImTe/z0
aN8xy7AZsj7SQKD66RdDko1NmeGY8nyLdCIAaabNDz0PYJCU/tcUHNstf7Vh3qka092TskVJPfw9
hv/ROR62IXQzMFDp/x+QkK1vXiOfO8W3Z43UfcyA9VYrl7jzmOshn0RH3Pa80n7Y+KKp2vGGa1K8
AuX7kg2Ub9mLo7FGsVQbKkp8aonfKJjmJXmN1L5hP/n8E+9ItsupMpbAERpnGcmpBz019LzVuoQn
vLb6DLXUpIlJdPCKALCxb5fCdOdDxajqLN5YCUn2jyHC5BMNd3Qje5Z7sPj8kybmagx9Yfq++xqE
IeDRhqk8ydPyq1M4OE82SL38r+2BDRXP+FsUCVQ0pPp3UWgdEmOP8/S5Ci46ziBbMO+Hvs/L8aGS
7Pqj0toMDSSd1r2ydIH7IBsAFXgOmUVmmIQrFlcG4/WacbRUO+TqD2YC5yOeQoph73Kj36c0VZVY
GVf8AGYchN7K4sWagLYY4yzbfTuChGOqTXRET045YqTbJzWKT0H3HAlW/IpCxBO3RLZOfDt0Dx8a
PW3cKDMUG83A/wdXGvY53WN0JVqNK9H0VeXzHqUKNU0vkC1MeOF5YsCDZAjnCRf4S96g7ZiJiFbm
Qvjp+tXRXD/o2n/P6Gi/k0P1T9yTmNuiwU+alfH9ygilWxF1V+5CiZiIEY+gmBmWYpSxy3BX5NvM
wW37+LbzvP065em8vkmYu2pv7RD75LIrswD9kXkBVtstsi1tZLAMqt6TRJrgxh5ICBMrzbdI4xf9
bPBtT+BkdzdLmkNRHi8yP1VRHCNHAXoLrT6/+8ItCGDZoRg42PeXVEoguHWqmn/Kts0Ke7UOLjhq
7UWIQoT6ouo2sltMWFpHQFLD46msXKgd1jYVpn5PK4/pWuASQn6vxiFJuH7yuECmWkOQ14eCypYb
70Sam/GsW9bzvBNgXMtUxFz/FJh0ZSNdnR87gFX+51ZDMxZy6B+EGCjYjineRyuYHZgWCq5MuLIa
9D9CmWVkABz+Oy1K60yMubh/P2cYY2U2anGRibcLM+3mV2vcxuhOYlkEVNheTOgIfqBCmKC8vbca
uFsH/RcfuGT4J0yepHHnU3EXHnRMCS13eyet9sL0fdOmZpqeJ/31YCgZLXOoivnq6AsbtZGMBDrz
mm3b4yZIuBaZLph9vzsj38svqclFmBlYI1BGpHyqd8kWad0OwNAdosS4Da/pHgJdRmzKCOGdoQ2y
ykboAMVeViB5t+Xhh2EyhmEGeolaTmkGh6TSPdk80RsqW/MI9GdMHszKzdUxg8s2aqskRwox+o7d
jBpfP2cU6SiaO4Z3BlkhL8S3hFsjfgzcj2zIgd+CxcJhzAo6PBVmz6Ord6LVEvxZ6NsxHP7wZFGx
sLe7sxU+/u6WsdxiLHX9aJ4VySCEn4ia5Nwh5Mz7xNFZ+XoZMDIB31SyWUohULCP9zKOfFGGPJc6
7Gj090LnxxWb71YaO8mIvGHcowsaya38ogrUIGQKvJNrIXqmg0cm73bVKQDtQ+pB5LBTajUEoHmu
rpi2+N1gjFud4gNUfAUMLlNfHIFPFFl0amUDPFQ9KqtHt5wAb/FuW5xvlEDuTN+nYGUlDL5aCNC/
Oc4Q95Bz/XDRZ2uIu8HV45dF1WfatONp/vR0i+SQlzaxc+WnbCcYEO4vYehAyrL+IHJMdeECqIit
m68tVeo6toJ6l7aga3l39o1ANZHLfLHxQE+JN1+uAH9yCkfTAEEi7ngiArqBW7TsWuccUq5V81hv
yK8ujSagj02NhI3UdWs7VE13bHIxQeG3AcXVyQBYkEYUB7tKgpuqeCmM1j+xARp9QIjwwfr9dXqC
wdMJ+mEb6Z5Qzzh36Cfmy+JNahpy4Xo4bu7ZTY6Sp7FzSNdmZGMT69F7OkApCW13IdRU6qWvtN31
kgzQOdcf0LEYo7jRC7YSiDB5Fp6PEk4swxToE7/XeGeqQLplrEvF8K0Xuhb0yqmRAbNBj3tQf2AP
hBgMQZa26G+G+FvP3rRbJg+TVvgAI+6SwZaIXVFFJoJVk40k/Yr8egUfAAK1H4rVA0x6ln1+Omwm
m2Et7YEW1ecLWgJ/bucQMQFcleaehgItddl67ZVx03Av1uvZetQTRoBLdX+tpwJQC6xQCPqCTHlk
Iu9UXuLtC/J8omeswZR7tVk0a3cw7Bma8apkxZkYFYUtqZNGl7cqPMVRcsssOJ1RkFcLt8vEqJxf
zvLfDV3eibJwHc/ipL4iiqmToXTy/Sdqi/eHKFPOrlEduk/3kQ8vcJYp0PI2SDpXXek7rATdtqAA
e6KWZuuxoVGh9vW/2596rqh5qFDHdZXvD3JSq93fBiCqNPgQRlq+PWeQx3KCfS6bLrlKC1KgJkGJ
/fjkPLhTHVfQp7bblubk7fQICC1FyN5M/NP4G+BvqkEfIATxEBhUVUbakwMVNTN0ANYCUtvKwNO5
Ugk+QsB0Efei7pWdLEnHOEcPl1x54Ko8ZfgaUW3Lmob38wPVV0ngGZaA+aiCRctx1VMPrz6OufuO
GwSoRyXSZtS2t+VDy0uc8v0uSmIIKXQbCPo6vHOCApfdibnoZdsJvSju+W44aR6NtJp8veAgl7i6
O+3Kzs8OfCUce9vEQ4Vgi23oH3eg0bJ+3T8RK6t0qhm0vEPMEb2C17FSazo7kz4EW0QEykN1Sk+V
O5fBgICkfteHvvPaJ1fuINaJvQBPPk9bLMQG+z3dFjvxTHwI7lCvA3//4sZLIOd9+28H1hkobbq/
IAQ7Hw12GHTGXaw0vU48tVYtWPl85/ecOuEF6iWXDd4ucHr6/7ALppjkotTn4ZVXCBt+xrlx8Fdt
Hp7j1ro3BBToed+3+ny0XM5bKVVqFuPv8RyMFwMHYKIlcdyborLONs0OTx5/y5Qjw2FgwdI/TXcK
6cyEPglJgEtMq2C4LCrd9QYXN2Jd3RipP2D775rVWCLn6miwT67/wlmn04uZpDzhgV2a7zUqVrIH
h/PWIu17oGJWmjl+BtZujF3mAFeeTLttpQzXqi37SKzB5gfdwsI8CHGiaR5mMb1795BIUJ6tAIZl
blpCWZE9rNkFnoi1rvdTM2TldrYAv3MGVFmgVI6JFU1rVSi2j1ZQ0cgOfMw2H+jeVbGhmBpoSXN3
9jrEX0pIUVHyV3YMmicb4/J2DlJ2YVx07c1QI/8dCyvKXD5RjDSFaKZNWG0h7kxFTL8aXm8/8H2T
RZFzu1ThiczRmKXcw3Cyrs9EkciNxq07ddmrPcFm9y+WZz6QixQnqdBDoETr72Jgj1V+7jB38m4V
ENyAfz+//USAk97EKEdDS+A9YEUJMxBAK8i5382Mz59Oy9yVwBqOx385bGl7mMyfHk1JlDrLwtZP
Q1X4P0b81dPbWgffvjka+Qa4xPR6/UZvU52wNVT8F5ISBIPsgLnwwgZWVp7Ad0udSnYGOGVrT72p
OnyUtBypyu0QRcgVtFjEIy8JQWcP4R0YWMT/CAK7YuGvV1PLPAQ/j78RIPFM1oIYVHn+U2IUWsxU
4xuI5oaDI+JtQTnEwMg6SJQBmoDjgKZiL2XegRtc2GYNjqLxGAhsSq5sPjeyXg8X+JHG8xcitiG5
Zx83ai6csLyssZMbYF6GCDqQ2vmvww314UP2UejeztNFJ+2fANDylWAA9UZOwJ+QnR+1QwtqwnSR
DcFTPdbdyRv8ReLxosR0X3tpTGFtBJNzl1MEFnhcGm6WuDtnDjC0TdJJ5n+nL5oMKJQvj+izRmbI
a3YxVsAj9l1cMCa6iAzm6zP8KUiFOikjysLPH/TYtXMZXNHRikBw298q/BJyVXlueY+gBsffAdS5
N87nq6OhOBpIc0nFO84yWPkW5EzCTY9l6Xq1QWKtExtfuXyoTP4+cQ19t/1C4tny5txsGLV4CGz1
RwL3DJIUDExbgmf+ZGU7X1ED9kAV6c3+eW8Y1ZpcAwjMM1e2GDz95XyGglYm9Tw2s3ggrAmqaq3J
2CUbvqSuMK07eN66dMRDn3t/0evuEizdMPhWao/Am7E/UCsBZxAGzof73tohXYXHCYiKPoSJGFlO
CbDash2aXSmG+gdnUkUDJzMSEdkngGZF0Yku1PL6cR5Bn0etIQRA14ZnnoCo60jc4m/Lb/ADYimQ
rDzPnGMu0vnHULHuAsFqneAHTw89Mqec3gnI23SgvmZSqu5BbKPK0l2npl3EWS7u1SK8Vp2cUW3e
+YK0/EaFNTn74ZeUQHUtWGP2KqnRz1djKpDQTrldRQdHBKRQMpFf6ekbKJCyN6zk5+HueVHWki7O
mmouqRxbzyCbuFqRU3Cp+PGbcJ2HjUbK/sz7mDSAMFYGupSdxJD20p/RAjUox4W2Fj2Ga1PXZKjC
Ftwfs8adplXFsAPjObheZr9ccNcUKrTUqXx29tcE27b16HPptxupqFIAO5DBmhgrr9JOWkdhrtzG
/D6XCz6RCx0Gc4Rmhn/1lF4dtWkORxRfQUxj3wblWeIDZ6f/cR/5rGiiwgR6WY+7IGaCwM74yP/U
3EIwTl/95WShwuSsC9tnsc4Xyin52igLQ5UoXjHPZssq+yyqLXKFLZP76E0WdDC+XUXaWkYCESfr
wAoEowUDUGNE+YuEqN4JILdwUQJALwPkPGawx6s0x7Q0MoB3MRYLsD+gOpEs4CjDtLrpNKUKaGqp
WG1TdHLoszwkfTIUSqCT8IQA4N6dMIKwaLWHfoDpwqxDA7/5cf8exs6vqT6eX+WdcGXmZqbuZ0kv
EroXyFFQ40JqE+Dn7mchYRysN19XRHgXXmnVxvLRXdZwiEoiJYyekGRJHlbItH5kS3Ps7qP5MEL8
cwtrxbWCWHD5r2FNjDR6Jla8f3lu1Rlq46jTTEyneSwXqhUPmuEjZRpIHmJnFi8k1DE864tWcuFb
Y5oVY2gwxQM7nKTy0LrCk2TA26Momn2/Nga/D14T3ojsiiivZVRGgHR7kMYK/f/zVj3R9VZBT0Am
POVEumw5OFDA/j1feacGqHkM8JwOhEUooGx9UPKiK/xR7BC0L5ty7ZjxBxZvReMBT5kkynGqd/mY
8Tk7XXm6PlQxYDS1xHaKPfG/tA/PwI3ViMveIDeCkHVVq1dY0vzsd0hgWfurn+yDaNzgM9g/E+0f
5Iev03qB3UCnMxWSJkPBUHv1YB4PJnBDBwu4p1aXKnl3EAMtj+xyySnmKkwzZ0SgNuUTQvak4gHm
Bf4D+oslc5aJuLe+7dRS9mWgzW9wHQzzsz0fji8t+J3vfunRxe04qJDlh3U/MRsg+NrznVxYp2t7
SDpfUKb9WNzaeUeyFVSBDcCHaPgHH7pHhdpqTZDk7u1NGYUru23eoKP6N9pwBOImtBHkbc5rEl25
8GsvyM0/CbRAJ/BaFStKqhI1XNIex30C7Qxazl3Um5A1gW7Jbz6C7RMqwGlUyIaXLLWDOHuqEpT2
Zb5SKau3w5fXZLUCCQak+N8iIt2/8ksjb8xDDXDEr/EsDEPWZSCfxBIo0M8IGgxQrvIzWlM5lbB9
KSLgwLyKaPven0kY5nZvGn7NDS+0TUiAEqTHLmbyNQV8OXloGKpzP+qqkiCx/Dyqe5Pim02UrE5x
4BD5tv+cqijQthAE9lnS7PhRDluFtf9kPqOVxIvHAlBL28XG7bmeiF3jRapzBtQLnUMAiWlFa7KV
MnvsruuxvOil1f/2A9KFNAsn3HIXhvKOOXS30OnvsH3pis8z9Qq2oL2o8xxUUytMo3IzDNGD6Ygg
F6llGgMuaP0JcaKFOQq5YKitNDQPk85sy3OdMU22MheXIszm/zh+WtgjasEcbnbJn/YRu8UyPumE
X7/BNWkDaNEsr0EkwSA9Vd3/G69ObFEWawMEaSgyDhdCOCilXqWmtiu7pvSqFUzT19FPyXAXCgGw
nMJtn1JbRMSsd4ZSOtn8APFGXMpWenxYm0opT+f6hKCZ2X0BURiZ3Ijwjz3iDv6fZ/Evq65um0Q1
GjzJP0E7Wm46U3cy7FUFWDU9SIyTqxtbSfZtsgUjCyzJ5q9nY1A0dDcA+2z7dwz3ybmcWqzGJZbI
HeYJQcVQqahIHFgzdVGPwDSWEMMVCFG/JpzIisexbOYeUAcuQGl8wiHP2xQoTUIgHxLd7tQeCdkq
Pb8j5vFNi8Q+n1EQwHiUPayEkXvs80jNhhYkfUkx/mgDy0pese2ufMOr2WblFcnuBcBy5FEoE4g+
kQhrTsry2Hb8mC6wLk+bXba957Rmpaf7TI/2zad/0uH7A1qYyyPW9RKb5bOK8Vy/sYxCUnLhUcpC
I4hMmu6h36AvIeUgAcJbbaofbKbj8GrJUQgh2DRNTQDy7tDvM8qB1ENIUVZhh8SywKIsmvejfO1A
Kd3glh0/Pmby/mG2Z+5f3bfJeR6RLqpD+nu/zUXeOpg7d3kdWe2IRWI5/uhHxLLig3P3JLkEwJBU
WgykjEDS2lajNhJDfgQ9TIT/psguWrAEFkBf0BGB1QbMbH7+r83K993gMgAsKBwdBI3wIJT2pHHC
LNbqkmXRPdAl3cnsAZKs3/dTUch07a3zbR2WX7jqypk5GDp8vjd8Fj5rwWaMzCXQJs+2n+gGDBhd
6U8ToQXE3pMD/RBk0yMHlQEB/FZ5IqmlRlBl9nBHZfpr9903YbSYy5dgaKn/0RDUEZ7mjF5Cziqc
02JRvX6a3r01WosrR67aI676TitayVes7Wg4GIjm62bsh9O5G/PEcAGcFRiFiH5ecCnvQ2vF5Yhh
GIdTfXZKkrvabHJ3G8QgXFXfxB5GwN5pfyZ2Rb1jfNALiQsKN5O7l3QAUa6KiZO3QO4VUowj/w+y
TMlh1j1ZfwGjYr79kRCyykaBARmuTzDULmQ8rpEsf35S731S9Kt3E2nsvBuMAVL2Vk8oGsKD0Jfd
belONVgGKaT8tUzth2TVT1ojvnL7RD2igRXWKH/jNHvJV6zL7r+bKSJRm6dz0yPvzqWHb+NLv/ut
He9F/WlelLGldaegdkrSC07EP+XfMzeMGcDYZr2URfBqqjWzSbDqG/GLNMF0nwie5EBBV0AsekLY
UIxF7lDhzoMQu8v/kWWwLgF722Exca9DNbzyU/MgaZ2clXsIAof7muN0iUS/Z857uwj9YoiKtrz8
Y7YblClcsKtb/Yh5uFuveWMgEgbN0iXftcffqFPJQXuNJ+AlcLVyRTuX8FuThZNQUFI5rippIukc
mwYQBR4Ko2CCxQTNZy5g/h85tpRVLYAWY8TTkkI1kRyOcdMYUDsTFVXwpJ1y3CJHdkPkUlTj8tb6
G70m9RXnsHpMCwltDpyITd1wqTiYAT9LtnPD1pGXq66SAxzCHIKwPgjRxqH3XeoPScd4u/pyMA6c
/Z5pOsSezOT7keeTVJ5BsJFHSnDrEXn49rayeWQvaQjsz9SMuU5ZpyUA5QVFnlwqhYiyhN5L64vy
liVmBUp6ldXKFxYEG/Id0RA7grxQd28+h7pcN/aVHw2VahvD6CGHSUbw3NGN2Yfi0E6yVqWi/Xb6
YXZrcZlBNRfvhk/IsXkN5YogcElVB/w1hhqmOKKoCR4s3msrX++3mMQKVkTtAk8n5TDNbEp4/hAp
psrwO+c4FS9G4b7JiBUuM6gMr2aKNgbyt8Vt80iBIm3gu8rLr1GuBXIweTfq5Zo88vIfI46tWVBC
y5AI0o011gMcTWtN2WRp2KU7QourXKBBZtAgEWy79KsFemd5/quFs+d+4O/jsRrBQlyOeaaiED1G
JlXjRS8f5lqak2d715wzModD7n57gQ2j5vzCKBpZmynkPg5Ksa0/3VovH0nNAcfav/CZZcx0sllL
h8xeCNipBHBjAXRgXevGXVilF3JveWhsmvSXbKkkA6a64IDJVb3BhrDe53eS1Sb/wRMoo96Z1cHF
OzFQNzOz0muMhxcAXh859fUnQ8StRG+p31a+k4PQEOoPAKdMmUqEQ3+/O16iHfa9o30McY7GAtsu
wMsUvW7AjPW0BNTVMR6JyPMpVLKoK1kZVluzsf71s6xyGUEqIuEULChczS5OLAZMVXYoFiP5ooS8
KEyj017Q1M2uhzCWqN3b0DMAGBG37xiiXnsSe3aXJYYVAgT+DwO7TrN9ZtcbfuWiiKbI10c8ysoU
JQ2WLT337CZ7/qlZ6aFaK3IecXSbAs+2qsTpDceXXDeh8ALOp+0WtFRDaJBUDT/3M0/+8M14ZYWK
iu9iBxCSMn30LAI4yA6ZwpHKWQDsZp3KiO//Fsq67ar75OJcMXXDqQcBSF37Lbsud/703Fs/0apo
Qo9eOzHNxtQcNVCNq2sDoZnFftLeYmUXTNdHs+utigadoHG7qBNxlNoTp6+BZRKHlrLv5BmujXWH
AEJHMv81LTCPAfe0cvScIPgn4U7pB7nHDmZJbHkYzPaLl1qqMDOS1FIie/FCHhJilIOxerUv052C
nKVLvjqBCnyxKWeZscrzHU1pYbcj48NWBEZuHrW82AfMNZXTUV+436ok4KqhAoknWkkkA5sOW1xT
BuJxAxqq2LdsMmO1egxXm5CyjNMb/w9rqD7bTkNpXFFRjG3LwrZKUmWIkDehFpJ3k2eaWfSfxrJD
qBojmDmCBLvahNBbGx3zbxi78v1g6NnUAcqUalnXjGukOj9Rr/cR+tnTBky/8o6kwPAG2ab68mV/
PB+AM9dAcqkgoRFNgECsIqCY4d289yBNTBrPeuqP/vagZD17uvPchyN1woYsiElMnBYPJSJ2c430
ZT8q8VA1Cm52LeRV5jnPbuAbFbyhloZfGQ+1+STYW7dPPO69OYeYaUp+zUbPpdhRf628dW66Infs
PbfTWA3jDPLc1jpO82uYEB4hjnQzc9xQ2mFVVNbTjG7Vn0FIvmLe6LTqdB+2SIwtVEjGMn4urGOF
LOi6ZQK10GM6o7lCa6hShbD6PvD4zysQVv9wnWx9z7zoGxxLb5ro1j1LZeO4LrdLbFYsa4WIai1e
w23GksrbYXzaJKebKli1kkJNrJq+N3pcDIlzEnvR/ytSR38z355sd5YYRssStnx/T+BXSgAEpQo3
t94TAJsGrqfGdj6fV15CRjxG7qtWbjRih2pYzjfC4AEriEFH9z5OOXXDXIUvHYauZ/IhHhP+E7OF
hFyg8Cl7QxHkd+X5BFOI56xCEo50g35j3h7a+hg6hq6xp628uOmQct/LPgT34QTdYubda62WPDwW
He5jHmwQlpjsMT3lv8t7GYC8QoBVUFz1xCb3oFsy85Zb5Rk7a8kysWxrIulHJkn6y0oAZg8c6zFU
b6op8nIGjjWZKBgW57D8mezqLafFxelwkJPcHcSDlxOoR1pvCBTEN8qepPPRFaEir8O6wZETq312
jto39Tz/fZIaK0aHA41vHZLlsBkoezg1x2afYy7hkzIrgFeSApWgFEQvqyav+qdIo00FfHq/+CmH
xaFH1bpe4SeX5PxPo7nwyfgRm5k1MyzmqdJJYaMdGeEwYLE7NGXfvSNhx9xf/kNby8kWwLT/RFRB
4URiaBeIYGDXLMruVVR8jzOIpdwqEyAIlGsf9nC6groB5hTEdMNKCuJ4pnmG3qiMEUSZI+RxvZbm
g0s4UY4is+ilZP7fpUvLxw5g0OIENH4Fv7jKU4LQ99zSdWuKZ8Bf2s0sWPO7A+0VDauYQiWB5SqX
t+Q9wJmta8FBiivSybbphApBNhH+z/PXF7DekuNzTG5lnGbtpVaOR+8FVOYUDkRmKWrRBWSWXS9i
K88psLs4qqWulDHRPIuIVN6NTW/LCpeIp6CWqAQwsPTP2RwCWg1sC/+yPuw1Ypzdy3RY7/HqfPHm
gzwr+jtOwHKVij9yKrN2NcEEyxAG5un75ic4+EjTZhSQgKDCH9lTUoPfmInUPyRu9DGyWVu7/Miz
rHgtQopZeh5Tt4AOxl+PHt+NuMzJO9dTuSMRvcPWapXfkbDyMBVz2erTwpu3pZsBdKB7MuKy9prp
JAqrGWbalFb7m1BmoGvj1jGwohbEPBFYXVAa7UFcmXgHDzagPZ3ZBpJP771VHWuNbv8iWgNOE0fE
0FCJgXqXPQTCL/Hwm7ZUnFBoZjifFlekCTPZVlzlgMK5zoN82rwcNEcy/jeZukw1HnhBjzpgeMhP
BzyikOpfNjb35/6Y8XSHznVP8d4j5Ki0x8+ym2qqhm6sDMBQeEteqOKyrC8onAI7d5Ij3eu9I7bK
XRfiqTyd+u6YtWLb8tpRDWezGUhgAYMPRsSbg2bfbkZNcRC0iNxxJuRCgt/1fuu7Vf8I3kc33Tze
47KCC9qp5Jz6i2ciTxsm4f8RWpVc2wMaGizElR6VcSSovdMdmsflFR633o2QzHRka46OZ/fVsnRu
1SbYcx2bxbFOPTERqUgzZlMOjsBm6ebhCc3/wVieknE3kj5sNYJWlMt0UNhzCHM18qvaKb8Rtolf
s+Z5hmtQ5z7Z5lmecWszdHySvomsdsE9kHQ2E6wcX8pnVXpDzgC4+FHagccQkx9T/55ycNQLMGR3
U98lgMupCbjWJUV8Vh1WOoVIcnIg/cRoO7O3U8QP3eqPqTTg4VC/e//H8PxYjY2j5rlI7Il3/itB
4Tp1LLuWM9l6ME4cyXOLwDUf/ur9JPlBqV3e4Cy1j2H63G6GhjJr+80ihgBW15p5mpJ4l1hg48Ka
euVl2YzN8fRS1TllA/mUuhlJp8NQM8xF4Fy+gqubvThPLu5gzYxXfrXtAB/OfZn/36GL+pbvj541
MqWdABhUS30oBcURg+FHyBTyxRsDR955BZ2vD4zCU+73NJXx3FXeiB/lCfDNa3XcW4jMq19TCWLD
f+SwsKi+bbkuMQOAIkxMfEDRJeLUOu4SPSuacMVWh6iDhyHzlD6HeaBwsg63+Jms4TJJY3WHviYa
+NQVInZR47iv6ASsUhz8pSh1E9a9uMg+ich4Re9i99A1w9HdRs49FMcIYV9L2oMQc5J8uDqRn/t2
1DrSp3RtFLbtDevMrts2tyBSg7sFwKs/YShYJ3wtLoehldr9FJX+gtznWx/pkPB/g6YRjw/mHlBt
0MBpNwrOl0GfPaCTJZfJU9e9tIl33b0VCuCaO3HWVE6c+vyn96QVsiLx4zTElrbZwb3bkYezHlou
FO8kGMEbOYVp+kbUsdt2oC/zLQvbSQ8nkWUePcMsVrGcnW3TzDbH7syNU76H0ZWgCVi0n7OeVDZl
upNhHW8GmpcbAE9f/Da0KJ3H5bSZFsak09XqzBvpwL3MtlxlWQZink9lGVaDza0sHr0wt5cLkUqi
9VuPJXg+N90OGW0SZjJeLAnvwlCl8wfVqsimV8EuHC32LosmGhcW3VKPWoh+gOvLju149e2Igh84
uBfnJN6g36ocwseE7uV+vzmq4LOIR5zRc0hYXrcc5+8aiEjLY/tbPyL6PCTMCwHcKG5Or69b3y/l
fPUB4THhWR1lC3IuO1Pp9B0HTP/JfGqnCYDuZfPz00ZTI4YGUd/0Y8E/XGkKB0EKQvsMrLZCzviN
jgwmFKHv7u6w1g7fP3el643XLnM/it2Emb/W0LB45AGsWiIm95OWNSWiVw4q5NWpLmdGkcNBToJa
9+yHcc75Y2H40B5pokDBzLHOJpbO/gAoWbqVd0IHY0ILjeGbTXjUMTA9aUOdqZTVA02FZs2srzM6
xvcES2SJjiz83f4k1DMpf65ogOT67eQ39clGAh8JglVUvXScj281stkp59FgVLK0vVjP7Lydj5XX
55KmgWqPFFqE7XaANaFWHA53poSrJqgWerYrHOK/8m3CTiS+SCV3ioUxU0bKmF89I87TQVVQtx9G
3mCHe00RZ+/9Rjl2kiQaYZe3AmytJKlf6PQTIf5yPyNCHw4L/6mei1M/soAwDXxsV/dvtltssZEs
i2nChdT5UjaOqdaGJLTGZq5hsganlQy1ummTqTnw5KsOUe0T6I8pNrdEpQbihg/sJ9aSbBNa4l1I
hmLuOBKB6e3Ki5Y4fTAhZ/prhUPRuXuc11xzBs2+5UhcRFyey9JuifGyhxsybCVXVMmp0YXll1XS
SUQeFcShacdbI1MINbPvHhPMcUvIw7gfGmhZVbjiyQ3nKfkrYXiPdVuWMLY5WtaswvoB20mVKikO
+/5EY16kw2Bpw9btpKmAkKDbT6+Q+zlhIKqHm1HIWXZBcDqiBQezY4g94JXqD5WMJ0j9a0mTLzau
lm0WZ2l6Z0I3gn8D5IyTwC8Ab53MRzdlQzDNsvaU/QaZhUseANma0jI6+flgXGRf/5gOsbZ9p0N+
gcKwLxoNP49qq9efxKife5Og6v9O8C6E1ea1P2CQyGoTY1mQW0ieozwPsCyL+pDC2WxwdtH93thP
C103hBaqvOLyXvSlGkGdVJZf2+4aengI7THyN9i7UnKQpWHZgi5CHnCDFMommeuT8NUIeGmgIYy6
9oqBLdOlwGI1tSMa3O/1lkqEqfK14Qen9eGX34W4lpdTyVn9TkfuZQJxuZTrcQDT9gldsTrf/pUO
haozOLH87UwN7Ahlo95wzx1LYiPFZcgl1cdkJpxqSujj+UZcvX6J/Gg2z97k6/CYr833BysMezgw
8iIoBfizxaph+L1J/JGgpaArfVrC0A6oeRUy9xLOEXa07e1jyEkrp84C2PIMU9UQDWa1sdzAy45U
B5EhptOJa9DWghrsGtHVmLAnadxNZlhSWoJB29zqcnu8enLwsCA2m9zuHwh1XAcGzY1rEUlMvyK7
C7D8p+CVIls1tNf4FYRj7vLmegeE7TWg3RhH0Vaj09NXs9aCN7UtXd1PL2FToZaZeB7F6UTTgEdC
PUzPwz0AiudtqRX0sxTNPUfj2BnBm9qnsLQ6sXm/398HqKe7deQ5vfvC5pPK7b8mCa2ytOPo9SNV
xdbsah1bBM98iqf9CbmTt/qTNglQLBlREEJej/tZ+MZbvVq8xDPxq/jf+4RRv8eufd4lfR4XbuWC
23M5Oaop+yGiLh6igBPJYzQNYjS8GJmw8jGhHn2GocuO6AhOAZHS7UauMr6i2jjACgmjPmlW4aNU
RrkqbaD0cv0082jTp0OcxVsQ4VSk2dURd8MsYpvZsUEsjLtj/MTzEqOmqPO6mxzMGcyA1ei7hO/n
veJOdTS8RuekCPEk2r3Avxgyau4gWJGeSkceXissC1QVCZPy06lulXm4SwN1lJ3gD+/lh+aQGP9K
grPY60IZF5XSW7AS54af9qMvEt18v4OMHvwa+G3SuLJ6mOjONFWafxSSkhxjLPoGWwOuUkomPWbC
HjkPumzsdEtzl7ifHhYz1+TBIxakaL398HlfL2bGKC1h62rm8O3mJDt5lAPTtldOMUu7l1iHm9VD
s5DCM9mPMDWiC0wSSSDHk6j848g05Q1zSSpgvgOjBC3WwVDmHot9yN3gGkqFk0L2gLPdJ8NwVix2
OBVwu98suCv+eVWgib0t3nA2t5h6tNNCpTrBwk/ffmx1Y1Fzk/g0C9ry12GRSWtO+nllKivVNYrf
OQTAuDOSBglPGVPFD7zzlzsTa50aKgpiwTOXryF1l1m18MZv3xxx/kssS9hLfMXoelJH4xyzbhCN
Xlb00gOme1ZekLpYj61uB+E4Klrg18LRNlMxpFAOao62NLfs2lkrjyrguzOqdQMKlmSEApg8CVeG
q8uXYG9YJwM71fnXCsrP5w5kWvgDcZTl/Pb+yznQrh4uNj4nYedd6Bc8M85vCXIJefMDWCzf4oYl
1w0MTok4wHZJ23v+JCsLz6xuqAWWDTgqXgm9QLUb8pLBY/XRJXMZ6W5DLLRdFeCfyrdi1OXZhthg
IGUTsg2rSGKE+BipmMGQKf54ffTLXGMbIQz/5DXb0c00fSFdEZaldvlycyzp4HxEb0C0R8hmGZE3
s5u2CaczoLSXT4kT+wlvZn/lBFt8LgvpkdUl/Hse3Ec/
`protect end_protected
