-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
amGz8Z7CvEw7kB8uXdtJNRb7wHIPfZxvpuNJRIfxRKJbu1e8CI9ryEqj+oNK+71qCrLeFFlPmGmB
ofyfp4dBiBMZZqB3smU5EZtdZ/gzPoXYAGm9t4OlMXoJSi5vXQtxLea03g0GVL2uicE/CVPCKKRf
ZLDftk3jZjheUDIgWmL46UTN1QmfuVZbVabMuD6EnSln6NwFVFmAADPhvVyTJb24XGUxNZIbdMik
CyFNkKVWKX1jhwo9aXuKiuf7miQD1OqTvTepL0ul7WIcWSy/kO9ydOmgeUCN/0b0J0Z3tWFXXEj2
qpOmlUiqHe1ne+5Xp5Rhz8EQr8R1ZLIuAIsFHA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72848)
`protect data_block
WueafZW1X4mmou0UAwfXd9Ms1QRX92v5u35KNTE+rTeHS1o/xjX5cBf9n49bTLahc63/7T5PcqbQ
N5l1WeDhpldPTw+oA8/EUUl6w1VoQoxnU+b8mD1mw9lksRTbsLhAwxVbdqbH83vboT0zUdEcXy4m
v1LwM3x+SSnhV3ZbcfqRVu1ZURAmLAhUTYpAdjBWxunlxNYKJpGTl+3P6rZOk1dDs/LIyh1xovVR
KNz2fcyggt6FJOx0V7YipTVgnVya712t/cUXGBi+agipeXuBwKexDM0dvd3m21KSaPS5SxgHmvEx
2ahpNZZPwnNnmf9s1TcgT0vllEPVnoHDv0UYRDswfjq/6WYsvIdXNYujCip1bDpmmhhWGjAxwpo3
EWwWknJ194/oBE4bhZ4otZCXfZYPN2W8PI9laLkLEdKTjyDFIIohS9PO0IyGoGMk7Ez4kWhhKbaL
okZriXie5pTxUk4V7S1L/03yYlCCkPaoHWXaWW0V+RyFJTZOiRIEnkMOCjfqS02Nwos7EcaXX3Kr
1mu09Jj6FwOHJdiN+MOrw0bU/T/kVw3yciH20DfBPkTu5ZtetukXzI2D/Dqb9Zx+VqWE710pTrXZ
KrA8aGEKNx4z5P08VScsT4h/6DMGeTlQ+miVk+1X3s07YAIwzuHvyZhCPOcnYie4mAO5nUZIeTUR
9EU1FDjnMvORX+WwQCqBsqBJy77NZWnlHUwqNrK4Wyu+p1hZWPFmtMSyVbJwerpOUp+1JPDXfVf/
Y19gvjQgFjsaWrzS7iweMq2JTfwZXCFtE/eNZCqK84R/pU5TZr2UMYBdm35qydQvD7bK8+YDj1gK
lB7U9w5V5i4JYNIJWy3Jzy9OftcaXMVj2gN+7FbZRzsZ6s/JFUMFybh9usjD1AHV9CpcMRlYikvH
FkBIttylOf/qT+ekTuQbtCgbrDJR5cqp0EVGHRDVUAfGTtwWkOrYlnKI9kFwyPebl2Y+cHeQ3v+g
js/Q3Jqi8NNEoZWCW9aPRAzOQzxxF1ZSMTJodaqAPRSKsZZaee+973zueeoiRXABLZTp2CxcKyp4
gd+2d8VMmnr2vPvaaQ9wYsWW4rX6RixP26flvHw3dtdN7rcwm7syqx99hU5GzTAIXpDyY74Yk9M4
kIDdjYv/5p2bZAMKqEpP8pD2FBu52mjIgE+lRTAIf5QfB8AY1YeatgFddozswpI+mj2DeCXjKqKx
sHMywwCgTWFf/macNTdx1P5R1teLyorlqsdmwMQm32pnYNh77YdrqHMwp4C1jNLGVYDbdyQCJWA2
Mct643sT0eZMfjQbm59yEF3VkVNY/FDMFC+hB1piu+SCMyktJo4WX0b1QlMdqbS2S7Y0GcP6dBLh
Eo/O4PcbSWG4TO46MFeKixMIaslrWZl66w7x3AJ9QfJldrDeNnqFFdb8kK6J6cupS8OWBFCOAdwU
TdJiPuuGsCznsLvrmEiIfi5SgtGK2tWvolM873rSqrGspuccFgha5ypzEh1e4gtM0cXhll/IBRr0
JhOxPlQpnkHouIecJJWs5fSJTlS+vZGcLMSui5aFptEbaclBYBtxBfM3BGQfbHE0MdJPJvimilp7
nKd39+ailr58eGdai403umG8c14EG6BSpVC8zxHM0v1aXJprIJHzXhr1Qz3RRmEODwIvqGYfDZFa
YeHTIVymUo7Ntg+pqdnSqf2mHbBLa/G7q7F8CrAjY+bgv57dRk9JSK1Hbsnx4FH6TJziJSrXYWpH
UpR4DtGi/T4nu1C1ljf9TQtCBB8uQkGI3SITh/rQ3Gdrf0u+I48YYfkCRJTTEa9Kp3g+e/ih8RvV
fGOkt+MDr8i23T40vKk8zhy7IFlySYpCZLTubm5W6vAOPm15kFayb+xPSwfHupHODl/n0fjQyVAa
0ZcQxBYJi5dxLZkxoDb9mY5iO5NMGWGhrFYuDycWbk3BJ5W46WSYgVG2B+Khf08PNjuRinwVPe1w
WbElMqsZVCl8N/Rp9xITCKvEfEA1JHtyTGW3h8PflkphdOvZ+tAxgfjIONBac0NZ4DZVy7rgo1tu
jqa0vk6gqOgi5yLcoFgur29NbYlqTAmZjPlQIxQh1wveI1LZOWoLiJA2FabEOpz+VFEHo9Fm245+
rvFI7SHfEA6tqmqDhLlEwUx4h+sAamVHQ8F+wg4vU1WwJDBN6zLSHYavRfVlla2SOXjKcLyFrAlL
ATyYZW7oye6Vr80NP5Tz1540DEqF7IPrmeCjce++vgcfIlDVMUeetj+DGVKH9Sh3Su9GtXDRlB1I
UzwY5LmkRifcR8MXuI6sU/6qau5ZG6gJDLWiOwsahbRUezjXLJx43At3Ow5pG4vMQTrGXeEMDZDt
bT4vdhrZjtbd0D4FRN4czqVunPKGca7d5j4m7Fg3nmUySKeP05wTHdOUxvKPWFCxENWynqioVvNf
LyhYPOYvWhjJgVDfSm8IPzEZlaAcqLdr/Knpizxk48xAhYvIGyjd+mFjnF7AXNK4J+doQxvqp+uZ
PdKjs5uMrcb82AlqTvSaGEWizg6U9yLrDb8yJLFgizWRifEqPjk/6x9+SrucYvnWmIMi4RmTLP+Z
WIQC0vLDIpihhiroEVZqhEjCXFnw9A6xKvj2XP7Eyj4dSGkYq0FcjI/Wc5T419wsf6aqux48BRFn
xUCVQJ2ep3+gTDBd+sqUS6vJnKa7GpNppQ/CP9kzjN49CjwvB0gTz6VVp+V7H4xHKYyeoHkoKbGx
sPBPyk76myXc9IM4r0/ke9qGfKFbH8STg0FQvNZssf2AkpTppeCerjBsfm2ErQXvYf0mcqcBaSrj
cxD+L8Kd61M7sE+aEFpqEfOKNb7KqTZd9tpV6nCQ0ZswOAxcOGEqafBDgQYCSw26zz6ORciyoRQV
OYwLJVEyz8mPy9FFRwYDDqW5dYdE0V6k7tsLkfREWPcnZeLMe52CyNEaj3fLZ56+3JuwhzeAcGx0
YzPzCIXL7uv8rosZFOCuJ5VDAxSBb3ta6mHZ6xhKLfFCuyPZFo+CEpXFxSBDXAG0pCXPKd227v+8
A+WKd7uktyButtwKKA8xjCH32VpM7I1il4lf6QeLlyx1AIYkYYoZo7NM7WL/zXTdHC+BcCdrsiPB
d6X4F8O74vnp1sP8QqUfACelnU6mDV7sCsCBLVo3YHGbajISjhioma1VCPjz9xu75TOvivDA9Y8x
UFUZXjgxgsfrKlvUj2qn/hTHYMex1368WfcwMOWLhGDrDrySXRjuD2YZ1/OS+IwiphM8WUNr476u
aDqq50F1pCxBpgPld7uUgODEFRW51r9E3nhcoXIeMpJwmm9KH+M5Gz/tW/y30rTuO8lHVwTlrOIV
zFirA5ht20GGCTjjJMyPK4APBHh4+tqGqpbOnvBU1c7x3/gKo8qB7eZQn0nf5YBmsfGK4/FUVJxC
JoYyPLKwxDkApMM2j0NmHZRSGrLdvD1ROSLIRJm4koLWWHUhp4iOzpC2EyqkVy2VfZD7lYYNqFdx
MH9z2q0VvYs0GmolMxGDBqxsuW7sZfVatPbtrTeurnp+aZgaOSk5DzbYtgV3IAqboaKOjpXSPpst
tGnHzHJuLAjVegEANmP/U0pB7Uzq8i8F+BIpFtvkg7t/PD+C3ktSZTgZp/qUI9avIthd+XHBWtKL
VZoBvG7jtmsyLGXvC9ENzkeyDulWvqWm2Vx6Cr72DXkt7CNQAKrpyMNFTQhyUhZSGajUDUPIQYwO
4EGw90vtAGn59ocXFv01MIFRkXdfjNrhBvQp8FBNbiVu0O5kcaeTlPz58hUb7tIdTlBRj7/TJswA
wa6Eho+Ux3AYsLIL2PryQnj7mTZzE39RcywxPeePkwJHlKjArv4Q6At2HGE/6vyrCtTC1Gu9WI4G
uefv6yRNf03xWUU2bOmczvEAYeQxS4v3vbbUdHwh9/4zAAshtH00+OQpw+maj7d1F60O5N7246kE
hurM6kANHyfkdJOUUEzzHIOPobuCMLImIIss3DQrxS9lWaAQxZDtqizBdcigQwO2IrcvKx56OU+z
NPRgYxyCpJc69mK0dmkSLPkdEI9SDApHODp5f8PEBlO23p1sTs0VLEMZK+EkWPXE7i+EyyNxqAmp
eEmbKO+CMIcnSqQeyvN/2k7RkeNXNqUg3Pf8wwaKot6gCajHtO/S2WniaxinJ8Ov3E2qStBP3gfq
h7BG4NXwWxpecNHiWZUp7siEWTg7vYk96PhIV2YrqAL5gq4Z20uIS/nm105AK6wRjlHAQENg33U2
ELWQX+g0aZU0M+LdO39biwqmco/J/ade9yJ/Sx8S4wGLlZk3q01SBatkkmXkWxHO7gur0P2o1sL9
nirV+k/vDnGz563gtKnktCZv6QJcf3Wq+3lSSxmWaNSxGzGcNycUc4qHlQ0x8oA7PNOhwAeo83zj
UWBklkMcazcE546GsAMXoBdHWhMb6Yfncv0eqRWlAOp3z1i8Mzu6RaXmhZ+l9lzIFaBS/57STJSO
pA+iJ+gKFM4LFQyboOS6AuucwywQkWjyt2qBBETg6maieK1c48pGlAMu+4g/4X42+2yzl2Laz0Bp
krHTGabVJIdYf7Sa7uRrZkPG2DsTFmvC0bzFzS/QqxP9C+j3SG6ghQW8zyI/n5OJjNalVsUnNk1i
6o4wzoNTgKSsfRGlfzogSq0hGqlcR1L7uQpy+cytzkT4R9HOfLR6x/D4H+HtgRXHZRaAlt9cVqw7
ssPNhcxbU0SGbog86VSjtr9XP6E9iYZw7ikyFuA5+npMw/G6TXSNlkjTE8Tr1YaLEonCJMQcn93U
NUD9JB4fyxy54YN53Qgnbv0pV6Qek/AKzm1tO5/0dynvw3pptEBJMDgXagJtQPgzbDXnY4lZsZfn
p2js6wg0PBPlm6WZwm7fD7+1LD2FcyFLZoQjLbNvhtFB2iZ4jA8eCp2+rjJVCkvC7axB2f1l+7Mt
TyX/VVsIw7ziTgsuvijIvsm1P1BjxaNZzmMTBj+ceiKoxvFINb3aPh/5P6RTtUPcD7x9LGKM8l8S
DyVFJX1uq0NKL5/OczYYNeiCWQnMriAvvpR/g1svzj9uOZuV401LxUHnbnnWCYFz/3IBKBtuV/ed
vVx8RqnIfskmHYaJtLV6poXMlt0zx1/gMWCecbp0zMeE5mxK0j1TBqK9iLwpGJ5omUFb+IuwzBfl
IQzYyhSiUohndzk5SwQ8LmEHMeNfkbJzgk//VsSQqMJmOtOAl2ZyBwGQMenounPPrQqflw+QcG22
kM6FPJN1EJa/kVcw0nG+r8gtFenGu1+b9OfGfOZH7BH6nwj4qbkBtOcC77yV4/Wh4ollT+r3Uv7H
GbWK2AHstzwk7k13FBHzzEUcJuo+delpGL991HhhFzqhCCAmto2bksS2BW6h74jqzCJR1a95TXVT
mEyF/nxkXJ21jLgLmqcKBYp+a8kxNEzEIDrpvXbbvOqOGBWItVwH+BpHl9q1m9nUsMcifvkqDrA7
AdLn+5tg8UaBAg4gHQWbM7iUZI+cmGG4PFr3HEZnZfY3bxZmSUUi77fkpQY3TSXbiDGxWjuxaokM
XOrz7GcJDxC+llFCcvaBuw3wxnCLDPaYcS4IdW50kr4LBGMqjNIrNmXBzrXIvV7LkNKwie/xak5n
o2scTS78l8rMFBY86cVlNC4DcrCuTvGo5YKgAzNPuSbLcACQng8yRNNiS61yG6XFLqe0e1aXXaOj
aWwBWbkVASX4ZGM4KgTt1g74ghf2MTangUmKTcxJ8uHvNkKhwa2rxtYFLCikxL+5yMTtTbAIujnX
uuw8UaR7nBk6O1EFuHfrdl39yPFCckD58OC+HHuz3XmQmafFNAL+M8u2a1Tq1k5gKTw3vlt8HK1X
ln674n69bZxzeIhBinBLb9cLPxAcCsFVaiAcv+0Wm1zsmneyYciQmfVUcYG4x9tzKpphLjRd9W8j
0OIiptFJREQl9ssoPrOTUsf/QNuCwqvFJXG9WMJc3xWh3fy/nSCvl0aVlI16OPSZDZSQzyF3zBHn
GEh7rbMASu34KKZnU74X6tgzEqO9gc4LYOY6AQhXmMNsEQTr54Row48r7hfiPAwLc9GvGehPiEGs
dWCbbYa5MAdm4pWkM52dAZY1YVnsn7tvB/vbcRML7+JOOMoWJTSi+nyUTSALVx3ipC6yKWgZ4kHk
ox4RzjBycHEIS16sk1EmxlXAg1f6XgB03jMW8yWY+86W1RdLC2OqqMvZiC2z3lgvO8jCMKsdRiEi
P8vzG9RofMDfR7dOr9A8MTg6wyPATe15HK+MeEp6tkdjmjFkH8XhXH/XCoCATKp3osXEzCYwd2su
7CY5GpB1ctmyOdX3/jRY84kPV25ZuCN1O3ViQ+W/rrjxd9Kr1RhX0rDSnMe1+yETegyTBD6aULeC
QrqsiXe1arbsT/k31QY0KFYqc1Uqg70x0Med4ODzMJV/0gg3Mr2h94oT/p+CSERdgAS/3bYTC92B
fgqXXhi9RvG66nF8kU1YL5zfVdDe7mqpgOLZWIwZtgc2aSbv/JSCAojB6FyyCh6oBPul9yUPsRzp
H405/lw1dBAX6t+VIKsR8Q22ScYL8oAMgvDTR3TjOsfcHZEB3+jE5CmNeca+4ZpYhvWdINKsYVIq
abeHJPBhhfcLJKXgWMFRHJf9h6UnnwHwfNXnJkOQIipdrKHyYQZfYcsTlSSvId72D9OyJiJweDZw
3Q8ZCCJrpdnEl52NLyEzi95tl9e//oIVAWfNucXoDPYZzbDwdKo0CY21EvS4ZtXvhJVe/Fg4SY/B
5DVKTGqKjAuyvtZKVBnC1w95bN0OZ6fVr9YwiPR97nFO1oys7bxv3Js3h8fUSg5iNVVheU2SUk8d
EXDkCTcgDe4yyZVzZeDLOcxpzRGlLIHtaYKb26WmSD7BVRKRZ8nBM0xZs1xK8vv6WSAlTqMbGEDe
9ZCOFYhEiJEj0ROKYqsqCDybQE0u2K6MlrqSGCsenNO3xyaoZy5bxPEkK2wE2838NqwlTSvsEOFV
Pf/cWAJ/i1lSQ7Z2w+y6j+zcmSNsJj9GpMidiIv9ghQpzHv3MYCk0mRAEvvtOGXqcfuKx9Ub8twQ
44b2z/PvENGp49/WUIjMwf/ZXl3vb5hblO+Yo9FMW+zg4t7D8HP9FF3yOZJNZncUFBCPncXDHK8Q
/9LQS8hx83GWPyLH1Gzp/xaEgR2GDnbYjwSDlB6Hz7TuqkdF6dbfTVA7yoU6LxH7u1pEHfZheHkj
r4FytZ6ys58b86bCuo9Ho+x/VlomSkt/oYz0GfRJqZcd3b88nbsQwahvEnzZ2J3WmKFPbKUHbjHB
r/XZ56L0S6EuVb3mUHgvOvCs7+EekG4B0vtLR5SsUuNqSKXhSWD3/lPC7g9HaE0X6fmtPCOnQLeG
sesM3cr9lj9O85usTS6cPy/qWBTLWunPh6ONYzluZFE03WGRJ11I1v2ktasTtx2GA28eDGB06uby
dXoegec1SI0fIvCdtyMPzdU6vsenhnqbpX0XdaSnmS/1ENcSqnmlK077OdBa4RVuDi6G+9Lu0dA+
Rq31eioPH67hFVbJx/mIQh7jpvIINu+qbugPPrf+DsGCU+qtxLTC5Nfierwz+phxgqY+4gL8QCkR
4oHGJ4Hot/UvSC7MMq9bbqPym44Pt25P1bs7bKos0tk4bVjkQB9LaNkKLznwoDreqwWszNyKjjL7
u+XCNx0lxip7GHkhHVtxQQrPWYk8MtEJ0vaje77PXvwZNWYmVKndCDphGjxUkwTAka6d70eQeHP4
APHwtMTLejJ57ZHuYDdPtT9YgTknIJLmVw35Ixx7yBhrlHO7pyRS4H7JGZB9RtutmI2No+wNIpdp
3YPFgifo6vBHU9YJcLXu43DSo4XIm7ZHJ35ZpEECtcF0SEpurwUeS58HUx+qqm8we69DSC9StYxa
DPR5pi99b8+Sjk4tUKm5xtqImCIWlndP03r/57fKkC3doLgq5ytOjyJMs9Zi9puaYb54NC4aznLG
HzX1rjq3JFseMn2EnmfoLwTxZ07yBCQTtxsArC7ucJOZCFM+9U/ciazEcKBlmFu7Ow/TF1OBDKYV
ON0+SB5+hRQ5XdRpuxogp++tRqdLnrAwWu6G9LGZLNKMooxzeYL9c/4JDMT/bOM7JvASm3iuQn8c
7XyT0+HaY7hfXp3nIQb+/4w9MLq3AqJFKnaOzIIkiUCsdMt4K7ak9vIzcop0jSD2v7lhRjMWG9QK
yJRurAeoJd1PfiLUcaeh7gIg9UKuoptmsgdzO5xOd8yDPiWXdPYXl1eZfOYddSe5c2KGH4hl6evf
RC/BSkh8/qHLhr6vHXHjUsfSMpeC6aVH2D9vNUyTZ79zZvxzX3heonuCanfpDFO+wBqEGEh31tjS
ujsAahSIlnYAeSZbIlrmvMxcK78ODiQsDOs7vLEnTBdHni4QYolrJBf8nua2ahP5dvW1eWERKNHX
EC22Ftfugg4ZqHLB09EOhqM4vpOxeT0neeLQBgMsZ795nGq8pCgUAGJYKJ63Fk9Ny/ZO9XPEF2d0
yCWt2Fetq8IIC/Jjr7d+siCsBpSnKENo0NYZRYSAbAT0Ju3yCPDS7OmlZolMSHYztQKFaQ/poUvi
tuQ0/go4Q6KyJTnmdrb8CkoPQI8A2UNbA3OaIUEuIuIu9wny9U3mhNhxdox1USBhp88bP8oReb+b
+p9QkjivcufYti9LuDfKBXDiny9b67IJ2fzoyI4cHdbfG5FKZ37aiIVobu8FygnySFpiNIl5Pcf5
kG1CG9yofQVnMId6G/V9QO9n2P795dnU5L28iTTaUqi3EbsTTP2T/jE0IYMDL/tJsWTSxJt4nJKR
99etlJ6OquP+iLF+fF0PdDN1OilYGyxG4gCOqF7ZF9FEFMx5khG1WodTVrFMf2Sg3BZjnPYCIZlX
PdN0bdgieVQuip33jiMurOtFavt4oD69Akw+/ulX+O2P9YED6Wry6KESBf1CcltdXHQbykNH4F0x
fVDqZgSUA9Aq7iJ2PCo5GYHFO/zKTt1UTuvXi0Zu1zqKCmRoGjc1J+eTopBGtOop/bZhpZGfn4v6
ibQSc2LGzEMFwut1/fODsUtAMO3oTYDUjDY133TCqr3hguPqaVArQ6A3O6+j+I4w99EZihzhHq6n
u10SFwzwAgJO9xBO848YRlk9T1B0PHw8PqL2mkZQWe5x34Ov2LyA5wb8pev01Jjk0xyYjebdEicY
Ml8fGWHletmc87yXE2BO8i7uWRpeECcytRBRe7Q7bv19Dm0pLZWNxtu5rs/sZ9hzLdU0HxwXIZGW
O2JKUEM8+LlOIdEz7I/eD5DB8zVYRd8PqC9Vp19TKRqgROkLcALvLxZu8+KZ3rnfG3hQWNH/HMtB
ktb1tkmgUeR3oOJgadIyNOqiSFrvaCFovLrW2FaPdeHZbThxG3TWpol6GlZhxKxKbDucwleyKJuN
oxTeyNtRJjZ6xV2wIVwhW5mzOgol3XkDhdXp7JLR2ZYS2rg8D+f0bh1DVgefxsu6fMJNT9AerUNd
3E/emiWbfbzgXl3sjoFr3V13q6PWCjHo6s60NJ2SxRUzxoC9YZq+/Uey/P0UMV37SIbJLOPqd1Ld
fz9i8yQy78ZP3J0I2UMK7fQyYDTcx0hakc6Ye8KPZRJe8iSHaN6EPmiyxliYK4s1wiOVNiEgPEFL
jmvBKvyJ3XdZkao3c+0JyF39UHV7BeCwwhTisLvzoKlx1+t6/D+iYx+Ivxm6whauq9AMsuhWxLEk
swg0Uvk4dTlPprSap2b+l13h7JKwDJnlxDVuuyoG042FZy3F1p+YPBE1CT2UV58LBIoTZBhffxsu
xUNwxGzcD/0b/gYpBwPYf4wijtFlH1JRC26QYpWJGRELOlGk3iP/6PN2/bX/wJu6LOS2u0pkxWrO
Co5TlPv/kYu9eU4Nc8Wtq53MCiIpnEAjQTlLbuojTNKcFFKjcacjh5Jy1l/hr8awEZGPriSpx+v/
g8XDpl2Md3yE3hVT2CPTc4KfnyZ13YSO8O3ZlYki+RlLtuUTAyjNaboRlSu9L+7/m/0ljib5+ZWW
fqPHlu/Q8AKZ1fc3DyOu5ThuAO6wFeFGryNdTmgB/rmgdTlZyOz5qPm+TZq228VmsgixuvPxR3D4
u2NDJ9cbQj2nPkLr7YWQkMdhOocifIwkGvQm2UW5WjXWkHrpA7xGP+ZSSG8jmRgbWuy4ynrplaWv
oRpzic5NRSFsDQS03nL1032/jraIdlUcRAqMF4xnC4MzLNtBzcCqTV2QyjYMv54OynqQtdd4oxI2
fGvpvIKlUi3eManPCZ0AAQqx93H2PGL0mPSAzeMMskECN76zknrj2sU/RvOJ4M+vQIGqeapOrqSc
CAjfZCNQgxdcMJSHA47XEAwMOSKn7C+4AyFWwiFSzOf+MFlBxatIkO/NUTpG8FZkuhjJ0eXMMZzP
VzMXYjNP37deqUPJDY6eVxEzp9YFW8sn3v/qasHA1oClJm4imhLSrInZ9WwsgV7Adlip+E1TTAsp
EtZNIXKbDftshGhcMSqSO2cdw4CpP97cZj4wJZiGibqBS8sMz4lzYCZoyF8oZHYigY1Vw5dwDEww
z6M+lnXQZaud0LbFZXhTK1Vl5llwfQ1x46Djv+sbTqGhy/7uaRW7d7EI7GmEc8AGf2xdSZ7QC4sp
4T/1loB9XOg1E6yaV9c9A2GSwabtmvlMe5w+ml1rEAbzRUMD53wQ3DlOtJphLNioTx2EijLVbCqm
vjny7nyG1YxJgCPRdHdk4MqvA+tuLYIdLp0q2rahyZI1GBsRnlNSs3r00Os3Im3ScJSP4xFFL0i0
XcvIbxsrQNHgdXLrCrcr+4y2Zrv7vuc2K8HK/gfCHfYJAPxQZQqUbZyV8vn4gMoR956+bE7w6hJ7
P2Cb7/omO7M0MNQ5sCy2npNXcrUqT0Rv5EVXMOZ4yO810msJvnwXtZtraa5Z2yD2+JkTfc0SRtsm
crjs+UjuCXWVsa4Xij2IhBPpEW2VAP0YCjEar7y05AsOVztnr0OzypqM4nJBv+Kmqlq9L8bzC9H0
d2vO3YprAxHyGGEtf1pJbFRsaRSYMnLmwjkerjr1M7+jIepzTVcZJydqDhgTUfDznrxwJjFHslIv
AidO1K+WdD1a2YtoB25u1W4P4S7OZcAsq20NCmyvsAmj8bXXCtCU/weog0Wzva7BCF7Q0xDbXu6f
sVNogYVphC/E/bQD6Q62FuQam20OPJXcdlHyQ2TGBjn/5R8f9hCpOrG/1HxgNVWKD9Om6hOsaMxK
QcAStGSwh0mTO/2aUCUic6bftKunblXQel7WwzK2AWQJa6GBh1eFGxE4B+oNazOcysLpob7MB5ba
i4CTTb9m+7rwXxUK0i5SXq2a2BkI2pjykf1+9A9vaBt5QOwJmEeNXRQ9hP+DoernTnahniSNaC7X
2fUytdJH8cpwuyzySZ32oF0lrbz0HMb09Ku9MY7JiHRd1WAv4LYSggqoLPZaUvN67nNDwYI5Ni7I
RlXKonNhmipLknfIWR8sM8b0i3UpK0oBz6NNvr0VqDzH5G0Mq3vlX71QjN4EoPdGcKdDkYuC3tf6
5wyS8N9w9smoRrBk/qoUAfdlaNAGnbI7ln2GXYV6l8WpU85gO+q+u1+zX6i5maROsitpxGIbBwvr
XCaZD5vd07sCeYptlKkyHlveMf7GAGLwwdzXlp4PnAMnvoJBDg4yViUWD4Q55+2rkqQdK5TouSvK
uCqC8HcidMUdKmXKhSGk2hLuOm6qR/hoXvdzxTJtOMbLLH4UdkhzpmCFYr+U7T1ybeXksr5JG96T
+5CCTXuhziI0+/1RiToPpGPL5fcSALHXdMlKlO6MNs8GOrLLoSdTdkODuai4Plw8CmCTydWrtliY
UGzxfs8fPM9FUm5YpT0jGDFXnHAkZG+CQiX6qHOq3yO6osaLxCiSTgEZLPPLUniy05ORRY4/GkYn
Mrv0hRhRd7MQCr6hx7VR978i2kIted+PnHrLOylc5KmnJYR5eyqwIVyPAZAXDjKaw0X8VBd7S/Rb
bGTE6xT67EFf0cDH7LAIfjS+jEw3CrI360ObUGUUQEytlWIrOvVFs4a8/nfnWJuVOdjnFsEfK0X2
k20abzjRxR+n1d8VXMJ2Lz7sGCtBJVjRpV3LxJj4zRk3SAbBLGqSjshI8CrqijP7eJk9AGsON9WB
4RTxKy2B51XKQVWkcYE8PF9DlQHThH53fCPBdp7OMh9jt7BihyRGW8Rak2wInHA5VbeTm5zetArl
pDvIqYV2wMyTPVjtFtrhkd3XK73qINgB3CBPUdzUJum2rpHyeJa+SOEIyh7/gITlKsCbds9VuySB
VLnxNVnABc7eNo0gV6Os8x9gr3uElriW3wZF+qyKn13JDr4TuiXpbXDFgPZTj/3y9/nVTq4Gof4Z
aQUELo2aOpTNzug0h86msyCIobfDLwc7uIPNHG0epcbRZcABV3xVIq8+UUw9OjLApuNtZe7681Wk
WM69BW/cM/jsdjQ2XPiSLe9MH2osICQJl7GlniaTGU16vxq+ON8Xw0P4I1VawYYUIxm0ALzofvYw
tWl2YLCSBJcdCNeVV/TUnBg3zaURQeLfnu4AYqnoP26vRRD0bKxHTo+LVkRHSc/bKY6SbunjNr9r
6r8bQKHpIkmMm80pnZrfrFdNRAA6fKP3lUa58ACIYV8Uu/yQrtRXpEB5nXI5ITcjqTbgIiTFz/Y+
IVi5Wkrx0RfzFIc20L/GPTXXB/yAhNL1oQkWkk0HO8YM1n9p3G2gTAfkjAG7wauATJfOa+G/QevJ
JDImnY+gn7VUkzE4pOv7pNyzi9M0+Lv0wXwtXuLySvCVbLttYj7CIiyOmizahEXcGacrcgtmeLGK
oYWR/jc28/VIQwx0JzNZui0yK3UBHJmCW1D8j0Mbh6V6BOYpCN7f9NJQkDoZ1dShvgyCpqVf8Jei
/hMnc55DFnbMQxPBJI9236hWQn0i3jIezkzwv8FRO+3QGLslnIb20Sv7lMVuDr07ZqxDZN0l36WE
CQYOL0KHAgaUXnDkuqnD7pFqSbMXuKDW3pu1/uH+uQqJgMWlWbmPDvAouWS5kgIYGpprXBcRW4gg
HSth96SMPYPuaUfvXwwvPaxOAoLR4dETpbzWb4FIWhkZaHCzSufPifteelo91eCH/CG7KB+MiW0m
RjITa1lZQxLwgUV6YwOymwG/iN/Yk4MEbpGGBTTxV8AEc5f4tOaUR93D+E9GQFvEGLx2LIecntal
ddSbDySL1PQ62rvhTRgtu7JTSW4V4dPfXh6G07D/JzBRLKCieWnWdGGHGdReB+NqvQllx9bpkGqR
5K2RuvfYdT+VypTXSnm0kTdevmkDgT5WLixhSXz9MUTCeh5aLL0r1b0EEm/ByNTisPFfWlqk6HCv
G+PKyDkxZuHagihfqWNHyhVd+MN2zaZ2+w1eqtsUvvWk0h0BPyvt6jkxVT0PConp5AylaBwXRifF
i9QLHtp/RXuae9/1Pzt5BAuZ2fLMPlnWbncArAAyUEtWCPQ6vAWpL8nBftH5vm+BEGL2esqeGOu6
s5k67gOaEhx0ZEojEnTR6MJp/riG6252shM9oquxR37N87e5D03dWpQz9exTkFPUCk55s6wSRDYP
HApjuUm7AmbwI161lkTHICQYtDil2Pcea8/MBwoQkrEvKR1I9Hk1XedlvYh1oqXdPAmLoalykU2P
U/Ggov6je5XXwf18bnEEcF8iKSR6hxFXpsU0QMP0lNMlP24Ew1X/nOw22L0TpgqDyXuuOrwsvquV
TrBNxZxNc6m4T/YP263ewV7AaotB5eHP8mYozOLwDVuclCCyBVUBIGIIYHHTCEDyi3mnMMADY/FC
L+fGbiEnNDBfdKHfWXQ+hFm7tReKRZcyaEIppDmcHuHj61I5H/E4FI1a74kbmFSzoenL2W7vSu02
kiogKETWoMCPGDmE05sVc31EqL9PDFUemHYZUvEdkDohZaLukrP9YB+rEwaq3T1i9Skl8Okg3Xqn
Hw6R5UmVxylK2oh91E2IFq+fmM5H2Ca+1+Bivc8aCkws9io9GhKFcOLhctk+xfPia/VYE5MI6/Yc
COtmfFHiQ+qLnP+Ajko2f7V3p7mC+doQ7poc+o61Okp7fBf2mysDPzCwE6o69ex7h5o8WE+tI7HW
H1PpKssbgMdeCzb13MPzf50Y/seY4yydCg2PNyPEkPS6NTRtM7xJu+nMlMtDF5Yscr/l++YxGGw+
ybIxY4B4+8OGiqQALs4TAvzSfMjZksdUVQ6qF9O6kFVYlnP9z5GQ1SE7vzfrVgVqX3Bxd5w4yvDF
Ab1Bhq+M7Xk9oJKSxweYmpfeJhud72mnniDVtIC4npVAain8+Nv4JyWwPl5+/oXP+j5SV4sqDEYX
XAVDAIDCy9aHJQmywrBajan6cmZx9m0G14tI4HX8kIJLOYOfdtft5K7PwKCOCeAGDeuNxleXcBI/
ySgWQfv5HHj3WyUXeGoKv5Ja+XnI4jzsI1IhI3vt1Gau3W0RzAXE0D8bmb0nkibFRydgG4HlP/PT
ScNA+9bqhkQIMEEwl/eihmGSWQTElpMABD5730Lw2aAXajDjwmSS/SZu9Lk42+9Oc5iofMDGDirL
04DlXXXb6LR1O2Blp7UR4fzhWmQnqahsJufWkVYFSeqYZgr1tpTUqgZLY7AcRigRK0aVEOnEfYvw
r0kzEgJIgM/q2op4Dqe0+QWrlhR1kD06nohWlM8Zm+CMOiZWF6+e9l2uSjnh0aXZ7xMxCmk1DiuT
9iBNcVLRgqBM5/UhcgQGCrvSSYklwgZf3KND5tukPSPQjReRVekS3Y7iHzuWHWqtYaHljoB1wepe
5m0QMO+Ly37WvCyfeFM70MeHmLXKOiAJPfTn/pYMbaAzBxqtR5phu1kx+s6OHQkjMQAQI4hZHawP
PI+a107XY8UNn28kHLMxPfR9ZvjQWVoPVQ2LP3J3KAS6lutFzbc7df36RzNDu/Bhs5yLpdPvAMC0
cw0SKa+SydWXfVKzRx83JNhnUmsplv0BRTsGfDPd6FfqOnmc8dOlt3xcI6eJEG5EO4NMfir/ecyG
JFAaxQnxo8O19nU8ttHHcP8XruTpZ7R62OO1u9HT5nBh/KtV8ubqXjWTPS6viHSRSdkwjIWuhSD9
OnjVZNDwPIuLOFat3nn1Pr3DwHb5tvXoDu0QOkZGsZcbqvqFoMfnLSl/vnnvkcHxzNqtbvT+CgT2
iYYfN9bCfl+DnUq31rgE5Z1XJrJ+8frN6I+ADve4w+gCwyQSx4+njrdNhEcFwkTRN2JsGRYFCzBU
hs+55jWWAHB4R2VRsYGHceS24jHm5WAggnCHWwyZrfUAOVLa9DO3yWEIvp8Ffd/f+z62neCtxtUo
iAeXVXDawzKWe7aUO7Ef/4Sy/l70sVkJhrJx5ruLen1fBhKVWQwj87sXMrH+FKw/TTaCm60ClVj7
nJd24RgW7h5F6aLGGyL7jwJ8jDwTYgkoFbPbU+G0uq3B2NqqQMujtXFxZ5yf6c5G9SbwwYpiUmuN
6zKHDrmJIfNlkhk9fGYUx5e7bAgUT4gwuNIBBdhC8/GqCg7OklLvTiVpXc8y9eq6iYnfRZo5ZF3o
chjV4xX9uBHPJNhu1gh2NVcOtJeypNYh4EG20saES6PXE0muM9Yuoc+ABELwD0EfJclluzuiFxz2
9sH9F/aasvzxNU0rutYpX3dSBwcFt8OHsNdx3X1Cj9YSyS5MOgS9bC7AE6OB3BMHtVK724y0ssw/
/TRXZdFwLP3fwekK4Q/wVUDttW8aaNw6sDzJX5GLdUV3gsQHSCMIpmb2NQATHw0NlBuodIpYO99y
RHMSylSl+DPIa5Y/FPq3rDGO3B2pp0et1rACX7EAxNnL7odBxegTJtchvZsOU2XDNG8aOeFb37Un
sSAgHr54X/gH0bK51l/rAweTX6oCANSP+x2oRGO53O8gUe9FExmMdxN6/Ni2+56oP3WWwkrpsfcH
rlrHn6MqUUrUUIIbXxxnqMo8evJ4DGsuuJkTQSa2F3oirKl+B+zcmoKgUw6UU3RW70OaJlYFbqiw
e5YqJC1w4EjORPYI0hnLfgM364BfznscLAlL4eoZZA2wuAN3MA4kUjRWnSStMXaB76TtwQecNwp4
qYU1hVWQm9o69DpXujU2XARKET5DDz0QTLw753B4kd21mbrbLGnTF15feqtuawkZ4wy6DBW9amrA
OFxw58ROW9lLl0ZiiwidgQ2ucRh+F2clDOXLS5w8vR7BDYCZJfqKm546lzaGDB43vEQHFpi9nKVW
oifQS/USi19xwoXTjFXKAZBkNpTKBqKyq5Us1nYKJDKNBecZNcChTi0lGJ9hRHlz/ty37kDUZpv1
cZrztoI6l3sX5jgA2YF4Pq27soztL+HoP/bjdSEw2FmVA/trIP8MMBGPgwjYoYEggF220eB5d2x+
h7kZkl6zDJ7yrty0gJbiPlNkRdUtoRFeYl/UWBKlm0Nr1IR29lCSQIbhlMf66D3DI2K6reradoPv
gACLlRbHJNQt+Ep8duIVZvKOUz07Fmb0IrS0JERHZ1gFbS4cYq7h6YFJFGK50WIYTGfiVrx1eb8k
qmNfefMiWVPUxJvBGe1DzLna9kxZkzPBuxZXmSY7huiK6g9omrXo9L6X5g76LbAGbt39k9qIAdQL
kyunY0zBuOQvu8MMn8L9lBd+aU006uBM1se0RsOcCaJoF6w8rWAqV23iKqKTflqokGwLQz7zjWiJ
xjtqZQHaAWONtgMMyx95Fh+qqfjLARRVYHbUdAxOcP0N3GZN6qIm/lUg5xQwxHZACmmRV7GpnwF4
w91Cd+FDjclX0Au+z0IeK42379u8nPvYdSBe5fWyR3qLxPSxb5iDaAJ7o1kyuGFn8qe+vozSQDxu
G12Lalh14TQW65QX5bDb+3ShLL6WJ3JcrgcqjSZuLJP1tWZPZThATa/gzgKJNJrqD6FJSZF+iZTF
CnCWMwS447BDQs9h0KrX7vXQaO1S7Aieod//xbiOR3ofTdL9oXZ6VMMDTSv7Z1UqcD2G0cGQgGBj
R/43JKTXL759S/jHlqWcgtnCl8QknJ9l3vcHCBKyaZFHp3rHd+I6Zi9Dmly3LojWgbgjnXnhnPMb
97rhTXMWL/2WiAO4dcPV/ddXQoauLormcK15XFmEfuPdA87yxyr+ye3+fVzu8ANmc6gbRQWOmYx7
+WBHm7EGBMk6/P83Uf4gRwluZyQUa73IwSN8+c+ChcE2Bjo0op0iXuPstBs3ZcI/6fh8XPvkZ/K1
MCTafDMXhdPBIBcCpAmR0FYP5t8Cw+jEJkfttQ3h3l0IXbgLA2tFnGrKHvS4U4zRE3/JDlBrKuku
a8kncywY3brYd0Hv0w6nIf616Tb26UaV/Jy3l9mz/6qsX8YthwhUcMVjsS8vxvjbsJuqLIFs3cHx
mRK1zMLvopaWmrYDvEwDaQ8b3iVrKA6gci31FaXRir4fcTzjCKhz33+6pOQrNEcAWd5EF5677TUR
Yg6uX6bu+O1eXCdXjl615HtDa7b1WwsQAFNsaxfpVgPdpO25qjxhduy32f/cXsZhexdaAlcr3HPC
isSE4rqpidYYILwUyr2Q+JwVAZZgkvh/g+yrN76K7sN3+GaTcSqO921XOnRFdO4y/qCxkYlaYdmw
lmmJiP4MIAxpMphl1s/2/6PzJ8R8LzvjSt4fOLCP6bPUUdwjIQOk1oCy1fLz3kzJZMAxrwWDEVml
XP/T18PudMIhvfgcAPsbvTrzJChUoeGjDLGV0kF70hqSK/WDVCq0SiNuK7uwnhWsu0KYh/pv4Gyo
f8SL5ETAVtdVWqQbyFYD9ej5bLWsIMQJXh5+FG6A4avZCuQ4VpqBU7AzO31kPDK/pKU1Vvu50Tos
Ujap6DI1/qDilZvy/AEdCpG9cJ6KlqICN7ltcwSzAP5m9MxlKPEQHS1bYjIJkjjwTeEX5hC9Io+f
HkCAcXuGLY0z9totIDphcoIWdnp7uwLC3O2L6LSbwWXmZbalo4bJ+8RczmUVycT+WJcTb62kL4zh
62ZTLs/zIzR/DB2mf73lHeLOwsE5WYS+pYeO/IP9hFTGv6Vr3DexjnFZDzD4uNwtEis3x0fzLna4
Xzpn0tcnVoyeaUNNtlluKntvQ9iJMYoesZiNib3hMO81/lD5GPurdrXApIxcrO86wS7+xftboeHV
PRnkkIFl0sAmbVgHW57tqukMeFJNJkZ9sJVvb4dsnc6fnGNcibofR3VEAOrZXS5yjdU18CMz7qPV
LQoBUfOC0svVzVM3mUZqrt5QH6EsBct5Hij5ehljQ9FAAiKXcO6mekK63PAKHB85dzrMISemw/6v
/t4fIEer57CeoZWRkJvOf1AK18Ix6DwrSqAIHSoRxLfm1IXwApYd4USNnX0A4ZQvtl78yKWOEuVw
dlbQZQEr13D7AJwFD8x5Kk3VHpBvPV64nnakrmq8+cE5CHljgI7yQ4/Jfph7A0eCpDieEBdfJrOF
GOuEPtYfAsgH6/r1OW41hmd3XgsIO605nag3iQ8qBx/pek/l4K4b4lP82WCYlRWtedeXFpe1h51z
jNBz4/T1bhrzhs5nVoQZLour1iE9TTcjMsrc3QGgmxZf7HO6qxbdiNY+J/DJWMw21x7PxLsHc42P
FQxJ9f04UXKJhxxNg3KX3qL8y2VC7HbtUTNOxPO0vWW5ELak/o18MvmsEqqqMgzjidBVMARTgI5l
U1Tr5TWeQm+DpipSRtOjBn5QPW3Whgn6651Id2fGp4G+JcysqXK8yLITlrs2YpBE0KURNXuBo8Vp
qu/UP8PhpTKdMBuzy0OZQDRaaSSHI2aeWYLQIJ8neVWDhQlJ/j4WUY0ngjmkpzDfJWoMnc3s+9dJ
HkVLoZtkhSUBDHq7aPiHuEa+smY1sDYVusDk4CmaMIiOeAw7zfDnTHRfGnrDikwO7Una/5IGggDe
xTT+Q4rkIKVMZUwHWBbLHmdeHGL1+l52S6Q5szz6az2Mz29VJrpfTMG9O0DANXAp93lDcLmFPI4u
DpvfAyjiDZ66J393Bm3OfbdZbJS6ESmYJ0OhFS7GbjKPWOcO7/RU1zUvBwwRJnSKevE0niaGroxv
aC2+IKIDZmKKwWQO1uIhfQesuFavn9D8i6NArKEABx2BhLB53moXxgDNG4dJ9sIfvInwcG3scCEb
Rai5adJrYADAu0pAuq01fu7GKVA8RH779d/Sz0wIXi38xeMLnlHm5y+buxMycMF0SRTAyjdcQHgO
K5vD1xAns1GV8ig+VbJ+I5cL+AzrTLSrZmNDXCr2CUXMr+F0CKx/x11+y5SOp5sySasQ2goHOzck
lmr/37zZhRfyv/fXLrluNELCWq9AwgJ4nqWdYa8j0jXwaTPMyjOVwFk5Ppw8ja2gv+xS1j20r0NF
upIcpMxyHVPHb+aiOAKDdJ7uX7eOcLcJJWcFjgTLXA8QtWn3qDB6EYOszs0WfOqda7NFeI5ssJ7A
35O7GLnw4w6qP/OtwPmAKhezL22jKgFA2+3M+/VEkdyt9KmMSIybSW560vDuEhwiGeq2L1+bGzLR
qCpBniuxuKhNLNpo/XdYJw/Ogsk9NsgYEGCN1NJWcTDpZMv8J7BClF16L10oya1ScuupGWy7GpO8
/sEIE+ypDubxtEX/dSxbH7w8VbBhWkBXQ6Ikk4IDD5aryABGazUcgN0Pyiu9N2PfM/35w/SW0wi1
03RU5t8553Ig/Xw6mcXNz4MhEaa+RXPrCjbII3AcjESl5VlvwX1lrt9vwUBtN2GLro3JPl0ku/1c
46oWXxLajdg6R723m7i1Ni+6pMAyB1IlVwTG2WAZgKl0aClfnDkSzL20jxZgWKGOT4JR3JTUdlue
YJ9tG1xt7INLblxjT0GFqdMVD0994S0oZh+R/4am+woy8lKa5wjyJr5MnuRuHZb12V2E6wtKerIt
Ux2VrSlDEt4LLEucpWHporDTAUfE5IKRzBqwY1Ig6JxbY4/Mco1JH6YquFCg6AAX22j8jEO60JaB
3MDCYdZiMDctAUJtIpeTgaKjydfGWPdpv6Hml3vTona1h9w8L6h7kDtIuSnwhp9CF5ppB29f8+JF
aVnX2SnUkFauYw2amPEHTKQ6AXZMxFjtKvUMFMm4Rdrzgd6gd9JmRLEha6J9aXIKbjunjsvlpMj1
mw+8mUwZLD1PBBZSzS8wG5nQIPhwwD/yiZS6AnfdqcNxo95ytkE+keInSw/USl72XzbGILJ/BdjF
QmAP79N5c0uTAZ90qGit8xD0M8WFIRHbk60ya2jTAzP6DYI72qV0pAY7E6bOZz7hy3F48v8M0Z+q
RnCgZMTrkbchBeBypCtlgGwzpFmPer3tQKy8XKStymV8B9CF2l1+7naMXzMsgrfZ3tJMdSTAK8Gg
leXNTE8g+QFReATZa7qvOFOFojWc7Gxs1q75zcaz/pMK0GbK+1VKlY/zIz1GDqzlaVCe3k4OTLyM
CfTDWMEuqDieNFWu+5/m96z8ET7hpPw3RW+o6mm99SjwvEBF+hOGVwk/WIglDZ/3+mg5ZbUjn2Ld
G98K3S/XNFRttfQnSV2GXVoXBZPQPKfTMH1vF+Tka/RK3nmdpQcaLtuWIWvWI9UymVXn0umhG5Jq
8CsJLQ5OVBVt42HfDH4smtYMpy25DNDoOCFdhgitUlqTyF/oQxFXVpE4t9IeB9dX0iK2oPfPoPki
IYWFnuUCjs1T71bzQgO375ULn7kQcvIM4sdG6bKRGNLSu4YkRKBJ3Nb6UK/T2hpBNg9YsKcbEbtl
ki5TdGu+hnklY0ybrN1vcnwTg0Hqv3EwVBDVvaDUyMMCdY7DI0Sd9RTW/FtU6gasxMEQIqWZ93yv
qIv44W4MPsaftrAjDWP/SQSLy8lqne3lYHOzmbXVEc1xiB+9/UWcq9RLvAlTxzHn3ntcggYmsryL
AWuI4O6PbPJ6GaBxiAGsrjWXEqi7+FlmcZTN20XJovpXQM4wnYtFMd8wVeQhDtf2NY0Snw/MWyUM
C99/Gurhp0yYmoGIsRoiEqjMSJ38FZ9tcSq3T33ipmOZIbFrimqz0yuU2pjANqzxUtBbwtFV3wAa
gA0W6fd1dEj+TM4JHUpu2wfTfISxjMgS5hu4RoU2Jlgo7E81YbVbFwajK8PkyuLUm6YfTAXojgDy
Zb7kY+T/6ev2xypjwh16Zw0MOThV/tF9x1r8QP1l/ORj+zgM2VaK9pQeolAtEjQgKcUUy2xBnPyJ
Fqb2f89dzBJWrAB0U10g2yBKkoqndJ5HItZs6UCeiep+VXyrm+vjDfSLa3UBGGnS50JzFxELvLSA
VCpVDjYEoN0nYdPQ+MDkhytenfOXF8cKDfyi9sf4RmO5MZ6Z81PolF2UChicxwiOwBUTWNao+3Mw
V+/aBl9BYQ3ca+kv5H5Zf5/3I7q/jWZhzI9xwP6s2aVyLwhvP+ed0K9mcWoM6/9xX4U8s8udWxgf
4RaTO3wRudZncLHxhcKe2ZWb53d/OFbnC4Lnjvbls9owJC3ncIOP1YlYgDoUY1C1G7wFZUsV22Ou
nOUT5dnPl11Kkzo8i/Tsy8fXJZawqGJ4LIwwSmJ8JgaTSzIOw55Q5w2r8M6uaeWYlOQkPW9D1Fgs
NPL8yqbmw1qRCBFkZch9dBndzh8Hnd5yaLc/rwRVSxctgl3hfHYNyXh+0xS9GyswQS9t6CJQQn92
lMb0flXAAvJiITsrdq5fv2DrhojNmDFe9U8KBAjd2AannmwVYfqI5NqmwieJns62kEnmot/0WXcV
fkPUXvoRzWJuxqSu8NE8SDtC/GQSfvM1Zhn2yThMYvAJAPdcmeqJycNrgb+/8sSH36eCUF/G+E+n
T3r9f6joXexn8xwEc+j0vg0Gyo8wSX48KZzPV+6ZcTL5n2/rII6jqRRaQm7xnD/kzgiKaL6w1aw0
G7sAAGHJXD4QNgfCf3AZ0YeX/trqRD3TkYleLKtKhRQIjTBV7EZWjDyA/UvAma2DhLdEJrAbNUbJ
7qdy8pC2kUbXaDbvDEMc4UbB+J8gy5Cvk+JyOmKB5x4encIaW0amNq/xTT+Swy2qEmrivl89wUgI
mLGt+0uHS0sQyIWdHNxu3SG1Zieq3Sdr26TpAr+rvtFpfFCAyW7+D0GxFuekiDN98G/wno7XE8PF
UfICIU9h35UAK2+r2T4l2V5lHP6CdpQ2qbjRyrYiEakDi6zolKjcTmVsajXNaHAzDpqA+yUnI+z0
sRBIubFQ1A2/RA24Ni3IaQuG+E7DJzTVF73asC65r2ij4veizBRRNfnt82OWcYCnCb1GIHsAsHPe
mvHFv34frzIZex+fBPZxEST8Zx5O9fL3UTKWXFt2cWc9LzUJddfErp6DUKQNlNLYn16+dqdRV6Lp
xp/0Qbrn0Ob+7zr2HkFz8Ozvq/Rc/uQAQiUU6+PJZiWk0ODei386+dozlorwOw4y4AbxF6UYmoFV
YKabVeJrnCbzjd0FtvdcXYHoHQTQJPlj90Xhzr+omqdvDmnSQupxPeFByOemv8wjygQXycgQThmj
Yu3b4kzvUE/ZNsT1ES4fh8J4lMz/nTzcR3OSZH1sonpBhuQ1S2M1XUO4aYRwgJtqhcKhIMbGYSHj
YIZRBHVtMc3uNgPuEI1BkfPk5zwn0K2UGrAsaOSrTBiahU0Fbjw7HluXK0M18h1b+jqShFCsxkMx
PkxYdoFYzt2qMObixNqVoDh3TS79OSk5aTxfflWCNrnNKRxCmLGVM7uqdLfwoOVsEv51+X/eKu/t
nVwF3T1/OeJIHYDKL3XjC//PZiWh2ZpsvfxfEzjkelyePJ1EvtagsDV33ATgQcrsWsQ2LBqrFlbO
Tg+FY+Wf0T8wFng9FZ88NeY6KRWS25HC5cnQG3hrobMi4pNevx4a4+kH2kbVWZeMIwgWcxZFxhQN
iIys03H6zptMix56QSfvM7i6b7TbXUhXI2GyempuHl76Er4FZGp4fbaLAkOOer5uA+T2p7gXMKf7
p08P3+sG5ndwAYG6WGwWsLlWt52nlLGJ7J6QQGxVmreXQSVcaMfwVUum0MRVjsgHwImhuCAb2LOT
3n1A7d8fvdXijaj7foQZTJ91HFnu+DUoXqb8N4OB4AmroewUzM78gIJOHtjoLECkXOyYCU/dKgSI
sIVMZqGXcmZx6K6ihw0Dts+1o8WU+0ODByEvfeK7eknf4WbRLvR8Cn9hvzAqnijtDco0MvSBNwlz
Ms9hoDcIz+JEoKzzJfMVGPAFRxnBRhmT+LcQfwlX5gwnC6HIky8PPQ/+2UpxOi8rR/PPrCuwPRLz
WEvypJJc7T17bFqVRFXuQz7UCwqJgJ99pCx0WupHocSVIKCz29ZtgXRXftO4WUdbVhs+nr8oSdLP
zk3H+dvNLDogr85PvAJ5WZ9hlpEb58XcULfU07kVe6ecf3/Em5wop2RgpJI1CnqlkXH7HTV1SRjk
HyqJ1nYppIeto1MW5EGsd9BI9TJ/DW6A1epkx4EaBiHfOgYs7PpjZH7Tv+phYl5KjwvWA/qGo1y1
utl9OhxPx8Yw60KXSx9y8xeTGRdGYc8Ifo7VvBSTNGrxkfnG6C999tx/AbUogRHwmDs69X7XaOhD
ExqChAj3nBhT51DcW2KgVY/cDRbmCzJw7a2wJ6S737MpptHMAtCQ58CqhsfSr31unrhSPfbbb/hf
PvlpJH1xwQwNUIG3ArSd1P0XjJo/LUBT73iAU+Ch3XjUPHu4KGE9okhqJVTE6IO8TRw0zWR+q89L
0BNHaZBiyIJ0KnvKH6lPz5DX3kquv26UJ41Y0UBiOy5pUjpiApOnixobLulIqVLbBqmm33/yAdn4
S/dAjDLE6Y6peDcQEMtc38VeacggzCA8xPU3SKfMvmxmSluyV71qBOORWp9BrhVfL3tkHFtWNanF
reIFZe/KIOn/Ws6fMEvuFlh0bTdcqql2leqfj8X8RqVHcbOk4dmZAYd6r3ownVbx2VXo2KBh0CzX
Bwzkx3zIEYP4MXBetAtS+HckECpUKOfFfwUjyvpVedotk7AZZcGgS9tY3u1DBjUU66hcGiqrhLcv
5JPuMYct3wJUosHI8bPSC4ckAq8kBgVCS14KyS4IDEUgZ2kCBTHvYMpR6V5/szC7wnbSCgkKMUH5
yoqwf8CjagGtOBGMgHkPPnE7uLEpFDlOearhFMO8Xz32D32e1asWysz5xKyfUaedNVj+JMlehZd+
iOAkBUeR9F8rzj53etrD6ZCcSIRa+G553ALaZkCuvm1Nbgr9O2xMzSXgzGKZAPI1BhNzIYs7a8l+
nMqXfec8ZU7dGBiN77ptwnRqZPPf/moEla4FS0ZJkFhTdxSQ1m1kKTGUqlRX3aw7nRV/y1Gy8xJl
B2UogIlKjuOpla3ETNnZQ3jP48bLWdKM+xCvVbh/l2/gTu2IWWbb+UUInfcvcNAKG8ERiYhUzyjo
oSMGHJNoAIt6bknKtgoEHd1tf1NXLkZa3LXkYEJhtIuurv3/R0Yl+W7LvJt736Uot+X14/gju/jY
AvQ7sNK9OwcU7Mob9fwsALow8JmkcrxAyoE6UfG2xOJzjt6rdJVp4BCjTivlj/Lpsf6eJ1qO1WnS
2qdzRvHUtxrbjk6R//pSTnR3MjIBCaICUfV4JpAIRK7k5usS4KeTGRYED0LJOWRTTGXDl6CtEedW
tozX/zEacKoLocMn5gRGxEqVWaXBXLQvx+wnN2EnjfkPQWoDzRkJUtPb3tZs/qDRw/Hb/7FfIoOc
u3JI7O1fiKmGeVlR3U+222FScAOWn12HJKSjGIL2GdupTSqgYsEDycIve6x+lB7FY9pBiYsvdH4T
fIr0ilRwHYcIHuteAyE38m1nDOx2l/QLcmtPg/OEJHg6jmgwXqHNoWLDrv4LHJFk8hoOEm/km/JV
O+ND9cjadVa60Ie7jMVHfXMz9aqk8RptCXKXcb4OHEJxds2xPP31uMixLqN6FoA+WnUFoW5XOIR4
wYjFBa+MFUMizUP0OGVXY9HIFUtKpOdvSyGx3zaGfTw4FThfWDn54ZyuJJX1T7OVWPLocZ511hET
QRN2dc8u/P/RS3MsbJSDKh33OT0KR9DojY/22Ajxc5wGGIv3Jm3ELnftyHH/V8OAj7iyrkU2xZ1y
CVa5v5HtLLhQM0q9/amtw/+uj4Sje0n9KnMRDaz2fin8rpbVni0DNw0tK0ZaEnfVSL+4YUzogmqx
pvwcTEDHstJyqXWzsprnQmrwjaehCNPTqqjiwvGGeERuwsWgwETmRUhVDPTgNfTMaIRnbnfsyaD4
l+xB7R2a8B23mMyWzStpLx3b+QVcvDrDphtiun7FbRbH9f/fLTLdb0oE4HaND2BEQma2W5gyek69
LNjtxwk7BOBxwJlVcsymtmP7zJlox4au1ESlT1ikCXmL2Kl7Bn6zaeGmOT1NmoZDHw7AledoP6pw
jxE84TUXSEZgAhDtk/UMUETF8Z9jQZQpQ7VLsZA9ojii+HXLZGmHs+CWyxSPorgZII59oKxGZDE3
NvQZ0Y8QylNL95cosWwHniiln6LXLMCex2BqMGOY69FRvh4houMefbp6khmUqHPej53vQsg+cmuK
ohYV3tJfKN9HyIEFcAYnUu8Qde3kKBkHtMS+j0cDY2pOHAEV0vo2ABx+C5XWsEv4KMV2wnCz3Cia
pkmv9sLrr2baP2h3s5FS01jkqbedZStlOTZE84QR2yKW7vcyv8vUOP3V7SYXj1xZ6igJu2cc5eAX
yN8rW8+LQy+BswBe4cCyMqm8820QfuwbMw8ICbzglFEsCOV0wRhto6hDe6Qb99NwSNse0zkhXtve
7mN3vPgGt60H11Drr/mQ6ZrFF3/io2Me9Ii0teNr7kszdpiwOUW8Gb0iHBXxdVQg55/F6QfVSA3/
MOTVHOJrWbTOVJa4tCL/UPnQ5A5T7Qigm7iXCQVI5PCV9MDJpUDzK1PSRjTR2Ms7YOWX212gUvDy
ukVQPHCnVnmRlw+zBAgND7pD2A5zGv1q7NdUUgaVAYVKf5Nuk0vzV3QNf/sIxqXQMnYNit8SRAZl
C68XCIh1+JioGHqiNrhVL7IrUS18cekv+p4qZNRXKSj1WSVnnxIG7hN3Em7ich3sheYV2z7g9wKU
kQqAPpZhjFfRvNH7vq9nrfx1lCnEZHrLRdf2v5aWB/B/pG5F/CrLVMBCPPcqVdwp1OnhVN3MJ55Q
pOw/TJVGt1Q69OduK+3dG83tQ/RDkj2LVqDWbEiNQXOxBPS3Z0YwLIuHCE+Bbpgrcg6MGRSArCwa
RU4fLechfvZIMbewswwEZghGHlnuGMLAAvEZ2D/1+kI1gPwAWSGztT3D5CTSKJpTNcr/kpwDxmMl
eEMq5Ns85rj4JXytlVgRHxXCrXcovYNdR6ZpyQ1Gsy/LOHLwPKPJm/6IcDdRYCwAY0uGTk/m40JQ
Ysx0CRkL13qnPC7e9ko4B4QdooYAGbwvGsNa3RbpIP7+1NsCvajdAnmn6Z4ljbUw92S5LctIE0vi
LRRkH+Br3IURCa66zYiCYS89HyWqpUrECiA7BLC8Vqqpe7hMnRxHQgiiPFnkncfApakXD8drybua
Y7aE8NHo8cckTQEOpwtB/RRFCB7ISVq2KvslSm+/JoWGVQNcixlnudehnYrvmo7HTOy+hHLig8aG
1PyDBd89llk6Ur+zDpLimzfoSo5QojShUqJOGRwvKx3dMmqfC8XzaLB/udVsnnrg23EXa4xitM7j
kGHE2lgWkYFuxkOeXC9ado0NdGsR3fnOS2iWBlyuhifiAMvrOivu0AdvOCFnYEM8C2oX4A8r6MkA
ldhKjAKc4+guuTd2ZYy78636bsr9kQmDFoDjCEqyFifLPo1FHtC9J2X/sIbrhnyFyB3+6/NS6fCk
DAJ0+a7Ha4O29+NW/P36LYGpmkWmhPcw1RWRagjUS7BhPrCw8ujLSHhZGf+l7+3sRP0Pk0oQWsUw
E7jYv/S5nBSfAA2vy15JFgnqWWul47TQC/2E2c1aEOH0YULHVZ2CbPhPrXwv3lSpH9mrJY0dNpbS
y2CM9pQWEhx86bMuoX2bBC+30i1E/KVHCSACZuEA02sPjRcP03V0nBl/FKstJCJvnjHWj/8Xshnm
ZnrAmuFZR7BIBlexW4FvPOczrhZ+6dziE71d3T3z3bGxTf/6A6KAJ2QHY61uR75Ya8OTVYg2BgQh
V5ztjZ0vfPrV3rKUpIIVbKuOc0fAtde/3Ugej3uG1vA39w07c8IMM4OXc24enUD+WManaRTrdEor
rYtjL4iuec7/6npLCrM0vFYQW2rkM7/Hgf52AbepjUOekEntCkAzYHDOqg5OP4pVJ6NbgsCrLwM6
it2RdPzMECbuevVRZenyIqwcknpl0OmLnA9/ge2p7XkF9RGtgHDFyKfiW52dBrruuFl6/3+NXHLx
AMdstwTniG2G0cd6Dby26YtYna0RQ3VEDIHinejZ30K+ANTfNkahh1ngdCVNUuMU+CuH5RFC2tiE
cCZa6fQw09cCtbuMIYFM5DlpDwmpjNH3xnLRT6uZn9YLV6ljZkjDCOz3jLKaHCMzl9XKFIdYK5Vp
NkbcwwumS6ftD/9316zXNjmKJ8hTEZ3HV8EQKyPRjvYKu+KgJH23BLxGnMDKxGsiQDWSjGCylJGA
HRKLrK5FVRn5nqhd3rTzdhG6PemZmHpuNzI0LHtxgdZBs+ungxq4oDd2kRKE9iPM6KahuCIvPydz
CdAtLpgTrj2QrBMju3+HGgKrlhXQurmNMwpYHJkQrvOthe/cHlRlyM4IXz8x/eLKjtrTYkAjBFyT
6FaP/qizDE5GovlHDP2814B6qPc+nv1bV6ZGZLX4jW33tJzXdkB/feHRvTpGsM2mKjadOq/YPf2s
bwsgXCIESBc1QY2WACFZ8awwevHEZVdhmFSY7U5Eoi21jqT9HNHvDOHp8uRozZoQFsJRiq+BzDvH
6nJUpi3o2Cx9xmwFGyEj0FWdfeAGmsto7Jom75p5MG3xW5Bl1l6jzJviu+EFIrcZ2B7fvgbTAlW2
pC3z8MwIyZJi017lM62TLXVx3pDoic2lXqifvNBEZkslTs5Mw6b+LfRO4nERVKCBvqOMfMEGIq+w
tS0dvKfd4FV8aa3to5wxH/NYZ3OOr8z49WUPprghPjVSbTcfI1QUa4LvklpSP1nzpR8x0e1tDf5I
dS5dsDzGJqWLKb6GSIdqkdS+T+HHwRWBzeT7q5KlWc4teGF5udL21dJ5UkDHd/CmwK8M+gOMqVEh
sa06E4fyfDRVsyQ4UZtyBhLDvXpG6YOFgjWfgNWqgElLQjZf7DUqFM4QtCzEjDsZUs9lTGk6O4RH
g/gBfjUWDfVpjz9YDwSA0JO1qA0b1NyrNWPaS69WW8Gpjts+bcR2YpvwXtgKxF68MTCJyqy0WNJ9
FOOyxSXPzj84eCtQ8hQ8F3qUdAtjDMlvtsd5l5ZLUCpMwEoeQ6DteAEt2VlPGykRx9hsyU7W+Hto
4F7ziStVUpHaoOLsItmmNIBBK4TV3dhbvivXoEoHIsr+mRMjbfErOj+N81arR+IYMz4u7CDyFPCi
s9VpCOF3/T7NOOVD5BbTxd72BOgVqjcY51H9gZvWbqzeUBzsImZwmhb2oR5d/xSVIeSUNHmH7yMe
ceGovMPBkifEQ1DuESjA66hAtsyCEiAWT8+Thfb7SZ10iP2S9BjbL6Kt8RTeHYoVGX0myLgtMPmh
YVW6WgvcQQ3Y0/DW3FENDTZtvJgdrguoOaGWTBx6iWh0By9g+jXK4CC+noClMCbdBT1/NoDXEOr/
+QRqh3kQPGXtJuy1oP+OVWKO2ojxMGNuBITR8MyxRu3nq0gYjeQ90yZu2b5dtpOTdXWJtY3F2oSi
gRb/lUAaGzf1+Bb3jifBobKMxvSQg5pKOeTizNk5oyS0PLse3TxWq7BcwXV2gI/w6Y5ikuMgUzfT
TVZjg9HJhEFPMD0kKpyMu3BL/1wbxGuOB9bh7a5fecgtabrMYJYwOJQ3qgw9kg86nhtkuGyY7IAU
l/tDar30YyyECcITMjOf+e69/blZVsUJXG4aGddPULZb8fs/2vR6q5gJe1UEB9UKvXPJrUi6ox+9
FlWmDVRSvLMYqkqqBo55fetUo4bVyMEZeSHebTNCiLPFEwMli+c1QQh8ltGleNpNINoKZAMSlTpO
IPuZAxX9/KKycd4jCTgHauKOPRc2xrVdbHupR/vR9W/9o6l4jMJezDL0PoHbonVMDCqjxiMyZb3j
tGFOpU2ivmSEu8Kt4tDPDns9gfKejNdGhxj8jsG/d6AGCwd09gBseQeqAep3cFnM2fgj3Ul2ND5q
P5oFyU72WmCa6s7P/vhchIHQwws482uNrhsUp994FTtshVb7qCBXHGrqRjUbcHJj1bYSdAsTICr5
XudRbk8C1dfi6MWDPNn+VpVDZuqi7o+NtmHzJYoh/m01O2IEWftFEiG+Ok4QyVZiaads/3MRyuB+
ze3r+ekyFvt0kpPyg7YmgDDNb8wkMweo9WvOAoU67kekTypyY5uLhGT6RJDgnG2upgnMSD7VTgZD
TJd22fBalH2Zhcl1Op77FNSzXwgSyqUc8Q8I+yol9HkDZ7z6p/OIPRXFwFp4Mr9qZP3/FlTby6xn
mn7XLufShVnVoOW0qSrJLx+QzejzwhNORhcDYL614jd0uAAOa6r13aKG/f/G5jb0GUPvkJeIQ0G8
T8RfizddehDKqb7HMwgqL5WywsKape45Hv6qemxTnvHf5vpRGyX8uOMEZkT46eXWloACRMGluf+N
qt/FFzH5SBvIZGe5xCc6o3jLGlzoP4SD/tcvba6WMvdIH4/Z+Hg3Hy3KwLnPfIsN4X53qnvr3REl
ayot0hY9z8a2cPGqKyIUkDlE+rvhhDVU+HFwLiq5qtJ4XaIJ8bQXNE/kf/98zVFcPXUpVKanIg0c
BQpdv1tAh3GLRF0GIshenvwY3J6DAjeRRr1Enxk4D0d3eBQPqRCiR3uHfvyis1hIjj27LJZgJ7lX
LJErpcCsVDtw9x37KMR4XXCgvDBGYaeV3clVkOiib0nl6dO4qLD2JLXytlzWLJy2VmLXuwGWws+w
1JrDpfB0sFTABYDetosaA7RXTNawCVvJNZE7u3nq37Rw3OO5z/FXd7tft474dtWEDIKpPvC5euBk
sXlYBD3fptYZGSiEut+ogTy8z4FkxB0GGUYTsDxb1TuZ1HYW5BArVka6GbQf0YGXw270sria7Jib
rLd2S+bWPoHgHzFoaTNlQ1vStzTqgR+Zz7WfeN1XN5l//xrxA0eDnBgyEwXOW9SNxOF3zOklepSZ
6eExoExJBWD6p/mXIb9p+xjsVSVv2RerNj6rvQOTWpT5qfyAtcjl/as4avX/HYot9MQx5zVscpPs
9t+ravnPOgblyaSX15Kal7lcwiTCQQXfIVHSvfo6mbQorf/EUTlzs3YL164jAXo9U+y3g8M1FRQS
c+zjvZUiLClouxjXEhc8LarFVYhXsrRLzJdCx6OvQ5r0fbrDMoZV1SUYW2lkSeDVEzoPBmjC32w5
0gXLPP0bOiPqx9xXBO4OiJ/MStn58IARYpVfjjDRFd+gJtgpgdyPRIaXuh+PrXteugPc9wVBNnt3
Yjn6r/b9IT41ncXXUoScxutCpvmuBTDF8ffVZ6QQLjMzhklR+7yGFbQzfHU/8LIoXCHWi9S4zi6q
r7as0bbo9mm9RJmGhe5B1MTet2JpvbrgtlQhhHstxrM7aqn80jGsygknycx/2sKHrkPiU1d3eMDw
E5OC6IF65fDVzWldFno2agQXJ7Gx/ICRfhQK09DP2WOonX+NtYDkJxK/H6FjfmHYUq+5LvwTH6Z0
TM5FDkeCjv+7SAUnuArHsESc2wJKq3Ke22Rzr9aKa+HGg36+g+DF/M9ceNQd8nasauaGnF2NTjt+
P0CCKVFrh18YfVUMMnVL4xdOKDrFPw4VVhBBaKjo1VFoSZvbnxNTRPYIJA9QAkuO+XrIqkIJRGsp
q25aeHhjvdKWcDArKCTT1CEG0mNFw9Nd5Hbg51PshBaOflSocQoczwPoZCCvs7wVzXC2e4y5VZFD
yM3IwjKVYl8p1eup5ip2R15bxGHBgu2v/GDCZNZ1NxqaCFwDVchnxXMQBNy+ME6PkhDgMGbguIfk
G7WTGaWseLYRUV/34HOJtpfIfm5kEO6KzurA1VY0YNeOsOZhA5UiRVMRvemyxVh3z0LZzQ0Yjykf
kcWxcuJIJ+IZMuRDO1A5Zia2ZraEbnoESSSymwncpmy38S3o/ClYaH2dREhFyzL8PZZipFFBnKQp
D7gBVcQcuOi6Q3QqP/FWkT861c81c/DyTtOZnLPbMRLncY0Dr3Wxb87jNI1GrnDp5YT/I9Os5wts
Nmj4wNqxgMA4adUyKOQ1kMBn7tKQXRlIlftZIxfDT6/Hnvq1wCfGVqZXUkZ3WlBL00ysD/BHOEnG
APcen5nj2sPYOOH6BLqJgiG7M5JItorXEOZFPEXougpRVAoOTVc1ANq7ijjQAKBBctqN0JgXfrem
gNyVBWLF8PPPSU2qXspUJHzMZFcA32eaaQCUsgWtjwT8hauMC6jW1hTsoSGAkwztxgS8Fv+cLV0R
+mRLDBUDtV9riTsNLvslS8OFxn6nBYr6L59PJAsvliOtFV6tEeV0paC7Dm3HYC3VecYS0GetRb+g
sHQgzZ3ff0ou/49BKaJJ6dvHb45vOvlHc39+crwWBrYE/tr1Bw7MzYyK0yq2tuSygZ17BRqHU4Q/
G4SgziL1BtauhscGixuwJTTteMAyRQMvIUUdw/IzBCTq+LohlH6AsEAsR9+gW88Lb7LrHKwaUXK/
OvVia6JxOoBQIO1amjBTDPL6cIV+nnQJTwqiuD9+dHGn1gr8qg+MYSF5z+H73c3nhoTIrfmeN8dD
b9ZNIUsP4i3CS1XZtLLgqEKRDtMQFbBJbJSEK86pXmOUKVcCYyOC1CfyoLFTaTwzrD4FADN7UwS2
LHopegtgbWTrmoJihWCDs4l7PuBoeOsFBFl8Gv5D5O9uehnzuhIxVZfDsusaOR2MkmvuLZEth5ak
6xSL+WK8AwVkgg9yFAGSXyt/rItSLQENu3p08+tOc+cbg1uC5AMFnXKgcOi2B6b6jK7TwjC08cIq
YaPFKx7MKUsioUFzYIsHZmglrfmWye3rxRQXqbmioNBtYx8t62wrBa2N5TCYBfXBhbc0HA5gYNH4
hG452x3A/CkRnx/nMTgEeBGUdSioFc+XVw2DRXlYgmIleAs0SjyGHfr8Or6xEGMrt3VVAhiWmhib
7o8MMW8F/TgAKyHj8sHQls5iyZKu79XJQ+w62gihDNvdpOZfO50kScuu/nM+b1VMpHI+t2OA1oOs
k1xape6TN/AW6APfYc8Lw6o1D2Fi1gl+94X6q1TaoleIuT01ChK2yeCiJfbd1vR4eXWxG0v3gQtl
sMW2Gp0v3BZTZq10vQXCopNarmsZoJbWHeJnGiKB/v7gPBqPWUMXITuUsH65HRcMBlTUH+De47K2
mW1XEKaN2ztDkejLCLpcKDXV0OPqPUqUMmCeTPSpomT4Hc0Hc7x1Jy610vdRK3oGl95TPgEUMaB6
51LFiVLsIq4wvIZJX1cSCRyqQiMaVSCkoJJB6vCDiIBqDNwm5yPpmaZXWQmSR72C/jEvongPrSE2
mIrGFmksC/Oh0l6E9EF4l6W9a/2tpyVq5C6a7lXuoKP405MQWlvtmN9WmRvPy40kfwxp6KwtRHdi
wNLEJ17UV/dCMZsNj/zUNjrRzeqSRFwA9N7Ml6FmS9PNShk+3O0Qy1l7Jc+tB2y13pf7eH5TxsEp
3LCJuY/YkfGhz28EBp6FTfGapc5wgql4kI0nr8IDDri0e9oiYGDtoNFaiWLolsHy1eg2eXnKLVua
uPVdZzIG37/kdCBkBkNTnHX/FA5HVMKxa6lxVZBqr6WpTE/KDn0NTTDzFPiDLIr/hkvn/8H8PkIS
QF43n/VtemDcP+Qn/D0tTo2SdowTWDW8vkhLy3ZRspkdZKTmx8M/tCN++Vlgh34Sr/ocJe6cZAjR
y1zlpkdokm2JVbTMLq+l4kHPChiSIw4Su06QsjiHUTM3pxKix7u4bYcoTvSsr27rUH6mKuj3dFBF
MNcWlm+caEs+j7Aqh8aRN2vIH8kdRJo2RfFpYWLc/CxnugbXtvAVu2o4b6arZTl7ZfecqRK/KDJh
d6+WLSHiKXc5WxVuYXaCbg+kDUaIeR61NEPY6hnmQMSBqxipeCAre0BUB45YphFnjPcqZ8947+U9
rxxEPrOn1TPI9FTCBwtggJJtCSdIErXgwDZaUI1UcwlvcZOsn+nx1IHq81klXJ/vveZysdt5mQmf
MYY3LzteG2pc84oxbu7ve9rsV4T4Uyp9CtwkxO8Vv9Hfye4qTSyT/aNxBIcLqCYC3NgXoW/mxIw4
VyR4NUI3otAsT2ss3ZvWKgEpwZcX9YKzit67mnQ6z0uI8oXCG4ZZ1QR0xGxrAOnMgINHTI1kRkD9
bW3jR/NvTKfB4+es+4Vj6RRopX9qtNSip5WmBvlL5Pi6v3cl6htZpgzbf4UWLxGx1oMpJMJgeaV4
hv5BuXbzrjR6n0dFhKPVMVTuxcIKe+rEz0rZHlT+ZHpLn5StJLqH+17ie1xVKn1Q6+7dUV7mxweQ
1x3h701tmC4KLWFGDMfRWF57zNDxqoZWp7OOxU/aFcUhhRR8PwKOAERTc2mqrUthEmtpgWb2eepI
JNe0L4IJQhKlmm3cQ+0eb4IzwKD3PsLPQgtXNdeTjFs9UMlQeLCvmtGnEgQ29JvX2A2tDHA1b5KG
U+y45pIA6RL+zTkkJFXDBeIx3A/LGPm+NFQfGN7vSxPcyFhhlG6Tau/7wB3ciY6PRDW4CZHJuY6m
m+eOwlOTfjkO+HPcEwn2TFOMY4qeVHy9oVZGvC40FVEtvyKUoy4SUAlBlITy399nNijRi2/Z8aYs
FR+sJlMdrM/YV3ibl6wmCw8pLrO+65Q1X3m6jrGNjyNbGzVISB3M5f/JOAqZOOvGN0fLgMTMAb0c
CCtBDc7XQ1Yrqy2HqK2618ZVHGoYXCjdgVVsgi69WqtTazTmBw1yWg2CFFagBGkmVOnG5YWxlHld
G5t04ZwFcyO26h2ym6k39fk3/984Fo+DeOeA7vjNjBktpWCuPRi6T5eloh9BOLZWZuBamO+PwCxc
OotNaZC3rj9t96e/cSu8rLVYmzFuUZxx6BFTwJOh3xBN2CzXzf6UYfx91jV+oy6tQRWSR+/bIDw4
iue7iZvuYOcMHtEJmax14cO4Km0lcZDmv5e9MZ2EJlG4cYfk7hF+14WhZMj9h/j1LfhixScnWGps
oxpEf/hDadlzqDrwF5h17m2J3e3yqcLuAt2Xf9Uul+EdrcfE6HYUDkHMsYp3Ym+PYm88iLC45HjN
w+JFROL0pMtWG5rcCnsKtNhFfoPBeiIAUO35Q7DjEFJTTYyd47rSs5laY55Jlo7MsXwS5L6eAwAX
f0IVi63DbOmCDGMiiwSdUl5xQCIW6HCcWUS8S/TcdgwNHDRVDco7t8dnl03/yg3dRpoWnGcD5OmE
gYRx59qGMO+ht1hAj4INSVUFP2oDjUktEDYWywXV3ncyYTsrBY2XpjaIMMx1NtmHA42NqVJGSKWu
R+G6F/dSXdPrY6VF8NWVtlHcwfroJthhqqMjVi71ZtpC7kf71ok9Co13JTUqmlOGLwRBJHeWi1bp
MY4znV5A0BSJRXgwJn6cAI7RaZJpmkIChFZ7g6rTuR8w5zTi55HHHK6MmJ8YSPxbtmKGgQ1gfAIr
vkTaEugUIRhuQPfgKTr38e91gl7MOz2Ij8V2pNkd93hd9v3WoMDREbkne3i0vuF4dlvqk1cCK7D9
bp5EkygXxBI8suGY6eYkUVqgtuOKYG+kPYjO0v2uS51D50BoOWUpGSyiSRgUxeJ1MPGwhPjRR62v
NnOv2FEaZt+UtE1l57Fz9ojnUIAeyHp/EgZU1i8KixwG1LnvKkSAdZJogrh2wKcnE+7HUVYbm895
66CizVHuntvIioH8HZT1Pob4nPYdXSxWH4SXqNTHDMIucYn7vO71xM39AR8a49FCPCy6K4xueAfh
2o4vt6rQvAEmOpjl+wEWzYuix+cG7x1c8hw3m8gl0qIpBuDlIO1dqxyF2XK9rYJJ2tRGLHGBBwcj
br9g2GbUwsDXD8isncki6vwTtiFGoiAWLaZNmd3GvT/vpkgWoViluKsyZX7mxUQl7Rt92Io6iqkw
udWrw4h2Y0yZBNzNMjUczmAEWe54ocOAVA5G/nqQV5/mbxvWt56y3DlabELimOqyYQkn9Ld7G4qD
qTrJEPxFDdtFXk9YSxvF+LkmVY+zOhJ0E87d8NOrWKI6Do13HLGIc0HSuFtkPHyXbO6lVL9HdcvN
UFHWAcLj56slWv/LQGHQgSJ8QjMCwzRmvg3nPSn8NwpzmPA1HmZzXByKrOfDWr3Rp0aTS5WnY1Ka
HJyi5z5U6QSMnUuKMhh/TL5u76W5QN834Rk/yPi+zL/tU2jXxJdeXyW1CVi6RJ4i3y7+bO3LhJBl
Todjul1wkVv2iWMNyUqsq2ooER6Fq9GG3+W3lqVT5/vxVZrTb60x2NWHOK7NGqfJhtuf9ewZmYF1
POFugT3rWIcrWemb57vJ7+wS9b2xJestKRJ2qPmZmxvL/5bCL7DY3eNiWearM47EGDZpowT9BpM/
xcrqv9CbN/8Ko/8U/n4u1/WRPUVV0/yRcZ2ripvwPr0jDU4XgTZ4SaVeZivn6FIfFMOQ1UO6Ip6p
/9yLRxNQLyDvOAW7XhzT15U+5h2Pz3/251fK+YnIn/k0zgmBZ3gEn+3CIA9yQ/20JfPpDnEPW03Z
Or6QUk1KMK+x+VSPBtMy0KBYlSAAdzKt2SRUXyPfMNLDj+B2v9Z+9TrDxwyL1HZ0C19oRLFNWtI4
KbLY1nDd0P5IGwPkypShzQzAqim8Kr9n8NEB7fgqJH4nVzkRoafUvFGzLSSz0uGzdUSnn2ALsiNr
27Zpx1YiFr2ol0oKjF3xo4/vg2ORV6IqaqN8LgUyfsA8ppOf/fj+ypZXmCFdfGXUDG37BZUzW03S
TPqpdSLrarzolj3Cbry5mnv1QpSzmVcfbnvdRmDjc0jc1aBuJeQrejPYlnmMA4BR+eK8jCpzDIEI
iVEvW6guuO5TB/W04crzvB72ZB3cxiBSj/VX4RHFl6Yznagn+N3aQ8rJW0T1EmKQfP2UAQvwODsR
3Vo1Uh5+ZchrhADB1bSwgMjOdCmREY/ZOhQOWoGZT/eQgcJMw/I0YYFhJA+XOsSEMMFB7osDNR9g
BveTckY+6AlT5cMQGI+GUPbks7JAboztnP1T1LIuJz0GFjq98kRxuXbzCgqK/if93VmZKL/CchFo
f+0WC0WlPILjcuKw1JOCa5sIL1b3qbYFuQ8pjOfrJyI4LegEo9lKNqZ5h6005g1ztzkBHqhgzLfJ
jCy10O5N1mxD5n7Aa8TIMb/ql0kLJmT+y13mBIuXZjdABeLj4B3ppeVArcwpyDlQOuqeDpUy2RCV
f/b+vKFYiwF2xDKIRNpXUAe86nwk1ZXPyKSq5RT+QBMQR4hNztbJzq6BxZLek9DwWt+ut4H91vmM
9DXisHFuOR/y/M3kUUDzs8z50WZKE9gPz1Ia0n4hlLCTzpKvmqrgq4miwlMnbqp6AZCE9A7sy7D+
30ob8MhKL99VJ07sL3Q3DgpFkPxNxhrDISgwLjWIIC3tnD/sr0OlgE4ooT5ZLdCNRH5DNxCH1im3
JYM5c6c2Yk1K0+RXEGJ0O1XEaQqIxQ/Lo3k14B/dPFaF8VqCoDrZEhBN4zK1kxPNzzSPxm7ize2u
HYJyQn+u9mZtingGXbrB9jUoynMGrpZ7ni7oYHu1vJ9BLMePNawdI7akC1ZGftZ8mVURRJsyLmfy
feY+UmUcMYtcutvi7QCVpnIqVg+r4O81KK/t5rVMnR+kLE5zncV7CDld3asIoCQV9vFoSHAK1bRy
WkQ0lgSZ6BZCoqLxRN3QlegNssYZ0iufTNMC/QT/cP/AazxlK7mG3Vc2kWRE1PjYDxfzehrR1OVV
IixeE3k95VWG+seRbRz2qkuM49kKJfjD12CIJHeNOM30vvXXeAtW5SwkN2/4WB1ciEQnTDRtjC/f
ZQwh1Ju7WcgfXS3lgFaUwsVEKW2uhUWjzg2Te4fHZd91QX/5Cxj8s9Fvc4Gb1r7DqiguDpOHu2VE
oXtgnF+7jJkz3DeAkjsQYmmaG6Xew5DD0PP+zOBIcDNz0Vbn/gnIEYO7j0X9/FmfRMWomNfkiqlt
M260XqzratxIRAM/RN13l4er1uSIh4L+sxrxbLasFOp8CKM+Qk0zY9NMhh4CB8d0FC/ad0T//82l
TVOLpXP2yIOqlr0dGib7QysfB3GevY03eju8O0Tqhn8bHh2+aAkGUlmWy0BQuYSp499Y/T0AnVvK
Q6FGV4ExElN+uCh30ABLdoVfZNgghkWzx7+699IHGcj1tzQd2C3WPT2CGW0tZQ7hGAfaa/Eq+Jz6
g7E4nRED4vJtmb5soQbJtgbXlJgzebfLHgnNCuI9+2zEP9LNMpsiUbmduzXnUy7SEOmnYqBpIMrJ
biz2fKW2emyt5jwxoxfGWtMIdeHP2VpxfI5GC7WgoQcMvJ2/50Fq2SXF3RccwstIbihOC7pOHPWp
c8OOKAZniaEG1nxTJ+b9Ep4MSSubrkNWCyK5+hpzKdl01eDDrCn2v2NOSCA0dZ4cPeNkP8vhoE0p
2SdnOLQq17pwiIuvwXJJPH2CinOEoqP3LuUT2WhDiyDLDjWAHy2rqdtJL/aYKvyl78Hz+pwj+J0u
VWvP94YCrHpaYhUsUsl0238IVEbG2KKBdIesptFY/oZo9/Kk0xXm/lUw9KRi28ycCnSOxzf0XNqY
5OOkGDBMWtB7aOwNYahPXqHSGNEG3r0UzmzuvKyY1H1UYkqivDrmfTKCqwKEXtAVonEpT8fT+AXR
Ch7mFqNiGKDrk88rXj1BpmV3Ld87l2giymRGbPZGNxDjjempbGyg8NrPuz6GjcEJhYHQZR0WXBdM
yOCB+ycCmFIHd8ESADrUVFRm5NJ55JgzDXlK8dTDnWL0nZfG1RJXO8ULfMl/PN1PGzmvT8EWhXfr
sqZNMAQkD7Pihq3BXMZvw6cspNFvwPbpudlIcZ4cCGVL4qvnzlEI3LOzHWPbQI4iPupV0S3aEocv
13cgC86wq6szCmsafi2wfZLyTFxc4ywvvwUyK5FFPLAK8q+sZQk7gWZSvTu9okHieLKRjtmvpNsh
R1mz3ZJQpkgQgououjbT5aytV/aY2YinnmG8JPMGn+uIxondUYPDNpU6NApYQUamkOG6MMPKn+Wa
Wb//2NuRujaYjYDiU5CavRcsAwTNjDbs79gkoEdSf46DVs9RYnpr/5y3+WqkEN8/ZxRcng+8JOBq
OMANUmrrIX/C1Ozr5oEZVBeTKPReC6Z5ct60p+nRcaXIDHd3705F1TGVTiXuxLciT16uQ2+3Ndwy
d79C6ovj5/N0+FnU3P83QM2TEJKhzUkKemWD0rzaj7w45TSKcttnW83Zv7g+k0NIHRCObIJf8K62
2rgVnpmc2udaSvkze08RNMv3ef0r6m/VTLYvozRGxabhB4TmWs7FqZydkrdsU6Uuk/RFSTJ73AlP
mzYQTVDcwUkqjMQfUAJmFcsmh9f1WB5UKss4wOP/QA/BkQsTHR/kZI0FXuA68o7kS92B/ABf/Fuh
3f9DsR17hf3bUjZsN8I/mjx+BxeVXjBjdnZa/RkWbS/bQWc8TK4h0k8hqWOUf7y0Uusuuw85DpKV
tkFvlP1QZ2JNuszauMlgOf+NOlT0QCpmlSHBXmDB6/ZLpu7QXziVKH2lT9JFP6wn6/paitZZLk5P
dSCcUvgFcP5elSvb8/C11bRUBcsHVP3yk8exaoPqdRCkUkJS6EUKYwdy/o1WFwfW0Qc9ixwwM5oE
/Nu8XyvtGzlBADHeKmnuH2PGroHr+zw2lddAyMUQcaJDj/kBQWKei40vOMUJtOiLUBJamP6UVQQV
Cp551wjMo4BftvSzjrk5Lgm8lg+BgzeXctdiBpiU+ckibUXfI+zMWlzcirt6AqLXEK1uTwo8yJ3t
mJo+5aAehiiQ5xdOLyA6/O0TAEtzPeAoYup64GjyHb05iQYGKZFgIpB1xKFFQVKOZAAcesG0BDFX
9fdLXN2zVeID+NnjZPDf2s1bqBKqaARZce7EQjuTsZL0tGWXixA4szZ0lsP7ugnxyyiac/dRkSGQ
wkw9kyPyX5cHMu9Dv3stFdjZEqXG0aAG/+fc+yTwIdQ7mFmiY8K435cOCMeCECk38Xs2+qdgYNH7
fi1ztCVDsPzE7LDgRBY45h8NKaQ/aEWdsLKxkBYvgBaquu9ZA8P0ILlKZ+0ZzCzZdESOAtXPsu9R
SMB/eiafG2I2C2S64rmDcot3ILQazY6oQlaMhiF+8puatsG1crjGcYveWcXhN7sGfxZFwEMyLbdY
6r6Dz7d+zunKLFWzQE67UfqtmIjLMi2tYWekD7bpFDVlOa5TGEfTsWvByRlHJcazQgorz93sWd7F
AOAypY1AmN/v/BOcNB6YR9awhLSpbG/kX12CuXZxss4BlzZllbeHY1cCweLZwa7KKCPvdFkLgYsG
oNyAmihxUp5Kp/WMV3Pa0rVjgDsYqIe5DjT+yj/IEpdSGXb8tyhoZyT9GXTFpGOPkLNpzQryi0gr
NqfaHl5c0ruWU7yp1Zw5eCwwB5qXYKOEcN09CYDDGe0VoJG9iNSScz2Igp7Gdu1w4L19pTCQZjI5
ltJdBS6QzHgf+08dB7h4reXezFPJCb/tQPtwDkUTd8o8Bi7iCwg8OYwa4sakHl8x7ECFBLtK80SB
DF7WzbM0NIXxenCgJjFIWKgzGYRLt+a7qh3q7FNAk+Sn+sHzU2aDu5cXgwwSVEaAu6CYSiyoizFn
IIyFrz4AtaP5awRxseXRHUV60yc6IxfydH8PB8Yp0r1Y1AvcNw/YDQSJ7XOWFyyLWC1sVSwV6EB6
VVF3ezRcMj7gzxV6v29yh13p6+aUESzSJc58Vjo+rBTHi6MMXBggz/gIQxgRVIDBGw3GW4NB+gik
ekBcAOAWIJIMvebDQJG59lpvjjFvlEdKNf3Baaqkic09Bwfb4fiNY+c4wJ5tFYRNGWq+Vmbh3Efp
A2rsqgI8mWNsXNtzs6ML4URbXD6bAMTvlr09ZjlnNbp2s7GTHjKC9HnhWn8zvSZjEHQLEmCYbG/e
drw0TkMthsT2mjhnKwF/uoBBpABC1SQZgRmv6wSj9ykb3pdLUUTg1fEl0L+mqAaTQOxdL9nVaajT
0VwCWUygrEmuxveFI9o2D/uf1nfYWLYHIf5RBuUXr0mMXjmW4l30JFHSbPPKAezYEWiRsS/TtNeN
7fA2lJoBibNHS2uLFsSRK4cKsnoozUY9hSYSl1btXhzIVEJhAZrwsAkJV/gDeYYQX2v7FOZztq/Q
6uFb4I4bBHJ9Y4i0DSqoN6huBRWaMlwZYtehXIX7xuL0d2VBY5mniccnOHoyhql5gjb4G7LVJ/9Y
rQyn/24s/EuMOn2prHUrUSYrko8ouu1WZfUWA9V+YM1rYfPdDEkS8iAX2dq1kt2s1kPNFrJVgTP8
4f7aZU7KvyWbJQ8+wYtjUF9QDCU2kPT9uZzpD7Judoq2nrB2hWVdnzj4o0hjRl752aHD27s6vMyl
yFtlaShsZt/bURFVG/GaSP0ttOxwjl9auWkvmW4fhYvw2P5x5rEKxXWI5r/21TtvAdpGwiqwD62q
nSo1Ag8a7TsUsFIF9Jw1sL+DzXK8RUsnqkqtR5X0HDTflutP5VGDq1zKodkQYxwjjF1jXiDMVijG
lLpt8e+3KucGuTfa3LREMbaeRvvjDrGd27CAnCJEngKPLL3otZKlVFGF/GfwoAoGNUU/sQcqHVjc
pX7wMDAkmj1u7oyDcsZQCjLgin80oZz/GA8feNz4RVb2bD8YGwWgEHSVKjzSPw9I17oN5ZB9lxBu
9UMgmk+xucE2iVdQovqYRsFsfU8a7pF7PZVUgdcMr+QKAIEFCfE3B0TwseGm+yJ83B/dKZavRYqr
cnmFIhUNTnkGgvSOPf+LfY51LHM8AnscdA9TNRQW3wwFzqPlvtYtwks8Wps+/DOK6FdjDzKAtFq7
YhKfZK3seA0bLS4jLsZO6q+IxjKf+k1DgBLPBiD5gdIXknVzkgGcKv1swDu36gt+tWWs8kYY8Po0
YStUJQyXf4D8z/ZWhcxxACtZbZWsPoV6a3vVL1zXYoMb79jNrZqqCgNUKz0/0NLn1IUrgOrfvueU
YF+U04HBB56A/0dfmR8L6HoMqmpwRXxAxVWny8y9MfAWYJR2R9vUORtt5WxFR+NmD+XUmna9haAp
52wdCF/KeMWHRT30VtT8ntj0zf60TI5G8kpozHRJv6TUqAZ06AkOAPujSlUU9tN9NrxmufQJ0SIo
Ez4kKaDDCU2LUT5G1vJCftFppCYixbU0PTlmbci/Mz/pZTeHQKc0QkJBlAaP00mN2uSijWhtoW5T
qxfS7oKZlbgikoEK4ugs3cFgmkhZzqJw9eWqALt2KxuOdeYS4R2k4k8hqG9RyCArahjJVZVwCRWX
JB5ygtnkNhFLbvjoZ8G77ruXvD198jssZEeyT2cyVYKCgtC6fOTbU6yzTNg4jVPHNtCTukRgZDdb
76eATfTNe2grjsiEG5+bXjxxGIMm1EdVzFBX3sIRX3H/dNY03U9CqtwxWWNHo7ialHx5R5/EAud+
5ZLIZ3vejS9EpdCDuotAmmGb4HnPTgpAbrmsSCjfk/88yCDvCVRy7aD007+UOC2Kqvdbe+l0XV68
bQjxblpb233i4A0OPHVWgG/ofrRt0TFDuX28RCxwxydfjy9gXlzLsE1+MgndZM/1pmTfn5GfO7i9
smV2NYgmbYqDWSMwit/7Eu4nQ4X9h/w+Sne/jajrFldHfXURNvD2anhnqHdGySk/O0JXZMJ5DKAj
i3HupkLwzwuPHd33K6sJ77feEMh6XRwRl2FVs/jht0p/178KOFtQ5aOL/v0bejE6vP0eeA3vNLN0
U6cfKfCinmBb2/KXUxptL4U8hu/45FtDcmQQ461HvntTrGggBaIg8SMGcjUoZLhOZhxx6Wu0Cn+d
hceMb2iQvVBYJKyAyCslhTH2e4AjIGW74pK3Fr7PD2LHYDkWyMYt7MUv48FmsjUMcG0cb4Nzo2my
vz351UPDtfzJ6K04KqdkjqMd52CknRAH/C+wl9frHXsRPFLI0ZeyEr2Uod3ZBBkLMDo2xFWYcX9c
fTXb5c6dlwblMvjgV5MQys+7e1jwowKs5g8VeNp/rSLjCZRx0+EStXA3Qy88REP8TuBHq5eiHK73
yvkznYJbG16vcbQKvy7Mj7xYz6FX03tfZ0mD84sFExfzmasE4L8RXTUaZwhuwgUR/Wrg77foSQl0
EG4CcHMWbSxNdcKH9gGANgqknlPoND9GTrFC1wW3o3DBGcnWGHRPz+m9GYr1lgoY3jrG8Zk+Fs8v
CvmMOtywYYjXqCx9MQ610XwKC1ztbnDVFpkQNvsfkd+oDpy1cv4kMDyaIgIbpJC1GcEw60uj1hRt
YDYcwMn7KE1Wg5xM270Ebtt9Ud7GzRWSTEkEMcQRnsYgSbJQzz+cDkRe6KjMyk7wffaCocm3/ROo
UdfPNW6p3eSxRpc+HHvqj0jwcqWntzzYZRiULB0XNyiXoaAnRQR9aME8+EdGcbLg/DU1v7NTIdjt
W2T9Byi3jf95K6JIf0aYV01FNu4q0IWss4/u2r6KLS6QYBcwtnADraO3l9PlpL4B0SA8XWXQjgA6
d6D2QYyF5rS71IMcsT+FvzrFlKeIZy0B+BQ1xVQr0M9w0yDvcJ6cN+G6/mXKjbIXzheE6NbgbiVd
nSmmCxnf2rlfZalQUnWHwRytRpyH/3zvhBd/s8XtKIa1Y4EwwSRpzqN3oxK0404wTaFfQc3Hn24a
kSR4TTvj7PltC7rKCdRn6uuNuyU7OE4qQ/BjjS1sMVHnKELDW9XHJBBawCdI+L/sUaWA1NKULCm8
1j1a+3nkIQ2dTVtVxqEd/KeBzxgLFeA/wFtnXhhecr92LPsdVeZCJ1amJ+28NSpZobJ0DKukcY5M
b8iExNXT56GkhfqXxatNRm4K7VndwE58Gr/5k1TcKkFVFbonmtmCCeKslEFAw2zGqvpfKQN8haMB
JSnPwyZcXl4dEUF+6ILX/Lh2Z2Qemis1gP+lMGzJ+/hpe2i1tum6Ah6wuU3UCyhZKTzO2QEC9vCa
NH6Jd+fSABh23GeFwDmnAyU+tFHE8pe8+jEkcoNS2wsiOBDYUETYjPc0UiqWVS211gK6a2ZG8sPk
L/es54tuvIS06YHScUW2easdvZoMVqnrcwh0+4yFliGu2mGOZR9RWLJiLq75Y8f+j2r6rjAi+2Xj
1ttikOfOBwKONUPRJCzR5uezgKw3dghDDnT3XTApibq8xF8ZbD3+LwdXJ0OsoAgBd0PEIpVyC46V
mxg8NthW9WU+P/Kj8M8bDxZnOqq3hmws9gPH5KDwHeS0SQEjMzUsQwtcKJAiqeMC34qRjJR/CYgZ
7jOhhWXKh3vwHhIe2caBvo0sPmMsqFD8GlKoaaX72ZWF0Z9MXHh11JbAB4DK8+aGMBuSjWj2B/KS
hFnK08WowfZPtyJyN/7TnENGxVmdUDOzyFiyNjziXHlxwLcTk4ilpOBY0HG51v755dRDLAs/bzxe
EUE/oWMRQ4nDBmqAtCuTQs4zVNULLI5C8cAUsb01SW/0TAeJfr8d0tHWzjqA12wwajXDRs/s6tvg
uOvS45RXTC19Sd519VxeeqOzmMX3sgxOJqovr6jJgCb4I/BUoyv9XiudgxuclAKfYyygkAP0Ev07
8KSg0oQI5stDJqS1uJSyyns4G0ICfh2qq4AkDhZxHkyZ8aoFQqz9QbRTFJ8XoHOdRUIoNqbFq4KG
NFF5u0ZrUBuamtwUkn6PY6Y0Qv3z/9yMhb2fJp+L5OBcGLhsZw2lisNaIKYDURzvMcEguCTjOBMl
44FuIFaPg1fSPMw6xaDfcJNZOreyvqL19LI/rPWMnL1tDbrmVOgJ5GMuiANHY3pRMhK7AnN2V43H
YaqXdon5+IXefQ8l9F0kRA50ugu0M3XAIiVZXK1Ym3o+hLJ9XbNTpNlV9FYUu/aTFNnoRtkAefLp
0VUabowsQARPZuQH/tmeMHCZuJe/aUGnGOvx7vayPOy38BJcKDPTe+BHxFc6A0YasmU7DOUKNM2E
4OyK8CyqexNtgX/pePpGsgFG9Ef9cbjNRGks/tzKxlHFZUXjaSDY6nZIo/tI3oiJVVQWGNV1/lKU
ggStbVKLRkxTfQcsEFlz6aqBQw/JeyadEwbNzsYq150GkFPLfmZmhdqbh9ytmMdHso1ltz2FD29W
EDxDIkkUOolPR//T0xmIhW5Nb/qR55pIq9Vypen7UjadRQHpsId33bess2zPh1W0RYXfb4Aj5ZcU
4LejTycL2ctz8GbQynbpweTOlvr89tJekwGUSOEqkir7yMXzK79SBIeHAmnZCOKl7ceQWrIZ5hfd
8bVkY2QIJ4sCzA2pZ2pkU/DEd9r4Lh3Kfgilq7kalwWYMKwYIh+zJK5ihXgd416RmRufjGSZ5g5V
sfwML0JwbAqsrjXOCSdizRvVTvzBUd0KFYYNN1fzphJXYH9pfLkeZ2EZMKDpakASUSx4wzAABUV0
PnEKsmdpoZ49jBs5sbduErm2PdRSQikz5plKNJZv5GzpnuqwaknAV+W3jTmTF5b51Tmp3OS2uU1v
I4HXFqxZT39z/uGcDdsyxIF1ScVho/1QyjPr7SXyiOyyi2Njuzn2yWA9ipBIS+vLx/5SU5yzRmNP
WiO+RY/Qnv9zzZYS5KkG9iy9QS1WfVBUx8Hay4RxjIMP6+/j9eo+yVvldzyhx7P6fX93RHdsNVfZ
WoWWUzl3rp4Ir1ZwMQoFCr2qggEE4j7R3a3ZqnnXN2pHeXTE3dtgevRJsqlnT4bQqgBPWJrWJVFS
zFuWtzjhfeISlOHH+7geI+Px+JAEz4n8vFZdtm3eY9L5++57F/ZW4mun3/+rZXUaIjuEujtcEtSA
i8eKepwMA4TgGTrnXs+HXmdqvTrvh86j+vu0p/2596UU41PZucx/MOu9DVOTTsLwg7MkBzCoY5LE
M58DwwfAX7kfT5UwO4LgyIddG0HqqmXr9lc8m+eR+B+gqYbdbpjFOqB0MmW1sc+dS96G0hXFh/5y
IbWRGhRuV29fkRb5hLztDuq98tIEt1LJRI+BwsCX588A1uOM35J9urIxV6azqcgu7t1W6jx1E4GB
wtvlVT2IAZ1YvCF1ZUgBHyvUnK19E3Hgro0z8lRspn/h1XfIV2zwhq3xEo7uNySWW7uhnpbYFXS+
6wukYx4G9xK5XBmXgfCZKutr9BC5XXwJiTOQbTlNXO0rLL1jE+5AUP9gR/JbcpVUy72fEfAPZdy7
pF38P3anGx7zcgNXb62xtolRMji3rASMwSrv6CsTz+gNs/HN8H37+/zgQE8+mmQ6HUYPjvxLepK9
48mpvnV1Z7B1wnR/dCapgHYvG47ituJ41Lf9M/cqODPPsi0b6Ju16lEc+q8YNiXLSjeIfsyIFXrj
9Fn1CQfw87t6HuHJR2VzX3XHxhB8xxSdPmPfxcgSOX9AgBGV+8kDXv7P6m7BE9gy5ilTaYsU4zFP
D8N0kU+aW/BN1v8feb4651BOEsJR0PJT+/j5mFTw0WdtyFUazboBF8cSIyEQR8qxgscgREAnIq6h
LRP8Bgpvr67+f15gehKo/P59jPhlwE0QGX6j9uPOgcG8+ooJiKA0deJQtBE1R7fWuSoOAi3AHS+8
YWXTNF+wphn7KW2aByMAZKe4Zme65HWzpSvBw0B/ackvyLvRYvqm+ME561cNZv02+lqHoNz6ON74
j2P9Zi6qZjFkZVnJWXAfNfHE7pp12pt4T7+ly12xuTH/aghbZqT87dgny8pb+y+jx4VVtw4bWHHZ
WQI40c6kX4LRK72u2WmgZI5RE9y5FUxDxfD8Uc6Ce5WxuTWigxeaKKPbBrzps34JtkTYRm398IiS
nCOfwX1nYpne8dl1/NxUr2HBdOwlA/jq/QimQfwvFyWWC6nZHNC97dkaUwwnkjXb/cEjLVAKwnfI
2d6W1xGg/crmhUEfgB/OVfHgQ+R9S4yov58l0InzhUMZthVaW0wZDwDyFx2pjJjHwUqhG8ePJ+by
opJe/IGcqqy50dLQZIGcGdKkE4AaV9UTHGfqeu/UvvUrY5mIwuhf7M3xilgQ6L+4lfTGzAXBIS8D
72lRf22/TxXcPJeYScdCKYTRW2R6P826+LiliWS0AbcpRrCecsOcnUWo4YN2DcDaV/jSsH9fhzi5
OGpTVaOMUVF+hnkb91KEKsATTjDmSzeRTYtMv56qDu+EQGV9UoUvIkrYb3FAly7qxsflUwfJ1/iz
q+4FJz53Bf8Gsv4TPmcUpSMnUgXJHcfM2bDojzc5qV1nXvRGKr7GiGY6tlLz6MFjbWkk+00RMyFY
/UUe5EWnwobEjQlaleOi79GXHz8J0pZ8nb75Z79hiUq61ejbh48NWKpfWnQ6f5Eac2UxpYNyysIH
3LZqODVdyWgwiqwxyGkTe5ZIcJ8Yegz87KXmc4A92s83OlbX3/R/SRdynHKQ9LKBZoJd6614gArD
me2myAXowPKQUOQFRArizSfVjd3eYU6ESbU985AKrEkOCFcGAvLKYTdPnnrQESHGnsPlmtmH+X4H
iRc28KNwe6okNxuZYKQLeCFF4ZWZz84e2vuQg6ppy2QgkhAO09I/Af2f01idsMagyVTJNbo0EmxP
NVCf12ttPliyCeaby60d/9hPVnQcWuJX4NJjJ5+jmAJHpbGNJLUJTRrP0qmxmCGQ79xV9wSsmbPv
m/8SnlJPIl9HzwNHtdgpRSnaQpM0k+IsSttdbSCYhmvpXXK0lGCCFdkbNTYPiGMGKzG6qjvmfGCC
7U0D0t0LD0KSfYf2sny+J3TP+dVHa2Wv+jxW6AzcACM5DwL7pzsbERy0SQombTjQRr0zM0+xgmlC
HC6OjzFpahdkanz9nnxp7mwozBRvgfxfPc2xtlN8tyyTZc9ngpFDmw+08deMziz5y8hAm4bNyJe3
ZslePfhY6lgt9IKbKF9E4VzaxOhx2RJGMv2NaovgtWlL5/QwfcAAEm7p3QI20lsNeS0bLlHeMAnS
Imw2gmjJt9FKCF3HyIajZahv76KDNVY8L0nFHh3w4yfKLjz+9R4Z0j1mGf+Ye4+tNuGu/q0DXCUt
sDEsn0qmH4u5edQps15LoJ6hE1JSC7DcWNTU7kguiRQcmFKAqKyo7GUS4dejTOXQcTiUIfcovWfw
DhEct1KZQ/Erk29iVkTD1DegH2Ia8qaii9lsyJuueAPsaOly7+/qMEokzekODC9nKoRBA7m47gDA
109/eaHF/wbFtcQMB5nUkewP745u4OIobOGPLQ7I5JC7L+/2Q20wm2II1Q1S0Ag7E6s3+M1SMcBV
cYj+4q8NGX5Ly0EKtJPO84cJdWFd6cg875QNu92uF4UYPciGmgRAYcWEM+qxSQVynVxlMphAWHNW
2/uBVgyGPm2QDLx6rCNIjNWWpQ0RtD6DExCJMPZT0SVm/FJ4uybsf8VrhRM9IjYbu0y36w1VbPen
1IhTSG0IuHSQmlU8Y+oQaztRppTBKuIBCCPdZquFrgPDW5rS9bOTfUQaMkibBH94EkNe7E4UE0PP
DNHzOodGLamJ+hOk+xim2MzCSQRdZhw0DpdDDM6krJgHN5liWm40hqvsL70mstMv7UziSAj0tc2X
UmkO73zmVAKo0n7ExFkKhDJ8xKy7ZVRx5JP0VDSldR9wV5wE+0r7pPYtUa1kBvHLRInQDOOkugXF
72Ry9du6T0sNA2a2HQWAGxuEyiEeCxaFjM6Lt9/6sBizeyXYIlE1S+RmEAGnzGLT3F8hYDcRB+ga
zASQFHV9TCddXcfdSdxY9G29mnPHifkAEINU5rhVZKKb9M6yeV70CVgifoOp5X4CmLMnp0qBZHKV
XKL2HvfLOsi8BQcG4QQpLtXBaIqfHgPZ8J4uAmQrxr6wtgZh7+3VVpzbxrBY+Zbf5eirte70Z/NK
swE2B6WBFHgXrAIcUhb6DPFuPbntv6vx/zUE+YU3AtsoG2VJdxx64aXR2qgymB1RsXE79fvIDqnm
yUonf/hLbfXVnb2X1Gh2e9QAcDE6eA2FizSe63tv0MoUpWOOPMfPuRhxqOhH5fB9aQ7PUQbaRZfJ
h5/C/GnYBKZKuFSFTK6aZJY4sSo8j3YQA6DMH/6Fe4OanTllwjhQ1uPmbuCZX33d6+byqUoJoWSh
S99OsIU/vXmO2junl/o/smMPlv5ztnuBjop2J8o53rLhKysWtxj/pvbER66JdU57uu9gVXLYEV35
lePe2H5RGsR1Q9a9goaqtDhY1d844fE3J/+LL5sJT5yekvDqAEU4GEHRtB2bnfXFUSKvCoprEwJA
rH/dljHa2uxDQ9CffS5SK6rmzXt5120OYIZWElnDDfSQkRYhUTq/+NISwPEEHawEYVTZEc9Xl1Xs
U2ylocpt1J+mf3GnZUCk0fi4u/0lMioNe+6uTWu1q1poI3w13w1FSeVxLPqAxHQY4zQjonXWoggO
zGyCcQOwTVzvtwYR5+FARLS5Un/lMQENIygXTWr3d9Sfpe/6SNfI8YjTVSziwyWPUoeXq26WsuhG
sBEQJw5W4ziN3v6Pl3yzg/oHX4L5aE369BjutagfZK6w7zRQO+sKohKgIl+WzA28o0e1DvpPtYRW
uKGLH4B5GZG86h0okwcuDRxLT3KxD9Hwe6HqFO/rT4pWc4fU6XlH8yRLr0iULc86kA11jxEMCpjS
bnBS7MTyAVkvZbT+j/C+AGI28zzV02MaxmGznB5E0Hg4PTOO2Vo8wrJxFRfVfdFqw6I9JP/UlsVw
S8TklU+I0Ey8fDHf21HpYSqwQMbeJVZ+miRACY4YJLo9BouyCzzWwuPf7OZpVhEsQrc1CduJDVQp
wmX/7dbR1B3n+OVRLf8S0osSR7rqBbiqZFpdAPyDZAqQTmz9gozGN2uyCII/bUQkPUt/DFYI/Caa
OORk7c3l/nvacId+sy8ZS7KmvOQcuvxaHDeQtj+XFocws83tluNZ5KGcJrjfKX1e9AshSCViv3f8
1TqXwPr1rWVtQZ6NNVCbnxYNzfFg/Qh3Er2jMshFBmX2Ab2GFvoBcWG6D+pFsX5vZS25PSqb67VV
P9RBEpC22iN1jXCSv1UA1oQgMxNakOJ02jF3355wjpeU4oeRmM4/wGTeswna3MKACWJr2jAg5wmd
G9eXBpb/cKr/yrkpfRpmu6084Rt5LmXekRBDEyOF7ItNjShbeYf83e2pexuoyA6sY6dRSp8HlFsU
YG6yB3eRAi5uhf2pEN0VId3s8IrfCoNLjZyjGv5sneVlVk9P1FdMJTdcAwe2OSLHrr37HU0btoAY
Nc+am2r4NmTqq9XYMA9mIt9g/EekVqAyV/xlYa5rwvSyk0+Ru52/qmnlqBvFSFOLJXdBAzA4Jj78
Pm89iPr62QYsCMGZrxTTX5JPAZnk6ohNJVvBkKm8c9doALfzpq/ez2iqXdgsA/FPWDnuq1d8HOlH
+pTz+JgY1V6F4asP3JC2Rz+/iecYJ2i5IZxyVUv+yoslgfF282GsKyw1TQVx2OLUfq7sgTBX+AhH
jGeVEp4DPrWXs1M23Bk7W3UYB62/Ps4kbVvaqG94JTq39eVUDlL9kF327wRqsNCIMqg3XoFYameC
HU1nPWhXv7YVs1VlRcHUSYenU6nBy4FUCpoGHQs3BcfWjD+qJ/iG1vqiIU3xnjrXYIbKe1nDx1lp
M5ky0LJ/kelEFOESsADAz6fPGHbONRqoRJB5UsqV1PFcDzhwxVUrjTr6BEkvMoQ3FcFnrPLkYSGD
qbpkcfVJZbhWCRs1MoJ7lg6PSHKVyEyRXbx9Be2o024orkgfhe0TBm4XJslDDEUTAHTfjfZUWUy9
HBbza9T98wkWRR+jSoUQS5ZxfrrqUSDxmx3MsokWOlj1SyKwH8nom7EVvFwF/z2BqaKpBziKqA2F
yOh+0s1jY4KSe6WTD4zsSu1StgoR3WtLw0jbrqFpUJ20xGnxDKPILyHCFAWlmiUfRRLofMIAiu6p
bq/OdENCoqqeRlX88ucpMfXP/V/Bw//LpbWoAWxlzAt4AYWYx1mK/F4agwYOVy3hs/b5b0mk6kM0
9FkjKQPMsa6Zse7o6/d0jL/R3yaYALCK7H2rGSv5o7LHaPtr4LQqqp/2e2UvstkYgrjmCse5TMXQ
J3FZcY22doWt+csoieE5tQR2d4qxsWQx/f6S1gstSYgGWJ1d9uMeKjG22DhQMAFmcL8B2P3KzIQt
IpsncNhffAIiwTI+1eHvXPxaP1/rlGsRgTH+xVm0GjN75h0PfCSPd9lPzmOlHYxHWtDuTEfZPYIc
g+SARJtDivBKLMLKP+oJTBydQpXPaEFwZqDHjeD7VMxFz0YylGwzohe1CntDAhd0jbHhV99PwNmA
dvRHsG1ZtvKx+GsFbogAiBCFA58vKZ5NiIs5W8HM2xS49W107FxlFpQlrn7iZ85Fi2TwY5CbSM6T
50dBpXctlsPu/1Kgt2dav+30rIETy57sfv4+NRk9cOWR2Yh2KvIV1nlhfFqJTMzRpltjChskVi0Z
LjWgPgJc0093Ma4TsrXFBpbRl4J77l71x+pdQylTTbYY+lCzjEAQnQUdTq+sQFnbejr5gcM8iQpj
//e50wGF7WEAw8EzAtR9ZLklQMfLYG9D/evhoDq0gEdG6qr6IvhhaL101X9Xz+2kcMpncvJjX6Ki
cFCMWFcmUP7+egzyE/f7IGButtasEN9Z2nlzJQYucwjsR+MWxAi/SzwUetyhEAZxAI1S7jumJY8q
6GdNNhB8SjkCEUfkNEArbXF81cOW3TmrzxKjW2VEDq7vjDU/raTtYgHHIs2Yi2uMDG+XreA7rZQv
/i7WmsSWSVtjj5OxmpChUpQoDBaAeTXSPfl8pNCP+TygPTyxXvvdciI1+mqRpspmxYJ/30lO5IMj
t/Wuk4kWQwts5Q9MISgJry9JcV8dTnhi86XHG9QMZd6pemmCk88tZVb8QyNiee+baAAkv/y/ftuH
Bp2Ia2hS9eHGO25FDAnX4NC4UhL+Rbre+LRdP09tHgIXZzpXAm8tQ4azYWRKcn8mWJzaMzrM8SI+
6DkEd+s7Ycz+y48/X+ikF+kCJOmdUkP2YvBbqZTPXHwp0ii7Z6tGtoSifRUdLANhSyudaAWHIdut
CHgbPXpkGDPaY+FrCPGbtLhZjUUdb5enLrRNU4MuQ/8td2VIkDXQRMnZh/nVrGUCy2G/QM9vRVir
W1x/6E8ZlMVdRpD0mXJ7EueiqoIKoW0vFEkK4z89GlE0E00ef8RqcTnRlow1LMpmQlZpfyF6JSi9
vuvN8hhHYMEPc0JKPYY7Eni5SZ1eHvMKpRbqQVh12DZeM+GuPprhuFfkHTfLKCBNCNv9m2ZIGc0Z
UPyRrBR8pT4j2xeBBlgQdaoGmCeJiwLTBGoRDP68JrOTMsj2xOdg4g35EY8bh9zZGNNueh0ivP4H
ekMjrBZZmTRtjCl8pKxt+qcRNGDXPFL1mgFYvdn5WZsqgyAhwHr8W7mwYU5PQrqDmJMZy4PaqRG7
kmXitac7SEpMifD6lg3xbjFC9X0VnV9X+A1XxMa7R7SrQO6F+g3ygVzBKspLf9djcJLYcgM4BQEE
eqXrqaBzo37JVpKKl2JYCH06HpONSz3HeFBsdX3jQZ2aheCTtKM14sFe/xv6J326xhz+US0otCNs
OvIXsUGV46e9pfFyHODkYxO9pl7+16iMIz2MVtc9wpU64kwNIdvvRieQAoTgZcU4MTqLz15VbAYW
8slL+CpweKfu+T6Jb/nou4+nK+fPwXVExzfGKeV0iuRSfXdyjMypOz4tXgxkzWGEHRgq8+ibpGtL
IFwEoMMkIHG7dPZZfLgH83j0V09v0JzZu+brsuPiWgguYiTCfUFQWzAt/A1SrqPi/W5G9JrgLKOy
MYIkgfqmqfUc3FW7/UbLLPfHmqVmBVEqB95k/idDx8o5/Hr/HTGlF6fR8ykalQ8LA7oDi6xlBph0
qb7LbLsbae9a9aV7Ev+ywESRtqKpT5X6EKKmpNIZAuleKZCj0wxrghz/TdRJyKiBPEXbHnQRqFDI
btgXNHPIwgxTFJeJ+54jk/PY6Tuwhh7wRIprb4/4+/FCKCR7JPhYTAR/I0LCGKL95/Qxoys36cqC
Gxyd+IBw+8cqjCzQ4bwyDYK3IQjDuTnWEQ1TXBgs4Z0bZR3bDw5uvdwkl6bImWDc7P0V+Yg/pnYH
Pk0bCS2HTUdfd06uf0pFNhfz4BQxE8wEXZeeMJVXGV0W4UCd0DOJSGoWZNQ2Hj7uEtuQ+SMTlywA
7f4WQj+dzbiwHP8cpiXOp3H1mEvhG6sfIJoqjaw1EnkF20GDzl39uiF+sI5xBkhKPBnzYWQ51yyn
FzFSSwQb6pkGVjZ+fm0J9LCDsxe9++1FcQ6E3uJO2/qLiLieMFkJQemSrl6JilPJPATbFV+R4nk1
22J0AK7zBMXtI42VroeZmtrpNqxTaRCHqOGdyPe8G/UoDSBoA2gTea4zjAGF4J0VSBnPbqU4ipN4
lki1jTwHCQXyQ4CakCGCby5hG2jkSjK0svyf8hYRhPwX0WAfHLRCVCoc1q3L35lz67KjC9VXkVEP
EQ3i+eDHDMhdv5HPl/F/jsECXWKrFKkxhf1NaSddvNjkOShjEhIUXZrpm1dptCpJVB9zcAMD+yYs
O/yIKVjfH7/Cp9uyOl2gHBs7w6tOJm2RqkOH2gia79vIS0r3Av0j56kjovGgDa1n6pGuRVDTQxJE
lmUDg2qSxx0EUQZVCBzfjp7VJEijVFvCswCzHBr+5SGD1fMCmut8AdQBwmJvxLKDXTV5xhK59JQG
yYDa13W3fJCARpCb/m1qsj9m3whEEdgSvx0XeO05QeHDx38Iea+kUW0797vSWhFHccjP7HumlQdZ
oQ/4lVAGBDFJNS5G7wvda0YydyLnxGTVD/+zyIDvizXVjBhyhtPQ8bNthvWGwjzArRFYzHVCkT1S
qSLJmw4tp+xL6XBfmTRRQr2cs5hOXRSQzkXu1Fv2Ble5tYe9Tq99uEzb8X8YuAenLSUU9p703/EP
G4JqV3cxS3UZ7HYwOCJ+5kzmlUBLS2NAuhJBi3JI9ghU6aA9ta76aWgmBphvFmT9RwzWwihlxS+F
Zg5Is/0DdNBhipOy3nEDFfclKeJ8z8nfHyQMOHqxahNawSEJFiqJHBKpAqEJJg14jeJtqwRNk5CD
9m5zYp5MPxriXMrGdf4wmvcWIhh5rf8UAlqT4ZzGfgSNwL5kuKA27JvwC2CgeCrgmdOMpOEWsZNW
knWHFjtH74AwbssCkK1TmDpTxu3rd/wHZezlRfjP3Nxmk50aZqVFRWo+CIk3C8d5GYlbi8JhFO6v
hWQGIK1E+jhMO0PQiv+sJYPt4JghM8G2idtPJ3cB238dfrkMJHp0Ilb9GqvOu1/ID4EUtYiKcO7i
RHy7l3WihvhUhAuuAdohIQYJU/t5O+z7BKYpXFpADTt9pjyokU+RTHBjxPeSZGRZ+0xpx1/cwwuc
bzy1OzOWdDa78NAe/5OhouIwGq/QAg/ROUCw2Cl1DsYybTB3h6kR9VV9wBguBWEVQW0BIk9CYEz0
i/gGTr13IsCxqljuSfX8q9GScN9fxIHrfOAMMU5CqwxuY/hG7frQdov2w0da9qs9hc3kc2b+ZS05
f7HTDVxe3Gx4y9BAnF5z0SAL/XqOToSiDWJkUM/LOJ+8gRTVeghL4NQRa/eDAQnDZbqqFK/fWdNL
Ebbfm0cf4DqMOwqKThG3BtaEzcEblv4GSfna8E8al0lIgTe2l0YGUC93NV4MeHlDD120/BN/mXha
HKAEUqrMCEfWk4BEA99jCbInRt2vv9NQJbt8CePoO4kXksB7NnicyMsJLrKE0qxL/vWafJzfU0wz
0MRnwx8hx0Nxes5GrJuhCpklyp35AjnCbpK1LP78rWwB9Qyv7l73ZUG44dvNhMHazmYl2hOMSArj
inWoUn/Q0zMNELCyTaUC9TK0smgAqW2w/6QeOOlI9EKS5dHvIVoCwkTDWvMDvhqgfeQBE3jUAgUk
P0BBQPL/7Z0nBhvV3Aeu6lPx053umcCMdzEPYmzAVLXu5WGCjDZn/37zcVqdD8XsZClm9qNO7dGQ
x7Wncv/xKiNyfp/K9kXmeqNHm6dMmcmX71yksOXV0ewKmYjmH7paWd56vctVCzioCaHvSK/bNsv4
sFjDPoB4xZjO2/X1zYChCMawqDfo8htrF8k5YU6G58D4e9vqXxWh4+Oyeu5YUQxVn2dzzHB19jsI
AlnHrdWmfBw+hFJweZqqst5KIUFnDmtz/BIKHOj/D8R53vXAPQQqinJ1iVTyqp19RHl18CLlmeRu
T9D+oAN7Qy9PbRlxElGefMKm701sISCp0Gs1h4kIKdqEKCsZmdFrCkj5xQgkgnn/zVe1OKr15pdD
MvTfMMiQqwR5fYQHrZKdWL7omiO/ZJY4mR900p2sCMfG0z1azB9SmfDcQrPo3Gf9PkNupGfLeyoj
6dWCnONeFMxHE7C3InySrZQyJFyiVTbKkA4VuI7q8yIByy0l3ryGk6TEtpV0YnICO+y7BoHVYTQi
Vh8D4PElJ0aqqeNg81+kBeZ6VPy/VUdoCN1bw5WtIcgRK6ox/p0w75x5i7bULEuoKcuyczfXosOf
eWnnYuR5RR0+oHjvL4XfOGG19Tu+jd7hxpNv+F54DBMMDNabA2fXzrBQs+A7HsbHk+UzkBWjC+jm
vJkPmN2VpfO607PSkgwKdMSD7xH3HJAzGTfXx3TYx4GUcKIZGuZeQK/sNA8nfGGvraL1vCNDNg6i
R1Q0ovtOYA3HakKSS9S4x+ai9Goxkz1YJ/N1viSZVHfxKKJH1AGQVniwgT0gY01EaRs3X21IYzO8
Dhlq3ABfMaI/H+z1QRgBZwn/JXTPyB7/guvzrcXs94IUatkK8du3ARJALhnPpZBWGjp6mn03nmRN
sdv+J7zjCZv467QwYnLZg+YFIp1lE7mWpBrtuNT9NiT3RCsI2O1zDK5r34+jyYLUPzCq7O/wEN+c
sKLxBH8Mrv+wUtEWQvk7Zs99dvt0VcFgYr/ZkiNMYMG0NWwuqmaZE98fwUG37OrfswWM8Wqo31US
z2LdJSH95f6SApEp4uMGZQskrHuDypLx4wD0ZJAcSln5kkkn5JNR1S2LJ+Nidd7jDmzeoGRqvZqB
5Ff2ST0Qa0lBkZ9CzVsjBlwil8XDuft4e4voIKlKMo1yFx3Zi5NuQjCvxzSLngbva31FjjjAiyHH
sFd6nydvL/agR4gLTUgL5p+8yi24wMTXxDq+nMHSb5ZYGEtU0mJhSvBQ8fSSn6jpCUA/TZnr9XuK
4qjc4b8jLqRaUroRyH7e5Cu/gxKGCNWM3nC4+Ys4nC8/NPxNqai/5A5NdHZofn5bOLdno7MhZa3s
t/4X3ufTkMRgF4ZuxqB4gAcxk7N3iRIfvILJAvtV0Nzb5wDe6AkfWMZURSZJg7ugczbqU4gG0S3c
UD+953M2TWzR+GuJYatqaECDlrKQGgNDFQ45Pp0aDobCUl5n1DwvRoEzDn6PGR4mKrWC220Tg6bo
rvDEKN1kZ7Pl3COdjpRvHykYz9OsAry3o3Nrz4C4gxiRltbhehvT7ZaWlR57iWVdwYysh6ka0GTl
r4hL1IcNCpp8dDIXNHms8flMeVfmkyQCQCkwuEDoAlp1ZszVH7P7jckOy4sinIKCptWWt2SjtP1d
G82N+NoAOIO2lg7Bn1mGydpF/xMys6sCLWwTcMDa8RP+PQtIhMSSg0iK/32Ctla51n6AcC2aGm1e
n4e/QK2FinSRsUre2F4ByE14c8RAqaV6XAd/d06/A8m53TtAa4Yrct+25A9qqQjWkrX0/v3eOetY
gzCKI0D0QXv5e5U/wl9/ReP6BId17UAKDaY5xGImVDKwsmKMoRGJ3S2xmJcAP3RTiKIuXYmBljpI
K203qwGQDyT5Gw+QHjerCXvmUVsiNjuaqxnB+OenBn9A2BHkmV7xzFb6zwSpZeDwCix95TFiywa9
xSylelh/a3iYOpXCXWBschB+32AxJfbDVk+8yAfnd+ZJdc3Duz8K9tCkQYYIG5rQ9ZcJvHHFVFaQ
GnfFK/GTpT1NHxFZ39hgmPYvippYgQJmhhxCME+17FklW3DSqqdds0Qe+n+NwMGgJWhbanGXRhST
u9T8/UrKoKhiFqUjQijqbRB9g6wBleJ6a8ziADRW0GSwPYdl6vrPB9uwoLOcMrLVs/PGZC1BPu42
3+18ff2qawe2vInB1mrzx13dfA4hTwDwzZJsqrFFgAE2R6QtZbpPM2zSI8x5nbMvT9+1mqNhK9MU
CFYhzuadwC07ap9+K38LqzvWTI3A0N80hYEfaIO6S14GAG2w8SiPNGBEUcpdCLlwPkAwsCv6PjBY
n2/2js7VfHFaH8pyhuQBhAxWG5nJILoRoqqJ8dUDDfo/zytyO7o7cE857JjhPvQOsKetO2pfh9vo
AYgj7jfHfthzcbQaqUVzaw9Huu91SRaEtV7X4nlqUQaZ2VcEhyIx/jySDiuw/HFsZvbi9TyygJ5Z
t9WjBkTJm8iWPzXHlwFV3OaFIggq3zLcWRzDlPjCb+dAuFJ/RmeSmxhcZRVElN2QUokR6lVncgkp
LYMjlt+kyRXbiiHX6ehUzsXloaOBx0iGLJHOHu4dO4yiEvyMTjvr5+Co2wcNCNP5xOPkysvn5ojS
ru0vxcv32e4JtWTDj3kj87fY5wwUhjT1ZQQiQA8xU8dDHDdmvDsDh2cOUpp1olmja85WwKx7RhDY
JYMnSx4hzR/aCCzRc6VpoTdPQ2sao+ol+gjlCPpiiemwAp9Uy9LygImjP0QfBXeuuILfDIzluy4n
oP2XutTgtd0v5W3UPTdK/zVh3oPrvKbJX1+LFs7FsAL5BBZ1Gob4WSVoXpCKIw+6c0CMuMyauJhO
n7sXz5V1AkMN3JLxGG7zHapDPQpnU0KzuPyYI9h50PriwfQTg7ZNIh9RlPXyYmduTRCC/IdolrM2
93O/oPvWNBXdiDQLxfJ3X/90ZQvrni2wzd5Wxo9h3nCsmGrxs+mAGRBbr5J2V/RwlYxqNs8fAKPX
0PAKrvPdyVqwsEaN7r/cZD+wiuQuXy8v4M9qJDNV0hS4EhPKTZ7FOwVllxoprfOsxpLPSRyckrwV
yQAYi2fqp63sCaOU6hSYMr5mRaakCSxSC48fqzPk2R+ooRFKIvs2fmB01OK07RvHo2T8ccZBI/bO
1HZ51Iau0RwDCjVKgM9qKBPoJEc7tkwUJuAYmjNloR/qoSLs5CxDlSgj0CDAoaKxAfaXCbQHKA1V
JzbCkC5DOUsEZtELp2UoKQ8LeM+TZVKfxUYKu9cGDz29TSQoeGjs3F1W+4Kn1c5+BFoBsRc/bfLO
9o7SXf3XdK8SxrCzhYb7zWRGUQYATdtL50SECelxo4HpUmcRX1mFTigvmMH7vt0NoXyz1GLZjuGh
Ydn2uJ61LnReaQ2PAmy4dxoLjQwIaJtfyKeTe81IzQhtpz/5U3+KrtmLdmElt7+xWZGCj06Lh6Kf
h55rvLdkoQ3a0M8oqOfwKGwenWsvsKHw5NFRfWkHBvPb720yhL1qIe0qEhfzCittxDxZaG+a9UQG
cCWAtaFIeQH3VX18YNE/ZwfWHeC3nuCHNWnqRW78Ce9ftOBTikRMReccY1vw2OedfMiKLekLQa2U
9LFhvX5njCU34xcIY8RK3oXAObfdQFCtB+NzrZiiRIPge6fIers6rEH3b1IUif0d9mUM8tgf5Ax5
/6xJk3gt/aUzFHH6CdLwYL+JFYb/hYdhINKOYtYiVJnmx38d1mv+9pIgDuNhXYT66lsMKeDwLkwM
ZqcjKmhfocEfSsC99MobVkyCUAiZuFfdROe8YOrQtmxW+vbh0qF7omk1Yk/OPkIz2xjm43FbEFMO
xd+xE6/YnERprSmGUcHUSIb0dGEyIxHusuEGuXkXwU9O+10JgpVJ/zTMwO7pn3FeOx1ncq+Mw/hh
yH2NptEsz2aZo+0M8cgbDJHidNgIT62uXUkDf6Nzndm9e1pgZmcuWTgMPkyb8ZXNVtvoewwPQjfQ
kygHawQIGCh7aQp7JTuoqUNogni7PyZNrtaTUQUpelIZUG4nWo9Efs7LC+h0KKGb+JGD/xfnUPVP
LMgc8+Zr2vraXSi8KgPwRk5/vMEb9sgNLVbhbv/fGkdPfYOYHpCg89fHNZ1rnE5jzquV8XTRaB5F
5IrNrGADArCMA51UK+OHG4Qvt3gHmYEMv+rihBNCZJItryNl23og2av8yzYx7blmxVmtMCyXPf7R
2eHuRBvZRnNlduAzgn/UaVpME8vde1vD8weL9xI1hl2IANEM6qqdbNNLZuqfs27FdrtQlVif/voD
YcavlFXFluHsJqzxHm2NYfbtwS/EbOGEFKAkWfqC5IR+kIS2jnveVzwTN7JXWgclrSGc1t3lwnH4
NRG0FRvI6Ax5J1Efxk5SJ4ytlXv0O8xmBRA6o9dZdwDNV/uNIqWp+qOsFcUJMgVxYHABG45IknFY
kZSYIWTcSfiOKfbZbZCm+UKi/UnnM9NrC4iiSl8jphSdGobqqf5LlvaoObK2nJW+hfGaZKK//a/6
G1AARX31oZwrasFGB1o6D2lQzyvxUA2ZA3/0fYxnJq5B77lyEXjIuox1SfbbmBZhCfWQqJ5mjZx6
Y60NIoHPb54DPMEys7IrRKXqxf8Wh4523z0FMQYUHyUgDT1j+rL+yroJkyGurACMJLidSYYnh25h
t14L7qy05gBQtlIfv2H69FiMGAYtXrWK4wL3sMM3OlwsgyAUhUMuF9cc/5yJT126wDlKAQUKZz32
KKaexWHUcmjJfAr7Odk4QLt9NZ12hT4tkTNLOf7Y+442O6ff+TEdBt4qg8eJhUG80qXbKHWYmm2B
uQVvHtmZtr4Ng+BsQdi3Jd2HJADPG5do2B7KO2rySoVh4eW0p/SR/iI3V0l9KwLMpvWxwJYhVh2D
QP3uuvboG7d0K9mFn4nRF1BpvtI9+IDclGKyGa3AZ8v9muc28YOjVG3Y1ZzA7pxnfuYncKRpjBgD
O0uaRnsGlY1TcRfwggzUSOhMyMbllGt/1VpZTUnXdtV0JOH045ZRlzOTJV6hwOYcYma/7jLoyGuv
bTpKtQqEswfoLqfUxwwfF4nl3S7+1Q+RS7N2gMbwTvO+Iw0w+LPFwAksrxyda9xFxVqR3+eai7cD
Hl7JYLxXZxxE0Gvz0ciw/V8D5lAvmti0QxVl0aZx+zV29YPQlnN1Ea/i0vU/1p9ac+0+8ROXleea
kC5ElyIN7X1QYn448fxuTqrjUm6V4jVSm1tqANBhz4/megJKdhQe2Mx5tS+7AjPFUhJcI1DFmDC2
XjfH3WXpnz1gO2Vi5qnkGNbupR6RoIQ4G20k2w51dytIf7HapmwcNZiXdSa2824UlshoJyY51gxF
rE9XR1QGYdHcN1qGFwNrwr+3NLSTjuhw12xiRTq12Pnl3YXxG+nnFlixPfN+EII+MgX+QAM9f2kV
2U4t+uHOlo070VurpjoU74OtbMfgJ9xo5EnWjlicFBipa8B+mw1I7ywIV9SdDSDQnkb4Z1FUN86Q
fK+Uop43DLYLjsBBTO3biKU61R3/P+sHgiXlPaArN5dF6kDVJA6UYopAbkBwNdgKqKNRgcqax3RM
QdKAzBQ/7I0+A+7BSJP5DJxpHmJfJRvdPsxv+gaUfDeqHsgydd/+A5Se3XcO+xk5SLfXtWbB0q6l
zhzHL08CfeD1RvqNJgU+2iuJg4NkNHf3syefaV/5k+UzlwsdR5fcc4wtGnOP8Crpz9U6DuM0WUhQ
sTINXuQSP9Raqb2h0k8B070LPGfbEGYWevwNGUV0bd64PKOMQ4qvbxadiUxrP0FnJqvjyTi86ybi
IGnMxQiT/Arns5VN6WN6Xdt+4Xm47bmu9oGESidt+dhQXC6gfm4+mRtDT7PVMd8FruL/j6wLdrqD
rX5uiEpjIurYv4ZYLnlBySnvb923AOg5raRKIdktVAWWtmQp6U/ovD9FafkV77UzsMxGytKfiRxB
FNJKD0KBJH3djsZpP7WAOlJsVsWKew7BBcwdgrOS3sTOkSIM0kXutZabw0OrT1EwONhcLEzG+I/j
eSmqDdfyXh/8MIM0ySu2n3n9Y7whFZ32bcc7sGa/FRFvnI/cLk/jJ/bHJUBRTTRXYhqiWQEdANJg
1ujGv3pnTbeO/XFkvJn1MlEmMYvu+IyYRR4iuqnmZb5pXepfqnHrCL9QHW2IZJPVzPBzRJ0xPkqn
0FNdq1ZfAFoAuHRCkcPNiQrLsOcmBtPAwZK4xDlYpUbmvtDYNT5/R2tP5O3JVOvcceIJiMW60clb
XkIZ7ltstWx8DbwSU5lnuDyU4awSwNODQD6zffnymFcUoCCop49mVsxIiO4QF+yle5m2KFqP9qqs
EQxg/vTo0hapEvXs+iKLs7V2k5kItfVwZCF7eIhQorzlI0IJsWYbfsMPNI4bcO+6K6moJARdBfpt
bWBhTVET6YKqyeg1tzib7XD3WKmNcTEX0og3BTiqnQR1hRiMIxJVmSjqCQ1q9SbC2EYaifar/7YD
simwfw7wFPIdJlPhqTk2SuNYRp5I6qsDHdK3iVzB9gfJ6o0PDl/nvkdWjijMllj/yMY1LY3h2Z8E
XZwaJGuJnI6rw/5kb+m19JJcGkhxGJ0STiXpK/X56Y9U4yTsBhIhbnJGYykxjKEsUImhUn08Po97
74jOMzU8TJfX1/LLCFO+LGboRhCvhEA4I6KyCMl7ySHvFbD8rg8f5wyJT+RuGTz5emQkjbCxfW5V
go5M0gK5nyBX0f4xrXglD96rOaU+f+wEi4RrBS6lhBi+gNtvQAzAOvR0x6y4QkoJofm1gOBpPrlV
Biwi15GfPtOma1Wt04H5y1nl4LPAalnKs4x8iMpoU20M88+KgdCtI4kdY++HanNkvo5BIcC482+P
OmI1BiKLrappWCTsX89d9htl73Z64gVltgp3yCrJsNWPYIhKy2N1VNXuVXiYNCw9L7AKhgyGWp2I
SbQcOGgi2m3btqyap/yl7F6cfIWmEKpGGgqVAQ1V0TBxxcmh6aafOSXJ17khMeSaFpvAMWpECHUE
pax9QOcnJ7WfyFx4HvDpDQiw0tni7WL8I5MNu4Yc1PanplBFlkGIsVwV4BVnFfFuwDHhtcMqAMnT
Amta02R/v66CYOxGjL+9bB4zdcciVr1FV5t6yTo8rBPDgEbbF5RTJ77bXXktnxicyysVZuP568hu
1VDZD4JERi2ues4vewBpJMhfdWtpdOzVxST8nc2jBKjS+afrb5DyRdcCIyV56TPd5efVhOQFqn3H
x7Oyvnm+tLgwM5SyHn4lWOAzHFPs1JWodvh/MrnxetXJ29rEewZoh7EM6m3W1cA+a8kojuBVgi0a
AkrWI+VjCSQ9ldBGK58a+orcURrmysRrexzRlubkfzS0VyoK5mrjdMwJJDYUSOY937zPpLCtLNzu
bQfWzdH2bmJ/q9lRxCA6zdpFU2JYhT2+kcVIim2aKvMa0g9FndLoG+RtLlifAa2ZrV7ZPoPEW/lQ
W0xkgoifij5h9BX7ZnADjIgxVtM8K8xGim+613Wt3BB+HScL0Mg95abuGQxozQ2Wkq8CaYFDGr77
0gg28zFeWQehys1ZDL90xiQ9EVqNG7Yqd/WIA0YiSSDd3PAtHWLKr0+zA36uzqiZBH1hWZaG7Q4/
/FXi4nMgtQtTKYlGdNGHqzCY/hZ8cjcvXHgHNZoi0LlZPmcycwRnCqh8rPIRNgRjPBHdQIAGFbb1
DjAXDzSQ9/f3U8CqzSfZc5i0kWlTE926s77812yAE102QgXDoo74mFK5Y3rI6OUf3UtYIvMt28EZ
MWjwDxyuFGZXGjKEVYKi4sPzvNFdBNprMmEepNXqE59+bbErhvKzTnXOz29FMO8urtPnXqAOfeca
zT19VE9vx2lIv0CkTBtpi1m2pLwrm+LFTgDBs/jH1RTELtXCrlTJd2NB15LdvAtTzyTA+vsYDJu9
Oj/vsB8XG46Onjqq+yVBCeMfagXfUZspQaIm95i5/aC4zBECu3GXC3bo6mGQZ+IHt16wls2f4U4r
kwyzfJlAtYpdi+X6cm+rcyrc4qniM1qozmrtfdhTBkNWi4yhBqSAONX9crVuhFBBdCtSq2MhC5y1
ssiVv32u/lgHPhQ3t5pWKT195Waxj4ipIR9DO1hkpwaGMY+kXFU9yctSPrHNLphYYZwKy0GvLY0s
fUYLoIYOnklFwPaTNYGnSk0KaD/4d5Xvry3GX+HDXoBlmkmD7yLcgApmzJIe9gxQ3ntjAgjL9kyA
stE/fWjjoW+AE70aq89NLb9Zp/GJm5j6Su0THo9+XdqLTbu2zUrQAFQWI+TzbGNh/P5ltnrnk1O7
3ayClaZ9rlKP32y4UT6LQYSFG7XkPyntdV1j7wzIA6cPvvjxLYVrkyHK9c6++i/fnOJFNmE+AHlZ
1Aq/ibi7Img3ynNVcVOWPKlQWJmnNvXwtm8h5l5Kv1I1CvEoyMOLytM3YVwIp1S/vLxuN182GGO2
4i4qXprgUZ0Qw2bI6gIrhkqMF47A5FejJ5D8pOv+3sUO0G9LVqCj5I6HbqqtTGm7mKkr1LomQRbu
hRvdEWqBCcAjmW1i9fOybgkApd4kSLuIjVeJXDuL3g7BHqu98aq2KJu4JGpApdL3VM774RfsCU83
FuoIlv3TPOS0lHIY6zTIVJungO7lmsd+691ycNijyK7tp4ImS0hJiLGxv7FIFaVcMKbmNdRVsUnL
+6vBq6MltjPo6/C2EloIxLWN9RQaviww/X+TwNTYtd200/kq7hhSfmr5R5IduJpByPFX6gfHPT1q
vR2ZNFq5wh7FXhKFiusU17NYicpRM0j3Ct1cYUqFPobujZExyKM80aIQ9E17cfCEbtglX99RAt4b
F8tUNw/Uzx0e9dmRKkD9YU3RTojO57ouOc4uvz3sjwb7v+ArwmdACtyJoxT0XK4bQi5mDIvRWCYL
Jsa/AxuRCmCicKQbav823mpPnwDDA0bzT6O0le6/dCQUOziwSwjbIh8/b6W5+3JUNoIQJjF/l76T
puC2cgIu0yhbr8nHc2vzWO2srTBSDwdGLnS1R5fGb130THbs/1E3Y1zqrUz5/SDm3IV8+pmVWjiy
1LY4196MMMGniJZp8L6eQyxK/inU13dJLuVK4EgEuFJJkjrTpK0Xfay0HvL2mcFLr5NtBJRJJHDU
tJNylg2wUzYB0gp5ICFF+ALwcSnyNPMwUjETRvNfm4KHGLcAR/ikmf3epLP3bUUG07WlGgALEpJh
pUo+l+2sy5jt3wfTxerSNpHiDBkU14BcTFv8yDCSsf2wQvSkjJwkp6w1cZnn+6Q9NXpxPze/uK15
6vsuPNbDOEyc3Y1i9OPk0OtaWPgRuCnsIdNCP4qlf4a5ova05M+8uXk9DuVQEU6HBmR8bPAgYIxl
x4idjoH7PNKeyZd2b/DiUIjqhISTDRR7fWZIOARCa51RWQ0UQucs1fFZfhbBC9v9Vu7ZN6sWqtDH
GNnnN8umfodndTJBwbr+KqryKKeeAS/LxM1bjkPoci8ZLW9apT6+dqBoLw+Tjr65llELGG8X/DAP
H09io256JQ5eVEvcmSHQxaJOMsHr5VSLxT8DRGyORdbWkq5zsWsDhKvJMePadFXftDzoWWkVpXX3
vXjxMAFm6IKXx97C+Yq97YrElGBOxGgiNZql4x9BgsBleYkqCtJNDUeU9O3Ewt4NCisoWY9K4TjL
2+Ti3iwBr4v+9reDjIaQnxMCev2lUr0W0gEppzsi/GDBijUI8ziNBMVRNaPn9EZYkhVKfwpsniYq
MDVq4JCFituXQYQwrxx4u4aOqkKFf9MicwLtGRJUBF2Vu9rI4nwNj0RbnpvfdhtmFl8t1FQsz5vB
pe9BBEx/wdBroNOfLqyt8fzER1ZplIL03F+8w8PURZzjfmJml3xKR4upSkOQCZX7adc54+m/3cni
hQpqHGL7IRQWHbFxndMOstkpNImNlNZ4Mwc49pfAjhlPZ3U+XDNUvnt/oDcOMrD34zl7xFIQtIKJ
piGiqWTy1jqkbmYkU2huWuQcquCChmoktrjsQzgj6LPUeIxKIZhhOnecrV98BjtGZOMUrDKBcWeN
WJmjdrQ60ZEntKb3R+xgzXslS33svtLSGhoR+Vmcx+icWkEG/JuuIRiMPOkKH2ui53OXMwLVr1kU
HJExLFU5Y1uD/S5vledhXu102W6vkpypNYLhQKQ1RVFT5VxAmedD3owRw1edG+cJBjnjMDBWSdpm
1OrodR/wKEFCd98caoAhbRkRfFyOYQEkNxYWR298hU52aheWcQ1jbNpAk7b7WtX0acQG/H1MH3T1
IQyPDN47EqM44PFfSO+JWFFAsdYwesNBR+rhKecyKZlycqGS468LqWobljFw3yCLV/9xan4ItV3a
ezUCCmeLFcPLkjNj5Q+2fdj9o18oVMzDUhsfmsP888+cYhj4aIEofj/GUVeVmAuUdqLqI2yBG8H1
CM03Evqxu2e/RLrKMGRu50aeMCKhtL4Apoh0wdulJoKQmYHewwoLiCRwkN/0mDNJoU+lqEueFrZi
JlZu+P9EkG0E1+3YaKgYDBDKa0EWRrXoEmmZANBeluoKi/jduSvlDGNFP6jLRfDKUSLosFEb6fdU
tRck9CQ46xjm15eRSHskHeXkU7gu/BhV7BroHZ8g2Rge9YKcgCy+j8dE05IrZijD6MUMJkYqsELU
Cq/nrvCSq13SJfii9WhmMBhV7usOJ9v7LPyGt80OLv1HBh0b1noac14JSM7dvyYdGGv8X0j9fXWF
lbb5qs+6ZuSnLTQnODfRPTYkdeXhPMHRiYF6CL2o7RRO9ps54mmROXsQImDQHJb4qfPG7S4j/P3x
MHBmzFwdEvxvgRcEOLU7vExH7ojoCrar0bGmywt0R+5p6YO/+WD2XfX1ZooeflEBeX57s0XZIVOY
0IfdOUMUmdJ/4hcIMqDWDqeHSms2NquCjQIoVv/t+Qfozv3grlLwe/fjHNxgtdut1ev3GEMYJLKF
l/kUy1Iq5b95XfhdrubGUcrPhroCbweW1On/RB56DaYK5D2Ix2VhrrS0M+p+7tJhzgnHrjlUTZTa
EKH909TUEqGxeZX7HyAU70ZDCpfIdFeqd+cljj48rYakcbgZ7+74cvwvGQlnUlkaIW2Q7yXHVZBA
Uh+fJwETpu0Weoc4OzgZM6HPDN80Va66ZVm6S2zEVpqXVWM6xDQO549BwEYk99zf1RrNVhnWM1QA
sMFWZYSZAYl640CUhmQoNY/1Wew/8a/w6vvTRaO8183fohdQR1iDdhG1GnF0sJl8xu8zCb113jcq
9frHDuKug5yrcCd/utNDTAzaXQSJJvLraOh91SOIeVdOI06ZN0PzTXJCY8HUtz9jvO8kK+4Th1gU
ll/+RXZLI8I+oPJr+2WOn0ZsaJ+cSL/9a3EdHBoinej4fWBfMLaMXK1afUjnyG45TcKhhX9mR46k
uekl+YNFHfaDi4B0wbbKhM5UHZn2VliX6daa76VvniWDFo/7vyHjh90bfK6REYjT+l6E2a1Bu0B0
p5rZUzEzdaOgJNBGKCN/tu5daRDlPW0aq9lEfY373MQmGFBHYKZLER3zlWjnWDLZU31mvUw06L0x
NiAVwN1CHVfjSyX05tf/y0BMekAt0gG4GtNejXeR7kXE5l/o50VzXQjgR0Ywk/QHUgbtXzc8dseJ
P+OL2HRwSFA7Rb+Ii+nHiNRRvjyeOEJMapK4T4QmVbZG4TVCgXV9k2TKzxpsaBLp5iTBklfIhfFg
kqOYpQKDlq7JO1bY+yf6jdpS94eb3++L5r5EDVpZZvtiJ9hSO5kYwy94w4fG04+4q4uw8IfVX6PJ
8fsX/orDwjii4QbolTudTIOemK/QsUyCqZZri0iIm1PQJU36mplmmYnkbxEwVxoutYcGfZiSAkZx
AdoZ+q7T8qYEy1T2bEFl+kA2Xv5U0pgRH8xDR1o9GKN+xdOrVxQo8pSqAyhCxrtMEJYHenW3Lw+U
bzfZC6gBaPmzK9/NuJlCadXKfWpsuc73M8HyasLychhtvkUkdJrH2I2VnDQ7wBdrLOpHXDg0ihTI
3G/PpIWHuS6AWaVw4VJiTzex4H95mBPzfW3gG47euWpt+dqh+Uf3zg/k94rgAyuUVMfQFwG9wHP+
q/zAZHOkoo0X+wUjFcPo3Bwb6/ylSDC8lEjPTRPYCLY18t1UuQ0g02Ve3QXuwDjBPdarFoG7oe9i
h1Ag6fJdFfkqYF0Ts5htX/urRR8ulT4g5v8bCh7RGrJeUvRSE9u9jUiRXytDAYCYxvF4pFRD7xM7
jOJY5aMnpNKyvKX3+6og2lKoztr9tzGZqlgP4FkOOra3TsVDgcKhyQYS21DqbBTnp6DE263yrPYl
BdK55O8fHg9ntC7p2F+i/Lag0PdLBf8N9IFrOuRbo9P6zLqrqYX5yhavPFF4ywTuP9fgRUNs1lNP
6icWhfd8rvtHAAvTH73+L/s2tLISq7ML2av+c0KulIrquvZe91jLn1kcZ/pBakZYUlNgp6tBXnai
J0U9cCa27ZF2PaJcrDC5A+0w2xO0H4PIgx378LW04Gx8gSstK0bMKwRaBC2J5MvjoOBL2rIBZnFv
/wBv9CInpkOJy6YreWnQ5fT7nmGoTdSK0BINVYLL3+mTBz0MBPWrGXGRYx8vgtnHG6jEeAFEePqG
b6YmkOESQKUQuEZ3lc2HGAQDfLff3canSZHnoQVe6cXtXbzUDUgEdfNq3IFx+bNPhLKSuYlEiClN
gB6RvlD0rCh9frntH46MP4lJA/J4SdcWHMtg66Osk+Wk3eLHfOjjiL+FdgyYbAtB2/+1gYa62EV/
9moDq1GAS4DyTDRx0chp+kJYxYKsQrFR/uEgnvqJnu/CI5P3iKoG7peXS3EXj1HKw67Nkqkl11e6
KZrdogjuCNy4wfILthkVNwbU7Phe35QBvBrJAPHHOgZXoBqFQy2J6YoyBeIoMGITNwTiwE5gQIJX
ScSDdkw7ZQclEE87C2A1KicGHnZz/XdpoIfEXPHh7AVcf297nLfjqHNCodnrFsyBdE8RZhp7GJ2+
G3saZrgeL2tuQ2EDjSSZTQvXnMqXWyhL6P7R2zaXmAzmkHRAxcAZQNt6FiT/RsgcloGyXCWNhAp2
Zv/SlJIaqgPv4BdLQXDF6AO7/vncCVJ5iLRk4iEIgPGlAgNdZoOhnnHNS94cCy5cBrggEnN68R6T
RW7gd7jdi6ABunwA0AvLY575XJWr0P/bO1Z0sPLnLS4zJr02oUGM+sWyV4LUqQFq+ogG/QK3NkiF
tG2PYEC7mx0KfuxNEoRfeWiehUV3Gp9joR+RDAsPC2MFWTNkd+qzpj8Ewyx0Z/pxLNIR0ytiuLTK
R3xM4pn4g6MVHShsAvUnTr0aWsWv/tmpj9u/pMn87nmq17QlvJiazWxuQz+v904x+YzPSUaY7TTP
+bQa0A+jFItwJrkIlVwLjpnHR5z1AxNLRVl2ZUfTgWZ50uzeUOKXfuZtKGqcL6ea19fFwJAZgoAN
zQJ3cSkN0r64XEdBJKQ2b3A2mKn78IgKiKZu8zxw9EnaxSpZSVSAyOJOiYwSpaAYjfgd77UVOhbv
asrwH7g3sJMhrDSY9aesCtTn2oiq9tN+bLvJvTAJjavWmb1eAQ9LM1xE7UnwgCysK2DjekWKwlGk
4gI4uRcsmLiEEvy9I8NxarhIMRhODz1gikfQAxL8ScwwTwrZ0HQoDhtqQR+3mEy669XGEiyJgfxa
ivtcu9f4a1e3hs6YY0G/NwGTQQrMovCxOLERZ4ytJLAetXbEkSxSv5qLW2uqcMTaI56x2GJgcWJK
B1ZuBe7gnkSNE9Lxe8cGCvkPpG38tdcVaXLsp/J72M+l8nwkr0lC4H0oyD8LkQsiDsK2k/Kp9PT/
YqV2VExRLbceHMTND2SGtleMgl3AtcYY3HMHWeu5y0OjPAPpuGUTCz4BVkAd8pH8bAMXbuW8VlHn
0HyrKMwTSDQh4PsHCSKaPszdWMz67ZQF/SjA3FxIrX5AKEV520aDx+JjWIemxY+rm75/Jz9/wk50
NeXN1jPid+jzloRLoWwr4BBZY8XohXHW0dv0T02L/4G9G9nT/cNMwhqG0RuRabWllVXUxDNdGACU
e/eQsB1jBqOyaWKr6OcmaSbVyH0qfG2CbxtF7z1iV4kVlPcKzuCl9Fe5kzbrEAyrftLFpuEynHaN
7AH9ne/XT7ttEWvStJa9Y8y4PigwHDqEw6dS9BYdqR+7W8r+Ug04703WYOQPmuyvf49ifiFjikTo
qnf6PTUniMjyEM+kTAwnxOchnnZajVYjKw4HNj2NI/kERAB/c1j86+13eQ2k+lLGg1aHAo8J2+1s
W4M85coNpmNsLq/m+4JJvemyb9XKyJ3uidGFXLt/rShZqXy6VoPALpE12HGzq6MqZN0mB1rVW1uf
vNQtWlTsHxJo4PvgPZwWLUrNOLOVD8anb3vELMWmgJl9sLTfXjp0fwBtMCuJCM0K0TXWEiwEAqNa
WQuu+FAP747PFy3ZsH1kCtn7ZjNv0qZKOX/DBBLzX3yxhic/9Prg/ekx6EcB9cJg5ea7vMwRLwyV
R3QXcUTuuPxhDXw3TEMhgudQKpfmnvGnuizL5K8ged8GkBZDXHDpHEeFOqRJKN/5xdvTFXdmDtcg
1z7ve6QaOUvYBnA6MT6CTqid/nOYSlIuDoRgUrGM20p90pD2o37Sqhkxodw4GRlcUTvXOm8UGQEm
d/yjcpqHbSTGygnrDApTaYY10Y8L/SFU4lY/Qo5qzaEEWo8p8CHuvCqPTvC4XwFfRxVeuS3ZXyFA
kdLGMS3XbfD5hpJhs8BWfirgsf5s+xgm48WwSnlHMfXP6FFrbJdGzJcBBFVgWfBSCJXhxKooMt8P
dhF8vQ5q2OAf/rvRmCdLK/kL51rmZ1h/yctliMyRhw+ZXmIPwiIJqFFYZstaxMdDkzRPXZENvcI2
YYCUYFpMSpB58/iTSSGjS0F7aUChV9Tn6suYNp/Ai4OVL14lRfDld4cI1Nr3LdicJ9FvYAAGhB/T
B5vWZapI8v8DbNKWxtkcLPebQKGkyDqIOqYsTnR/PdtX+h/ct06r/u3YSSWyFoORMzJvSws1OJLr
qlA2DFrcLAuhdmsqoLiya4hGBl4Hw3Tr09h05ih5zRuSmRvOXfxLxqzKcLDMnzE0VbvhpPnhqFpM
IU8+lT7fpgI1qS9F9zv47OxbvufEkXjemAV+VpicdJVjhZySBrpM4XeQzgVBY1Grc+wb8j2Qz3Fi
RlPGuv6rJchQbsgZJuu9u5+0w50CTvseGJ5ndDKn1WJUHqJMC0H1c6/0gktSBzeiZ/wMzn0wjzye
xlNcGEF7G7dCAt1KXpRojcayx24Ts7lRfZ1ULRY0bBpm79ZIo0L2OghztYmvcOdhOkg/EWlQn6YC
UzjDauA6QHwMDBfEP/nFYOo3kBP/N5PacAzCe7yxlcKrdAJ7GmqU7NCAUJBEbXJMOQPUK4Do9AxZ
CcDdU34i5FzyJqEFLJBQj+ixZLl4bCe+BrmHRbF0ZVuL90nLlydM1E5b08Ifq+uY2Du3UrzRsl6o
y6/Oqfahn9loaY9+xcof2aGjSnCuUZ4rWqgU6xdt8IEVxdicGGJ5uZAY+ZG3uJlET4Sgf2ewGFS0
Gklf4sR1e9WLsUChHuS6deRH8yrT6Fz952Mpf5fOTw/JrFK2aP7SB43++N839EakoBjO1omAJwtG
KpLutWoJYoGNht5ALlyW29KNfY4YwO0OH4ZqyR3fMmcsD33UQxPrbiyA81kqIvf10CY2knaA2M6a
yRqipfFU72+e+Q1FBZ23tDR3rz4jW8i9AInCmwKNy+XbcHsOAYXkog81WWNt9FFe2OzAMNW73o/A
Q+HAWcCVQP0lgvV6g3Jr7DqwP9Fnreir/zF3tH/jlkvn58A1tAJFwe23ayKTV0OLIjwSUEkaERJE
7fP2ZY+qwJZxNgoLqyZ9OFNoMhSk4foj6t8Fff2CwEKvwKtQdrY7jJ6EbKrWcdgeZw3xvt720YUJ
OluGfbJZl0zuM74b6YXAvsnGihb4IrMZq3WAD4lTPuOMJQ1Sr2v0eJaIspgIYvZQsGZkhl5l0+6r
tB3wOnboQ2NZRekQcpZxw23yAF1NZSd3WfO0a+ARoSq051n++3VIoqRW94787xtX5JD0u4+TeLh3
C4gjV1UNuq1EtSlUAy853z8qGLRCC0WAtHHrBnU8CZxoyrjVzwpScTGa2LIRoRJBq0mCX+x++qGP
Ct4/+d/CicAk6zgXAnpzVuVOaTnKPuD4ZgLOFww2kJY6pSrldcZW/fTT4blxt9QUXy6pVs9Xhzhq
PvutOXHXst2LO7PqNK/OttxjDpu/mSP/WkQaAgkueCW8/hAKj5EAX4dsmESBqK7Q3qtOL9HRtYG0
gFPYkyJAGU/dPRMTr5nyFIDAjcsjN3HxLlHCDl3GUEbDRlHtuK2cn6M8BCvmE1B5Aw+M4Yo7TXfw
xqc5mOGi9KPMYjjZ8+TQ/Qu3kTv7AFMF+i5IWAs0VplJxB77G3ecN68cCFi32MJYwTGj0g+rzdUf
ZbVFKCMgr+wjNMsGit7EHEWeD6sgPxWtWd4QtEXDdt1xLAOOVNn+lQsVx/PqVmE4jCTZR0Zrt976
ZTVETbHZ6VOaF/Brjk7dkNPUenZcBnQojYgQ+iGTikivjfn4G/2AOGfEo/keYbt+JiyFV9qStTse
3S+a4Pc366F8CHpeYqM0T60Ftt8o2f3kCDgEiWa2dmq0pw4d/7ahqXGZfJ+fAJ+hi/Xi2fAX2Y6m
gC+RJngrM3YRQojTec3y9nnOqRuS9zdpYxCAGbP2a6e+28jxWKQ02q2u1fKBQ9oPgD8zsT9/cCvd
zo4vVP09f+gcmYAvfqVRRpoPTPzU9QdfLCCYoAnIaVSCChEHYECIqwzfOxwVFkvLz4ezrAKvB3+j
Nvm8Q0BMm7tPc/mXyKQWqI4Uhk8aE3J+5n9ks9uSCowGoI7R0m7SYCyOcmcBAg5pTBUsbwjLA2LY
JOhbsuNQ8Dz2is51+nZEPoUBcY9Me3egk9yFz5pzWV82KzVR3BoEA/WS/vP+jzeX1CNoF3oa8TcX
RPDCOfVDwsQP7FHuDZFbsRq5CaZwzBg9tcUQeUfQ8/zHFhmMS8uT0Q/5NKwYfSuh6dxQqfipEMvG
zEFCfbxkJqh7Dr0o0AyODKeUFlOil0XGKg8NiFVAD3nXPaVv9Q4IFvkbHi3rro0MSUTqGNlIm7ol
7V1FjgqMVf87epbZSv61mbbOT2H34d5ozIXj/0c/dK+VyA6kYXmmfZWCnQG4z43IHG9r1wwlYEWQ
QM8+b7y4TDVtONGckFq6oRLfsekNy8wPCi1f8S6syWbGpdlfNRkEK7RonlrgMnqHf+2TbFg7o1YX
wo9fAYmW3e6vcHp8T41LaYGIzM0Q9vxJ2BnspFwyKwLz6YHikJGgDThcq0pJc2/pooDvp0rV544j
QeHuUn9UNqka/qu9nel60MPUTdC6x53urkcR0MeEHUHdk/+MAjc7hCcGE0K2r/5ji9skdyKixRp0
ZjgkovQ2D9R5sqfnnYn9aNfyV0F19R3y4LrZLOhJLABgC8oqjhY71+EuC1IznRAfOOWT1ErugV5A
uA5aCNRyoOjH97NY6vtMUzx/IMBIKdWi/x4m9yE0NtuJ2epoprcYfW0QFrjBiS2qIs+acx/t+YlG
ndO1gJ5hnjSbWrTNRYVO3y3AWGRyRX0jITq6YfQTxyDHelLvnPESnDCby+tJvLDcT3fa9Z5s3jQ4
PKm3tU1EWg/2Nj31YtwVBadxgvLHKRLG7docHKU4onoXFpb3D3ceGbRzrHdGKm0iQpDODmFFQ99i
qTdR/Dgk1cZDAFnQZGodJVOHsUTEu46ZS07jksQwGo6JfiD3iQQDB5uvlvsb4xDGK+G47ATlDdT1
QI6diT2/5mnPTMruUJb6YYKn/DAoK9DF7uYjreRUPEjZjD9x1vg6gW39Y54bhhoK3IrEzJCF0O2u
VrFn456ymfpmblwZ61PYKhFz9Im2kN09LpJAw8SSZ/s75dmlrocVsRPXXEER2X2YQ6bw6WmHkkMD
0F0c63LzyYBthcf+P/qeUNnnE5uMTjbu8hltCcDrcbRDg5zVFf+wrWxETGl/iFIGFtiDj6gst9pC
BpAXaKzHlLqYduCI/rDVoNZEv9CVcKZFllKr5MzBe4bqUcjcNdOo+VdeIgPXtzFfFJim10XHy3o3
vJoT8ILkoPUnpC8CD1TUUO7Y09/bCHfA36W5GFf0z/IvUd0+0RLXF9XmxLWi19fbutRUlUzzCSOB
+zroffZ7Ixz1DSo8UVmcSrjo+Nj5C2kFxKqb3+aHV5ptb2VuWR8P4eql4gEwzb32xRtPg2/JpLqC
W+23sIqiNtE+iHhsKg+3qO6vUD1Gq836rBXLyxSjnf0cT6T8JrV21t6p7LXUP7JgAuQM99qYELZ5
KqEUB0oUmCsQkYprV8KblRYEclcsIiqphPZSCLpBW6OBBRbY1qpf1HKN/C3Jc/nqQqfXE2+SQDmz
8MN+K0iGeHiRFko+sMzWce8pKds495vQehgDaAlRDpIl7r10HRwYziEm10NoMYo4IEpUTsaaNiGJ
suxUgD5huB2fJdYgcx32r7w2wFTpWKbmnIg/R1qxRBRlje1FqGU+zPdGFSs4c+AxJ2vvCW9RPbLU
TAxDwQ84brmNelR49JLq8t2f4NqFof5vW5ITTw9MkTnPFxTsjq5IFa0yWmw/vA2V672pN2oV1wv3
FMchFQAV108pmYHl1093ZzQIg7H5ooFxt2shFv/9RWfvpIM5QfqEO3hR2aRT94QFoJ4nJ+JJQf2n
VNTeyYeamjirI3ulZeZ8oMzztYp/jw6m4N78qHXFCqPebac0GqA8ywvZZvlas7EQ/PyM5huHQ8jQ
5U++0if9tyj8IBb5/6SLKh1zUKYquFUv1iGIil1e9n5Z1Ua8BLM+Kb0P8mUmD5oENphdS9vuJAwO
BZOSOGCr/VNxdxILmW/PRXv3uT4rwq+wLB3D/joBADfdVtQIYz6hEDA5PpYfqLW1uqt+1Aj7i6uw
yhotP8pl8X7DaZe+9E1WuCnad+p8CsATf8UAVuhIYE5qtUlO+viVG0kjWzaqUmxDf2U+LGWMkNxN
luofksM4UvOS3WcRrWOlDOvkDIE1LlFYI9pKAzbo5CcKbN6ShefiqqrEP9cGzE0GKqTIxDCYfvgu
PLJhT3PtLyycTAybZPg+URDpOAxVziNAZM+g3w38/Gepo0X0alaxtHJNMVJtnaKpVipkPfTw6Qh0
fB//gFpGXA1vaZM+nqoYG6Qn/Zh0JJZP/XRmtiDK7DN4TWd2NOZrRNzpCXG3T3/6H5BOLmygtRK4
Uf26DydhgxkajYgCqiYXsC49UAmziOPQnbcZm/Dkba3bAY5n7C+rgKrUBP6RNa2zCmhdOUsWfLqS
v16/7KXdmH4wWHkdinbSQjJUFpcc6gFpKa7e8K5JFF1rjsREMaKFWJJHgct3luIWoXu0wxELHpR4
zOHLl/QNYAo+qy7aCyob7wM0H2O4nL/4RNvlDiHfNVQusMbg4fFtEG+Ua/1jRrNhy4IXAuAnSAmV
nPJmYWrQIsYwUM1fEqzQ9wUj+RZtbYApSOVF4TWwp+5fIFwpmsjGWXCCMDuEP9DRSz4f9418dH8a
qD1Mv/pGjvO4KCziHNxx9G5wkx9q/HOkgLjfcnigSs07dqvszVvDipWPkR8/PoDedL57IAYEPJVA
rI1PeEE55AyTWo9+0TzCztnGmjHbicwldjlnCFZC764nVpSH8pZWrMI4MfuSQtb3/OMGozPGgti1
aGt5luEXRqBkFYpLbWPW6yWU90GLOsNc1+UEqvq7zmDhtOJG6m0hWp8xMZS87DxX7pInHA66L8T1
QyIk6vAChr4czGRpVkO2i260mJqmYLbxgohNrj2PNL8K0z4Z7GOqMKpOyBRz8o5jIlC3c4XON67Y
u1Ig6hORuPzyn0fQaQaRR3ZqJ3QzJsoIUp1e6iMeASct2tjZhUiJ0XyW36TiKE+J8p6mpCIHKAzH
66Wtjm+5iSs6e/kzmZgPZV9QNVGzfy9WJo8KnMM4EO/TRg7J1mJpgcnXKWfwc/nclx0y8WNErdt5
MEF/vNtl2YYitYR8MqajXM1Zgte6VrVlXO6A6Fwp3tdgdLfOT3Sd/1fqA+XnCUW7MbTnIOLmoTW+
L+vUGGKbp6tup4xdcy9dlRLjpgL+ptroA7VaDHOOl0OxXfOwcxCDckiN+Anklmt5/LmhqTu6ZtaP
KvsfFGbyF6/RUaAKxfguGcx0xcQlSFTIz/JHBDxeyTV6Tu2cMMVFaxD0133sTgjZ5BMQ2M7tozxZ
nl0BHn1/2nOOaSrpvlpG2eZ26411h6HeEe75X2Vl+Y2yDitB45rBO27fHtYVz0iS+k+tSc68n7iR
zv9bUK4rlDUR7b+Lo+UPy62GOZe+7nRHP1a+5u9VU2Xr1PQNIr1aRbnqMVTDVKp9qCJiyRn8yWDv
07ma7JdQlsDA8sS6kU2PVqXt7hTdaNzgSUtxKESVjcrI8V0DRVXQ2ibk7QnAzYHqlHOR9Z2b6MD9
+tJkKZN5DKxmSeFdb/MSznuzzmzbDjlhiVkrGdKkEbJc8T85ZteUuyARbNcZUwzHBOlpN9ZjBqG0
tL31RzR9MuykgiKfaSVf+hhCA/IwB9RideNHNwR3RigswIormNiBIk/u3BsQDlGisihEVA7TF/eP
MSt4N9czKPM6obZv7e7eao7oK8msruHAXqvNqJuJxjc0lEJmsQ+Ql30yjYpAdZ8ykviTJvpLKb35
G0gphUapAkBGxYd8tsk+qdOF6Pq3+lz4dQUFkrpfVVp+IZk70cgN8TfpHIriQ1fNMW05boSeu+uJ
DhXBpNyFTetyoKsLcLckRJAT3xKuyghKZ4DCLrSMHaNTa0CCNw84U67W2Ff/vmzqzmSnVLuWAl5Z
wwmMIqG4z/Lme7max6uiKKPOJinU+CNbsTEQULDnaMUew5tKh84ABeqPWWuNvS59EELzRKS/ni4o
0nTr+FQ04lVdQgid8fsLcIz3lc6WdEQC84hzMB9uoc2XLN/DTUGVhgfM2neHYry7viKzGZhxnc7p
EBldLOieAMkl6pik8MooxgrodmeFibDY1aFmvOOzDdvtvmZbRdnBfa4TrqSPwkJByuMESuy5ynce
jjgh7uxIrvqIGzE4y/nGECEmg58KHdfdg6S1Fzzxh7muiT2yT/Tw+sPcov+j7/eyrVPjJu4zbCL3
J17Sg02/7sT7cLxiEU5jm7oRw65Si4aJHJiaL+YNJIBu1TZ0eLJYFrOifl70tSbn1rYl31yxrjtw
oE29qLRnpV2ZSN9Jx+HLCzDIwkIZ/sM3sgNYUKbOScd9w3zXTsBE+0Cd5m+0r/ociDKJl7CAx/wa
RIFfYdX/H7xE0zcwHBv/sG0wWJ1ukpxaxs3ZhM9njsiLSaWFSwnP3QUItdRsIQSLoTKLIsqHhl3A
NAQ3pl4ju3FPjm57jome0XHZ7K9vlMnQPjCbiAwqxP5wiaEiyAyfMCmkUmRUKuCaFkPwEH7rTnky
lCPiGT47kD1bM9iabq9raCSfUANOglhgGOr7WIuibmfDQ0Ll4y6MsEb26AZi956QNDiKq+LhFh5L
fyhpQUCPMCTMs7OkDENNFcCYUdVbh78N+wyJf2SmSRjAXoaH8AjRc+FZz+TovxziKd/KKJMDwo6I
GkdW0Ad+E7oFIr+RAf5KgH8K3wRuyDJOYmhdST8UcU4DTUv5T+/BRJ9XTpdSWJuy0ty/CGH97XQq
WpzoHoi4xcxfG7Yppxv3DI8J0KYEmnaXsk6BvtMZ/vbs032AjTGY3P+ILLpPAtYASjetffMiqoh7
XaK7r8gVTKk/Huw8bzbliwABWhCaxv/W7P1/Tp9WAbCJRW/uvFJ6vJRFBl+1X/LLcAHYFMKZYV0a
oxuCsNMlM8f2NQZ6cXcr/qU9Pn2SP1ZfwqExhye54bU9GsaUw29RpT0/5Ptb0WyWfWpDgt/6HQrS
xsWTu0A/d3H0To85LyTMnnFAVqz7wElRaLcp+xrnN3S/PNiBSfs0ng4VhaHB32oYO1z41GTFyTe+
f9+7KPksxayS88Com5OrerWVLhrNerNZtHsd3TQWQfkCFoPSUSiUM4+I77Y3lMtaIQAunIS7Euaj
Ix+IHStcLFYREYKrOHta+3tbvMP9YJA7fCZqtCxlmqTGaOD5QM405lwhDtF6ffOXfzBFenT6Iy0N
niWoo+zHlG6g8whHVIIffCSUHgBamnhhq21I/Uh3GI0CqPthRuEzKwsIp993rbBSa4Jg3g+/KSYa
0Aa7fcT6m70ANUmKjb3gF/zESCCPea88ABTsvuLWN/ITi8E71IG4WBZxjowf2B80I2GuqCJhaQBe
/gyEbm+DyXn9yXPaHokx2Hizp0N2gAvXFGaJpQAx8ZvGc482w5n/uv3Nv1NJ10lyH86T6D4KA+Aq
+FpI5qJtcM+1WpqF6Z3H1SBcxTBKCQLYhtxPddsU7uEv34fBdXI5vSsRMLyiVDqBoFecUJV+WFKR
niQfoYuW1+Yumb3h+Lnih1KrGnX/Vw4ztcfL3PsuFlmfZax1H4OeAz1+Ns40ZmDdYCjZVMYOBIZt
29JgSw0lhLi+597Hs61addfTQB4nJLoqhpRr2glUtnC2wgO5PTopYNs20vkzyiNE44rLAl9o+ihb
xwX0DOqClXU2D6EivpSaQSFresDN13p7K7s/M16rBCFjbQNe5ZwnvKBZjG3nNnWBjAPQKUuO6BWi
BotbuP+OSSXdVF8/+6C7hYCbOkdqXyytVVUGVi52ComyEfmw6skNGzuc9c+kkglVcj4k3gtQ9lsQ
/AMoj2aN5g93PFIqQYdLbZwR+r0gwVsM3aCoW2EsdLwY5YUw0nqS9Jz/r9TIdgjOkhfdleCgkYE1
F3gL2gxz8zLkkoPhqxDy6w/L8LZ6dPATBYrRP9NllmrhTiYiVG44g344qyUIJRN0NucxbXtlK/Q1
rejt0EYUu2ONu+MfX7j5lBeyujLVyQMe7xIiB4YpqoODfuj9H03Wknc9MSdtoJBUFuy3E1kslncc
Vd0PAGrVFbrGWKvDgKSeJIzOfdkJKOpUxCezwd+pwa7jRTUz8H2PRC2XYGIfDWsjkKKoZWcl+J/r
PONMINR5zODRv0+68JAZNpH/8FrRf+SSHNnCaGOLGwDOVwBB6H8ni0BuQhXjTJZLCxYY/EK3/wDf
ctfOI9MWMWKb7QzZ0CSfv0KEuKJ9/WIJBAxrfZBH0qQEH+hnwQJVhqdNIUgpaVsgoU0fqDI0YfQm
Xx3VM+xAfqGmDRBTqYUdqcc0WquxeWZ68AqMb/2hkP2x7sgsaFDLlYPGpl9N0CfgaYDMxYsqghCO
Mvgt5CCzlUBdrc8qOqqXxbf5pjwWRd/XjzWwUFApRkFb1Lzjlonx/d9aUgiYJMSHJlqWByzD9ezO
1T6z6ZPUhGsO6JjU1NOrGLkY0pm/hrsR+MRcDyltgmylfyrf/HzrqvCIEZ6fhm657NdK2bISOrVQ
PVOd+wS4vPR9bChGY+82O+2wb3hrbT8D5LBVDP7Gx67NYIciS1twx5vUC/L3nRXtPQwS6CAVcG2w
c3NHU29toMXuauv7MTIhEuTQ9hnfeOnA+k+H+irKa94LRn++onKScl1CRZuAZKFUPgZlM3TTGFrO
EOJMhRj8HNOqlkpHIydO3z1Zmy+crB9LRbvbzxr9Zl2EnBvkknfZ2lNsQr2xnZH71acAwu6iNk7+
1OcUXzOHGaA4EDVIDl7Mawm06KU6M2vBpir1enrbc96LziCJIL6QR9Utr+RPWtt1Xhn1uAie+GQp
oeW/GN+Fc9SazyzENgM1QRrf4lfZLfdZRMu9uifHFwLZLRv7xICUs326LG7T7TnZAiIsXWUOLCpE
7uDZZTL0akcjFqOXQ+lxMTFHxKPb2TTO/D83UYhOBo3ywnr2tPiGYfzp6Fd77gfW19rF8Tcvmrs/
cYIYhQsHcYCeK814HBhTSJ0VCaAQ3DNmmbvGwnFDsKGrlXrJD3/2iak5C0Vs4vX//mzTB5euGZvu
tqWNIjg1MU+6n5Js/HRWA+kbV6UNQbaHkPZepaV2CwiUn0TjFQgXYS0MiFeqdcXrf/G4Re22Brr0
FowIPfMV+HCzZhZqISkAIphmWujDp5Nbqs/11w4dzxRj8BARGrzSCyC8FDK3X8udJsldBZaUHSgD
4ozLk+1IeT638ujzHvaKdtZyhN1nOBykJJclAM/COMM3XiQ/Cb5yQAq3ONkCVtSYAxwJitZGe8Te
90Jo9p2LPWDCcuJ176aV7KwkG+Ar/+jPqMNdLcDLrHqN8PS2QlWKtiEZZwppaXza1tO2PvXLNXwB
aFIyZiUQnCbhse8V0k/RBwAcIB3+tfUWSxtEiQSfgGevoY6gR3Sk0Nb+XUhx7xqrd7/7FVXY3Yun
uPEtTCfLH9AqiJQyk/HM2ZAjuQwjnGavP4gMiuXNKDLnmUApkR81rq8yFc3QzqLfqldmHYjOenqs
2l++U80JQkX1+zjSmQwfXRtfvho790M5tVAbNUW2a6AKvxxWhh4bv849Khe0fQ0J3SoBbwkabN57
Oox+Gvuib59Q5zyxaPoc+ojwsyiYNM5cCR6R/Ow30s71HJflrayIaaTgvEJL99cGmEC8WmBgBpAp
nlogSaRt8Uwwgs+svCHy96NnodT1LMNdEJNfv2GVwO2YBFMFsuSLueE1LLqkqPCtQfOKTW6XlUQj
KL1xnL83+aoC/D7WC3Z6vI5DCxCDYD3g/aC2NHVxe9SHzYOwXKo5Rpkxsxm+RPs4oVNdd0Mv+QRR
s6ACgtRRpcJ12OT9jikOFZiyb/DWQUaVbrgF7xKlh0I/7uUn/xJv9QsE8xTsO4mfuRwskxeWPo4p
SoPNeO2XZBDXnK6w0sWkk++PS71OfNUZWoS7zdS3A4iGK+n8cwGJhYTWGbjgjZOzpciZuXtcW3xW
7qBKGcgm+BoOvlyFdXQrCVMCSPixRtwZXuhhzD7Y+8baz9KZECnanx1qsm31D0K7a6LJ0FmYmYXf
G6V4jS8wFJZxGKZc5HlgPdf2cdV72PoSFxOg+GKsOSfY3YhdccdHlnUwVn886gIPjATqHVCnnRy8
GAtypSuIYE/Yaiw1lwxsGLEGNEG6XUbX34A0gLx/nG0vrqh91TEquTU1Upz0ZByIApdvq48Ko0Pi
et4jj22I+6X9+srJTG/j54ov1NL/pRMV4AvY0VL/4G8DSnEXZC/fjYPLc9C8AOIgBOrWOWVEtuJv
8tFu6LdeQtfYrOxpg7YtCYxYkSOReUFOivUFMT2akyxPOJZTth3AmYVWYvFBAl5d63pNpLj6IILM
L2x0puaMFvZCek01OVQ6HU3ssr1jI0Aq2YbnSHJ2O3r9DtpckeNFdQWiR+k56PtgeerXrTCGA+4r
BRzS0Uz9AdJ44t+cnQyKsWm1snvgweCVxQQIsqmGYDTDP7rHhw/jT65OPgMH0MuoJW76jZj0x/KU
n4SL+O+S5tbroHvkRlyChITmq4ZOvSBrrOQnkLZKZtDXcWL39mgCxxJ6Myjzc6PZ5ix4frRLtCy/
qaUZ5qoR1dS8NHUwzgdIszBuP6raO+m3kjdJ0NUV72RbLix4BwegHN7p61GYdyNdQpoi0VCRQIpI
R5ei09mFDXvUAr/qfdWJqR3Y8ogVE8NMJrqJ6KNuJUukBMUUsXvI5z+J2AXxlFFF2NUAY/QSMGQu
3dIYqPASaNfPyBQ1mgmNqcWiYY5gmpztaR65czfPhheTciBQ9qU6iEyVJuXuM0hZb3eFoBd1QQml
MBkHhfqEmcHTzvA4LrHX+4/lusBSwQ0Tyug/UHJ/cEbtWtf+JZ2OXqUgpK0ufa4guu4rblaY5SaW
ZwkDPAaoSVx8Y0n+ndEqBx0knRVfQauzvRER1siVdA07XNt0cTYOZRGgzNpfaB/GSPFqAxVDTx1e
NCaaN+Z1hPolRZuHjvcmKOusd5N+9vI8cooJqsGUiPY1eT/dR3aOImUpGW6kT3NpGiZWNLR8pvpp
HjZeJzjnAt700ZaV4AHxvuH6jxYS1toUlDsITjbjs8D8mKPKufO7cZaWkp2t2Klq4hw+TV7x9OFG
rSKoKghHwfvxbQHTy6jNZDxGHzXm+2Qs1EA8Y++kgfxHmWisGQaLpFsMEGYRRFZjkbMmfWzjZ9Tl
S1aSZ8vuKLhiRDgJfl2120t+bA5G6zXrOnq8ZgY4KUVBHbqmfx7qXArmMC1KSJ1KE0XwU8ZbNBZd
3KwcjglaOpD9jpvtRrARmgWxmkkbcwpOo1+W1w3pojMon5s8C+NfGk0P+fEd/+/qAHBqTULZ89O9
+sL7k5uJRben6Ca6Cp5z5cyWR1G+GuKOLVa77UKmLTKkF9dN2WFC6mTTmDxTV90cS4tBz/O/dE6H
3S76U7slDjy+xcHwphTuzGUQRe55SILsDjpLBvRdT/VqE+oWNVP1nXv9IcHRhvHayWEzbzuz6AuM
vxD40BBloDsUnDSP54+Y9pml3aedohM4JUmhovlu+0sAMiGWFTH52LTuMb4OJUSwDghL9Tx7AoXD
VKCaeErU4pdYye3wf81F00PfYMjxfkD7DKeZuF1whDTQ6i6t1GK//SE/hPTyLEbStQHJ6APcXgiV
AFMN+BDPO4jaDtlOecqByjFS0dus9Mw41vfoj9M3xoCQIyPEa8JafydtqFd05HcIc2wnAJnce1iD
Asey8tZW1hUuL0bHh22Wf/H4rToPfn5g/qUQoJi+s9tyUt9vGTMKV3eyMkIqVpJ8jlBH2ocVMOqV
dmgguwPJbvMn0q/oCDh1rCvtEKYBN6DyuNeJ/TwwNzOdqA+UIMlPOJpKVtQYEDvM2xRnCYAEUeV/
0ThTNZMBTK4dL3nl9TzWRf8zhI6CMdWMsNmloF+ZVplqpZiZMboScYtZYA3JELIpJ32iLmb+opq/
/EM1USQb7ImRPGvngoo3ldKZDHIzUim7TpFN3TLoBx/Kl44VV9xb2NQtvnXMBT1StDxu0RLfkTgW
vQsw0b7w9bpQC6itFiC3Un1EFo3PuaZCaEvzZICrviiNKczY6d4k7hMfw5uC4Z4XTiuZrRZzkNzK
imZEiJKRyknmEUcbUbNgHvDKfAPfwdMm/DvgIUyHAbNH/mKBP59TEvo18iBO3XMAV8on2CyZz+8x
qcN26NRXYo813vSvg5/5lFpz1fsePAtk4S7GhpDq433GYUM4SgmGCfUT/EpMaqqUKYZDPGRkgm08
MnzgixJkXaa/AmYO1EXP4fAtUgMW1me0qZ8kc0jCo4FeQqlJLEvL1FfiXUTNZBwlp7Bow+4W7nm7
LJHNCL9szkMkDm7MdVhXNhwoWJG/w8CjRrWMloQGrjFiQdTCMjTkeijTOPFqhtNraBioSnhBjP1U
4RAoEb4SvKJzqMUxk+/fGIDw4/UUhxEGL5/mJmq7HK7lbTltS0tEkpLwxON6vp5ylc7KzSbH/XKS
s6k9Y1gh6UsYxT8A+SzglI/TMBKinj91p/zlX7YKhP8Rp2JdtRGSNJ+iPX6HUZifRrnh7FRpamS2
kCZhNYJsQKagzmGqPTeMku4r0WA8W/twyvwLxPYc23/IljYIggm0WNnQhsE43DoRROXWIvZKU48P
cc40tLTgzyHKFBSenzhmkolPXvCcaSU7blvLrvA5u9GhqqYWIrOj9ZyIdAqCjwalRcyEU1McknTR
LWEOufANZ3zRWLwbTl4u+7Y+dH3QnwoAebJ8XtvG98M/uL8akI4SQ0fgev+02u04TEcHKd2bv90Y
hRhRI+pK6zSTrIJrofX/O7kveIzg7W40dGEQPUarFnesD0jxhIAsyJeB6w+uyivQytl3jYBx8jLZ
79a0qG5ls+ADMjNcBdBl3Qey94XkzyE9rkdHnJ4lAK6UYfjASYxihwbLxwvJqHuDgipZsTdGku5H
uT8GwQruKtg3x4j4G3nQ8ew/QekMpSgOEdqopU13WuiMNpog+aHcBo++WHr0fzqU4euNG0IZCx/3
psQzRE6pbaidtcDPOwLdRnGUqvc4/kpB6h+xnHQnbAuSI7TtulUwh7X4KYsZhRCNLhQ/ALh+RUJ/
tNgIpR/KaXPvCqAOWSqkFmQUYtH2EqLEC75CWjYreU85K1G44ylQEcKTbuo10a4awDX6Up9OS3z1
6TJWCCcvIVA5LlZDLlz8mrY/j15K55TrQx/XXwWQ0jLVNhwUAsOdEi3RU4ZL1rP16IX95L6FUYBy
jjxo6GxfCY3mcc2Vu6dmilhuJ43/LihQVN+2oZ1NDVeKjkCbVqxRaNtoxRlKPYa9FozLFSsb//3n
2TLItkvzxtDgwadCZU3/BXVPIaru1B2z09uT++Vt4qD4u8PCLsSMR97QSAOH/f2SsTQznvkjiGLd
sspeIGQXmleJifDbjQ6c+WepQ0SH3Gf41TupOGA38fNM6VjT7WU+CZA3/rinw+eqnLKHkD5RMEEW
mqlNnR3oz3Z3EUL5ARzY8QBSdY7iLyUr8E7EWNuU5u9sZ5115RHh1C/87VWwCSulHbJ79te/hxoK
2JC823YEPE8johrQ2D0Ho25aKaov4RmE4nAoQhWl9Kw6IawlDGz5wCRPLgdHdUBTeX9QdRAP2A+6
s9uEj5TEpsZeIQZwgHGdWTJRW6YD211rJz1XQihECfXD57jlOcpLg1vovcDceX57SR5ACUPG3O7N
3c6MNpmkWrfiXZOyd0v49n1EQ0///Tu3Bg+TRLUi+C+BLUZjTzzt0GAtVszgtY10rEbzaYEzQcVm
k7XfsJ9sANAJYtiAdyfl8iK/B9ummEW8E0FDNGc64FJq/9okzx8e7JlTVWaaKYsaTQNxvu5fWJRX
5uzm37Vsk7g+3q6GV6qI6IC+RLFZBD8p43wBp3yad8hjfgTGc+a7ejerbrxuz/JtUywUues1w3zf
PNg8htMtCUB8dcm3lg56TFPtVNt99PYamTvUJU4m3iMUq1eSKelkAqJHR9rbwuFSTgm2WtQKDvO4
0gySXn8wxAyez9bOtF5RIJGv4outLdZDpq3BnIzSzj8v8XMPZkREbnd1VVaCD1lfFruT0nbQSNZi
xFGEdqMHIkFBjOFj9KuoU25EbAa0mM5ap3cEiZhsXz9UK1e3tLiRCFVIo9QOzUhK2MxYIyKv/vRk
XEMsWgja7Y0BlTdJwMXx0YhcsR8khHo24aJ0i1I0AsjnNSVaRta1a1Tx51qcsilOlsP1CQ8lRPHe
qHpxPTLCtjeakKVsipdJeSoorRdVTtL2S1SP6VTOcBqXQ8VXEqwAeGZ8RU5Evdu3IVuKguEcxnvF
bByfpXd9cwS1nwXd+pyTfpjAXMKbvD2lwdNFadD0wvM6r9qPUE6W5/D3Z4Q5umHob0+oZVH0TjtF
bre53ee2K4i5SnqRb4lDyVOcd08d6SB7NhIWhFLJgdh4jYUyb50b09w2gtiJL146i4yG5DRuZ3z2
t6IbcfAnMm5XtRbAdIcJcjV7wVRleRe09KIRfGuAJFySe0qQUGJ78lZv2GOjq58wyfCdsvGyNqnK
g5Ktzs4yJlEVk1/0WznnZKwTMjgu4+FiyCMBvu92QT4w/VukF4cHcQ8XRBF9yKRobXVVaJdekNmf
0BdyTuyFCfMX04rs73hnj0imKO2jDNo4xRym7GvGw6dV6OUrVLTyVWZ4WI1HS4YS+H/qVeeVLQJQ
JYG4pQLtoeYFu22H1PhAsEsusOAfiGD2kA7pfTGbx9/xMG4BvZf78M7I2rppWVn0hOaCfavq4E93
86Jur4j60Mu99zobvjJjMW5AglqeiFdaoQ+0cMuPVlfDgULGosEuIpVF/8UpU7v/7PWY67oSP1YM
RVp/wXfztF8Jd1CVkKth9dh/G1JF2tuqdsKn8E2iScAwErZPpCyilHLqwvhTUNo1EKpcCQ6SNlm+
RYXfGZrZ3DQ0bd6/QD3t1dBFeYNQ/K/KBgxfO9WQGT1VyTYMb5mv0U8rPsRXVS7LE/0wmm4YCLNJ
H24S47c9kMoOykv2/7MnKbyZwFLIp1eFweyJksnob0pADZOXbFDpeFxbinQCwpYwr4ZtevE146EY
welhq6z6TbNJIHlm4y5ljBFtAOU3JI8j7T4vdhHdn9WJRs4Ncq0aukzV8dJrwKv+aGUS5jMLKlN0
NXudE6mIWbzcwykvJG7wlAxUVIVqPilfTihrbsASg7o5VbKaTb/9TO5WzhDs6ILDgP+NkWC0qrH2
8fpIXRmEZgBMB1J7TIAVw95H69DKFSkXzc6vCoQGq/zibtH1QhYMUp+HYwW70FVocKVizWELlSDg
cSEJycW1JH/1wjH3cdPssVC4FxOXryE/hCWvHjxwf/eERJzyEkdbs6BWZA8Bm+NM78lxO0A0HfMJ
2H9vZivvteYeEGPUGimdxi7aWd0QHyGMGM9LnEUK2ea+Bs8WJMLs5r+niscnD+DdVCzxqmngU6ZR
+KrD0056n6gnDdVHmu/2hIUBE0kHq3/7zke2PbY0pL4QO/ckegQovtylEEXCOoZ1ekYplNrh3KFa
7pvBRqjTQ9hlqxOgxlioHOp93WQXAjxsSnduXLOOQHwOJJS3Kquxq5776Ru/Ix5gJvUxeFbOSK7T
bFNUDShTNbw0+UGH1yFeqkC+fZ2JB8w91PYGn7IQEymaKoKvTLqKpifphbryKGzfnMrjHjOKmj4z
I78jludEpbdRDlqB4X2PwvxiGyYMyGb0ReNW6VaUjDqvaYsgP/NQKyyZNwSUAc+kmpA0U8Il3o/+
HrV8jgFdzZI5x7GT79EWr1O+vlG3heyDnpSRccskHrGr4vd5MgLtt202Drrm+/XKjlI0JMZQwN1v
Snzxc4ob0HCAKIHAvfZf6lFs5I3dcIRbYCdBCkdpdhCTiHweQFbK8gTmKnGz6iLd96urNyDeuB0Y
vw0Hse/MtIl5bpVBfXKAWm1ERR86fUYHXcMV5vpi+PxV996MyIjc0N3xDMd7p/wJ85R7Y0FSkgjA
qgAz5th9D7+fIAUpRaI11UgBqJ75uZm6tSebizjsT2H2wFKi2fb+WA7Y9S9bgPlM+WnpqHzs/qoB
CKJpKvDLT5TNPge6ffmIdkFtABgV7vRXb7ttRUM3JGiXMOHO1XGuLfdbM76CrI+XUzinTiOdHulJ
ZEhc0S4h2CuMNPhN3msUiOa+k1cjvDE6dxNHJY1KSKdGAP5o1QIRCMYPz2kxtyl8+ar/QJX1b2QU
K4ET5GDwLls8L7/mFr2jA5Atn/F5HTU+1CfbvXHE7YMonwwOWOp+Kz4Y+WApqOBe7v5KutuE+G+m
ET0KFmDnhKNI96eL2nHC08HRBj8QWjypBe/FpmvsH4t5wTB0Uv4KJP57Sw14zP8ne9zgD43jDNE5
K1pzatGxdWCO2u8EN6eLqVhe+a1TKVB5X0GZo0tItO90T4XYmIbPLWm0WkxvjTseuI0stE84mPN1
Z/KTzk1ruls6aJWij3UrMvhhveiSI8pYF7wIUfpn7POmZLDK+SiVL1yrMjTIU4L7n26CpzEhJJNe
H2NOGuUqR5VC/1g8W45AzBA51JDP36nb2VPJ0Yez5HS3o14vF6TwiTBFV2w2XW+L4H1eUjhVllv1
0Q4IeRVj7vRmAjcpcXqpHqBg6q0v+GVAakUdMXs0aSHwWbFy5Mjljv2IEnOaPyS7ryDagi3nWiP8
FMstVj/R7kCPgsPYhc+zxegbfs9C6YHqT7Ym15lDcANQgMknpvoH3ra1HISF3ooRIsDH0jvR/mRa
b65b3a8F08DNleKvdz1SzAYcxiJx9F3k8Aau3w5mRmQn0Wo+9HbiYXV1nSI7tZH/sBEyl8GjAbPA
sqr29L7uBCptBTZE7BXL4aw295r7oXlV85lPTuwBoV+tKHQzmeis7oyLmTFRZaGP0BJ8nvCkcDF9
o2sbdoQezn7h3fPey731YHMp4RTG2JokAyu7w0VCdnLwQOr+qkUTKfgI865hL74txsjoRB6sYi04
6mHgEqS/y26h2xrlDkF4ztpm+T5Q7ms2ZzvpuicmXZ1FYvGtevjS1RlczhMKRhh2wAnTgtFIQqaj
CiMF/jE/tVRHRWZgnmRf0WoSHEFdJ71RUKCfaZ6Nf/Zu8jnTfku49jR5c1X3P7W3nMBMsy2rzO98
G4ig8+rZ7qF+6H3iLjtVQp+39pwrMEHC7l4riek7cQNriPR13sh1vcwVdVi1HTmNRiJ0MDbzAOt4
cjGNhvjBNlFbtBZbOgheD0BBeRyIvcC07Ol7gHMudHrvhwDx5BNER4u54dU5dXaHu2+JELHrUmX7
7KdUHNnbZ9k1SMJw4//lxbE572cY/tyg8Kn5pi96moq0UEp17/1sAqrOkQYG964ouRKNV5/npdFd
qYhsilDMDjy3DbkxbRzdOk0OCHpbEen3OgTA1ludCOe3v8eb91ZjuM+qcEFN75Eh9etI6jyiswTQ
CEuhkgIpwb/Q/XYowAA23O1JxLB8X9v2tFR9hD2tv6kaELvDJAk6PkDPZ+F3ukRZQmrnGyvr62HF
s7xjVjQNqLlKVdeXdaItyJUMmXXyoZTiuujo+74cVQS4JR3yFlSjiStP5yNbs/uws9AWhACusENQ
zrMIA1wVurYDL2LNOl3Q1KzKy1WQhWuYEId5LhsvpYK/4jR59es9KkhYGHEUCieVsYQq/yoBizG+
RBD2twxJQ+0w5nsd3KOP7K7vVGuaS5xgLbNIoF3SCyv2K3BQcrONTbtmu/ND0MGPAvKIig/JjmGv
4/lIKVj+IPShPCUaafU6su6VNgm3X1KNkw9g94M4oKY6LX7LEsH8eHDCDHuWa5sxNklJHxOAkaTt
GqxsTsfFTnMRRoupim89YA1m5nNrn68UV4OVKmURMF9N6zcVKpHVQJXVokRmTgLdS9jnw3+pgUMl
O6PxAcxII5gIyVwIDzEicowqGnGyU+6I8Z9EnNA6VRzx3BkU+cPeEMV5Skuqe8rtf9ksI6MkZANL
Xzh2Qj9oY4a4Ys2sDA5VFDTRraMjqI+hu/Ti0RAkKcxs+32K42W7ac1AxSGrZHMXgNonai2pYp2p
0TxBh9vzl9xzRzNBnJSjzikNWDYRmF26XzR14lwEiIBDqIUuX9JdNcyra048E/umDL7kDCdzEPAk
SfEBYFZvXXJJNtpTxUIbnIRXwsddhX5ufYTIjtyxrp/GV+IA4EYnFGgjDn5H6LRrEAraPsOBS/Ua
sPj2w7QcKYh/6DA18XHyKGWFmOxrrMtg+sETNRbpSVgpJirtb+maoHhIeS+DZHdpSUvf3nKZUNYu
4oAOU0ISVPGs5StcR5ntzbd7+YOtcvyKKWJd1Ua/MZ5Ax90kA6FdBjs6yrhC2ux6JgfwsK0RHyOK
dCJPyDuVXgq59u55iHPrpY+B0VUCXmqjennnR+yLnK4qMyW/KFJuiYyHqcAaiQcVuGu2SazyqkK0
pMd88LUmbQRAi9M5D9osMCNSAjCopIFygKRgc43jrutmxo/BZzYx2ONcz8CaSazntzgX7t+keeTo
RFrImew+XXLYKMWVrhCdh4+bPX4e/psgQXH4yO8Bc1f+UaPCgrPak1s1/SqOEeQgrJsAVTF+13+G
dHjXVUX7rptC4rxQT7tmB2JXSp7vcWZOs1DxqAuVZrDhA9wvkVx4JsjQtK8YVlP1wkTkXEyibtdJ
7+hns77JP7utXf1Euu86p8XwqpFrvkNFbeofo8K3g08iRv48qo0DzLdubf/BsYy5jgQMTqGSI2WJ
LbXR+mk71dj6n5gAr9GvOG8MetQbdEP48gEpSr0htHcEoa4Q3KYmC45EWMKqEioMWpWsFwURN04t
agTMJGLVNPcXdRsuEHfw3sNVyW+abLD3gwbynfxiZC7F/t9qkAAuJAP/VaaK/ndmhgCd0BeyUWLq
YCP34vLU7g+7FM5JcPBuztQqAjJ4p5g+vz/H+MWvog9ptU4cNBdyqTVwl1tu2IlGeXDVV3b/eXPO
25qXj5ab2CopNNSm/ylkLhXi5CzIJknpZVk2t5LmA+te5T41jKkxRcrvSlc52fqv+ycuyspITFgE
Gwrr9TKPIulJjlXxIU+CofwJDqA44vO/2/Wu6v+yyWDlwx3HQYxyWsMXc3X9XUm2rA8mSWfYaTG3
BqaRnAXoCsXZmUtY2q3Shpj2uVBl60CKqYRDIP8JzHDKSPufCEaJjxjgaPHszL7M/1YPFvWfM4bE
G+7PP3H9byPKzeEmXI5DKo2e738/mzUdW2hw8aRncaIbQa6ZL7IxIxvVc00d9p7Qju6IBa/uzjMy
H2mleJ5LeJ+XivNlmx0WDxKIZWAXZy/m3IdF16dXbS4x3vfhNK/sFjHBVMTn4NaZA4jbClUsoLRw
yvvz6Kkm/XBX+6fpujHS3nWHoMX0KIXROGokHxnUhpkCJODEkCBeXRNk0kqaGhSDzFNa45JbXsVk
lyZFT/g1w8HizV+yQjQe8DBagCbT88kEl++tu+iYQaTCV1cmEJNrdRlQJt8mKTEFfex9F/5kouwn
aJaDNMxK/RxVUwNTTXiJdTe/GwqPAev1jVyGHmCAeAcn+PIXVoet3oUjq0npzrlIQI+fCfwZwJjP
7urD68La2KRZTIb1oiN9uiAaMNeLf1r3SAYmBpq/MQN6yXvwsQvEq96louPKotgDqAsUyQyf1FsB
YbyaiSTwt+XoI9Of2rAMM/MVwPFzHvJioYg2lxJg1uuqiOtoTQYgKwJHZTIkmLUcO59nNtGD9X5X
x2mU7UHhoQl8mfcynrhACnSbDt11MmxBcq5R/z3z5O4Qoj5R99VaoSGpkBuGPQ6RxcuCPtgNkzkP
WwjFD5uzapTdzmQ3XZ7xX+2CloTc/8P0GrG0nJS9+e7lnPRMOR79mXaORQ1ilJqoZDX1bwifipmf
3s4ZgGyiUiFRkw49iSjDUeQ+G7JLjYCTzWk6w0WqAEYqVbbSNDXwKQTvpkE7zMToBD8TAZzMj7k0
tdX8sWXNTL2x6+4LKWcFkXAnlyImjZDMZBy0HMWq2OFsVC3DfCB9wPbwBYhmSg7Td6q35zIFevnl
C197Tik50NdTDqGbF03pypr60tuWdE37Slsyh7ZGl5UTKr3eVaLFM3Px+1kLcY8pyLnLcnhztBRQ
CixMerk2WQqwSL6yjVtlw+V9atqHSuHV327GqP65/XiUgAsLQp1uI2gnwSkIcWGF1Ggj4sJBQHYk
0QmD6HYkFtZ65fQ0KW6c3XJdtm9SBIcYH5nUYViwG/x3vP7X3WJ/imCrwcKHn1ZJ424SzhUC9x4h
JFezEjaIntu5WOMrHmN1SCIn4cp+UtLGAfY9nU9ggUj6lvSZ88lyqF6EEUc67/sA7bvpgv0RycrV
IYaaWsw0Ycvxq4SHjg+blWKxb5BAVU7iw+0V337lsfMKn+ToB2s+pi4kjalnW30u9GD3zr8geHl0
kE/sfxS+LgY3qkOBpqYakZOyRkiQz2YqJDOFmurJhRsDiRgEfOWPiTXg19og9VfMJy8vCmfgDKH3
fFcNQnbRPVihnCq4KTewsNzJWEMEyw49siSQ+O9rlh+NwLpxlPqSBM8HYWiUyeGTj5+IlWOiDACK
SMZS6DfWzbiyKrdWGUoHwSeNN5Rp0wEDsnA/w8UqIHh0jhKBaIU+9jr3jon+FmYRIzpdBJyQa3lf
8FzHQENzDAVUOOWCxaEl5sXw/J6oqPFd8OQhhgfqJpBxeozdadHFEbr/R3VJAQPBZ9ZWuaV1mw9Y
lhVPQPvgCXkTpaq7geazRl0BqLdeUiGks2ta9L5JchOrzEtoV12zP4GBoA61FibCq8zHwuPBX3gI
9mGJphWogwWPUcTGzAjH302m/6egkufxYOFkmqZyonIaPD2CW5kb4bHPpLhJ96uGnmd341h9uDK2
QoK9h417B241JecXghYpBk5RXhOwq/YjCbr7EL78KEzbIOrglBbjdzvoBUoQOjbFutiRJtg9b+Vq
Y04I9Xt8Zr3aEhfMspw3AR5OdQ+R0WWTSGfCbJGzQWWfVHAVCZ0XcwpGu2mBSWc94+GRpfH7PGu5
aRvDcmN2BBtadyDXImMlxtApbBSTRJeOsD/1q3vgAmdi3rVBXAllYNbL6POC6s/viq/ELb0SISfo
U3Bj6F1cnBYrxxg1Efc86z5ByvUzyqkYd1VCCezrz5B3EGTFuH75OUZfp4PdrlFDyXDGGx/hVuMf
+9c3PHlMZ5z6vGCvgsxfLtycxTN9Mrnv+YFiwmiPPpKrKpW1WGJydiYDUZUZrX25ci5I3Sdm2z48
Al/bvlM3ps42aCMzi9Ajo9CC8GzMsBTdlVF4/hUAe6wYRULKoGTWeCDW/9pq90r2KxLfGijcjbqt
X8j9ubuntmCQcBMQvCrfAyVfXWRQITcFamzut5o7L+Qh3B0M7NYwhg/W+ZT6geUaqlrIUoTdliCU
w4H/u2+e3YDnvS8wTtAPwztXBmvWwAIlH7EyQoPIiTG0REEHxDdl62m3rIPkYaxYVdBUF3I528Vw
Z8KoscXltDVEZjqTzLV6o8PoPqYGx2oRSECx4l4Da1qw4wA7/d2WgXlUIO3JVVrXY4g510LIKK/Y
mqXOWgvCDpA0d+Fcs4KPrDT9gk8sTYxk0v5H9FJlWmRxP02wQDNLm+UC/APmahNz4vu9T7ZM0CWn
ahSPylP6D4pnNzQqo5ghIOpHnV3X1pNdonoWrtrD+7XjflbOWWNYr4pnmGY74qEKsUkACFB+yNp5
EpKeKvZrpGcpMEHzqTHEIOwWikO1cH1bivMEF/dugK4QdYlxo2t0oVEIM59u+zQApntT9ZAt2SI2
kPMoQE0LaHDZ6637sW9IgotC2Np1f5ypbnmmM8reBurmfDyerXj+C7uagHUt3b9UrWOgSKSazKB6
lcctkqI1HzMNQd7W4ClAJhKnIX6NAXjsOFUr/YxhEQF06/eubwIaPk2XOgp6DWjIIF/jYn5HAHFX
RpMmI+5XbAIUPeZ9AieMRxE0xOw7YPKIJyM/kXmwrx2/jCw4aOmlnT299YN7XbyVTczwshrYN3G4
NOoNHuevmyYCSLy8bIXKKjc+QlquIT4eQWChthwp5/2oQRPPpaDN2LCrzEJC/jerylm402y3nchE
YZAPipfECldQw9Aq5XnTccmdpqSUY0WRvbL07Oz3JbgeH4dqt/5OxhO0zASZPZUOLVCW1gIF4fXa
7XbIVCo+MpCI0rX1OO0i53Vs9+50tlrrvCmndLkDiH8Cx4aNOU4PpNNqsfJ/Hc+TESHm62rg1IbO
q9ioECbNV3qzql4JyLsNyhNfGKzOXmhBiBvp8lsrl66dYU3k64mrXC8s0POso7J1bXiKColKH/V/
j2DPYm0e+1p3bLaFKW4Qf/K/7xwbBm1VpBvDILzd8A+qqcgwB3RgkR38qCUPrCsOg6dRilsbIGwc
7EaVSaSRsuWBewLLe8UnHzoJIuDn1DT9f6EMIk6r6vdNvkby7TUL1mUbfZmKMLOat7H9PbAmb/IU
3Y7Ze2EUlObJerrBBZCsJ6vaTk5GLz3eTHmgNSt465NM8lzXj7zeptqppDPjGzZvdWvJZu3EIjgG
OdyhApDaTJAY+jH8xLOYEXXvSFfhdWdMIQhHGTyeRzxpplDsRy4y/66z73odo/++NnwfiZgOE7po
T3LbTD4wwRpTFKngeFTx60yKeRouIICZuFD2X1OYESqAHzI149VqJyR4bO5YqJ4q5iBnbDKxIg4m
MfrEWiDRyhmftBfOrqHLDUwlI/0Of4Rtq5MFV8Hkf4PPNjICO3i1SO6zpbviA6rxGsFNVE/4Ttv2
85u3Zh9a3N+w1gpMR+EUeWYNTZGc8QYsnSksgiQJlxXpj4iMkBix4VyHU4jDFeM1JywaHaVVyl1G
ixsNkzplqp3dw60MFvebAM7PipnNa3fXCfkE0gm50p9Oq0rouaRDo6/5NUVEHLPBMVh8i3XgFErr
tS6PPx6F43u3CNDXi7Uxn4MpAQZP07RDt65G2sPdIKwCcVmYAm0CWNGYohzra3o5EBBLXORo+Qb9
UTJlgUTlLipwi1ofJkDGxHyoQdGCAkjmefTbB0MQF4WIp/CBghSsSV41c5WN4ufLJBi9iUdsoeAI
o3YAM7I5T8JbExai7pnAlaWFMQAeuCrlOR5ZXHCeavz5Im1EUZOdKpbfoaSfYYtpQm17VDflio0m
p+JLFyQe8QOOzG4bmIzetK7P9Dcg7LtejFuby0MVDOx8bk01ImuqUrLRrcGHw1LFEwgHwRx1TYDe
Ofgxuz0lW+Jg63T0mgEDL4Y6+mr2HOFEgUYmCMNY8wlLyha5zbtcc3UmLKJq9r4utgcX7I7K6omP
dyUuUA9OKs7ZV7bu7IdyEOepKb1tXsPVWuPikxdIAcffo0R3jH01zkLxCo6huW47uY9c5T4dwSO2
Uch5mbWwiJqhkFCnH/129kKCUfDNz+FkouIxMy8zuJImmTsttd/98jHBAY0cUduN3Nn0DrUydAuZ
Qi1h79ggw6Mg0AwEgG/kIN2tx3ZS6JSPPlhtpWDQ2IA9eq2kMIyYu/oBzsMSlOpeUwZtQJdS67si
d2d05ZzVx9SkAjoBwz3EQm1xZtEAZO9grmN0QH8o1Sov2S7bifjT62ZLIM8GQF75IKNT+jJVQsgs
Ma1CMb4hoWHhS8Cw0MFkKLVg5TxVPxEUl8d/8B9VwLRysx/jCzruvi4j6ktgQA1Zeo8Qvai0m+U1
VRTN5kGDhQ6qE6ZdUxmor25D3uxcWze0zl7B4Pqu2RMBe1aDfCMA6QSMdVDgwk4uYHrmwz503NS+
bhSDX0ifMBucffNdz8bjP7A1SDEW9ihLYMzuKmQP9NjsEvg/RAvbHFEfiLpS0Xe/Z456mtMfJS1j
pYnHYu7gcx0psuPfk7w2792OPL/rhP0tqhqLDmRNY5FV7F4lMgtrlNnQU29IWX8MMY4oUv/UtID8
HUVYQIbiEImw9U7gCcUBg2nPWdI0d3g82X9BU9Eu10Dm+8mXj9511jxRzjLYRHa8IS4tdaogBtJd
o6wBjtntSe8WPyiI+8yKcBEVIfxbWbIAo1GIf7lCO/FuNsqora335PhI9oJ09630NlJoS4ykX5ym
efbeqB2dr5IvnhlW+FP56Z6lSIqEiyjuJsXE3ENhkoZDv2k5nDiY6WywF9eqwKDYpj3zk/6ZKpP2
sPyA4GllbXrDOM7EUGLTkOVhbNuTlU0zNVnvyc2l1TAZJJbo+F9aqTp0Px/D84JGCIBGtQs1PEfF
0ig8mXUXkqNGGWrzCzYzAwAd7CJl3qM6sKK46KTBFppu4Mh+ZvGyjw4b4SPWXRA9itXchXLhoiza
27xVHleSbCufHxCS0tY2hf1/B74aUTMS8YJiMCok/F7hgxroZ4fv5kajfOunCalKycAcI11do5ZD
c75qSyIgmR5DnSjTB3i5yzjsYtP0ACRIl8QRnsFgeRP5MhfjiDzl3F0zBvmAsJsYhFD7anBMMNL0
/HbXppzCKfv9wmwAy18jdIQsv3jku0hPcxDFgB1MCKLFVgcQkURdkfuxcnWxIVqWo3e+uPrP5TAl
Ql8R90Q00tm92BoSF10RjzVs2xd38sOGyeOOaqXabhyDwOq22vd7vHbfwAonGff8Nrpu7f2H7yc2
wMIbO4OH8XLckwMh/PWWE0wym+m4fXJvn0s/JVzTcMIniEYq6Zbh/jCTwB1noTxWQHBqwYdaBDN0
tAoTEQ3a0/yI7pvOCzACYfG1qEgn04L/ZCyYJrwxPnelp//IlMcuyWh+PM6jTXKYHFphIMl2zPu4
ibZEdTapIdjG7KM1/P6pxJ90FGn1qjHDdw4VGAYgyu81WH94j6seyAUOjwRUpBETVQcVTERZDHPa
T5VhAiqP0pq01qRHPTD2pSvvu5V40PSvnI8gzJ6aZu0rBTyUT4FWG9kA7nq3+zjzYwLrT+FSiDNt
wZKc6JEje7aMuBCUaG/8tWAOyU+ZRbEvSe+j9QlLOk5QkK03fIDPHtuX7+JOcPiWTXNU+T+1l4lB
2/EPGKF4wv7RRbJOeKZ0l8eS1FiB+2zgpgsjW+kCHy4Du3neAAGr6DPP5+x5GUYeVkM5tOLkDe0Z
AbZTkI1Yb+batmoAnmFrMg0iQsneGdhWop3PBs/5YxGt4n/7tVMv6ZMT3aOr/YX4hXJVIzeAbIZQ
LdDfpv0vbST0rjme9Cfik/+AduD6eV07CjGVrq3TYP+atahUdGOyOQVBTUc3dcmj4red1is2SRqk
oIszjShjNEVBDGYNZb73g0wAymZbM7S8DeR+Vuowai5d9ci+DUHflXFOCjZ0PbRaA/dG9Ohnvfwu
tZHFk04ju1fn+RxyWbllNW9FWcD/pwNVyTCYL4PEhjOhxUkqagRNu8bHgToK3L1bP3w592VUCc96
phw+4TmT/iX9WcyZK00CC9F0w+z7XRRyVjxY4MSTQmZcUDzT6Slv8EyyXxP8ChTsQa0laHEx2OLn
O7Pez8987CPbE5YMW95D+LqJwsoIVJuy9XZKYhG0ScEKpOn0n6u8jnLUilyCD5N60/eU8eola9Lh
TO+FdCzP3hMI/SLNF0l5oBiCAWPV34/+RD9huMwNrrdExbBrvpNHhlnqquG/mR4HIgQztduUonzy
/g6lqJZ7vEAfi2FOAagbYuy9V99zinN8rG2BZHhrL6ucfFr/aAOFCBcjtXp0ukoGO/K9sPgAkfRV
WHWZsrI5K3xjKQYeL/xjTQyTPG+b/OinXFwrdWbWTPbztcr8MGS0SX5lb9nqjAyqzHpDP3XPUeqi
Vdpk2FQiJJP+0/roPzKSvTG/csm4YoszNmkHfFkuBL2tXZiCJAraRtgga6AMo5ubcRnwnxO/mkHx
+0goyTsrgdDaZ3tLOEFPKeYPtw85tbFV1y1AfyDZ1x5d6hKkk0Dz0M+rX7XxlcAUaB8uO6RsjrXg
3sRAka/WYqU12/2wn+PPydQsdwxuAvUP6YjysrLi+/J3XUGB6V/6OgwJ5Umda3Xt5hpknq3BrWzG
IErOYtnAblKItQF6pW+f2i+8+YHHxzBXs896vEO3HWm+074GGJSfu09x5uLoQXzHueOEZ+QXKJpO
+VzYL6qo1rxRkpoQGQ1R0kxEot3PSyGPJOFZkI0VU4wX92quyndYtkhY3Dtl6mDrHap3EE0Lt8FI
eUnTTVLBZYB1IaaEoZvb8vOfZW3nATpidpJS4vRYPiKIeqDYGRot0u96mbvaBHhtzhZJ3vsOgsUo
symsVnjJVD3gC5b1DWZa3TyHSEvcPgNiJipZCk1Xz5MWNMRPF6fSg0FKVzFJkHtq0gx0fO8BnMW+
Mewb1J92ryravJc8r5K6wlCc29MRZwbHV1CmUEX6wpBSG+QIZeqTe9NOrNvT/vKD5IFY6f3tigPG
mdnHyBvZbMObmXDRHk0/dVU4kn4CWeU7ZRFJLkaFQLV97r1iiSzrZZK/U85eviROPnwyzB6CU4v+
I8JPlGBUjqYFFSzRqrVEUv1CQp6CutA+1PgWNGZIhrOAp4wkkiRTTWGIQ1gXMyFJq16UJE2UmvS1
dUVJ8wecgk3ejyw79MaYJ0Rm2gC9F4vFbesZuZIErao4GWLC+u9fk8JDRv4z1GhR4ZNowUzBe+u1
Vxpq0yU/WyshqMOK5vkHX6qIG+1FuXPy7WOfm8gjo5imA8mCT2bK6WaqJsPgyodag2dsQH9Npn9x
lbGxP717MHeFXeBMZpoz3Ptj9PMOPJ7LPb5OYUBSSe67YAwtoeW7qJnZrjwhQW65LzpX4xDxYLeI
0RbYs6uHLs4yNLudXeBVvwZsCq2KDxtCJOsFvx40tTNQmsOdh4sNX1MC3RoLR1n+G3PDP1ei8GA4
Im5nMrCjHZIkNYRbF4NheAZLpsFEA3xV0nFdvW+VhelQekZmepi2R4KeWB0ii2U2TqUEt5Rdi7ko
PjfszJMF/rKoQyeJrMdex+bfc7x1jRRBENbtyrDDfWiywwVJhhP6K5Z7MNYVIGb0tESPbJNi1w7L
hM6DGsCNOL0Dtr2r7G+x1v6AeoMSkX7pQsoN7ZJ5jWoHqZqFNMsDSM4ZTUzE5HxLeH6AqtyXnVEj
+pbBdi+BTgzo5uImx4rlaQYDt71k5U/3ePqFffq1AHlY3AqiY+9AgfvRTzkr/cd4JQdhWvQu2SHD
QK2D2yMyDmO5a3XIlyNrkzJeHkq54JrsWETGaPqskkQYm+p4LnUUdOx2AvsRgrpPcCzWn+nyCZnu
1qIhJ43C30a7DgVF9A4CicScUGZmXl9lCzuUOHq/S2VO4/9dJItdyErgBVez2CkHxNmlBgbhq4J5
uJakw87NZ2kCCxEjoG2vhbjJyj33b2LPMl9c2eroLmbfya8inommhH57pFU+CNORH0EA3VNlT+4I
qdPWA1ZVgZxpkzxio/NR28DRLvT776jJeiQBOpzgI131girjR5SnRHANGYmJx4UscXZDYx8uqV8z
LzUxM6SvV2i++R9PIbBKLfHYnRjLpb0g+Tr/62bBMMPF3yYcePNSS28zHgMZiciVOmp8Xylc70y/
3G0nsFa3syeAPfsJW5nxaYv26BQXyskeOBL4/Rbs6NqWsaCjf7dmRMlIRXxtoH7b7oaEgKUxwBC0
O9GKVRHkFHj24/97f9zt9aYzolX5zjOuoLBjvBXMwHy1B4t/LM2DRuw8yZgt6AbkRR0wn8KntNLV
zf7AvoX2+Wb1jPHIQaCNppwmIvqqC5ipARkisIFa5UxAi4suARVOYKgnGNONwZgKIx6rhUJcpzg9
V0sjywmFtxyxa87sJJYwFSH2nGRogNojJmPfIre0BNgUrVnvE98zdHnqruZHS6UhOOTnBzQU0Chg
iRL00TzyKXjfRHBFobfr1vCpMczuUG4wqxmCgaSpGTDlsHRoTQRbVRvnRBis4Z9xp/pF0/edChmm
DJXbpL1ySuBIPNm7E8RiF793dDANq7aFKl5goOVzr/G+2mYmw4zr4OQYKySxljoUp6Gj1TDFewTk
ZNI=
`protect end_protected
