��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�2V��QV-�T2���A.RZ�6�-�β�vJRI>�O9Fun��#�2���]������ Y����������B��^ /�����T!���iTGL��=��������MiO���>��XSP��*���M�D����������"b��naS�c��ӥ�<4f��D
y,c����EZ���[S/5y��*���L]����՝��7������Γ찃q s4]͛����u�\�ވ~$���GV7��T���9pY_�v���%���hjf��x���b��8&l�?D��Ð�Z�V�r}�����]�] m���d��^#�����$��'��@�JT�w����=�G�j"C�c��JцRW���?{�ۗ��-��\��o��/2�"ĶA�HBj�S~���u�����S�"&�X��<�tkLj�[UKg2��[��-�q`�Op�Z\Z��U����Tw��/8����v7�F�V��9��w�*�D\Im|+���N�I:��v3�N!���(�?O5��ab�i����Lw����u硃#�ȁ�J�F�2�����!PlP�d��9�T{	�L��{�U|��M���	F&OޠL��ÆiR�)M9;��%څo���5�&/y�x	J.���#�z�c|���g�0�oxqʹy`�PBLJ�+��h�oKB+.��-�;Ԯ�:Ԍ�:�#K�z��c�M�w���:�eXY�0R����bj�5�_t�{j�_�=s}@�,=�&v��u^��t�A��Ȉ�7�ƛ�����E	h>z� ��h����q���'�D��63ЖY]�w�����ݷ���.�6�e�/�<��YO�+�B��ﯞ/�)�(�ґS߮�G����0��i�f�\a7��|���x ����)0��л[�|
B��E��BaT%o��O�[m���0�nj�IF+=s�Z�|7ꕧȊ��֬������9h�T/������W�c  �eo���p�����%�D�qb\�k����P�K�Ƕ2 �n�B�KP&�ڽ�@I8��aR�Vq�p�Y{�:��F�S�j����������{'z���{$�w�U���~�ey��*T6��&��c ƨv�7æ޿�(/xǷMG��VPLl��u���G&�n� ��_�����hUe�Z�k[�o;��i5����q+���+��K]�O �����a}�RǼ��,oMh�%�DN���	f,+P��ZH�`�?�m4U?��}-�y����d�2Ǡڕma1`�Q��Z9M���=���ƇK�{�f�P���q�L.`$�&�s'jC��cz�X���t�Ql-n���r!��d�*r�3�����4Kt�O5/��W@��MQ����U���@�:>�� a5SR��L(1�|��T̷�@���V����fᗸil�"���V�*n��P/+���fT=���^������O͛��J�o2�鞿���;K�O�ݓi�rT��AR�o�'�r�zx�,�a��C�0�Q��cw���ˊ��#;.�'�����M躇�Ƀ}���t/L
ö���;W�� �;-�h�Vf5����ʙA:S���#(.1�1ǧ�{N%<vir��P��p�O;-��%6^QF�G�4� և̠Ss6_/9>`E�Z��'^ꀌd;>���vX����#�f�(Oێ�)W*&�VNӲ�B{�u��N�LRr�1�ޔ�����b=�|۷�X��a���|��F���wRW�>&ߓ?�����{����v]ﵩ`v�ަ�D�~ɏ�v� i�����7S�����\�%����3^0�Ən^Ù�S5m9�4HY�Ӎ�<�L��h��Rnw����>�j�N���&���Wj����3C�}86!.���1��MN�ph�����Qq �>>u�ʳ��Q�S�L�E~T�F�0���y&���j�L|9u /I<���5��K� .�٦�u>"Þ^R;Z�e���qTU�J��S�¡ ����@�	��V���l'v~>t��ʵ]��ݏ��r;�À�Ń��%wkف{�����L�+И��ءgS�}�&����Z�z����Ј?eP0/c� ���R��Ŝ�̌��E�j�0��
x�$�ΞQ��(�k�{b1Zi��@�\��6��e�q����V���[�i�xs;�Z�z�������	�ke������t�iZv ������m,X�=��@ ��\
*��$����>P�������Θ@�]��>ⓓ#���D�����t�
���,�W�e���V�̝�K��	nޥ���:8�*&$�CǄ�
��/�?�V[9�^obp�k�
��<K��`�%�,�_]���'J�O�l��~�Ĕ��m�=V8���(B�n�ߓs��2ώZ�a��f_�+}���t;o*�1	��5�ӛƥ�7�[nM<��A	H@l 6<��o3�|�ʐ`{�Nc��p���}GYЃ�������[qo]�)f߆�$y&�kY�2��j�G2|�zt�}�O"�\�<��O�C�� R��H���	?GB�P����$h4���q��ī|6CZa����:��ʔFt���0���OP���]N��=��z[�v,���?�Ǧ��YܕC�*��?��Ϝꈕn�h`a~ߌ;�2�:Xҩ��ל���n4-�yv�\�Q��D㙣����Ҝ)�(�=�' 86!L=�����#W��[ƪ�iW�*9��RRA��}�@q߉����z���2����SQ��t����b��z�s>���Yh�/�O�(�'N"CV�	\7�.ލ�$��ѫ����泏��We:N�<��O��|�-�_u����WC���	�r�s��vP޾vl1RS�����}�u�Qڨ�^"�J��4.o��2�9���kߝ�Ԋs��#%�b�	��UwRKҷ�G�4Q1��� �=�ɟ��ɑy�c�؋!�m݃"���)��;��U�/����QrԔtdf7�L'Q1��n<��џ���a���2�a�	��ު|c`kg�|�
���Q�=�o��S�$���I�7�y�l�3����8�Q���C���� K��6@�W*ۏ� � ��΄N{�]���"���OD%/��'�Ϡo�H��N��$�uS�:��$
��|L|��<�ٱ��JG���K!��I̿rtL����d����Z��lV��y"��zH鉤��PP0���5$MَE��=�@��< ;�4���mԜ&�x��<F rۋ�(a~����X���6IGΡj�:b��F�8��ܘ]��Y�:��i[�Nz?��� ���l̞��@c:��]ۗk-I��:(�?C��O�0���A��y��ŕ(R���5F��{@AEk�ju���zE��
+*W������YmF�}��(G��F*M^;6�T|�=���2&@��sV��|w��KI'[�&r���)���:D�,k��`����~�q���v�˔t�t$�c�A#o����<QOM��L����o�_����ǃ߹~v9������#^��;���lzs�a�S�1�B����b���*�^���ԅU,�Z:��5>R��D��Ϛ��T+ ��N�YY��U���8[Tt��l��X��p�{�25�@�nL�R�N��kd��[vu^����VT.@�L�Am�.�&���%:�����_�T!G����u?�`g����e�z0mϓ.����nl�>gI���c��tm���⢌�~l�!�ĬR��H�Bʾ���7�0y޵l�����	_��N���гE� ��j� z��M3c=�p0�|��D{���2甃��i��fMi��R�:䫀��e���6��S�a���^��]�|"QK�h/�]Oy���Ka��G���Td�rp�p�#_�|�ن-�@�%�Ⓞ�����պdc'�1�i�k�\R�k�=z��'�ݷ1�,u%L�4m����}�ˠ�"�1��!�I��[Eҿh	�Ex?���=���Ya���p�L��)��PI����Y�WQ���*jJ�<j�%44�gEJ3�0�M�����<������Fo|j��`k�e�wR�H�J�1?���H�Tx|�˓�@�M�L��\)��&W���K���k��{-�"H�����s�p֦�^�Ԇ&�	��8�ein٦M4��ء��f�S�>���;��[��`���w�z�K$�^�?�8�:}����CgE�w�tLӭDp�I�7�i��(��:���A��7c��N��|;������|Bf������� �VY	%GW�� ��#�����B*�㯌A�e�F�@Ft�W��8lQt&4�,qo�N�D2f�.gҶk���q�$fZ��4'5:>q�m�s��aa�5C��mN�Ca�"�����{3��m � �m� �A�=�K�"�9g�w'&x�Lg�H7X¸��R|b��x����C��ǻ�˗�P�'zK�̀+P	�F�x��@�W�1�nj�j�Z?vt�O��ey��;Nj:�#Z-�7��
��nH_���b_�y�aO��}J��⺌�&dWAH{�v�b��K6�H���{+�8��J�[�	�֘j��,*�K�>�.Ɏ杌1�������-@l��� A�U a�$�e��X��!�f�
���S 26���Sw�j�l�͐�D$�'�~�����\tm
b��^�R�㗑�I��X'ה0Rm}_O6#B�_��$�t�<��
]��
L�+�߭����,������'���?�W2�V}}�ѹ�E�6Nc��k�/j�A����{�%x�/U�3
h��p���$���&Gk�<)�A��y�f[��D�W�gm��1��� ���(���ŕ�!�P_ɻ�>q&��% ���hY"��d׏��΀�
U�Χ90����+��G�Ռ��Գ�^^�!�\vYi�}�tE%��a��ݧ&��d�=����6��^:Θ0��:p��pd:P����
�����oY]Ba�� �c����!K	N����T�'>ʩ!0(;�] ��3�Z�q�~ކ���*rnR)'H��ߩ����"gD��`��.�yɘO�(l��LQ��P��f��$�x�ηXi%w4�R=�n�Eխv�<���:Go���3)�����E�r�$�ȵ0`�
)��Ć���⾴6���*�eMv0LO"KaL���o�� K��ef*=����@,x�[�L��������\�d�b�D��p��Ī�$�z���yu=��K��Ǥg���	�����֌O'>7`��K�D���b����R=UɁt����m^/�! S�em?�fS���9��}�[�\_�֙?�LY�~G[���������UM(�R`�җ;"JMl��a�N�m|h�~�Q>�����iE�L���h�ul�R����X�t�u��IA����\�F�>^�#-�!�"n��Ɗ<�b��hwO����l��7�J��,J�M��������dWW�]M	"ˊ�b$����iݗ*;p �bq�qM��ʰ���(������!�)M�9�ÇlI��T�msC�ޝs�7׉3���%Մ*lA�Mh\�э\M�o�7��Ѕ�!Ӄq��K-�SY� ��7��N8k��+o��u�o)p<����J��Y.�����!�@_2��"���ˣp��^��	�X���{ru��-�H}LQ�	D�6�Λ�3=ɴTC�09�J��b�Aiv�c�}E�ލ�ns�C�ѽ~#<$�A�4�.�"�&�W��Ս�,s;O��;��o	�W�r�򑙿)��6�|7�o:>aG���7���'�Q�Z1-yd�/`ڱ������a޼�2��� #��w)�m̜Dr齅Y��O:���8u��
o��g���H��"�!�x�bzl?�I�s��,�R7R�� ����4�P2��,�,.�7nik� �����s=T�긖a���J.��FwfaQᴓ��*9R��`��xϯ�km����DI9=�4#��K�8Lۋr*LI�+L�|D��}t_�?lM )o��,�c��"�Q�$�0Y��~@W�E���p�>U}�ƹ�%RF��U�QAO��ɫq�%��h�-�f́ X\ko����L��a+���� ȝ1'��S{Z� ��=B�L�&�x��y�r�PG�)�S�adq�m��6�G��m�yF�%��@�=��.Pփ4A��S�M�:�O	[)�[N("GVr�bp���x��S,4 0���G`�Cs�b94��[���Q&��}�#����̉�!����{bI�	E�ES�C� �f����M�*���ͧ�1o2�B�m-@;��}�>n''�&Ӎ~�C
qO�?p�I�?ZRX�+O~�\\V��\�A����^�ͅtI��<����d���VB<���M�t-�?�5'�
�Y���pi6&��z�<��~,�<D?�b!��DJ��@�b��&b�/���|�sk����3��樏�j(�{뱆fA����J��@��{�tc�6Z?q��u�%3��\7%�#SF�r�D�S͚Չl-�D�X��X�}"Wۮ��g��8�C0�x�_ʕ'����S���?:����|�k�Fqn���
�{q��;�gTu���ꔽ���|��h�Ik�t\���*O+�-�Бc��M�7��k�dzhS��7B�ҿt�vr�]��q��w�0d��b�̺�L�Δ>��ۋ2�^xQ�kl��$���W;��
2w���t�����D7 .z����A�d�m�������b�g��S��[�j�$��ر�ǙK߲�_�/���/��g�!���8m6=4%�R9pu��\V�8��=sr'CN�������+���L,m�α*k)����O]����rėh�'�ũ�C�S?� �9Avm���`�8N�nz����[���f�l����4�]N�ʴ�Þ����� ֆ�K�Y�������`���a@���z���
�s-��}EѲ�.��c��Z�����ār���l��?�b��e�r��b	r���Y�� �Z�]���
��ڤ�~����r �jT��k�ݶ�Z��*G{�d�w�6's.= c�s�Mx��ix'�J�A �qzFK�8�����Ľ��5�e%g3�(�(J��K��ua
�w�������>�B�b��3 RlI��=����9;���կ���J7�~S�s�W~�-���Jڱ�%l�:�{�QYkҌ�g>/0J�~B�/��ʿ<{�p��L
>��<x���l�#�I�z̑:�ˌ�����H�-���_��UL�H�$��M��5�̄�s��r����I[yY�G���%N��m�,E�>�4��h�&�^��v�L�*^��{%����,�>�1�,/ d�������&쵩�"Ú6���5߅��0Φ ʬ�0b�_��پM�Y�2����AamF����}BY%:�E[H�/�<׻���	Lk5u@�v7(ӡ�~���Y@���f}�.��� �f�x�b%���O0�Z�������nh5q"���{��j	"w�X6
�Ce���_{}�&��sq�Z��E����.��g�P�i�4�Up�����R��R�*�!?�8���q�@=����x�"�P�e�K�#~���Ɖ�o9��6vT���AD��W�N����E�#HcL������z8�f��-J7�c�*��#S ����-[�����*qQ�Dc*�a)�6н<�qz�~  O�Wj�Ր*��;Jh��_��0�Kr`���h��34��j���)(����,5dC��N����޽�K�h��c��H&�)�fv�ݺ:גv��gîd�H*yv�7d���W�e K�Jk�m� ��x"k7OU��G�������6 d�1_(��d�Q��[/��6<�Kr�2nB�l��tIkx#�����2��K�3n��41Ӎ��m��\jW�����1BuXuSǭ�����&�ƫ��4i��f���<R��KB�$��C��:���HO.� �;F���2xq'|�
j@��}�=@4L6餳��R_@r�$�kpIQ�3�n;��k��U�mGh��K����e���m0��
Z9dj�87K�����b�}�Z�/��J�%z�_UW�^�2�=��=��&�8��Y����OQGO��0Pnwo�]+]��P��X�lN^G%��dO�?�o��ڋ��W=�	�w)�pR���-A�T�Ae~z�*����Yc��
���Txۂ��4r�[���H�2N)~W�7��D�X�����u��W���<�.�J=�\�<\�6g+ñ6X(9e�>i�bl���J�%���!��șT_�� ���'�~�D�1�W��a�<E�1vy���3�?��(���t��+O�6��s��f{ds��������X%�\�]q~hC�MrK-�H6��N<������"|rUc����!ofK���?��"�+f��]�I��C#k�rْ�Ho����������'�2@��%��b�:ʟ]��shӉB��XS� �9�a�.
��Lk��g��ai�ރsമ��U�"au\���ä����x�(�Ǡ���W�q�ނ>}5]��j	2���ˍ�T��)Ǵ|�@mV��_FS��m��g�B�K��$ry�ʔ�kYֵ_r����#Aב����*�2H��#�Q����(�(����z�t�7��֏��P�x$hl[w��FM�4C�][��eB�[v�W�!4AbҤp#��y��������Y����4�Vh>�2.�SW�����`��C�+�!� ݣ�Y;Aہ:݄�1�R��F���8�Us 8=[��~�朚�V>��0��?#�}�!K��N��JB�����K�c�nK�/�h�!��["���z�s�+�j��f�m�a�<]��p����~�K�a0�87�x9��,��F=�;N���/	L����|P�ףƜ���P�9������y���c� ���B˦<;%ާTC��I�ƪB�U���3E���;�}>���fگ�b`���7��|_
HVv�L� M�����B+0w�բ��9�N%��h�(�������E���"�|�k���m� 5�q���f[�cs�4�O�,�y��硟Q�Q��v�-��# Z�吪�0]��4����i�t9ZU�8��:X����OM�IY��[��C��p)q�����8#R�a#�,Dn���&Zy{�x�����pQ8{\F��6�.�8F���.Ԉ��	IȪ)k���k����Ko�^Hq7	pK�3�{�q�����*��ޏa��SE*�:�`�̽~�.���6ܤ���,AgW!3,���C��[S	_��*�g�d5 �zU�Ik�?��,��'���)t����!�$� R
S����$�AK[���g�(��*jJ.e�(�N=7���M������<0񎝡�ä��q- ���2G��&�]fjwW��q��>;��A�Jk�	V�����cz���z����Z��1�[܇�m��QNw���v��81HD�_0�*t4~��q��O���2�U�}�0{�6`�Kצ2��3������[as|�����w�?m���<<aw$� �/V 0�_�=�^�\��h�~��sK�,6�u1���^ۛ����*t�S�ę����_ԕJCEԙ��iRHič��e��F�x��N@ZY�{��!#_S�X:^��|(��:!x%�ʇ���6��lU�NRX�qa#tԄ�P�s(�{�%�ȧe%)RakR+�@�;�	��%-`e�]]f��
ᙃ`����������K�
o�D��[(b^����l!\�W[>�#�'4x
�H@L����j�s��z]!Qt�F�N*���D��\)V�2�U5�؍C�˔�������f<�ix#�l6 ���p��b���z��e$���֑�m��%8�YDW�@�
�9�3u��#2'A�.�E��p,��쿄ʊ©%�Od�ɑP�.��	�6 �
��K��@O���W6��4��c?�n�ða�rߏ�	�9�!��9�*�Y;ru�)�K�A���^��lt�4@p�;���F G�ԋ�c%-���.D�.ݕr.c������ﴖ���$WVD{Z�а�Q��a����1�!=7�v�ic]�#0�g����}g�W؅s