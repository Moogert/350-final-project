��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.hP�r~Jzܣ�JK��`�E^z H@��G�s5O���$u�ͫKe��f~HM���<��;��J};����Tn�+qs�Q��Ϫ5�JX��}�f`���C��k��{�]EǗ���g�٩���M(��f�$2|*�N��m�Y��J����7v?/^L���n �/-	�р�Ag�d�+	+�KcrLt��#�_��J�ڗ�g�$>��m<b����T��-	 �R�8�f˪�8b�N{���B<N�R�Ύ�) � V�Sx�Ʉ��%�x�yU�k �㐹}y�d��
�y����SM� x\C6My���d���ЁP|��d�Q�q��M~�=�������\�Qk���Nm�Y��tJ��`o5�?[�@�}�,��I<���m;�|�:DH����^-[']�c-=��C]���@���1IP�K��Y}l5�ɬ��cf.��֘y� �Y7[����W&k&y�)u. -w3u����-��n&����o�z幛��,��D}6�9�؝?�t
�b��7�"���}F�s2�p��������_�i/�i1Z���5Ш6�T���=��X��F �p�g(����y��"�S���c�T-����{LD�Q��R� I��M>cӶ�exĹk���<��
�a�d�֝��QZ����5��B���p��A%(���u��2���4V���㺆W�<5�"�*�٩��΁j�:_���|3[����n��)�9��1d����$��$�b�E����{ U��
xt�(5��/Ҝ_=�ᮕ�L��iQTF�H/�N���9���OtpReJ�#	�<������L2Ҏ�8,��
�Q+�F_5\9�|��a�T���U��[���
jaJ!o���=4ǐrNV�U.,ɜ�#��M�p��vT��`���v��G=4��82�M���'W�Wt��{��Rm�W�"z.D�R�T4�4;E�$���Dd�F�=�׷�_y��>���	1��H#6��ZmN��.��^���*A����i�Ov��[~�"sx�i�X�֋��3@P��I�R���t�@[����fV}�޵zN{���7�n ��Y��p�=�8�=�ꧨ�!h��oL'�D��Bd<�4�=�"Q?��=�����Zm��X���F�sYa�������ǥ$�[�&׺c��b!c.E�{jf���Kj9.Ɏ�o���х��x�����g���g�JHh)�|���>�W� �Ǆ�WbFQzf;�d�R�O2�Ƒ2�;����J�J���K�A����ݺӻ�~�1�aS��p�fMXda��D-���kiP�Y��hqȳ����Ԙ��$�uJ��8%�Sh5ٯNy�� 9�QQv !��W"�+�M�@W��e���S��{J@�7m����ԣ�zi���u';�`V����#V�1����}0,C
X��� cp>����Z�>c����ʱA���d���^��A���]C�DYJL�'
���Ai��5j��Ս����?�cp^t]]x�6����;"�ӪT��Ey�ɀ���W> ڃ Xm���2�	˜�� �Z��fʥ�"���f]����lfNy��ZG��!wp���J��Q��9��j~[����iK�P]�Sa�TF�����=FdT�
����;��YZa��77ND+�]'�7��?�VX�ΐ�w�S�_:�hH��y�%9��pP���*њT3��	+�P;M;O��Xx޳3�
�}<�K@�8lm1p�\����S:�(�>yh��3rջ��m����NdD�ʭM��E��*��
X����j�?���x��Q��<C��(�́E�4�p�w�Z�\��f���Rv��I����̜���m)wՔVt1�`i;T������,m#���a�n��)�eDF���&)4˒d�8���K��*Q�\���zkq{�z��v$�����_�y k\�����y�~� 6��Т�׀q�S���}�.IV(PU8i� �7�SK�7Hg׸�>*�!2��dL��羃Lʨ�t�>6��9DW&����oy�*c��3WEݟ�n�s;;���Y)�;n�2�l�.L����Q;J�)�KiL�"�c�ӱ�d�2��A��q�S�K�"�d�^����НU��?�t�d�cC��~�&iι�Q;إw��`*g�6�E��W;����x�1��
��%K����qJFS��-!�?����C��.��2s��Gto'�^01����*������!�u��z��#f��30�O]@�l��1�z�EE*6�zfN��53*�W����:7�9��M��,��O�a%�g�4��i�L�Εn���S{i�����gN��L�N��m`���g&���=�}9f��PBy�5V��u�H��3�fGP���թ�*��@�Cr�ِ�P8���W?�w�`����W�����HHXm�`�EQky|���87u�p�7����r�R\��t���9���������
�
��fjɪ��0� �1���#,�/��J��^�vє�Ј ��O����z��%����F�WI��_#����]��l���$�j��˻�7��-��vLj�l�-�� �t`�%��8l+D�?�R��"��A�l"�(����	�`(^U�y���k-�m��8FVP�v�Y��r�Jf}�t�0�A�VpH��ERẜ�W~��ŵ����%��GQ���2dr�`�U@~1�|_�n�i�d��TL�#tX�T-܇>@�Z�$R�po��<fZ'H�O��Ҋ\k��v9ZI �-+8��<F�,��e ��m�&w�sL'_7��=��?�j�٣I�? Ɣ�U@��x����~B�9sS3 ������E`r��[�z�=ws.�Q��(IK���;���;=M����C!"D����FK��(fn�_ڻ�
 &�~��,<Y�k��w��Cu7���f�[Ȏ�G&�o ����[�(�W��/��Z >�
0_C�N��Ģm�-U	�����&+O��D��^��TY�PY�lT�4�u�e;c{��u�>룧��u5l�Fc�e-�+o�y/���}v���9K=aoe�6mεO�p$�G��p�\B��M��'�Ȩ�W��hE�e@/_��������_D�Ha�<鱷f��f[�1�~�]uU�p������9�p�n'wk�?kcRB(:�`q�M�2�3�j2KBڇM�|�լmR������P�����]Nɠ4���j1�}�%�4��ra|AxvB�l�ѴJ�f���^j�.�7�ѓPV�O0���쿘��c�G����F���D5f��Ͼ���;��MH�F��x�ZP���B&d��]5�O3�-�����+Z��\ ����`�k"W�0��r���{�n[�>Dԉ�&�p������tK�ᙨKu���͕�#�ớ�A`�8���O󟠸�>"f��=�sY�o��/���� �������rգ�[$��(F"N�$*�%����ӛz�"����S��+����P��,Vr�m���Y�T�/:��М1�;�P �����_%� )�3���P��7��Խ��td����mk�/�i��PB��l(��C�C�N�D����q6|�����
}i�m�#W��Ä�|�\JG�T���݆2��5P��kjז����8m��'�E4+Ě��Ǘ����\��[@V^�iF_��~��9�:^<��v�F D
�60SP�����/�o���i������0�sD,ģ�NTޤ����
�)\�~9�������if��X�%�����l
�*�Q��E�-��:�eP,�p�?�ɕY�o�ǣ�	�.�9�_��O���z�v�u���2?|U��kVhN|��j9le7�x��i��drt�%W�5P��QD>�M�.Ye��������׬pp�H��P*E�|��)٠T����&�(���7�V8!��\<���!S.���2�=�M읂���#,�P�P0�TȪq`����d�#eIq��g��17��*#�wO�>�.�4�8�������|��"hI���|6�2˦�����^��x�ݼ�"vI/�Q�|�M��G�d����Fi5E���� >F%K�;�0�����CKTKJ�փ��3�D�ߋc����tL�p���tS8 ���zT�}਩��평]�CD�G́a�Rj�ҏ?��4����CXmJ��U@E�'T�'g���M5�
���'����ܥG�'\��Z�Վ�3��rW�
Ag�q�S�p9�����\d��[��3��W��,1 ٯ���(������N��I�o�kG������F`�t��87��E��N;���j5顰���˰��v��A���o�*��������K�&��Wj� ~��hªO�ôW�5�d0VJ��<o��$mӁ�@'oc�����*#�4�KF��Ɋ��ðn�{ux|s�J�w.[J�:O�7��$�N��qo���[����<HC���ڵVU��5���X�!ɋ������{N28�����xL�~:70C]\s��(�=B.K�`^��}^��,����Q<3��b�k���:	�>��h
B��<�Q'�YπS?��/�l(��+�B����oW�ͼ�$f�M�4sd��O�P�'Jv/R}���7Ƞ+�����n�1ЂK���p�y�[#x6i��W 6����Q�r?��i�a��F�q�8N'�>7��"T��)"-����D_��T�������g�e1�)��]�;�w�Pͪ��N X�dS��ݮ��;�wq�O=�uF�xoc�������Eo�5�4t�mT�id座5�o�7"�5�&9D�-�	�э�O���]�9zO���)��|�25A7]�� $�&�v~�t���*ːL�h��b���M��n��
r�緃�e,�1G���4��Q�=��D��3������kf�C��ն �R���������7���x���"��f�'w�#B�Y�N����9` S�Ph!jB�i�n�_*/�H$�İ9��������.�ь�Uv*9�10k{��N���k��<��d����"@o*Z��rn�]��D|�쬯��I���8���/���x���v��ҘI�v.�h�{2�������#��O�R��&���)���@�M�T��Fh_�ji��R�E��9�G$��e��8j	��\:ʷ�6�w�ph$`s$D��iE{sּ�P �^��Z^z�e�ٿ��<����XP@^��:5>���ԆF/��T��۟� ��p�h�;���p'J96��-Ĉ���������*�j/�NlIG��֫Fk��'�V����O���"���;s�֯��K�K���r\X�U�'�~������Y�7�yFA�mh��%ch�V-�	�w����	����j��:u)�σ��G�AAJ�q�XT�������
kW���+��7,�T�7x����Dg��ކ�;Ȇ�'g
�b�X��	���5�P�-�`{�3�
F"���������4K��w��v����3k�5���wC6oCLS���+.:yF�
��R��v��" V%>�UP�؞# � ���:i%�=/�rxʻ�o�'���绅
A�U�[t��p�C�8lMl��^��-�OX�t�*ڱ4�ū�4���$�j������!���>2�N��d���{�A܁&P:�����f�����G����t��S��!j��A:]g�z������;��}4���W��pK.�7�YÀ�'���ڈ=6=�s�H�$�����=���jOǥ��48
{��z�vpS�|}�=aj�k�i��XH��%h�b��2�B"fZ�c�m�N���dA������,&lti��F�n��S#�p��R쌗����dCy�dXl��Lor��\96k���j���^�1�)�W�Dʳ�D�	�L�u�_̧\�lF�p��7�(g�AWe�
ޮ����և�;آ{�-���z�H稞D��������u1��ΪM�?Y��%����N��hDl���v/�K!O��~��ZmS�m�CW�ig��eG"L��l��U������WXEWḘ��f�EN�!��7�ʘ,6����A����+k�mB�w�M�8< ]��HM_���j�ir��CΨ�GSQ�Cz	��/9Wk��ʲ��P}�J�,y��ky�q5Aiz&�fv��c�"�k�T�+�J<1�D^��}��.K��#N��&�eRfcp+S��a��I���x�o����$���7�-x.K��k��o}L���>����eej�̴�W�J�bnW�U�G���Y��m�	�g�
хI{Q��l��QNQ:�G�؜x��ʋq
�� #�u�����S)�h��<�J�`���8>�q����Q���y��K�b������]�r,�gdw�5�6���}m]����b��3�����ӊgu����7��*:r�$��+����{פ�f,¥2ޒ�|v"E�<Ik
X��`F�֐1C�����Z7k�C';{�-��q�#%��4}5��K�I~�i��/�y{�4�3�
��?~�jM:�}Hu�����L�x�7�YП� Ω���{��⾥*���;F6s)�q�ɫ�=x��1��=���¡�Du��V�+WI�!�X����0�\A%ʗ�"she$	�sh�fd��Ln} R^HȞ8Y��\��J�$�U'�y�ʓr�G�~g��� �+AO����}-��1�`M�y�~���%�˼oP�,�n�h(W7�~T/���[��g$k���@&����}@U��u��k@^��tTIn����la���<^��0�r��$��� <���^2�F�7O������BD�HMæ!T�����4W��}q�b6!���	���t/��)V��݂'L�^n���ݴ"�ۻN�����J�s)ca�^�M|���vttt�!O�Jվl�om��I�]`V��DrJ-��d�ϼ)���99E�*���60���8����1.k��ʭ���l��`�~��3N�ނ �/z�/T<C_�U2
$cN��c\p3� �A2j���Q��
5]�o�i��c�r����c|�ӥ��vY ����i��FzO����Ѵڋ�F��I"����'�z��>l�p���d0*"��Md�>*v��&�#�Q'�59�>�=����4��C��[�խ�Ӗ��� ��XM��D��#���Tq)	F����:_�_k���)e��S�:���\��*3�b@�z��ZT�':@W@?�իd]9u���]�l~͕d��PkVÛ�2@�e�XNX���z�s�C��?{�j� Q���k�{�o�r嶗�U8.K�41�����g�;8h�o6[8�Ĵ�,E�Z�w�,������h�G���}r?v�cFjrc����g#tx5!�}v��"k�?�G�l�l݄����k�'5RW��� ��d�p��3ɿ���-�
�f
�- �F���T��^[�/�,��j�T74�E��P[Lx�OҜ��F��>��
�9t�5_!ؽ�=�%�>�pn��X��/a�`��Š�O��xOÃ�����3c��_� Y[��>��.Y�:W~Ҹi��e�f|j��n�r��@ڋ^%�X��M�w�J-�=���E��#�W�,��&���Ǧ݂.޿�{����<�dqĸ`�7��ࠜ��7XH�o6U�("ѱ��M0n���/����'Q��b-q��Iu��	#1�L������q���5z�+IH{�rR1x��(3 ���lag�I���^!z.�E�~����/8�+�x:Oa���xIq�[O�D��;�����v5���g�s8�\˼?��۫I��,.�g�^�O
���^�zl$��a܉e�͞�1�8�[GM*o����'CQ`��f���O���"��ЫU�R�&�B�=�d�ixv�6�;!zx��3��XY�Ȅ��l�B3�n�h6:Z	�m���N����������"OU�~��x�)��d:}���IdfF��f�}��=�� �疉T�6jM��uW'֝�:ڢж�zq!`r7��1�.���FBs����YDqr@}�ؘ'-E�ro/�hLZ��Ȋ��*5)�`��O|<���8g��s^R�~�[a����u�d?�I��\ed�o3��'.y3F�\��)��6A�vۈ��=@|{,:�	&�Q�t�����@,?����@�*���h�2FcԖ�т5(2�Ӧ��j�͏Ծ�6$��V�JGI>P�V�x� F�T,��V�w���<5f7�U���+H��`~"5����/o)�)��n����(�� iÕN��*E�gWZ6]�}[]��-
_��D�-4�ИFO��j�p� ,m�L{n�H�C����b?1�)^߰M�ǂ ��	nQ�*�Zs�2��*iz$Q+���?7ܬV�Y�1Oqz�a:;:�;(5�}�t��!0����tx�|.vś�yֆ�i ��T��2ǜU|-�e�>�Y`��#*V�]�'� �O�!4	}7N�{���ʨ�u����yD �1t.�m=�����[� ���+5=���,sIgw�G�£��>f"=��XHi}�Ѩb�`���%�Ձ�^�F�d�>Ն���,�k=��S�s���ӥ��{{����LP5�p�k��%���')8!h��^/�T�\��'��������4� >�2 q��4Z �Y��R���f���핻�����&���<a��J�����-���z'�p`��ʔ��}����OI�P�����z9ٲy�.���}���U¬4�!s��g����!N.B!"�e\M�#��G�7���vN��o���S�-��Do��T�XÄŇ�%�XIdi]b��""��:�2�4�xͻ�<��ҙ)l�w&J54P;�U'R��� 2��=3��qʩ�0y\�$ �X<pyw��Ӡ�]O뇰^�}�7�����l]6K]ig�w�C8�!ޜG�u	Y�ŵWvs�㤿��
m�Q~ؿ-N�T�n1�0WXZ���+�܎��M�f�p����(�߼�ؖ��>.�#&����k�'�9�^R��%K5�$�q�����z�#���@D��i����i7� ���S�t�Of~�RJ�V9z����֮	��A�Z��� �M>7	�vk�X��P갅A|-�ŕԃh���u�<]^;�0��ʃ)�a4w���N�$Nc� %�@8�;��&�<���f�i��QU��D`}���ܯkk*��RP_Xa'�p��4��;�3f|Ik�u�I����J��;$�t��@�ÕVBChEcU��y��F�=�h�����a�J��'��K���TQ`���cD#���פ��G��q���<&�Z=�M���6/�ȁ�� �Nu���+&��H�p��P#s�L3��1oX������[�b�/��Z��p�1�,��TƉeCߕC�FN���\��
,K2	j`�(�u�hXb�����k-�Pŉ��$0�!�ޅ:��J���4<B�߾�2�D}���b���o>2�͝�f��iJP\�,PhWZ!�;HǠ�fƪ�RV;9(���,(,�<t�S\����$~�O��D�e�Ek:����mC�hވ���8���>����J��j�S���B��4e�Zh���	)�ED�(��8�{M��gK:0�7E�	�d4y9:O'����[=0���S��\ . ҏ�a�2 w��_�z�5K���#b
�aknSq��c���㉙o�o_{*�D��CI!q�4�c�]�Q�i\߾�sVei��&�=qy��|��0�� �k�H6.���Bf��*�+�o׹26�0��|����H�y7ŭ�p�)��.D�Ǯ� u�j,�׽�r\Q<=���@��!6����	�J���u��~�ߝ;�\�����]�K��D����IjVN�d�Q��!�5��#���_�-�5l�,7�����6�1�{�Dg���d�z�JH�(��-:6U����x��������HUg��EŇ�ϴT`��92�:��s��E� <�'���Z
���8�\�^��%|���?�U>?,�co�G]�F�/�{,X7Q���}��b�nǫ����d��Fk��޿��{.k*��Ezoމ�X�/��+ܡ��k��5���/���4ѕ`1�|�	�y����Al��	�/�|*g�v�W~tc����rE"b/,�������2J^��㳖x'�pwީ�"O^�"מּ�R�Y5�d.Qy%����Ø���{u����)��~c�/_�^���,���U>�"͞��+�-��&7�M����F"����Zu�cv�+�ĵg�t��������::4�4��j� �_�$�8��
�Ak��g��µ�SJè����h�Ɏ�D5�ꯈQ�ɱtM�}Jq�ANy�{��U�<��
%�̓�����%/�؀�HoW�p^�TǕmk�^PV�'�?�9dX���u��0=ƪi�PW �2�]*��c���m�z���Dǡ�$tM�#��t��� ���A'��l����(���LA\Gs��50<����J{��ce/o߰7Ny:�+ �y�Nڥ��z:������$�Ih���-X��w�è�S�y�M����*u�$���H�W�5<غU�D���Ɩ�TG�v��� R6�=���Ի,k=r��� �ii�hn0ы�&:����;�UWŸ�X<Ղi��J�g|A(6�X&A��B��;�B�ћ����9�u��1~�����+̾(����,r�+��Xݾ��e"�X2�F�d=KH����C�]�W�@5selމ��y'��]z�QTR˶�� ��y,�Z����h0i�:�6����x�U.�ԕ��������D5�O����������	b��T�gP�u�Y�)݇��H�Ry^~�^y��{�r�h����4}�fvF'U�c���jy7���1�|Tɍ�M�Cj��1k=p"FT��f�J��o�rF��<���Nq�3�&�c+�øh�L���Rf�]��<��.ke	K�D�R���̭ �K�B�����膁�O~��q8`*�[z=�R�ط�)ҫ��yK��1�@Z�M�_,vj��S����$�tc�=���*[��>�dogbXłL�pz�]-)�G�q*٤�f��SE���?�`�֍"�ԕW7��W����?dQ��Y�<a�0��5�8�7�6;������X-����0����3L�������)�%LB7�� 
5����j!�j����D��Bmd!�tC�����Ǖ�)2��S-|at��pA������3vӜ�.��֫W�~�4p�x���֋R�ī�E�����
p�Ȭ����6�������
-Q�J����9��UlgeuuqN��W>^�jݵV� #���"d���,N��5�1�N�%�Z!A���'��z��]���k��Q������SH��.Ï�U�����s���ޥ������k�a��`��#�8ԞZ�yW��@�s�	��u��'�L����jpçи2C�[��SA�-[�L�3���У�Y��R�,��|��n��_Ř��Jwc'8,���=`qi�#=�T��F������_X����@~GX3��I���.��|��)=������T�(��}^�_�Z�_�<Yy�b}R�}9P�fS�J�y��^1�|�0}���8�; �x���l�]x1�������َˑ��UDk���2n���.���欀��_�$�W�Ş�&=����v0�k�AB��ջ������}��n��˴����S@�3ۮ�(��-�<_go6���>9����.��j�G��_B�Z�*QJ�S�B���&X��E�+�D��n�/�.�MlW��F�9s�[o�c��@G�W؆,���h�Sl~t L�	ZaE��}����E.;"+���?	�A9ѓ4R�����$�u�W.�U+}���,��=4�g�*ff�	}�(�)�� -�,6�\fB�(X���T���!����M9uR�����˚�8vꏐ��Sb� ���Ŵ��Vֺs`(��'5~-=�޲lD��+_��/.�ޕ�U1�s56�*��H@��&�'|�'�	%\���mw���J��I����ޒZo�^��Z���cQ�,��3��gf��:���22E����R��x�h\�q<�:�V`C%��}J'�\R3�jdO0H��%�=�,�<��?�����SAe�&�Do�g]T?��~Z!N��د��8�b�����T�W>�)&9[-M?a�.�Q��
b��&�`[�����n�2�Ak�,��ޒ�D7$9s7�OL�Tz�}�ݞ���h+��^�{`�i'�f�x ���ñ��r� lLk���ɑ\m��3p��9?���.����+jj>��^*@!N��qvwt�!���t�9���N����5�V�`��*�64�x�,P�;@�lg�D�.�g�OS�cAx��I6��x2X�O�LC��˳���|��!�T*;�BV�=H��F��Δ˫�#zc/>;e.J9�Π)�� ]�ǈ���W��	��lvZ9��\Q��p��{��us�F���"_��^pf=a��?�{k����	On6���ϧ�E�&��dnws^[�4_?��@