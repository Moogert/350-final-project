// audio_config.v

// Generated using ACDS version 16.0 222

`timescale 1 ps / 1 ps
module audio_config (
		input  wire [1:0]  address,     // avalon_av_config_slave.address
		input  wire [3:0]  byteenable,  //                       .byteenable
		input  wire        read,        //                       .read
		input  wire        write,       //                       .write
		input  wire [31:0] writedata,   //                       .writedata
		output wire [31:0] readdata,    //                       .readdata
		output wire        waitrequest, //                       .waitrequest
		input  wire        clk,         //                    clk.clk
		inout  wire        I2C_SDAT,    //     external_interface.SDAT
		output wire        I2C_SCLK,    //                       .SCLK
		input  wire        reset        //                  reset.reset
	);

	audio_config_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk),         //                    clk.clk
		.reset       (reset),       //                  reset.reset
		.address     (address),     // avalon_av_config_slave.address
		.byteenable  (byteenable),  //                       .byteenable
		.read        (read),        //                       .read
		.write       (write),       //                       .write
		.writedata   (writedata),   //                       .writedata
		.readdata    (readdata),    //                       .readdata
		.waitrequest (waitrequest), //                       .waitrequest
		.I2C_SDAT    (I2C_SDAT),    //     external_interface.export
		.I2C_SCLK    (I2C_SCLK)     //                       .export
	);

endmodule
