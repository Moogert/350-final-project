-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
t45QDhyoitTvTjkQpG/BjtzMEkVDhYZIVihiOdSjD/2QyO3vNr47hzegm3ue92GBs5A5gXnIbOjJ
2yNZow9v02apGytOE+DmmHO5oQJkpxC32L0Wqyk/oJoyN/AEC0MtZ++jPNYnPHjVfba4/Gtg54Ny
zrJI3Eo58ZLYJyiXkFpzXcM/71C8ZJJUHk9H0U/8r8jo7hE19rlTt4pgP55aP5nfgikwlqxwmpl8
s6syPurAUwRFeWADHITvcbHa/Y+Xq0CBoW9MNH5g+J6R7C4/BjgjRZkQyYJhh23wg3nLB50v2Vnk
rRwweXwqkV2G1i0y/Rm9IIHaOswMgaQvuWAY0w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
NnX46T5/aGgWFsNA5uHRutnU4sAf/DhpJySzJqA5Lm+mL5iUC/O1D0wa672q7u35TSTwklAwHBwh
YUvDcoSQYgJSQeQ7jpx0dCQpIb/3HRz9/NPRT7RrilWbHD0RJt86/tQ26W4osF2oiZ3TsIAXlmA4
Wib9voB5g5eBw0Bja5b8EgKcp8WZpL81AubBGhqK/3sKmCnabkGMoigMSnKZT1KsRsKGfVmmCpXJ
U944EdL8X9Dd03+N4LHkv7MRY9VlAcGuoSX8l9q4+zUdwxW5gGSpzzMCOB3eNkpcc2S5vlC0xqZc
s8gCoWZe2fH97xOuNFo2P55xVXR2InbDcXO8vMyAiJK6tfmfcH3kmJi3H/Nxx8KTr6YWmoPzXrvj
RfRs0etRw5AoEDQhSoJ6o6Dp88bTZT0nTk+hUjkeUnvelpzy3eHxCO3JGfh0T+dbSdVQRMRz39xj
Y0KVbh0GLxsIVlb91vu1DvL1WnqQIaPEoUObZP5lqy4iRkMJF7sBRF97gyok4wNmBN5hos0Lu6jh
Qt0Iqi7SmXNNBgVDrBBF0RJfgfmshGigmg+pr6Eyw/PCl6BsQyN8wleFn5xneFRhnRx1S613vfro
ORSYMa4p+BWZ6yKLedE2r3va/Kmyp1U4yMpPhwUTY1leoF6XyGZj+7/JM8APvvLBMBLkIeLt/nMV
w2L1/rNaJ94z9j2jUbDAbUd6H2EFaSNMsFAohUyOK5v5cigF+X/R93KX0XcslFLYfgUdJgEm3Yof
DWWp/9lq8z6q55je9vBdMIQpRVT0QOicPYtP4GzHJcyoxEz8s4RsD1M+8C3IagZPz5XfcMcZkT1q
8nU/Iff1sdhnwA6UrOgM2DrQ9UstSHApsNBisG4McCN+H4+F6xrwHR0OmaIn33eiLzQHJJ0m412B
corUIAjvyaFcD8czX40mDDOwY3c3an92fPyWmKcHkcqh+E0lqIL+pSFmChuzrOly3Cu5Gvcymtp1
xhjIsnDtLNP2xlmHsnH4erJM+OAKii9VuXZYxD8UgKsIlIwBEtBRomrJAO5iD86ITYrA1mmsumXM
i8xiJqj4OZ5VmO0+0OcjZtIPKKDmL5hVPtiRL2RH4KQQMFy7q69Vg7C9nF5dYXiycXyJthgc2pJ7
R3dOeUAkn5nUlg9/0DwaFc3eGxW4xSwZNRYUtWC623hOm7om87LeEMyspwds2b4/aj2SDiiwp9ut
2P+lWzmF1W28Vl62ZtVsG+d0bcg/orkNlZPaoRbFT7ZVJIh638P0C/Qat/KzY7StRHxOy1hvEBPX
C49/MuS5iv3KJLnaSIGAOJgseAcMWOFjg1+CETPbrOt+0r17WDhPBdqT+PQuh3OPPvKGn6yYkVcw
IfQ+Wno5NDqDa/VuiqpyvgoEiD15PscdEe25h2P7Uql4C1/+fWgLkGDmO+1TZ9IohavCHOQfUQpL
5eb0mPgRkcU0CiGfUiCLrPJ+l96SA97HkjgZ6ixRoYgVjEvEpa7pG2MhrDfoZjqafRIH/9o2PNvN
AseqzaWhfxFANJ0b3pjiQv5l3dSZUMe0I4n9KqYKb8dkWbuGU2xFW59wfMG+s5VpXadiLmdggNg1
bwqUK2dnNBBQ/E83DVKfV5ScceFt7BFP28uHhArSLLd7IP/8NqbY37COg/ztNYGSKzDpubwbncsi
oBdX7FH8qK/89MX5GMtoIFuXMP08C8IlH5JVLiQLiweuB7ShO2GAJAHLGgZoBqmGqlvGcAe5Sz9r
lnndioYXBf3guFEOjknELelZdQQNC8MzLkK4RzJxnC6cqR9yv6TTOfkLBrK4tERM9b9rbhHoAEa4
4VL+HTarbTsOSEJoduWln3CrqzIUeGZfJ8OM18kMeBQm4yFr6YFKAbXBF+iI6cG0DKc5bGP6S2Ri
anQn6fMTUO6wrQjAf/HCCzsZa788pZEDQepGugLE5wPeDDKDzF7pXpuwCsj/bF2ShlDOa+WfCDhO
u0o+gArnHWItt6XRFCRGsIv4JvkNlp+re9rt1XOLZMgV+todPV51cm5Jh3ykaByaWqmFENaDQ+T/
IinL495epXNnx83gDlpbu7fBkTj2eOBJsqERnaJodEzDKUp16Ltl3/5SZyGXr0gx88zRN6FrcySN
Szq8rx6C2wDNb6wYooPAecLsUf5Gv14WlfxeD6ThzjMM8QQBANyeZsRhasJRO/0JvxggqHTU5q74
3s7D6PKrtm+zYfijHAz7Xl8icRlpXr8hUujb3uEA+N3GDIoOKr4SeECoQ2bGVgfvVdypnbU20MRt
D0+/U6bZZVOamozRcspvqrFCOjl24HaAc/1kLXTOaHocqEZnd7IcoV+A9XJUemt3XAL7r+xiCVx7
ixrRJtUWPEyPEuIRF1LfQSoKnCoeneTlfOkLPvG27ObOtL+7/AGgWljOyra3NRs2Xb/h52F2+uQI
c0f5x+c4MxYa3SsE2xiKA5vrXC62sRxTqJ3A1lujn5bfjOdB3wj2Cl/9Lq5Nt5DxObj63VKLUUN/
nFBq2XD1OsAj6YYc1YWEHbUkzu/VNzskZyPnSaAx4ocod0JJV72tre0IwsLnJne9DIdTRwQE8ROU
Q1w2ufWqsIkZisSqgm2UZC39H+RNjZNrSnKWo39GREo0hq+YvV/AlIkGewQQU/lNs4i8hQLi7gAw
GC8LduktiAbNbpq/+/WGwwgzwWfGW2GIGsbcQUejc7Fae/lA8KKGTJW2Q5kOdYidbP6itBQNz5AN
q6T8f4IVke408pYmid2f7c9qnJFJbbn28AGlDkvVGRUXwogMAeGLx4vLehH8I2Cy3tSVD13fHPtn
ueeLtMo/avDiyLy7Cf5/BdINROzPLP9vIfcW8WBtT1FOtU090Xix0KeTyGAe7TxIDghcLJ3g0kfp
MqEBZ5huudF5TxUVtpUACmmBHovTpPNBwAjkCgcPcXlhaeb8R2Q8Bu6T+V5ghhnSTnVInMqaes6N
8jbUybUWnbNoDB9iEY7TYRNLXMovWX8ffmpb4u8VmE+2dxLhGGOr/xJGe2lj9P5zhjGtxll2SaK3
5bFRGnmZasdUx4hKY4h4wLC+y7niO7RCWgdpMxvMMLmaV/aXkA7zfZG0pSu8zlTUkTzS6D6wCubn
mbbQ4ksHMsgBu4yk5ec0J3/9jSRt15dxzQQUo+IGM7ywMovegIHskYTb6ZqGBAed6DbNq29Jz7bj
vmHMOKAPocBEIKdxXMcLeuGFS+7BJbEzcvWKz6glIKReU3XJ2/BWUqADZMSOgGfNZ64BWtcv4ydW
h8XRKFedh8esGdaQ3o5zNiduIgO9tDeKZlq7zfVTlKfHGyEVOUUZn2Vi3486mb/tHijglGbqDWkI
qjJohC7lNG853aahOoYBAyWIVo8Rx7lPlK6v/8c/pFCnGY1u3hmIhm19CmXUDddxbvV13VMFVYp1
ItEs5pBvQMR7bUrolgVfIrp/SjJdPRd8Q+cjmKX//aNqlW+JPJ2eGypl7WYhZQYyfKXsF8+qaCPK
gT2HJS95YPCy3SIvbruxf/IElWurg3EzfT1zuMEtoQsuNkPBEf2pNW0zjzCioJMHitdQzZihB7e+
Mk5K0zHDi0TBg7pK9f6YrnPr7mruBj7sTQiR8FWeqlMXHwdUAV89/xqRLwOoGSUaJd90c2+p8TvZ
0JTi1gyR/KwJhCP2qJGcJypbX/XsQvVrMH/s28AAO5Gebqm25Y9lRR7BeogImtqnjF/ZvGtBdb5a
b+2x2fbpW9vCzgFDovCzqTmT/642Ozinj/aQ+rULV43cD+NY8BX6IT5T2WZE+/11YM+DGhdXpy0J
zvlq2PpM4/1ycX5nILp4tyrgHXLvztziNBfXnDksV7pi9gaRM6nGghd62xobHhgk0kE/qJXWy3lr
/I5iI8RWU5ta396TQVBoSF0AzCHx42g4nCZVf1QqYAsGMQHiNkaul0gh6iEHys/v7aESG1of3Cv0
o/kkITGfIPi+iSahstPgKjTB8ftyQ52RI12kvxCwS4xyjN34FLZqT/6TeKK9BLfRK060uknDY+Ih
DjCUzGSvv0KWyyycmMzbpaoUaXHn8rDGjq7pt0W1nXMJB9fCrsAqQAWHxytR+g/pUQWkE0+7xXWz
kjBsPoKmw3giSgAfl23jng8Hax5aDiAHxkhu01jAi7B1caYqK0IJn5q3bVBwRdhIsW1U5gbLcyqd
tGVOVT8sh+JmOQAn3bqTg3xX3TyKJCeAQ0DSYXzMRJAPKbFXL2AkqKc3VkrHEq3Ej6OioAgn09V5
6f8TfyUvputYru2oZM79CO3W492pDqWNKlnjfMKt/VQ9NkifrC+hUaoSb7Y/CTP6h5onzcrVJ9Qq
Zccrr08G0lSLH/vQpmPzfvHxSnEsPXCMaTBWhxTZjuP4tgt4jn5voetSFZvK7aLvMM+OsjfoQ3cz
SdDEv4yU5t8ETJx7z/uSYmL8ybcaLZEoQkAO2BXBrOiQS+RAOEDTMU+6AGviaDMPmexDOXL0ol33
saHQrT/8eL++1Bn0OyPH8SiKYmzFXr4QuMRDdtwDAjZEDYjRAPMb9Td4spPwyQXFYDvXux5fr4TE
u9pv8aENO//Br3j+Iam6ieyoIalnK14RFON280t+N6WwdD4Uit3FMITFAC+mpQbqMeNuOfK9RJF0
AWZ50TcXe9R/yKws/T8NUEQMAqfOiJ3G2cFVv2XHPLf9dFH/ov4q3fZCZanqV4CTE1gIm43Xm2Mi
yueiunktrWe89LdinBxAfr+l9jhaNddX1THYpMIyItpQ1SZr+k2UoiqVswIqmaYzxsrQA0EVL3FE
7rMZKtSP8lyaPOnp/QZVQOAnCwF6GBV1Xf9SRzq7id9PGTZ1pcLTwTVyd5pmeDVXMjEsDFn17xYJ
shc+OkmmuCzbAM3riN4EyZtrDwACUOKCsTixWc8voTaaGR3LFJlT9pUxctkTS5sKxAFOYeWcpay/
qG9glx8xwUOjOpKUrHfcY9k/nVoOGi2q1xzh2GZQc40wBnTfRS66Ne40DN/X2TYKoVg6S52jmwZS
tEb/CsPQZs7T6kLXP3HlRpSb9+uCccUf7Y7ckqmffkmoDqKazMJ/Qt5/erwJJbD3VXP8LeAtieNd
nKU7o+jiuOT1YFvTxMemK21hta1w79Le9dMkvNYj/Ioh4iON1b83f2QrqWb2JW5gIWD7RQW0dlLL
OcDCC/720+sz8zx0HC0Ld6Bn3gHZ0VhDc3J5DR5mf94WHxJ23t6IkFdLdV9mgAOR9heKFlHryQgW
J2U7dMUaTDk+ms5yzyORb3Q/8YM56y3Bvmfx9dWfjB6hB9mUZTyINxda4WeOXQyVlGir9xQiBsip
iogPIvK8XwnBg+bGX4w4MDoaadeq/L3oJyyMSliBNXPqq0p3vCy0GLat6gfq7VeU2O6JCOeMecV7
oWR8p5z3LTLZo5D8mpF6sr1VHUHWszVp+I56yfeS2ZXSvAgy2YmYTWOlVmAS8GNk9je+zoBMa3Sa
TTAH8SRJqq9USx6623nRC2R+oxVYAi0x0J1IyvI7EmjPZyFGn4NO+flLObdh6VYMbYg5oqMVM50W
8MCiDM3OmKu3aA+nMIzHEgFY+eO7xPPhcXziynNawCX7lBd5CzaNj8YLpaX3HGpy8Y+lTyFDC111
EZwOHKqCNZgnwtdwqxG8YXg3cpVHZZtNYAKeVEfeLiex4vJf2boEshMZzmBC8MinSy7XeqL6ogtp
qTL2p5Vww8WewCMBlRv1//IvJUnohnhi9ra5v40MS2WJEgw9GaebAN7J1nNujT1Mb4ZkL6NnXC2L
+8WyckwMJPQO6Tmpbjos0IKwhL86UiVCbpwP9nUKJ4dwVPvtzBPQxL3kM0xytqSTQEmEGx87dCBF
UoMoEerV8uK33lZ6Bk2nDSOPJAtiwSmraLU792o3/ByZ92NMY4Zzwkd63MSyDi3XGGK1mEgUOr7e
Ut0wTNUyramePmF2cLZjzt3zAohS+Fy76AVBg4ohk9OP8E08yANGKbsUTFkKJAZSxUpvVSnyQkD9
/jx5gEybYcljf9fUn6Hdwm6V7sB4T20bJY1ytyz/8vv6NVMaDKrkrIX6jG2vxOrrZTC7an4/Q4xZ
NR3MwJdLOnKEepRqbvwsyzfyvvP3eLjgWwN+V+a8igBHQkJ+kS81BkwincmV0K+RzGNL6XszYCW8
eqIDwxZ0XUGN3t8oOlCEpceAGOaP6jgNJe5ciSgL+Df/QFPjt/9TkfefJStTjAoSzXSjtNfaOjEl
5L4m3hFe7nh9xFwfXhqYQ2ViJoo/dnEuLJ5v/3Itt8m1If0nGcdamsG7fw0bnOsJjKZ4wX8uMpYm
7HKHDJPTTouFs/WogWHdMCVc8YEV6So6Zvk5fYVok2ODNSfeb7d3ygoJqgKobqeMjvbEUBjaEYxq
j92gaRhPk2Sdon3tguVXGnPpnrIB91adlDlJqo8Xu5rNTWmEY3XS6+toQeLM/oFkBvb4x2VqtBca
9GlpaHjdBo6azcxS1BqbAWwUQ3S5j/Ttqpt+rZdfFy+uKnbB+SZVwa7T71C8ao3WLhEu+A3DYlTa
ZGXfHuvxPAPpkJw6EugRwP6bXTrAMlKKS/+/vX3RbIJ02CX2qRVqRACON4g9jJ66NMHD5/Axa+ZS
iWJ1ZYDWQC7ExPsO/zllR5NbqDad/Tkv3ZBiIPyH4yDWbAAJnwVouREo2F4MIzVrBwCgLjCGraaB
FrrlKNXIHtJf+q8Chh6rjnJTh524q/DqWe2+jPLaQIM1GQDalHcjowDcdSoRfJcq7UijmkoM609z
UD3Rm3UdE/A0Hni9rfv1ckQrezCTDNRHZLHRbJT+5GhqSlCwMYVE3brMOAKw7+tsHNw7//R1zbdd
e3QcadjUfjSHAE2eyZbUSaJY5mgDACgFRDFb/chYUebrqLgZi5NanOxIe4pX2XvcScwxzIWufytS
ia/K+/dCY09Ae3UnLBUoXi6bxvUUQ08w2i4C0OGJXK/Dzyo5XywY+clfTmUCu9+QLaNj5VKEqASo
4lsDWImGihosQwpf+2MWmJhSkUJejl9dCRv8kLnsRL84BluHr8ultnZOIDxw+GRrTccgbbrDrK6A
T5Rma9tafAM6iOADVPSlRharKGsEAlTkp/KVw7iR4716OPX49NEM8Oz3BvJryEL+y9vbeHOqJnbu
vGxBL+apUyQe4Mh2ma5YoGJHacgRsnEgCh3vIbetntq/C+AC8DzHbtJ2fJA2tl8d4Uao6Qor97L1
6ejaCi07SvsTSNNpbejvqgntGc/jKmSmOEFixctqm2wLoHQ7aRJKMoikY+XYYB6/MWM06DTjBTqM
nvQBzmzWMnyJ0kNCtxbiXoOtQdWSYHtav4Vm7nXulkQzerxkWIdnnpJ2at0SJCzXk5XXjSV+hHbZ
owlBgsE6I3Ae+ZpZX9Z2eym4yQCy6xpBAsO/azwrxDrV8I2mo55njD7AfmxLSmTlrggoMhR++lR6
WnMui9r8CKRdCwHCZl3wsfXcgI9nLLdMXPzEdU1ICBtJyJCQXxvLPrmai2Rkyn+KbVpyzrm+L+6g
gSEQcCmXs/M48BZ9qWiLMilHBRd010uHLD9rZ6yo4BW8JKygGwd/DDO5JxS6fj9aYWrWqIrAynLf
3jpVlp/LMB9Q0OwnPyUKfr6NYzDRQ+R7ZjdabaW6N5VaxFreTPDXACpzXwOq3QX0L2dZw8ZX/6JY
ZHMBDFU3kLWHcM5CC6T7H6o3FkuaBT3jQFiI1dPg+3e3pWTSjyTcpBus4Y8tg+HBaneZYpXATWta
UGP0s3bfYl5c8lAR/SnC61od6K88Mf0hpBsH5jsrJQNiVGIRnmLSwFxunApdKGYTSp46XwKyv0Fg
AWYX4iJ5nq8tjjlW32aZZ7sCkktqVh8Ss8I16jBOaYtZXqfBszh9OurEAOZxVSSH7lRXvQB0CtSF
3+A5IUSOtt2CZz5r0dK4M8vvawPcyBOROjrO2Rj2gcOXSlsyjDBKdA4YmcNFuaLcVL+khTZYpNh/
az6VuqMzlgfgLjRT4/8FtVaPuVVT0Ytp+38so73t33IWv6DN9z5SD9LSqYWrSzWHeVlEVJ+w77Uf
VFYhr7frEx6bzJ9oEm3CUKrhElWiM4VUTdKHeVcIWCD1rtTU1M1NmRNZFKAQS48BtJwzAYdZCfo/
ZDM+IyRh/dA8raOSXHgBqqPTI1hbuu7ndLb90l6KQMRUytLEoQJmf9OSF36ani9//pixuXFXbgsC
f3wvl79gNOlbts0TEL8P7A6kfqlK6498NC3DCZcyBKZ2JWqsxBFTxN8tBvFOrNM3wGfGNfUGNy18
rhrbREl6KYmgo0EZq3s22h/+myJtlBqVQJBXT26pVFbxbi2KXP2dOLictZyjcXeSvs2QHzvj2YjB
iqzOp0jWRcyjwS2OPEFzK9rrtIbzun0rGuYh9c34cjpkoSfV4JlsqUlmfqnenOCVK56BAjR/GcFL
yo+o9oRHInHwswftxGvdXPuKqPvwB2p8jwph88lQEeQyx2Dq04DQqkqGjWEphxf2MJZIHLLLA/m7
D4n6wC5pzvTIqv4GTaPBH6blDlxBy998hwGEzigo30kFC6Zn6f2SKhZSs0Me+FlraHyCWSRbQ06X
7mEj5xp9bc2elVBxdNeB7axmHXpXpkiJACIJQio2k1Xjq8D73myWBwU700AhHRSwZ8Nc0p4ufVGl
WP8eK29uz1pA2q5JsBONtVOiFjawFz3l9n50asuHBc+ik3wkqOpXUGk0IgFXehIlmGI859FWKuJ4
AU/s5YB13ok2rhVEM7IuS0ufmou3i7KWOaq5qKJMDqDx4gwXkgYOgowZtGKSjfZUy4OwxFt1Y4It
5Tozqp8AqU634NAbH7OIcfpZKDlJ3qUm+5HXR5favWe2RGv6ovcj6KnXXmkIW1nH+kLlD8BRzFYm
Vk4n1qHV/juGkwLs4ALfLjUz1ns1Ra7xGUYFZmQERdYAsvyiorNeLlCRXsDzBceqeapto1FfvpGG
kx2GofahjJGaqcNgBV6bJivtxlDsn3wyzoF4bEOX3FPuoRzrENzF1HSduBDUTgyDCTFJtNxOm7b4
YEmstdokmtVrYRNVv2hXJ7tkuQg3BGTLmp4uXqYvdW35sYWV1kIOkBsFe98XOzgmO7GzlU5hklvQ
CutjA0Mp8CgmrnPhzSkjE4xviWyPVf2aobVyvQBoFKclo43/NXvjXBEPu2mIdhl2sWN+gadPJGQH
QDsEB2UMgZlRAS7/LBpbeRWDAecw0IkNXsyPnec2dzwruqzKqXWDbXRt/qA+OLDvhxc+qIQO3Wvk
2O6eMDJ+kWAMIGB9XV7Xos1yGTyzHDZ9MYw2as7JSLpELio5kn389W/9AEOvmcRIPJ1NkDumXFsj
yUFbjZMQzcNHOD5ODzuQgZrY7qEWeZvPI7IF+iFtOg/bwktzhgKEr25wEcwhh2c6WIT9FGjMZWBp
SmTcpb07JT0YyXma0potycyoqaH8HPkd8RRQZ9yIF+3SfnCHVJ191lEM7Gens/lW71Z8fncg8daN
N7+6NAwYS3pS3tMvnJRzmKWULo22tqvliZaW5vDYMbWE8O7/IrAdqK68OQ17dazF4o6H4bKKlO7L
JbzmZApBAMm3Icy5eSRMMg9UNhWZ8lnw+9t1eP26bR2cDX3PjHQ6EVSHHOZQNTPGVLvWLQbokYvV
BcD4DtV+1PJMd4CYGwcPw0wfdC/nLLn2t0487pMR4SF70KVO4diwvIVL7ptIUrN7/TPPRSgvUQGB
AV8ZDW4od6OYPWTCX5IZInxRz+Q2TmhZxlZLYA+8GCYLJqYxtcHqXVRzw+gyGarNcRUq4SZzV8eG
objVrwGwyoEAx3TyI0xYQxYYBv+wr59yDFxe0/NJjn3YQLnj32Ju2tBaeDKMi+/HulBcZcKk1yTp
xyIESkHx77oHXgRKcP8hY36IycQFF0BzES0Mjjsjc3aEv5smLDEZi/CUgQhXF/7+GVgHEi8iq1ET
3f5TeLUYNXwNQZ3IK0R5ZoTzdmzgPBkaj2FS8evbNNeh8qqiTlpWdwScIEP3n8YCBr5Wh0xgIW6w
zTfv26mqzTmXef74uYQ3mXgiEP4xmxxGemfMUo6QqDW4FAfXjG6B3VsLowpfPWiBRLnEt7KQokds
NkbpoXrAMz379ruGwchcPPAQ1j2yjTSMIK4EXVWCgu3LqJNKecsK2POOzE79DbhLdZQ/Klcapwv7
NbT5n0ai2gP6zhuvWeTudpc2yI8LiKOmssuJRm0alUO4Yoqj+ESb85QZPJIICxHdcIL8UWHQBHL4
OmV6eCLI5WaQ/x+i7C5Qc+Q2Xwk01JTys313Ic4bQ0VmYWELP1+GsBcx1PJ9W2QiSC2RbPQqnbB6
h1xsGoNtUWNBRLlLjFFsvwKIWQ1Vw4PG6R4qeWMLLoAmbmsWltHJ2TtFKchdGt3ZBqDwDVwhiOfW
xYdyoN9FW4dfV/XEbjJIIMNhScjV2LoSQ89wmJHL0t2RyVoQM9Y8+nfB+sKt/+AZccDYWwTSyOUj
VIQnPMmK5FsCLW4Tf+ICIEVCgfGE2RmJUinn+Xc+szs9zp4N1RyGeBWpR2K5lyVUCe7VGZN9AnPc
6JK/nqS1hKoE/md0evSySwAPQzdkdBycL0XPv0pUSZlo2KaF621Y2PGrTYCRxMWAuLfFY/bygivZ
wIWtsAI0ZBsg737gpObGYeCWR5+caPXh7qMFxPbn1Ymfz8SbNod7peV1zcdgP9Cn0qPskc/VxjxQ
iage5fnUngCtO+9TDMzmYYtw43b5xbI4z1rulGWmpEjRV8yyYQDsDfiUiGhWMMmLwRTVnOIVBUHu
tKe9Ki9fSfBKkFCBDo4Uk+uEV+MfBNzucmur2oCjKKPcy+5NeE0fKSgoDFcyjYOaK+nMtZszOeUn
37mXGen8TizSTjK7lyIQxHy9Qg/QlZsCJ4VOcRJgNYxng2668FRNe74BLOCwhergvw7kwn56HHX4
bblRJMHThsxcXaaf+329EMWAJWZqYBMylEjhiQhFF8cs2zihaPtTdNkYubx3hYksq6WsU76/8Yqx
R8DDCsoGmLg/yaD0waPpBFuTiq2Z4ASQK6MCIdrULieOF65/hTTyMLWoUy9fwHCqR4dwiL7Cj82K
w7uTkyzuyvoAeeT6gE42H/ObPyYVIg+cnxFA9Dxu+1HG7GvGzlO+q6iSEUd4HErQCHxhYO0il2o4
2yXkIi+SXsk9Qv0BX4e8GVzDsnsk3OEe786tLbMsSZNrh4K93syGCFEQg3rpJ/NWWAZGgdB/AnQ3
U6shbdS6DnxhKFRd2pvhaPghKI/D5/ADVwtJH0eUJh+A5ufyphQURQ/eNaNVV1q6O6nPsR2C5+WF
rKD39bBnaGpteVenFPZL4K9bXfloQPeHoaL4kJzcq4NlGRe8w0zogZlffl/2Olrbu1erp6N7pXW5
j8q2HSo5xLnOydzkgXgoMt42PlAOwfPj07iOr0MDj+eiRRysUIa5AADv2TfyHBSIIQGXVvIhlo7O
yeztxGZEd7nDuNfzY7GkFgo9xagI7LsoBdpLE71/DNJSpbUGxXF5bzPq6IZEm7Zt2P6/sbKepCsM
Rdz3erL4BCx23Dz49hvyhXke4GAZNU9fOzrOxv0tbvgCh2IyDPx0ZpD25Dtcd+XLizdb5OPmx0iL
3pvGC5qbaRDTC04gGsn8Mg1HfmXzLyoYt8BZmrFno6U6V/hwd/t07JMNKzjoN+UbktE5o2XEcMAX
shWFKLuAUChFs63HxPw8/Jrrt2PxENo6HAyrZRJb8VtL9TMQqoTwN44O9Onhslrhhg20eiPp0IGD
IZh2tsV8hRaoa4SmUMsiuswMswYdQIFOpGr6b7xnTHvWmYxPmwMz6rVJrUXeONMTafqe8QhP63Ga
ytvM7bXbgn8qjA/m2pMAdLwj4pN0MPc17LD5jOUG1nCQSPc+HZ9pFpnqnWCdACaMRqxOGRrZ8rDl
glJEjHLc7ugyqKhX9BWYZcjjfhLIolvmMmjb648Wm8hhv4iMdYYSuceZSoDRhmW40ZL30xnAg1yc
8gluidxNAmIqUS4f6T/GCccfMtv8yHIa4rGD06EDXycLxhZFAt3P5UJXurccu6BUE95oUeTXtuxZ
DTzXXkgDchgdfv6XHaMawFVHUgaSXLkomYXMcvTni+4xcfSw2sTrEbs2CX260WTNEjcycDTvNTdi
WmALuDEPhjcirVGfLq2qjGw/I1cKI+CZUIczfuw1bghF54mJ+pAfD+ilKa5vU6OznCWut/wUypcV
8dmt3H0KOLqY7Ngjn+BHVm4/QawFO+DPgwb97U6jCHiCiwuv0MlnbZSx12rMFyQ4qYlQqq1ua/dh
PcbfQjQ0efNrvdErYgOO1SMGnxO0AOOvj5fKXSX197SfN1wx51zxnlO0EYGFgXxusDsfcPTEjP9E
R+zO3xSFS7McvWPc2kVqT4iS1Q2TxobhlqsdpsNZWEPLnWt0eY8oOVIPYBh0KHUUM7mefrF7viwE
cM2SMIqv5oRjyzCsx/hHO3AnQI2BfleGaLeFw2hapDYSiIrsbSrlc5nmlCyEwnMPh25AOdc0+xX5
ZhMeT6//wgH6lbkqsHwS0neRNV3s7wM/yqrNjuKlYScQMYi2nrqXN5DIH+hCqSDBPzTgMr1OHhK/
F0foaBdfaTtzPAZRDzv+15HmCvyquE8uKGWeqjwQCYirByTuiRKU4FJWaX6tiiR/Ant3lJztUG+i
T0j38MIBl6rv0jhRA9RIMxZgU82W3yG0ryr3cHpctjirJATVJtXjsG97TQcOCbU0Ioa1/CEczZiz
jHYGZhBrhr5o3kJyGQ92nbW+PgK8p4KeCpNxsdt4B992ekotoNFqwl6P1+fT3v4P16H7iH8M5ALe
Pjj8USll4cHSMybxEZmw1KzR/lPdJLY9AyKji9LLDUywPRnpkdhnasDxdgxplbbkJsQPlxfAkO23
iOp8YWsFwUg0IX77OBZW8yZQJEuumwYy4TOQgCxNM7BYlLZ21wOAXR6vfRUAfWwlp4HNDMGmxZIK
Agh7X8kU/lkqqC4JEF3MNu3YOjCguE4LdKD4a/x89vv8Er3UsX164YVNqWypbf988EDpqZeHhOeP
2e7l+53AzUZcz8AZYQS7t5PZDfR/e6DE9Jzup1703+3y2Umk6R4ayBUnlV8zbLeDiegJAMFaU/hd
okBQIvUW0dWIMXkBujxu/jf++SmqCzO2j7DF1wHNcv960btZ2iMiQaabPK6xK5CGYBzPd3tBYAaL
kvl7a22S08gHvOc7SUo+o8G1VruGvGPoQ6uBHZ7iOL/TJ/3C4+s5nEIzf+Eu169VSupAFNSRzXFL
yepyLOCMPsPOQmIGjILS/ph9gpmuxbqtD1IwsDhBgYKwrXhH/jDIHtyZeTjp/AigtwiC9UlZh3Rl
pz8ByU8erj4WW1whPa21dIWljoqBDZE2q2Zfra2K6QLI3LCwp+rBF24HCOTq8/eC9/aT2Y96DEk0
851XceaAoYqFjIKOhoIHJTJfUupdnNe9SJ6oJYSz+Xk8lcOJfSHfOL2sqC5aU2L8E43q/TKBqs7I
0BLxy9CJD7oYtzfpeBKKW6DL/2EBXQcT32PMM3slplhd0kvXtiKmUQzUVsNstdOz6jPX9YaXVrOC
TlX7EXAOBrelK7BYJj1C63aCt6PXWIL6YwpzAEuPO9RMmaFXutb4K+G/wvCAHTeqmxEu+x3EREIV
cXNsTe+0GCr6RkuE2q8zunVzAXh9FWueGOwOnRRb63vq3ac6+rBXe7jyDAyzT7CLeKFnVQsZNHIg
hAYtnkUd8Vi7L+byBs7+EkDcf60brw3ly44effQiYcbNHmL0BWtSciheXODaH4N+QDVf+J+MeHy1
3fsbYSOLcvXQXKAKshymv08DfL7/Hx5TAwBfVkKIO5G06B2GHRhABebFP+5SXSNbSgWcnRvV2ZJx
ZrYmhOPjzQoNXnbWTj1J43HGbV07wqAPA/Bzrd80xO+JT0emXM68RKV7GsT5J5VhkFOlyeN+ubni
uOmHNMEIBNEaFrfD5lByeMOkX9Q8A4KcwX3kdpKRmIPYdmKDPYz9u0Vy1zp8S0kv+v0Ji+z/ztIX
zL+fegtDTCZmy3CS1AH7JwSU2A1Y8NT1Fp911zA1zfg7Y0iuAHeDQTtdxY5lMFG8N7aDsjemkD4W
MVVU74uiUkq0tYgCL53G5fphYckm+MRJ2puKPiH2g3bhquSFiieYjzzvvhVZnh0LNnk3L0V99fyw
A7IvNiMKjDNkQAr5eD4+tY5piWVOVldbSV7NgG5BWvyH34BoJwErL2yY1ipsWi1zPXUERxmMDCVJ
6SVeDD5tsDWJpKK9POLouWu8yY5/s4aVCBVYWAGs321scTho
`protect end_protected
