-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
w22dr/suwPkeqbFkzCl2A3qoZyImNIFh452mO5BYE2i1S1Y605sG3ah3eb9olGVgrJ2kyNduWyLM
UXPfrBT3A3QTH2nX85q5aHO9q+47/vKcvxWNd3lRh2qd60mhGmqZnyTTkKjdi8fCNRtEo22mAVe3
gmoWiCt0QAmBy8WMbYHn6eyUEe8eSpr36EML2L8NEbqaIt0Sg6LEVQeibouE8kCnNFiVTY9nJtaQ
IHr4xGCL07pFukHLbY5ilpad7mR6R7tQfw0/h82ttjrr6DM7k/EQR6kzuN26EznKhTGjk8Zbu0aC
u4e56bXNb6mM8f/SylYmk8HNS+driLFBQsHq7w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
w3+Z7xpKdGGxwZOcq3netGp3w6x0ebX+AONg1xAlSwIYwFgIuZcDBfyapxlBfBeXJ21SLhoENWku
JMGsPLCaGDv1iY+DH32ov40EvrvP9EyfemOi6fH/ISHxObGi+JX3b/vpTa5nhJEuvID+ioVmOAQ1
fgIKJfnHQHniqz9jGsrqz6GXoEL5Jf9QZ6m9M30a59xrL9kNv0n0e3GbDzRWFQdIhDkcatxqnEmL
+TKeRAmYBjQjNH8PLKa9/zhdHWp7UHddQGeWZVE8+naM9fKNJTCDUBGlHdQOG93S3QJ4f6sLw2HU
3JPcSeUzaSk0hLHe8oywtnMhT4e+hUqYp3CUBsS+dfzeHatB3HXihCBDIbO54cgxdv9gHMEX2/5l
o5zJGBkPI3CPQWVxo2uFYWa3VYIWtrmtzPfmko/qZVWIT3mz5yUVbtvLXLyoyPBYBIvW3LvYZvVD
H+QoB4mQOjiOS1y20K5ao+3sPZ2KkcnbUM1KpGmaGfxngMfHVtixZp6GfcjwReScZk2sNDxOFdi1
3xQN8nTFoPyXlZsgkGuuaeqbMkvpGHLqWECRYkk2BJwo67j+9napJjiESpEeDuU93sAdfZ9j0nAA
+IAqAaMaDPcXChi/XfiKzCVgrKheCN5j6d448+l9StiaOtoJEBrK7KTMMsUAt8tfHTVl7+Q4Oqpq
d29oWZrRnC+w/zfP3yz45K6v/pbE8tFRvSwemGhQxvx4lsPgomZYf5CCEqnKHXo/IbXq5qIW84v0
ikyp4iSWHBRby2qFnu9naBfNY43t6G5sObNftozYOGhU9aVzfFraXaSL/263YDgUcMhn3HyPAo/E
5jluubIbHst1rkUmFZmntLz0vfOnbjnFvq0F5++Od3XPRqnHTpSGugaf5K0hdbTa3CKovBlGH6f5
nRA/abbp94Go3LXHXhHIhD1GrfclkqIBb/XJtEi97wHJEqKb4tL+jHewoV1MNHxEYJgC36eeLOHs
sMFo9QhiSg4FOUbvkDioAsX+T7yajiWlO3GELyObntT8fG1hBorN/dPUAmqwkh4SznnXcnWfLAIR
m/R6AllH6ImF1Gdg9OpGvkmKW4f7s6srPDc17KWQZUOng8BYlKes6lr1RnHDBUGtMC7YHiO+ylMO
pUZ2PSCBdNuazN2SJum/ROY1ODRiyB8YQWitFN6/I2xbdMFJCeoSs4eHQdEJ9tV1R2nRWdoZrRTq
rR72OnlaJhOThbIFczawTKW2w9IY7mnGpu/eKpUEE1t3ImwT87pVrioecVYSu9UcZLl+CEOVCJeJ
BdWX2Iyctf00W0wYSnLHmRf1A9LEIBGyREVtlm1JJ1/+mlOewdvL5yrCBaJ9l1Miyw7Rg/nNkjP7
HcN4zFCfEDotIYerxS06YBXqLf2L3tlsKPRjpIn+s1RR/4WH6L3gVdWbadvvpCwb8MsWVcbZdLmB
ouZbCsND+cya+cFCz57D/0SCRMCWXwBLvVTrXdF1iHTWWGkMRFpKj2336oWAwVBvomcLOPd0sQfE
UFTaHYKJpN447G/xkYsU2X+jilPH08d/GWkFTkz3aho5/s3sHMNC/N2l0sRRcXU8U6lMiGjZSnKk
MmoZwJaMINy+LDeoCeuelMdJ0f3Ky5dyphFxu1UbCdMqHwcbRFpg6wCYFAzQM4gnq4ECt1okbz7o
LOZsDaY6PjcjNyJ29NLzIMpqbp3DdtID/IYokWfIVC6Qjx7R8yTUKHu98LXP8LquNiXHHjmDqZeQ
q3VwcXvxusHRRNT58b1n2hl7BLGg0D9rH1K3K6+EqppG3djaYXeFwSo0Yd+6Mn0ApV8ok2GQA8lF
Plnd+gUvLYCzSaj4oCA2MLdmqhtU+f2C2weZyrMOzt4+ftDcZ/s1Vk1i2YFIssNBXDc0KoG0RMxn
XI3Ya6fvgpseBaC9dU2Od6gnyIeTy53KxrZg78l4EwA4vcspU9AuGrAl19qLp9zGXPRBws5fOAlK
hM8RpWLW5pcP0unCFMXXcD5/IkvX1OyngnN9Uq8mHwK1/lFwZG0OxQnAGtzxQOYCWT6djOXt64Fi
GKOkZHufZ+TcLBU99ljIgQJev+XbA1eQ7XgmJQ5pl/LqUKaINkLCxqrfeE99QldmMjPojAruCsUP
2cKtUGQQMj7OpudIxXye4mhAyCMIeQdH4I0IBhDvzR58R6YLXXWCkWPfPFFw+RROECCRzVHVutM9
4fWp2cTYYfF7N+rIwCd/ruaa3sJWVGC+mqAvd85OwkRYBqfpPel5ElP00MQl474GxAGPUuDgL1KA
W7o9EeWmYMrs5x5ayIR7IRGVAM1hwDE191sosQgy68oCbqyo9fAfYBq33+Dcy9FQqSc98qCkADJ+
DSuvch2UhT8BGeBVoKtUXHcKfwCblSNN+N9wn2ABfpO1EpkRc0Wri3MCf+gicnm9uRU4Y4mHIqDG
DxC2N0nnlQPhw7PcO+kH5iykGkjCgw7l2Vm42IwqsF8CqHFGHvShZ/4cjCxsjtFlfpoB8OlB7b4Q
F/oQvsQvs9aKDbcJEOWrIw/c3OEiAinOwfw6KwCdMibRNfH/GTPdJr2dl9H2+6rXyjlejreiKEhQ
qcbU+frCQ6MYy9uhr9NDcNHFxMJfAPpV4jLaL5i3CL0Vpzy75N/3IUINAuH6RKACCc4+S1YTSB17
I7Sd1keazDs3yGpZHAup104/pd1AWXnrqDaZPhaJ6TsV8IckcM+Vesyb5k9NBWpx0lee505XY7i9
ANCPo+sPs66kjXSgo1r2EpfHPXVRvMXBdVZfEKYiJ3LiGn/cxHW6cSKvDmhy//pSGjdPe0jlGckR
vhCnV4A4kJbz8zg6g8fM4ZGgQ/zsk0+V95fC/p6aFmtC8Onp4w/AF77SE3/kuF+o6yJtg2HOrHLa
D558Lig9SxL5AHmnlkFk/9m1dCUSkZaYZE5rjsyTgQW93tEtwWXnvmW9XW13WO0VkPMyswZBoK2P
PBzHpdFTqnFC5toUSBNjDB7Vp4bjeurkmkpgCtTMJKYMrKur48Ef1kIJJWTodsyi6OrLN0MjSs1J
V9KpGwoz+dUxSr2oBgEwQg3ikFw1bpzbxoPRbm6kpEe0yEMWnKE5x0KEF8UqJK+wqNrlgq5+h9q8
hIEVKqxUtzp4YwfPDF/qo8JY6fkWmocpek+QpLIOYUfzHHb2Qb073AyiRnMUBRGtWKzHGPKMkgzx
8h3lUztpSj/pARODTUXYv9N9gI9gANCk1mq/egpwjnVh9pCf0/Ye10htMD/9TMAXeAY63dSFmIFV
ZMrr1jvDAloEt8VIzcYP1v+/hsjPtXSu+yYR41OSK9/Pqsh1dBLgnserHH8pauf7aKdp148wjciU
+wHVDn//L+p721PIeAVJ7Ko31QNMrIOef9vAVkOWFMyzv1Ic2yAL2ymXXKJtrezc6eDtYr2/qNET
NQuFESGUb2M8Go+9SBWd18MT1TyXKtINGhEILphb/63CQPD/qqxUHV5zpqgAgYMqDFM+BLiX1/Iq
nEPPCqGA0P5hknAegtS4anioKGVrPbN5XhaxZhsZNk2U2Fr8nQKsevS5S6I5irCKc40C3msjGiZz
9GNjG4viEM2Xv+y47ipkf5IxXVBdjkh0+WAtuO/kbgka5aBuUJl83WKIQ8LnudE2jI6Cx/CbEB9M
ZQLSZfEzj5JRtRx8dzkufZKmRH+d6K4mCt+cCHHjRoH0QxtojxP7jDus7DLLSdcMclBV5nIJmZig
CtNBJ4kRQp3gcmoDTsOKVHN8xUNisUFl3K0DKTyDmfjjGOUvjQWAGzOeJoi0s2jcPTf4VS0ONT6S
JPUfChAK1p1vTSAgdCLMvS5m5FsN7YVbtMS1VZYuQdYJbMkeDV2hdaOwd4qaooR7BK16/EDlPP6E
eN8zVojNE19qkhayQpCI38MDjM5UHFHY7JQTxXaxQ3BRQftvkxP1YBKiypX14hnn40Q/eXGCcSOz
0svCp0RcoeNczT/fCddQ7AN+kcI63J/Y0roHr8XhseGGEQ4hrwg3LcYO/SBL9BwciYbh7bFFMlQx
JKOlvVo4fDGRc0RKz1rAKz29ldu3FKfj2Gl+Cd0bkHfoGBfairs8NLrN+oVT8f+GxItexj83TUJ5
rhirgbkijtS11PFBEJ90uQQ8eB1XQW82qEUMZ0lbjuBzImF74duz1lYRvnm8gqhBWtJAX8xArYYa
z4RL3+uuGMLjtR5pisSMevEp+Cu0XGNHnfBCzbdKrhdlVy2tU/XF8clnHIbPxnCxZJkxBDGa97dE
bhuzN+juK0vR0Gxlwrv9iwbDpnVg5ILzQD0d4kcZWdBuwYxuH54R6S70b9kYAsMNBxs3ZIZU3eFe
q04ymqIkyDOjSn1FnmxJXnrCmjSxnDrKr+Qf2sPw8zBDXMM4r0GhvXeePlH++cfaGTA0M+ALR8KQ
KyUt4VpMMJgZNpuACw4lRmG/zdMWng4Mkwtc3IQ0gH5PALRmGm2SqCEgspy96FUUi4QK1eK6DTwy
DHazPjKcsSLzyQAyVDGoPcWpzIReAwMWWNN8fubsvC21V4husmIwBT6a3rebVt4AHgDzkt9GNdQM
46hDKWHpmKsQciLpXqP6UIPFrEMxTSQFRNp9hO2qBCJZBy1QI6vk5epaaXq0Lp3oz9fULJOXTbTI
9b1Pg38GMVovhIs6TjDMlEzTCFQtT/JdvRaNWkmb0RscVO1rsCeVmK8e6dEpKPkysQihGij3yWRH
IbkkWxSVd6bO9dXFQ0xASiqf0JPoVF296yRXZVn5aI4Ql1/t3LJ8Bv0cceMuQuj4FL+rXguCus+q
6gvWU6mTKcu3j7EG/aUdqCVYqVGf/rj64+sTwdxdOlSlyRAvhFySMOH7CXoMqIB2TEeeF2QB7zYy
RfujJG+yC9xZOFYYTaY/8nd1gIMKctcNvZNo71bcPJmsT5APhfYzqhZshcXO+xbYSBeQI6iNSLqE
sxADduaQRm3GlequcaDSpV9WzTRN7HKIFn3aXSioBDCqObK3lGX9V77M68LihDx4WTzUAUZYRsGj
h1On/6555LzLt2J1BJRxr385bX+9TpMT6ItUTwRTtgqMIdPt+JODGJCIDNg5mkRprv5Ul6ypcFYe
Sw3vx4Ef4clxNq1F0jjV6sBTifeiHRQ9J/FvxFkfesIJdEjlxstujy+oG4WPaZm9zL6uNecnwpoC
GifFZNnLD8va3on4BKnVXvNTUr5n8e1S5lxelfuG8YnWu4I540BQqXLWDHKfwFaBDWDMHGX7DKEu
EuQSsDDAx30qxNrYc5OLEpGyQpAhkwty+ekkafrctfgRZZZserMuDf4o0CPiykNeVC3F8lR+/wd2
iMFcCqu5YoFRtDaoEh33ZH8WLnhVzQkdz55ylZxDkwYjHD0V9KadloLQgNl653OCagP7SbZtrk/0
aggMHV2riIiuAwZcz7rUlxHnQ3QVRaGi73Syd4Eu8D7zbOB9tI2pL52qK69ZRvq6G2yR8Is7Ic74
smNnrPVz7YoloINZ49z1+c3+Vw2lo5Ff03sTA9flrMK7pMHscGW6C441sf+YfMedCMpnQI9A01cE
DBxl8NMa/DN//N/E5sApOB02pnJh+RNjiGLQydqx2sBfEG1jzN+VJdHlSBFjNN74n0qG6bkZxy53
0YAFmzA5kgl3XaMrP6oMGG7ixLBl9XJzcDoCLm8d5y8i5pzG286AKRuYG7h/jmpVX1whCRRu9fBG
Fltsi4MeGr5riKSM1RLZw5PWgS+JNeqw0zEDQDQRBreV5jl7byuyI6pzMkgRBtGSmShBOCEN4zOY
F2AfKTmcQmeTSQOplbQdVifiz9OQFDM938Aj+YRFxgBTYeNGpnFIkO73vo2/kAG54RX9Ufj3pfBw
og5uuNUrLD79o/lu/32sQ3/g5cJo29fiVJxmhgwL67t7RTj47VLnRhOdPs9u8JaqRRMnOHPr8nAU
DXP1r8rOZvzKZGcoCKTiA3kQuHttUJQfPzmaOEjbUmNb/2PXIBA9u3K1JijCr/65YYLcGNINSIb9
gtCc8TaDKzTGSIGg0ASJFujTtI1RJB0x/Sv1BvfgQ/YAJjmBOv2XLwq+MopucETvjhHbeRwe4d1d
AAAYuqh7uzP4jUz9HCm/0fHp1z6/gh1p3dGd/KtquQiIu0BBckrQMy9Ui0i09IzssxX2+Wt7AKLw
qgfrhLvpjLXAM4+9LVIfTg+mN9wUaClr6N3Vtnj23I8S3PO/YWisAseF2w2kTvZtGwUBdFmyT/Qb
4/L7ftiTHXg/ycdhnjD/HC6zbkWABs9s0b+OrYJy2lQUtmeKRpnrD/pLuMNn/TJllrGmySynHNDs
ImiCyem2bvTOz4GnU3upqDkUh23R/ZbquBpGgx+eczy5obfiilzhMGrO1YNjfqGuI77xNRdNZ8o7
CveCQoZeZnsuGlDYB4hORfrtqhljT7cE54O/tBONxRHsHxxTiAlVxCKYGgkBzDMdiLVIxGetPxg+
VCJxGZsiQ4GsJwC4CPzvZvXJhxda6eK1OvOFPq1ITrN7pBz33TFWMkO8KvxEYipDBnVZS8JWmOBY
vR9yUie9wgYeVToB85iz3ClN5//JcQL7LOV6YI5w1vo+4bL5pRdwYJSTZdWg3Tpza2mo3gopkUy8
eZSAsOtiMvQeAds7LLjtaAvWOTN/Qpt+XYjyRzKmJ84pSVZ4DvZNEvNa9KVWMefGCFKE0Hc5cnac
pnyFbKcyGK8jLXAhimKeUS6alRAc97QV5arqwPu/oiI8s+6H46kpYVFQteRW9f19CIIpgMj3w3XF
d0akvqvoQIP3HN7CF/j9JNElCXS2c3HuCsg32A3DjSwu/2Z59v3n8haqwRLHCAmiEmqRcz3n0yrZ
ERZccWqSj2HgXnwzlofgjv7lzW1WOZiFhW3VP6wxOxO7c6d95doJNNiQ7UCt+V+3Z8lTlKhmDN9o
OxdCZiGZ0rfLutWnGYK/N97bn3HEsU0e1TsgPl8GCK9GJ8QptzogvYfgLWsOo0eQEvoTj+5/WtsI
aBFZ/f2+iBf6A4A3TSUHc4RZ2cJY3RxTHedmvuAh7NtzTYt/9Ymr8U6cwn8PArZacCAcgLaF4u5n
4q9s6/F5SUT4++tr+yiQsR6fuYj1FmFZiAncGd1EhJ3RmZds+99U1UlEbHaSL8Mz7djfXJWc1/Ha
ZBhJ4wDV5k89R/QgwPX9PvM7lXYyqr74MJe9HG1WAA+gNSpxYPmFQ59pD1rSOPEkGoyl3t8j1WEL
2QIVaiW4safeP7Ey6huUptbDCphxlhmtQtCmKjUUiccssZh5yegCqZjeAVHBByc7WIQJRlhjomQQ
l9lzWQqjJ5ne7DCt3msLtD/i3zT9iP2PavBosUTDXc5dRz11qJFo8qfbBdjM3fTDQ4qCJpPgMyxC
jPMPRonruXJI/3y1xIM92BcKBTK7GVcYVVIReMBDcOnt0RZqZfzcnVm3RtvAzIVQCECSTGfjxtx9
xsIL+I3hJ0IUMkNqCi9XMjrVjnHdZLzQy0RB5v75zFLdVry+WWuIlyd7j8Py5DS4jmO0UUUBOZQ8
9NZI5/RQEGdFZtJE/RSsmTrCRUb6CpkxfD4kKw1yNhn2h8jsOeFnTdI36Hbms5HxfpjNUDMbgI0L
cbMgqpB753TSnDdNP9pqgR8y4NLl2DYb1BbSmAMo/IrtoBUpekc9isX4YtWpGJhG30tiwAcmqvPj
8PL/Un3xXX2JvMq55c+i5nXeTHKqjF4C84vM+/tb2iCyjNVWpHNJxC2R89wPm1MsnWIzzUyfIiBB
jZo7DDKwy/YoiKXy5TZ+bSlpRp0enyRNiegZBPzxPZwdiLwuArMbX8zUonx0n5fz0HHLc9YQU+mj
1aOsdXhr5tLFtNMFc+SsN89nV2ZaZsOD23IGtz2euWzm5dLiJK2WY3mRcDrFBAfTvK5xeoSSTTte
b09cptyIZ8q3hAeaSfngb/GZnVx6sGPuzTvim/M3OVuHYlnDS+5zyX5v7K1eZtSV4e888DY7fIq5
2NCnYFSCBe3YpiCkASBphN1ubCZ0M6Ugp5p54WltZWcNFecPWp6AIdTQkJ7fcskyPjlHMLhqk8cH
s7jyV/Lx7kWbZGidKMQkpNIgxTB11zYZIxQ0FCP7t8O9uRk6l6MRx3Uwa4AsRFf+jXwOVNeOF3yl
SYdXE6ZfcPy5nwvCsJ/pQmXCJvKzJvKUbEwtJg5RnP/TWHk/7tZlr6RhhAJEjif+m8xyHiYvPQkJ
+MfycICXaOwAchf8cNpEYK+8EW9ZFB9uNnwh9ccjrVvG3mfgeHu18YooxIJDoc1MWyaMQSKQaJpc
JRwBk7oaFjLXvBrUpXxwCc95rRSvyMzzp78/pmZkHeIlJnNb0j580cuJCuNq9q7N5F5TaORGWoxi
mpL4DMcvH6J+Roo0R3JoIx6QfnUXU9r2WScCCiwIOlSdQANjKEhyl6nITGUkkCTKDtIh9ySFUVBr
EegbobaK3f5kEizyuXttmgo6fTeh+BoN+dE9D7EuFlrGGYoCqp60PCU8YAPTIFtc5jYiQAAvvzvQ
PcXJXmbqHFEnocdgcsf+G6HnxaX1oYn7n/ymMC08A47ZAUABM4x6HEg2QG/RViYWJtzSUFsB1S1a
r2OvEPiqsoSfCkgPb05HTx/TIA4nA1/qFtNTUaDwI/8P22KKO6bFyu5MpcLryjq286KsYmwVEiM7
acARE83dHO/Jgic9DOWgoWA4WyV3/3wOKIbnkJvhU20cPn+nbylnk7oJTlEm5HAZ8FZ5JS/N/65p
OHP8XXoj5CJGlCaNMI1iXBC/pkYtAoU4Z+ewOjKLJ7eBppq0VMW7HlUHFbmN+DXPgBrHonsThIXG
60QmOmZ62kJZ5OzJ8ImgkUq5SPR4002bfgxVnIxEvYF4M/cMEPYgUPo3XGZLeY+Mhu9OsmO/cdqL
OhqCvShhk7xBVLhKFfGNbjDCuSrnzZcUHlOTcjT+sXJflBtIXjR834BBU8JPwMe3tBIUYZj+nReE
SPdGlSPiq6Aq71bQJEvTlAsZO/tP87mWSYDGWcwQzfr0WxochGx5MXRgoEonP1PtVO09urSYc/eS
NDGdPvGcXQY3Ka2T1l9ADhNYpkY0zdl7Rxa38dJ+uNkO3QjCUz+znbDBMlN6BSxzshT9HTNw8wEd
wB8yaep83H8sT+ryZanTniIiXHS6e69fr+/wA4CbDOzflaPh85/PCCP1VHfvBpXaGiV/drLcVCbU
3Ylp1TsFcZ6sSUEgJQ25ZXO/eF/GcIHC4kFXgytjSKCN2FTNuGMELC4pJrpoFBqRZOwj8mM10Bom
KqHdgto0qsRknI0Dug8A9pfUAEc6OnmtORAKZ/w2rRNcZpMdIhh94ilz5QJybfLaAlJ+caeClcck
W8PBM3b6WkNKXvNxFDl/vLcB6kh3AGGGVAmpXgUx/2EbK28iAQ+WEIlvcUXOpsOmyX7GWnkUUsUX
6twcSv2DpvU9lFbOEzN23Ke/li5LXLAKBKL3+9gUyBpozzRn1Kqr9NlCqMwKyhNmB4cBlDT6Oska
I0SbaTt3Jh8zgAbMj8qzYLlbLHFBOy1rVqt4zfpbSfr6vAf7uf1qC6v9RVplTbKYibdOY7Ms6DDO
Gcb5gTMAGspuPHzQVpqNNnb43B9bWJncFVzz391A7dkj3ttq0zc9VKehJUIYGdw7Fa94OSTWGnLd
ZrwZeN8WwmkDrwnEVM09Gv6fCZLGmKJ27j5JJYLf1i2P+NVIxQjN76MQTZe778JpsUckZi2CIo28
uokBHhghzrtogZeAb4iB1LQdWPRtIg1zQHMGN9YgedX3c0rZtbMrLuliCMu0akoMVTfhFdJWDcC0
vDhiAgtPe4Cemn+72JpFjXzM+O43vniqP23o4Uz9XDoLex4DSgbRR43veRHdvDAMRzQSgdEOoCoG
1lPzT5zBXT9M6PxfcyXAhDsawoV1bVSd2arjQt18Akyeywa5/aZ6f5wStZLfWBngmYhjJanpgMc3
Tr1hfiIIYm4FEbCD3zuzcuhzzyrAtDDX1AlscGuBP02fuarZxFh/7oMTEyNDyS9cp5eEuCTI8YQL
htWY8LyI6m6L0/ldHSW5mf8NYm+OKJOwQs8xlGnERNzRx4ZXU0N9ufu8MTUQaPhdRNAMGE9+nHog
f9ifTatmTs2ecXRnB3m4S6SMQ6fHwvxH8F8pgo148u2UdzfzYP8zwLyP4hm9iZRqx4XTZTw+U8US
RXAjo3J/4cMEFGgBh6bTkFHE5Ta4s1RqbKF+HnJv3PWWbAFjQidp1JUDEWYXTYISa+tgmIeNiEUc
Cvf9L43N9qXCeMUFd14ZMfoF2LvGgl2t0kZs78TsY4A7+10PXCejiiREDMlg4lJnNcHPxTvbqKDV
GH3z071KQgdRi5mK/bSPFUdmhxfXoAB6alh1r8Pbrs55v816+Z+gXDR+ri+FB+YW8/6Ctzq97Mnf
MwRMgZD1iT59KT4CHTO8+0BXfSGFMP+UpxpzjGgWU5pt9y+Q2Gbc1j8VFKhsPh0Ljn5x8jmN25dy
1h8/tuWzwH23iwJLk5EzPkiajsjINadYmDb67AGBBnGsV1xwPnCJF2a6YDqJZCEUtFI/zCCytCTa
WZ4MHjVk1HIscXZoUDzvNEBYLFPPspaXeZGIBf12SopaDuYv8wwOg7aqWvEqJpO6ylAX8IfqJ2ex
4asyymlA4atyg+i3KdQTEVh/2Si64ZBgllPiM6wr4lEMhzv2daa6z4tLpm2/5pX3dP2gdhYzE/vt
LSBdr1ysRuG7q4kSwrAPJLw+ioXL3CrosA7UkCdWfC3Miko3NH17kF3s1BMghGHYdpguBELkG42H
zlBhRa1TxHezhOgA4BHmMdrs5w7iIRvQF8+P7rQgYm2h1Xx0hrCu9c3ISw+mwij0WbmC2sOk/f1R
9t//eO2TpdBgfsTUGE7lHExFblMlvzqEwf3zJ1cIx6e2qOyKBqKl6am5vbYmYZtFcQbggP3xJEBy
QqxTmznJGfaiigl7ZabT/lJmeY4JrYIDmt3kOzL0d+GnUCRLQPV6YaaMdwkFZpnPE8/ZcTC/DUii
XyGE46BjrK6r9xs+o2xldIuRFXbDd3RrA9HH66QBopaNyxeUy0W7YGkgvdGUs/Ouoa9YNVaLNfKP
dd5hS0dxCRLX6mDLHtYpSYoEIiJ9w0WCxbGtVt2mylGIPR9emxwokCycv96Dvv9qxlweVQPU9cLI
5QF1VYaHDJijtDjzNp6J0cJJ+uRGIC24zr6sXij913rHtZV7z5bfcArg8NGV+yF5VkxalkiHUOjN
KXiLOtfHmytfOd9jcQfm8PqGyMpAJQDikHD2zUuqrgu5yqsRr/VedY14ve5rXHJitEpqGdAbiFnc
Dv8hBu78uQTmXdPA3K7yttVTC7sNX7OCVwWujB5B1OKdnNo4uDL8N1SyzNReR+s4k/5m1e+AAEBk
hR0zKnoV4FFkxsRWquCauEUAqu8m9piek0sqCboSFDioXTzgCDAWwrR736YS54epRhH6A6zFBJEZ
yhdrZiRhFH+K+AhugtTLkI6aCS0xsY++NlC/poV2Gv7xpRTgPFhHjP9z9xZD5fFqvsKO4uGO2cRk
z9sqqfONVd6Nf3NcSCU7w9dEGfWSwGj8mJ2PsGy5PPJ4VcJ8DK+i8/qab5ZiLnikS5xWSw0ytwbB
5axs4HfRU3w0qASS+ixpBqYqzELhqdkKrppVgqkC3JQQbyCx/Myk8DOwLLNy+HNbUXajVXjy1p0x
QWXSaOeXty25OLqQiyAmDJ4zVVYvRpLrgsyJiStXoanz7ilIE6aOvJ/algagL6t0yCLyySh+JDc7
Ncg0j5KPmS4/mtoAD0ADag0UV+KGodX1J6kRIz7EiDWvnPcUEQ0J6VixZpzAmfPdf2Lt2lVZbIqN
GxFNTAmkcNzccnrHtmVFvhpdcTGDi/MhoTSR/ApFdYezQcqMxusH8ormoxAa2KaOEXKxPDRdGaFi
EiQT+WHijREvWCmFAbR8uvhDwlaX21VGbhAMOuo8PGdNYQzUW8wdaF2nTs++OChzI7W9F4vvEfmx
fYBcHzftDzMcd9tBa0KifO50XB5lSX6g0xMDHk3NQds3/858hAOZojuxAnAZVckbfpa+QrLbupDO
wkyKAMVWPfw+iPSS8pIG3vDlmKDLag7F4scdjFhu6ETMFaadhwXgBRQvhvMN1ta3pwgbRQFPgkZ8
/04cKiEFXPHT6tLylcgLX3OXh8ycHnlqdQzuAJc+pMEt0clzQ9+CyLAN+UTSZ6Vt/DsS+IbLHUVc
3P6BIop7YqDGbnwPn3hSaCYtveA011YeBhDRSgb1/d01LZDAs3laeq1hSDiPDMl+VYFjpOfkspsC
TD1VHP66fFF3doVGUa8oye0JfRwhNdqVqIXsgjyc+sk6OBMdglZl6HTKlaJaFnI5UTSqHM1BZlsU
MsFWthZWpxk6RZZMLdyagv70XgX7gO4DBve/0fqz0k4VOzwyUjQvpPINELm6WLlYMT9et7fCLLgK
600wTJ7e1AS2+GHPiOzztoJdrH7IH4tvyYbx0kN9zTxAQOrHxPZfjqi7q5NhsPffXEnagyVRnIt1
y3pdr+ipRNSA61szeb6d7hcE+cGsWlGzaml+yI2svryO6z8MzmP/tnAU2YWUmsPhYWOLfPsgrbb8
E2dxWz4PXjqq4pjOdSiv0HuNI+iqAhrzyotyPjdHC+fCAb0fHoFVEAHSh7qBDDATaO/JGQu1JHfs
SGIq57/Ivn/vtJAxj3WHd9YnPSfShMtJfwrIY0TxfDGaeGM1eZmOB4B92bJjswIe46Boru4f5gux
3cORfEYNyIIauhIDErydPI8sGyPIOG1JGOQeCbHZr1A4hsLjpUDSb2C341QA2ir4hWuOMZc6m4fU
jit6tM/6Zp3c5MUHJe6BUGG3+CHD6PXM47xcLTbISMj9TqX/4jQcO2i2UJs+zm6sTWKh5POE/5wI
76cSSlNc8+e/5ZGRFn3V8VhklQwxCvakPjmiCYP3+Sb8gpB/m0lHXupT31wlv+hH3fWHssM4dr7c
cbaP0SVN/9hG+fVUF2t99fMnvPpuJ5bsg8QNqB/zIM6CDj8L3PXYI7nEPyVMNtgWeBDi+w3SkjgB
8dYJ7wQv1pDcFs1nxI1NwVVs4FzGMfPV5z2XoYGKWLjHzaYBPcj6xwrmppRirmATcuAniXqpRtjU
z8ByFEUn+pX5q5TYV4qRLH0btMmGq9rJEK9vuiXh2uvWdTsSQOgJzM7mkQt1bb6fyBcA0YXEuTkj
qE8A5VoHyfCpotzL9ifB/auhkQt2sFk/QugaO9jPtdEExQusU4lhjI1z3SncWzJriJo25ujCpa6R
/GEA1yoZVJW8mhpTT7f1ZMjg/rvkDF+/AkRpiN4HtQVzzshL/u+50qavKt7qVHuT7524XI4EwLxA
SyZS/Lufp0EQCK+33lNUzMxFhRt8wWKCnJ4DN2meXkI7bzmp1toCf+QwybdJ1YOQSnVOzKqndSEZ
i0B1M77FA4+wZhCJAdvOLq581ZG1wYoreB/Wjd41gnMiS+tj8t7p8kj3bvEJCMTCrdIoyP8esKoP
kHFzMbX+k3CfLvAhIrDuPJ4yextcaPqY6//e6RYgsXNLJzb20Em3j99kNR/evIZRbvpWJdvpztg4
nOhByEDLfVS8C1Xm6XPEq6tyYGZbYPB/ykNYXwlhtIAP/FF/jYSFa6pWa2uYQqAHNGN1bo6nM/u4
eCsZ5f0UNYzNGky4MdfsdnGhJNDLqfy9wpcuISbiBW5VdP9Fel6alMs1RMcgC1twJ06rGRx9KMtS
64moEUxxktGXGGtkR+xh7Q/uZoQuroRFdGq7IVgM3Z5/UjMHbSx93Ui5xdHkuYIDqb64Kz5Qsl4O
GwLKDug/BwbYv/EFbDN7ZaVW4Cqr3alFnJbtpaTiVXQoOuGfK/Re/I468+U0o746MzvZyeOxSvSB
rBpAs6eEUuCHadBdMDEWkJ+eI99jujiXxlf4NVRfea40BYmV/wRgMnVOOexXVmvvLo6uENvmIca6
yv86Ke9VF+vjzhPfWNJ7D1A07nwr/ANA5vSqc4qaiLS8cyJmyIKnTDTkHnlO5C7XxNI0OhYWONmD
7z3QzOa6eTLa9nHGhkUhr2c16z5/wuB2qVnYGkObQqJYZzdpjBwvRZmUaT1ns4FTAav79J0GdFw6
C4hxzIGKjiP8JM34/Q6aNxPi9CGxg+4/9EfOCgqKI0j1FptFF3YRTLZ6LOwuc2CazDduS6LZjNeJ
9wb93q0BcS2uP9lXWa/PIskTR97SFrymoI2nIJeiqsiNrz2DKBPwg2Z6YXXcBlhnVaDv6c0oGXdq
dhthY/zDuccXeWvEd2H9NDgM3g3qVAjRnlSGts+ZCDUV5/Osm0dSa7UrwAAdF0XxkRU5sDe/vpXG
1PskPwZem6d1I8BkucpVMyHfK2UJU2YWPM82flMk/TyODPNKlEEpFM62Ii7719hnl7vkqtE0I8fL
yCL0vTJgZ0t33z6gL5riI3nk0k/vzKJyU0ejvr++U3++9dM72nXTk4JQkKXZR5iytGTZzAYFe5YV
NGKewyGZLzS5bCSwktVh5x69xYyZCgOig+nzudtCU3vEbFMp/esvpA4jRh068iu1wS14L8cVSpwy
Fyw6nbujDni8l8TuxUDIqUrgAUwNu2/52ePsSbWqbo+46R/PRBV39xBSMNawOgTIKrVqhfrYUoDs
lmlNqp38G/8NGEB24Iqg6PY4LqVBtAycXznDrD6kMxDJQa/MLk5KaQ9QNJr8de/JP4PDknh9EeZP
/7k6dfi3uDhrTR1lBCFXZuY4FUHqLwds95PSZvUtPFnGhjUBpd9GeX5snsmRZg4D2FdbHmCUp2pb
Bvbpdt/jTlDUUHxToT+ZeUQrwQ4ifFPwZf7mIp5U8zBGevdirs1QhraBZt4I7UlZtP6ITHUJSmOl
sNgdLknGhk8K4+ouLFxtXfAB1a3u+rL/EHI1TjckBNlx1pcgSwn2+PGey8oLVLkethG8tS9V08mN
QJ7zdDkcgrwndR3tu4nk556g66n/beD4WdB4QWQ8JrTu1A4H8AAS/+fCuYA9hd/ZR8N99GAHGm+w
UOM8AGSt4v2TM4SgDgQCjP5yy2kC2UlY4PQoPqwtY5vndkz5yBhFMwgkVG3DPy8N8+sIwnHCZF14
6eC08OcfwWnoiIa4Y6UA4dQ1aeo8cmLgqARPuuTNb0xWuBRTItqjsdXhWULwmTCmMr3knFK0WUiL
FUkp8Clf0IjPLo/8bLQMDIy8XYm7OAvlSd7EPl5Nncr/sOz8vWokQ6fD0CKyXALtv1XC6wKsZ6HM
enuBMsU+kDgDGGQt0eJLcm9vo8tW0idDB81mjJ3wStcMFyx5QkLjiPT5FJnb2qc5jDvM++Taxrz8
kJ92RCeyaHJyFTxkdQJBqi15wGnI1l/OPRXITVvQ2IsBUrquvNR2yDLs9NWHfvPwCeL+yk0w8ogD
ecWwiQC7ZFoQGyarco+NaYbH4zfzN/L2RZ51xWEQLpVhNQ2xjTN5nEOG36vu+Z1H3vL+XbDfX6j6
L01tYFV8MKeQnewOyHe08AOxRZDrOfSiqY7rIYOBBRIVUeHzCgAqIQj2TkhGZ0VpIskBUagt+bbq
eIB7OjFrzAzWRYs5UGCUGMvJPMXR4scSVMXo+/KvabOGafv9MH+Ax/51p2GBWrZkK3FLVfVe2wfj
26R4+JZxuAI50LLdw60/XDW3mItcB94plHHBPjsAoR/OHx1MZc1ca7cf6YrFulUkF423n0xdZn0g
r/1e/5NY7IHSoracnRlh/BiVIzQ6IriuzBR0LcaaxSsrcvRTfALqZ+r3WONQgI7Xxk7y6D6KcCLG
KuqUfZc0odwBrU+zEq8BjU3cb+DeDckKyU1ItODi3ugPBIs24Vpd4NGD972WGw+o7i22Mgaw+zq4
r7rSWCI1mIZLN1nnZjxpn4sPNmNHtPw83P/Uel0y841iICVECaHT6rw9cXJ2uwvdZAqwLS5ulCgo
QSjcmQ7mp5PVilo1/akd4OL/yyc1leILHMHBBxJn3wGpWzmismpuK4s0/fh2HTNoCQbB0z97dWEP
kYEPVLA73xEIvwT2haLoPT10SVybqfjERDzKi23Kt2s9akIic0hufQsdXx3Ev7xA/K+HRYziRCO0
AxE3/5LiikVs5OPo1lz8ozbPFdUO5ZdUp0LodPqPYnz8SxRysCvT1lbkgY+rLZMhOF/NtK06Nu3+
XN9uwAH2tEIdcQWz0CYHKxvquACxVhLuAGuNoEBthDjfbQv9dbtbvFZFzjHb5dq+K6bh4ajQsgfT
sb7cnWxjg7duFJSvvG3Un8gsaaukwPmNMkukh8gQxLt1N1UnSQOIt3/ob/TZb6ejqnfg2FBzY8yG
7LDxsOReMSXwJTIOQQgVi+amLbEcazE9Le55eivleZQC2ew57KNAkpk8awNpVyKxSGPiw6xK5DDF
V99pHD+sSYJSzkwhiam1WcVXTf9EgBT2mML0zYPgIg5Fdp8iBbKm1zqCVx+KZjOExFmYKuJJzYok
2dGdT520bpbMKxkDzwE17qAD1ctE5H1CcUejjwaFyFANlfr9Tf2Y/VoHNUOmAbHcZ2gfnuV739vb
1IPOBpGvJafLvIydZmGuuqS5xch3y+hEB/DGE4uB7jwdUYwMx0Q/RLx5IASISnVZTr0SyHsOMyO3
y4P0AKswElPbLlFJpPAhuLuiZOr99deDez/xn2TXwbCuYLxCF1KTNC0tSlQpEyGH7vzDseGiS9P/
K7xVb9bDhA1ML5zFlY9MeniRaBv8NiL8dJzVuDd4BUfQXQbTMl+Z3KZoC87kL6LcTifzYMYJhZxl
6Gua7+jJZEnkTatrcB+8Q7pupofVDozaQealG6k8uTeE59K7Q53eM4g7n5NStYkzMhwQhKYGLj+r
P1uF6siXyFCRFJjEayP4GB0ZMNleGKrKqRozIKLTBJj0/MKgAFFx2Blu+R+l51rV+ClxkhsbmXhA
1RqNbRCDT2TsNd2SrXJH9kcGB4UY5PQsg5Zi4rta9uJzbJZtoAoMsGgZjgBc744fHMGNLS/NRDbZ
wUncSB4R5OUKdjSRTX3VG+MqanixQNUtjLGGlTjGqTi6t+02baPA8DmXid0Cmk2z5PUG7Hpp3vWI
VC4ds1QKZ4iMDmDXw+mwRZhjyhCQ4QldP/rOAoTJUC4uBr7HY5ovxKgH7Lm9iNL9XozVkRmma/Ud
znODoxRQdTJshzSngWns/g3OEBvtlz0C8V/PC1po6+xhkv9QJ3Um70GxjFb4Ok/orlzCrC9oQVw2
nUCm7W6WmsuMnkhV9t5qvE9oqy5wLa3E52fZAmOSfZCWa1t4dgwQf7cmaRCNFHN9sXJNQK35NVB9
Fzxbb2tdWJA3fZYpAEzb2ckvBZOsZL6brX7OLyfWz3WXUD4ngB9a9lwfhRjOeN8Yn4d0qkU6leqi
eTePeH2vADU0AxwNJERF7KXIOiESee6qPnMh8kXNIlK4PpNKdfHF4hoIaLqtmGn5FDtdAvz/Ca0a
LxiS7bSEWfQ3dqVYbz+YMiwbE4AikBLJMweAU4/pHoCvDs852j7kzPIAtdLlGan4e7nbcRyQBCLI
59f336suckFJkO7gZZ/09KdoIq1SgsjxCGaDz6FDW4u8Mc4kqL4g9ARq6ZnSejfWBxXxQgWZwu8P
nLErsJgg5y7psF0PHyqsXtOASIg1Oepw6tg6mXZ1WTVh2/jZg+7EtSK6F62UJQ8TJSy0k+gb3N+x
GGBTtyZT73gUOpSZpUfLzOJExxixJM1yC/8y+3tiaO+HDcULHuqKehpAATDXOsvUeds8mGE30m+I
YDxFEG3m2G7cinZzRaOd1T62/T9jVf+bhv9m6djIGktvYcYwCRmixgeXUHehAdiAFlBd3RyYY8II
M5SirEqnEfOB7JLXGWONi6G9YF8PHSseptp2wi147t8kE28z1gmxTrzVQ+i6
`protect end_protected
