-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OATOBFg5g4SuJ7WHIgbnGRs2mSzeWQg4MBYplju1/Q/Tk9GkyvgvKi80hbrDwjGtLeyFXjjB8e+k
U5QYjMsXZygTLOnkZ7r15jCcI7uK7+bLit7Nf1E92wHXFetzCkYPNly9uqHkeG34MA4UrCD6ygLv
DGxfCxdTHwkW/etXxVOtUfAcGoi4Bkkq24gEUqEnbiER6x7Uz+2R7pJYv2a16oS9x3zt0PmKc/ee
ir2/isPmrFcMNtzwWL8L22GHtO8ALkCIzEBd9RuJ3vNmuv3FiZwfGH0Rt3B5HhyvyX2OlghLDwHV
4F9MZqSEgKnXrjObBl5b4S7DFgiZlKKguC5MOw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
833XeKUtLS/wubZTBDkVRdA/bHvQhoeSs+/iZt6LKdSrN7fLckozw9AZpRccEtxMspx3fELuE66e
VDECTYxLrzmPjRvy9lBofKrUj96dbY5fmVcHY1FociA8tAaaDsRmtn6WnLGdAZESFNA2lj0QFaK3
TKUYQ7k2oTq6EPHUOx/NRjT8SxveBFe+2H+TaM16y53qZztfZ4xXLNJNnrEo4hsNQBKjiYgWMW5k
VaD2/cl1Fu7S3C5uBkmswLJjh/kg4eh89jntN7zH6FHwbDaJFHGIHBOMUVHn+jWR1PlF8D6Hfcyi
K0bUBk3yFKWvLk6WBEQMF/teYQ6vcbOdFPQphfBqvB8tziNz/ZtUinBUsIPcWxoMKC4bH+6Zd1/J
JuLo370dNyQ/Szq8M9pYSeCONXhhBK68AEdj9gjoeZdFE4ZNmzzFqQVroUAa3GIx2QRnELI7iHlW
hxtNV2F/Q7O5K/SfGfPaVHvY4bz2UhIhgX2A0JGLxa/F+GxLD1K+i3hbIqKLkU8L8QEtUbsjCOH1
Lm1fbG7zPCjVcJCDU5duEaNOEv/UP7Tr3PwnL2il/LK1RqaY5TWyqWp+wHwV63/QiNuC4882bRs5
j6KEElbwJiSbs7+1IAgEyMF7ZTm/MI2aASBgLhqsTD72f/4xFk99yhT/tfL+TeMyQ6vyJfzuR+v4
7OjVZUOtH5Y1yd71unBoGI+Ly+VLKvK6+tAyun3vfjUQSqe8/O3q+5qcVtkjJ8k7HvWEUo93O3xN
BT28jptLfp9dT4zqvc6iEVaJ3umVq0ZC2ilCSdwmFxajIP/RFddH6n2LNyEOlwSjY0ae3HEC0RAR
YTswY3T1+r7uga2c3uQRGiq6MsQ79hJw2aymGI0VqRG2lWCDTbeab+TjHXEbV62ZNffyiFpsHh6Y
B5EKTJaLViUpnLkg5i+tt7wcPfVw2iK5dAlZXKK0K6Ou9qDYfD1qg+5N8dU+2N7SzzPKT8F6JyJV
Y7yvhAObWa0Prigpb02rnXLDZo7up/8cUOsrH0YQ9LDXzEYgYYADqPCNipfbii9P2Af8xpKu9K57
uhyYFzMTE2Mj4aO/atoYK5XM02UqwA3KqePu6dGyKQd0vJMcsXWSkHJFalpUmldLkiFjHnubYkME
SbI1i1ofATn5BoZGld7w1AkMu5IdAUlUrBqVVcT6yVZ6/V/v7QgRUbKCw6MJ/ihRQoiv7h32yKcS
MDoDIKxVqXPIiYCpdEXF10ADPdroaTLIajxuKS8+Dk2AsMTqNCSKPwLCXg2wrBn2jYxrNSE4Chri
9SHIgAKPgImhkAFmYW4LmsERndYXasgHa+ht6+6VNFs5Yu7IjETenOjxuEdCu7IMJ6/qLfmEOtZ9
1+NkydylXmKZ3g9nrRVy0Xo+oGhE9H09H/0iXZYmTBe7uXcr7GHXDjygPnOLll6/Pgly/1/yTiQj
huz44ADITq6FLLUkFXuavcHU6znQ9c3YCgGLwqCKzP7/doe9Ka20PV9LfM4GAK10rx5DkQYkbngt
T9Ad6GnmqQGzzUGwP4cN90MiFs9DHKxfFFnfTg6wVIUTv2Hh4SDy2EJ+HLi9Z4fASlTaaKyar05T
NRKREw+DRu6L7nkNq1UUOhofDcxK0VirKO3C5IUVH1DVKKumf+UNi7aOkuQGQB/sXwXczg+4AwOC
QGlbKZxGDe+KcKzgO51hJNH4gZtapL2gN2mVw5eHNJQRSXY3vI8ig/M2liKGqz/WSo+/OXKr5oa/
Rwj+o4CQJUBdC4WEgPt+OsyAHX6NyfmvzrpT4Gy/hZqR+1QMJ6iCtDobH+bEoiL5Rnwi0SkL6lLr
GtHXWXMZODKk1SWerHifkDuD0oZw8WntJ61NrBptpnz02x60BsflDhwfGHvbPoO24ERXiva0ltJa
dhVMVekGcfXcSen5QfE6AUvdZ+q60GtgndJeHLSekTbqrSRyRDJMiAc+PBhF3hLVB406Z8lquA0r
j7+YTL+1z5F3Pj2b5h0RgHYwi1KKhX4gndl/LeM+5FbeUQ9uTSN1x84P0Gi1jvjvXboj4jEuBfDF
uxcj39mQaf/moWV1oF/M7e2L5PIjwwljd3NxXu0uvwFAMdgVQ9l4fp+Nv+XphjT/FwMFm36leDmP
AxiMdeUr+SJl+nQJ3soo6kt96xK9L5nPRNw8/m73h2ncvDw9C5Xm5uTTi+93ZBkALsmNV3ukZYZz
K1H6HYbd/5aOcaVN183XUBLH06kZilVSKAAr3zWHrdZaQAJdnfA7Aai3ufeDkUGXijyOqWnfZhWO
jnnqbhrsrMLFKOgK7nSF/wB33eU7ijBXUzLeApnXLfOeTl2BYEY8vgOTHOjOE6/S0F3vTGXF9ZP5
eXqggfaNgdD9jF5qKPxv2KOtqosxAeUltg22KUKDBGIW0fgcxOHxz28iVoqe7q2L+LZkWBUI0Fwb
jQFruDXGT3ZjdsgEfcVcS7bjG0LP0oWKGNLCs0yfY/msg/duUtO7xSZ12CInla9m3F0K3sTew/IU
iVCD103Wlu9PerHDrVTZ2RcO845XGdHH7AfheQHnuC2d2iD03XSPssbYOgMzxvp1bKT3L5xshqXr
7Gdjr/fJgMWfdusQ9CPnCuiZUlmhKDpT7Nq0u3raTxT6ZQ1rPl2rtVzsH8BvOECQqA7yPRgkvXvH
KE4QwGGKdaAtKHECKP/CHRc7f24gdymemnAKVeuNc1cAYHd3rYHyaGCkqtepBxYUsRzGyGGFwW5/
rrCVjPMnVeTwII5v5i5imPmjed3HcSqRgRo3gxZyjMJNBJ5/TJa3xAYzVm8s9JvXkpyEA4xGOorL
HXt7cDa7MZsgsXRkOuCidHPA3hW/MPCKkUEQaY17DLM6iNmcU9UK5kXke8JmlrrsPvEkpuZhb0tl
2u7sE/Bh6i87INyBh1d8z/IGpgVp5MpJDQ830pHsSdXZiGAUq1iipkl1FLfw9ZlbNLCQquBVBc6m
PTqhvjOU8SH4N8dFyA6AYSbferbCAbXVj2RHnZ77d2s36SwdCwL4mhLgD03whgD9/N5B5ZUwW8fd
pm+xhiDylBzAhW4N6F19p51rgKIDGhtur0scebUZIGjnhtJ9ooIUo1zTXPQckyO7yrJN0Ip0a5hQ
bqHehdXdVXO/N9UU5DC/YtDVPZrnS6hgvXXTLbmrgPS1jvjNgB2+NDRI7J73UImN0hh60+nlH+0f
OL9aqKtq+HArJrFj5sXyrZWzsxRQaevjpSd3tiwW0JB/ZTVfC2tJbmGlx/GxG2dn7s74E7dw3eIk
drae7rPFmvz//bYXISxrnYRpLi8zAEymMjV5RaKQlCAuu8r0hEe5U/1aMwkFOo8hKwFtuv5gPWfX
KublMcCwKIk64HzeXCntmvwPO7GpGqQa35LxjtBUwhcBXntZUugwGYbT5HgHSpT6ngI4cuuEuqIm
vXCRXPPzie7shw3hdXxVPP0CrQl9iCudwTl5Q17p1T0T8JlEVJf4q7VHPNVnzAAe5oTKK83DCHFF
MR2ekWCfOQGgP9euf2oOoYybcfEgTIu3JHfVlfdmlRB6p0WGSZzLLemB+aRbTMgXYrH3PTtz6Qu2
Zqd5s5Kz6II4cZ8Rl3fhxiNZYujQQM7db2cddGD4hFtXB5C4CKxFxBIx3SixWFrErw0c43ZjFdMT
xoRR86GE95Lpc0jOlRq6P5uPiwNWo/wydEosvQ3OweNxaGeHtwUmrq2Z5zm9J6UhSHysgwG0UVtD
A73gr4W2K96PrlK/RoXD5CVY+Qdm+iMJTnDbXLFM+QLzWu7JmWFvrFNOReo9btv7bLgFIyebl3Xt
97LH2UHbfqRdb27+q0QxtKYpvd0miOWiSqL3CuhgOeSXGnopCmiJMjo4s7DzcIzd+jSuoQ6JWzPM
7HgpNaeQyDb3ZK7wnl6UeEWqvmZ/9q7+HiLCMc+l8+IGnEYyK+4PxQdXnj6Chy0EuLiJeU8f+egI
quhv9vMjhk3PDrUgdqdAyb0z2qPy8kEJnLWM8At3DXHkdGTUlNmZE6yaNJM7qDnEVpiOpNQCyHHf
GO2Qe2+RY2Fa5W43jF2D3zV59bAAHb+0uX4CQVLz58uD8971ERU+pRYaefCvzoAbW35JhwGdQ7VH
kGZBbUnFjdhszkjUCR1aqlCsinyCSIhfoN2o0FxRJZQ9dQuoHTL/kpnEGKIyrKeM/5BhIGfOG0EA
qveUnhr3FTOZADebm9K/F9BzOaaluhUvHX1B3HAa8FF94FrBpqo47DajDrCCvhBiOizsf6hpJPY+
/q9pr44JpMakqG8kXy2oRY14Ou9RUGIHoHotJxpdVfgsLokf2F1Dft5Xg/YQf9VhVK+4MUqqgzwf
MOmGhAqW7w/IoZuSP9So2Hr3+ciiHweRxLRfxalXy9wHuzP1sjHPhZds1Z0Hi7rXLteLxRG/3n+v
ro16WFizllj8+ljta9S6jID83NiZF/OU0L6YQeo0RB9WR5Z1RT8urN2vmBPldt8x9Wyy13LmT/0L
TIsu8dHNQ/jj2QfInVBZSjUbWs1Mt+tk53l2NP+RHVRgaWmvOYHP2+VdVvmnvVLwD54EA/osmxBc
r+u6PHayQnLUkGUPzLOXMjyKbGhSCOiy9BrPbnohVqx9FaGZ0IIwJz26l2gl2h/TzIQO4Mso2y6s
DgUjm470Cra5SyT/TXgYwq17ykltKxCGIqS7Rn5mniZ1Cdu2dZ0Bkis+WlSZYX2uNwiJCbTAT4+R
uBq8aNQZ5EY/E3ygVDVj9GXi78ILbhZFGq4+V5VNn0AbT+uo8a0VNLZ+hQLvvFSK1EABwzN72hyo
hzvEHqIW7ZJo2Qq5ojISDN3VWBhFTFbaXSG42wUb/j0LEQ+m3Lf8chYU0DyJMmFAwM4SlwdU3V3u
792oM9KunvqyR/H2Kuwqb5uX1ODz8Lkol6oKW0EHZIRCLGDWVYblcrxAPwaDggyDJQ9DocnZ3pMJ
8PtGaXkzcy5k4nqM0mmjdozYWR5gR1Nd4cfZh1iDFoMvr7cnGvnHs2pQY6LYv/bT2mQbEWZhUZ1r
OvHSchB4GvdCVdVPg/0YCBGk8TkC0rpeCOMV1HpTjXyF8hZ2d5hRO3//j6wWqPp2qzNoaGkL8pWR
jhx7TdnKgIFAa1ZBkVUUaMFL1Qccoeym0azGJZRAIwS0CWQEagZjiScxj5WHHmctFjjd5+9F+soK
w+Puh12yLEsBu9w2642+aMx9eX5V/Qq7sX3klxj79ZSoXwc+YrT3lE5ipu8d1h4FXoWWqxUnX4N8
EGpYn38Emo0UII0o/p5TTR491vzXR5XVtda7cehqoHjrQFikyde59u5Sr4/iVJ+yPsOJz+FASQMJ
cGaplfDIE6K7PlV8h6q5xnAGqcvaWRiPEZDgK1mB2TjLVAiYA5yuSQTV7dqMEbzkqiAeeEFzD3LB
2U0fYJjBxrRDp8KH6Dn3Qqa/11IJvw+QvKW1S7N+0+eFklaeVeevy3yayyZ+tsAbFMKq39s5qIV0
YrTDuwYmz3wXPc/nKu+NIV1oCpJI1VjqRR9bFtpnyDYZfWWFvcEbW1OKFQzHK8ySvlD1tIpGlklz
GfNKUIY8aSwogyBZXX5Af2YZe60vXERZclRwX/7jMwh1+GJr8rP5kfAdmEsSizrhqCX4iD2x8Fd+
Lqb0xFxa4yLrLbZwRG1gnt7TpDpHjVTKibXxuYN7HZLXTgmIaBzcTy+0oEOahFTspzQM3wffGKpo
FJ46jyJ5/otYm/Nprjt5pS8Lv/zHVJ10iB5pFdXXZ9zTBhRw2ozga8WzQ0PQIml/9UHA1PjtTbcd
oT/v7slRbMxmYRXn4QU4pKu994ey5Xq72iDAUSlSMwjN82VLoTkRMv6/Q/aCd6DRwkEksa9pcVxY
Xqe0aGgXoJ7/mClnford62zX/nHtXUBOwSkESqEs0fQBaTlhpB6fYWHqIs8MdJOPy8XOomOv0/p/
omuvpfxjRRbIEj0NDxuxnxKi66yt20XS2lyRtXr61RFY3UYDzhdKKqMA2O1SreeM7WRI157DvCVd
xvlcRqxdptTRqSjr8TNNMH4WJElJkmB5ewqWsy/bcGvaPIc6s/S1U+cAZtwjDcf6cMI2BBu2eTua
eTweV9faY0L2uhmiscODkCqilke0LtPjc/BM2uz9rT6pMMhKmDucLk/9SOtDZqoyNxplC3gczT3O
0ApeoOHh10v/ezIKcWbprsquZtlS/Nsa+FMPpItM/JQmDtvSXV40p35mK5icWRE6Sc0j5kudl7DW
g4cQ5tSpE5T/8v79VvQ9w/ACaBoUPls7z/IhT24ReIShKeySuIQRIS7LtXqb6OJYCKskgN55znFB
woDI2Nw12Skx4I4Dda1bBRDl/FNCmZ5fCY7MSCD3YP3hvxo/sw16jqcaB0Cq132GJcOPbWDc5cB3
pVWAu8y5EHHJAE9PrZNRPZctTZGyAV8sU59ftzgU4WX3IEujoozni+aSykJxt85R2U2luMd4xGow
/fUv2MU5sCUIyKQ4ru1DXfx0J6EoAS0are8t9X4+nPX8l9eq6dnjXicDNwBM4UGXZPA0kGUXxV13
YlaEQ0caCJN+sAdaIygB2jX7dwmV/NiVLOQk51jgZx/IHiCL9cyb3DTOAqfwKVO7n9MUER8UpqoP
igsGYcyjOzbUKkZgNSBpbIZrw0rXE9qKDU9PbbTN/PkhIByfTZ5F07hQZqmFG0MsXMIpowA9t8SU
khh8QIwK8tWuAZ8N9r1alJcSX7D2GQPy1CKl9naJ0N8ue6eSTvXDrR0MkjcgR+GCFuIhaWXdgour
lbmtXyuOlkOCpZ521OxS8hOOqo5Hoz8pzbHL3jOWie121I55FpLx8VTRzKfqgGvlRqPwOCRgkgP4
2XrI6JOqBtTyGtXl/vErVJDSFIShef5dNd+JSxWA15NijpYemUZzO2gOGa2DKMlfmDFxWiDQni/J
0xVvucu7guIYeeZaZ2DFBnDR+e+JyWk3ppcKR8+6vwzuLsu6bq55ab5s4BwIX0JZUXy3WnG/W21w
/I9OsIVXGAN4P3iB0riwcBCqAUb4QLKPnv54KhPAS1oMms6JavvmYv2gu83IjhoNOIziYO50vodq
j3ybSo/sbL/ardQCv0aOV4CZPJiLTJsZX+/7F8VCvYPXPbyJkgd3E8XUTIlt2wQWZXjHhgCOgQIb
Woc+rkJi4tXfAe5eWLArp4w0POkXfLw97TuGNyUjS+y3/QcOvFSxfFA8FLUoEnXXB+ZGqIxW22pF
jCGY4AA5alL9eE6yeNIwJjG47eUWyyhZxPqn07h8ovfwf6Zw7FfPiDQCWgDKLpIzrRk/Ar0q9LlZ
tqhY+MzR1anxuqWZlz1WlVxYhABAwABfJBr82bag7WU0WqQZTLJUysDJ9+r82ygaHWlsOGqxG8bi
KB6zLg7rnZQIEvKFWyGdKSwFt+b8oJJ5WQgvigIReFa+bgzekDKisLLtMkRvX8VWSdZn9yM3mpKL
QaSc2J08pbU9UC77sddzbk5BwtJjkPeyfUJwhDXkKHoKfQaXW8geOplxGjl7+l5omyJt19TT8RuW
gW5jdT4JR452WNrIgAikTZHCMrtN8DQ4tB5CPuRTJQezsZSYPiG7y4vqmc/q7gMH19mw5fCtKcJ0
6o43ObWX5EvIFJli/2jLjm9UyU1KzhLRnz2EUOnr3F840pIDV7Iv0+lie23deShsY9ujH5bPcr9Y
su7dnQ6w4c9uPUD5dk9Wu/j/UY9tLJOFCkUNgdbpXy9FmNrRqsasLTXHpVpMWfGYGaD3K8BflcPt
oLxXd6reG1u85f6itcG3On2RCY4VGXF6rBMY+Iv7MYZuEK7wPjAXaF+C2ooD3SjdQ+YATEJdIoX+
A7lmDbLoSfZrsTws2jyaDpkdsH7DS8uvzIxsgkSz5uiXOCEyK4ZQVRdwh/t9MFXWOiQNakUkiDn1
aRjvdc1HXs1Urk++6dvxmCrUXRgqKEJM2e3+IQkdvPR9/zsUAyi7Y29blCS2V2R7DSI9OZi0eD6k
VyJa7gcw4YFqBA0Svr4XHtoICX12kATNWy59MAbd+5ZmSjIX44bHSkwrF4/1R95U+iEKa82XwlWt
yaZbVD166vTa4qicWNycn6rI8egjzEJfdI/GZnsPcK1ODgu+I6dGeRrWAi7+0o+Ga2JrivkYp+L0
lpQt7AV4CYOuzUDnmvMgBgWF7LMa4TJT8QrjY5Di2tDpk8e6tYdN+mT2VO/gGZooXITh2J07lA2N
xgGOCRBsf5fZ47aBX1tgxgx6xNIfBvSC5qhfb9h03JhmcCHfRhlIuW27vpYq0filWL/l8W5A8d1x
6171a6WFMYTopODlN0tmxtgIBfXBXSrVsVfUO66daWhIJme58Ic0r5uDfde9zPZbUV/G+1qv7TGd
B3v774f7oTqIIil+rGW8IOx5H9qjvXU0jXxlI/IhpF/lrnKSavh7rIfB0gLPK2movee4s4mjheeS
kUJipNZ+GWftJ6PLP42Xt2Pj6mLambHGs6xi2C6oQVXJeh6e8wa1BXmHvvls5WgCaf+NwlK3jKHI
D+A0hRClCllc2aTsDYdbnP74v16ITMCMAXlqLo7waZpxKuY9UaawkQOKXtbC8km/86vUx/kLNv87
V3J0h7t9LJfi4GcJ4+MkK5z5kGSQYEzDfFNHLUrUUma8OHqXGxadd8H413tuhvAWpAe03RVccoZk
5TOzvn3pguPsMWlbuBtbHPAS7a6mPXk7QpOZaGaCjBs6i4VRMtMzMZMBFV2CnZBV0GRh1+v3DP9b
5IquL4EFHPc77/QvMTNYZPd97bs4NS1yLCVpZKXrjl85DQqy/wtPlJ5muTKQmhMLE9mFoG/l9HSD
/VOKMiBVL6pdUpFPrAcAl0G2FVZB/eb98UYiOAqRU4oceC4L3KTX2s3IScMwhFhiDSM+uAS7bvZk
4uZa2+xJpef+JFyAotnMe+QcnBNgcAjNMxeYaB73mjwNa0Nb/EoZ2JeH134Uqm9KBSOJTKtHSJ02
xlcwYwEA35PcgkwfBkYJOw4d6e/x4XfSmMb31eIEDDLx8Iop7ktsqEY6fbiBvQ4b8b7rOGop3FdA
kvxVs7RX96cTyoRLZlUHp8cu+Nj73n+w/NXNlS8yXJ2DYZCAEHdxNFvVgEXOTdNFBUYgV11lBuPO
FzyZcE6tKSvNWMEFq5sR/sngzQw/8ia9dtO1KvTOCD5Ik7YW5DkjkCjVQB/kwWc1Bg+HbBV7+kd3
BJfnrKUBC/F5i/4JovaUnNYt/eHiWh9Yjpgv+BWDzFMXYeAy33tlOylefYBIDY+wIoaKSbpRKvKG
bl/3omA5ibtPYLNV8ZDYh2pXYG7TySxZRWGLfw2tp7ATzTjb0RCmIOQ5/HTgp/hmbVNuaVNJwbZd
JDSUn/FYWcTqnAksMffg/pMgeOCwQtLwHhtzRy+9+lMAq+UEi4ZE6/YU4vu3cMoGccWWrGp+EgeX
hLMX9gN9mnzuoTZx7tU/RFL+FPXUZfOYTLdYlqkxCbLb7Ny7lPi8wgglQjztP5kxfkvticsWVuN1
1yze23oPlSSmmy5QMGlFZqQXNW/D0RZgaOW1rbRbXnVxvQDVuNYciqd4s2r+pkNUuFelkqog8CPw
R0I8vXsb9J1wZ/LifAubTvOItqCnNT5D7+Pr/yHAlh2i2hnQD/gyQtxInbz0czV+58RGiRNsP53d
b7g3iU92ecr6lEp97VOJjIEDla5wQqB2aFMA5cashLT5G5cz4pb0XOSVccHarnUAHwjnUKBMn8/U
zUa1SDrsux2yA6zj3nU2qS+RBONjM5ljswtQNOnOsf5aDLUh9vlpCk/nJS4bJ7Iq/Sp/L73rFsBU
fu/SzAxqY1envQXRr3mkSOWkUxhg7mJHxbDna/EGR2XG9L+i/qWzUA9H7ETVlDdJN5kdYhyPrMJK
bszBvi5hXuZhMtWHnN3F18EOJoGJAH/HSkA7nGXJHXWjh/AoEezDwPRl59xm2sV/45p5/WxulMgQ
uL2DKOwhnlyuX37gtyrSMO66UYmLMeGEs1BG7d2OBace+zqkiUPK0Pc7GbYQgm+poZiPo1OpCcMr
I1Wxbi+CmMXSiZ1JrwDID7NoKB0pCUjuSkXqE3iz1i5G/ghKlqbdQsmzOGwyrdtDSVijdiVisFv5
2aIIklhqZHAzrLp1d/OLZTEOV2gVYk/IJn3zFcB0AeGRhxXAPuDcQtFOoFV52EjQcmTh6SgX1rAc
O6s5euiFGQlaeV1h+eiTBwTCyjnNcYMEVyTkXt6i/Vi0bsdxbSz4BcDk9b/xpTmTVPmARVF5NpIZ
ZAfuwbkKMIxWmUs5C9YQPBBFd55sfh3xwtbESB4C2Y4i0lvjF94i03m1oztOR/EMX5r3Xh+/mf9n
zi9xGMSeWUtb2/7EwvQuWxUkgDiyHRdyujFN1R4ZjdwOwkd0mniGBxuHoMKIm6iyRPIxZO3M3WJk
kuRRqgL2eXJ92d9mFT4fIymRML0h/0hbDCcPahpjiQ214oY7a0jIT8K90h5Xrsa3gCw/+CyR1ZwB
3oJucNWtq3Qeq6t7meR4OuUa5HLNIXBjUicYEz9xq94NRWQA48iBuBpZSWzZtx+67aiDdaseaBC8
99UMHknCs5fgNxYxDQz2w7X1f/S4+3MsSbaP9axmVNJtyH5dcMPrGcgZTMW1+/UJi/VRTBPNaB1w
47M29aMd2v3qK9N/WXmYfiGZbGp/Nxo3vLNqgroBQixTRmPH9jyf+iBoPgKS3gOPEgrakLSh1fwr
fMcISet31yV6O0vPZbJ/saxOJ9ZzXqtT3WT8+lqsMR0jGfGxv1R+vsSjqofaN3SrEcjKtqTBLAOH
5u9sfXmvYyHBmaYap+vaaUd/hset1LATaptvMQxS6OArjPjrFAxafDBavOskOlMfwDDI8DeGQDkB
6buD/nt9pjxbhpSbFhjym8epId/y0pQX+z2tJVl3gKx4be6Xl/VERZbAG2D1WKWvhSdnsgLTF+yZ
QQsO5NM0Tcu9MSo2xTaEY4r6NXqO+owZXXqO0o7v2Z/OeyM05tFTIL9xv8vPie+9sDbDCKgGc/v+
i4sBYq8Q6RlrO0W86fwWVBCl/HG66YPkvOKLNdynTrMGeQRWu5aeFvxcKhIEgIubW1x2TL1EOWBZ
Oh0k2HQAHNf7NRBGZM0jUQG+XzbGaY++6188PSlKvdQKHD6buFa/3j/q+yKJJMKCGtDFHcJK+3y3
5UEHoZub8oEZ2BwaU7vccZOXe/F8uW3P9F/vYipbxc4JLyzYyuG1D6F15aR1ODIot9JxMKIJEsNq
TZbNBhH713rRadrzJhMEonsfy1Ppzw6iLDRRd8BjvL57QMiqPVUSu1PyfnB1/puTdAXfQw1XSjf5
+qYeh1r69quhkb+yLPDbGfSqY3S5S3BAT6IljlSDGttoHGp+88YpA/xIJenOXAhT+kDnn77SGB2G
M4RYDz2XjtxoGMxZcTLBjx3mz622iRpjSeHTYkRpP0oEIv0d0LNGWx2uFjZR9Ts9XstCTG9O2Y1V
YLSUfEvnuI/svmhrR7stQmeZwxVUcOTH7sEZxpQ7A/6spROA5LH2nf03r12Q6qJKa9AkETrEm0Zq
L+lX5BY4ws4pnk05lbjpfwC3LhnCF2BTWnXnUEZrgtVAMCybAUTJml0P5tAbSeA5wIsZutaix0Yn
Nzzpi1dqkrqelMH+4OnEK4FuMWGuhc2wdtx/c5875c/3kM7p1jN9YhBkyV0qX00LGrszpCN4w49I
3IBvOKg8UjQAav98coR8DXwywEGfSKhyGdxVnD7g5UGyhXHdk+mEmYM4N8Lm1/sM38vKAmZUZ6ef
RH0/BKx4pZ2Gnm/cfutGDlFaabKwfqr0buGCtetdAXmwvmqZy9GGxMNwR4v55Xmo4uZxhcUtAUQu
awBtiO3vDsQH8pxkDQxZhjuBvodI++p1cjSAOZnR4iRsXW7QViJjrqC+Vncv+70/dWV0DLJpLIy5
Dl887LgAEPWjM7BsNLFOHqoqofkNb8xvunUD9W9goHgc2KYpk32aDvWdKrpM5Ek727sQONDUEXpx
B/dSCRXD33dhf24KLNbM48Gt6n9DrZ0vWummAZ4T0H3q53SbhZoI3xgBakZXbj0iwKG6/hbH/3ZN
Vw8SXVdE8fViVI1t2wCUpxYqnK7/SOvT467w7b/Of4DJUQ3IV1cc2mGdKt73deGN6n5hIm9HaUmQ
0SDeKgVVYUO2c9A8cI5COIH2uu8kzZkSHw14/2kEyGQcH4ckhndTmcDqtj4qOC6LYGUSXqDjOzSG
k+JMpNuXz2kGfcf4wfZAHTseCYEDvZVok6b+LFjrR/RHaIIZZDlIR7T4pnZAno3g4nnAsDxjE1et
/9H3IaXeNe8J5xyJah8IxKcrYyf/zl7jmeIAziBHE/sV/NBqL5wL23F7Et5+BgJonpDLjPbLMcjQ
4tMnHHxlT+2SeiJsHreSFbkldDxKqVhPQHf98uv4NWZBknXfqxfJRoBmYdYmae7i8zCVgwTptfpP
UCHCEAkzujfradh/zUuRPQJNJYWjv+14LzrtoG7C3uCf198uYPziMe4Av073TvUifn3BaRsDqg3h
U07bJaHxYGShNjE7sqruvtn/agYlhG+vE6LsD+ZSNrPG9xSBqCOZaPH/LXFhdlwyv7OVpMV/KBNQ
jg5kQq0qhLz49P55OhauWcKdkrYAZXtjwGtCCDFkp7HWaVYg30EV7brh6VffPn7MtANXTcLH1nVw
E9O2IKNllVuaZe9CCq3ih4f0MZCWHVJam8oR5aTWjFSVb/ArMY38MyVvIlyY301FWViu6nbvXB1x
wBqs0ifoFGeQpOnBFaeSydhZtsynn9ch4VQ6QLAPQvs3ddzX56RULIlzPxubd+uR9YpOmaAs9A9j
xt2lFzvlSVnQikSxEmIMuQc0kxSQwJW2feVXg5uXjF3Mg8eas7UduPi3PEeyDdftPnygkQvoDEx+
nb9OqblTKukpxamleBQ6jEbhE9LqRBc96x8f6KbKqR0olbGCzupinAoZDzz0AWLo3Pnl6YZ+tD35
0J4KtBV9ZGs/lFhhuAIA+G3Aw0bjc3bnXaqENKnNfEYOl33pQ58WK65exZE/UBuN8ysjlbQkcCdL
Sh03PA/KGpn/vRn3/D7AxeFA3t8qxzgt382v6UtJZnzK7J4a47RdF4VVP2xU9BPqb7lPcYgM0rDQ
QFz2OqvxQVlhoMtusgWMAtdfh1xIcGh3Xq/bbDiRMwRwGw36o7KWusP1EupBF8HF4lmqvuG8VwGB
aEYYOu7dFS0dIm4Hg8qHiKoug04+Vu2CcJuar1LZW5bYYqp7W6/i8RYV0cdq1j45gfRK5BsUJQi3
74svo52/Ch9KV0+fhULSzq5iQgs3fsSpFRPziEuj0oG9q/4Bc+JTtKPVnHG5Ceytln/9xG7n61qb
XfdBc9/fblXkGXKOI0UX918wHnysahabYjurw844Ua6BEtqfNQj6ndjhhYoZtnMWXdg+fhMc66Ed
dIvEh0tf9VJTpya5C2369UzY2YoEpI338g4FhqJ2sz9u4HlLaQssNyMJXBbth1GglOyThO6V4hxg
HJsPjOmliL13McaOKvA5Rkmh31UAXXk94+OGYv+H0EGMksQeCH1LxnukraMWRhCTrTrWM0MkqNRQ
EaVL1GXMJOZTrETZv1LiaKRPN8MO9JKlRq3QeiHTRRvxpkzO2aXugo7oSRi1wAUIXvnntWAlaE4L
t/sgQ50KROw7ioOKGz9+cWkoaCak+8vU72sokjH2nSSfw7ELRGrc0WImcuO1+3jg/uBDfqJVufHP
mqM9Nb3mdfRDZLLe7a2pkXkTyt5U2QFSnQ45Xytzr9pupvdthcmyCIPd05LD+wuqPrnsOTwRpPoo
0vJNXv1hTuI8Bs5NtR77wDGzomNvBx5ZVJtOnvOCU2uMLWveS/FvvMQV/LXfj71fiFTuAe0k+FiS
WJN0AjiF9UshPTz1s6qukLFaUfG3GkqH2oYkVMkH8fgICOl9FmBdPzyLln84DbW1i9f5P+ta15qL
IOJDM5ySVmf1EyaYeM5igCLASW6AiwjPD88+Qz7CTltE9gzR8aTNJcohRIAvalemdnOeNqN5fZE9
Q4zhSq424YPfyKjz9StNt6ZEjgefm5wd1WtRCYtlQ8uzLt0kBGde+tub6a+bebXVMnEDYmtfYUss
RJ/kEAzo8rPgjypSkG6URYoAh6OWmqYN3h7qAR4AuRCTSQIgz9ee5/B9O3pGK8lJuEnrtENDEUo7
HDB3MwgJkM1AbgTz/J5Z5F6rBNvbsJOmGWcTx0NVTNEujQtdGuwkCLfMbLkSqm/XnukTZ60razn8
d4tTxdQE3iRLzOoKLAjHHRLL3aaLkw2r1jCNJ41QKVkh3m4E7D0IdlL7q5pH87X3zHRKRCBVr4hB
BreUSt74/LGU/llOgTn/UTJxFnfHw6s08dXSKI5oR0twgkdYpt3c4VAJ3vshm8Fpc6nxYAHnCFyg
Au4q7gUgvqH6W0xYvOYsA4DQLdlIidf+tZmcqUdOkEupztV0IexH0Mhhs13YwS8rf/V83hz3qDBI
y5sS2s8JF08q0NHxsexZ0TBZ4JD82eQc5DvGl73TlV5VCg17qxenwMJMk5mjmqAXFhikjQCMaG4c
BMHTGJTkfL34/+/iPeZDMBklFTANC2wNRkqudwqVfQwP0moP/rj6t6MkvgmiBVFcP2gU1J8TIumU
UZBk7dZM/ZkwwqDYvpC1PQez71W8Yv+O/LnZTLe+1G0+VFjP47IW7E8VaphBDIQI10kebAiZK6Y2
uGXPLMGiHLhu6hbKk2SUD3moSCSYhXKRj8F8vkmcOv5vkDog9MEtCBF6pbD4+y2t2H5nxrOtA8z2
5avDBV1mtz6qYvhxaiGBkLuUi+Lc1UhrMhejm0754vdgajkOJqZCGy0qemFWNpmap9YBeCrTPH/r
2n0PEs1pIVgNzzFc0Af4Zw3oqJXH4n3J+5xohF5k2WkJ2GsP4tIQzFxviELuMLC80ixiVD9NhHb2
8FrV1S0368pbM/KiHpv7ysM1cof1S3BsPQdAYR21TN01jPtrgh1KpspzKKkx4tBSMju6q4rNzocj
Vh4YqwJslV+ctytCI6GqP2h9+j9k5XM/No3jv1AX/DkEnDCXF4g5J4jrct76aINdXnAgf7GR5sGG
vr073cPvvivCXWxuZaX1WZVI2OBzOP98oQUZVnkV5saYy94nUSyBt0HuQehwCouMz6Qu457C7wjh
jmRzYhw1+5qul2HHXcc1tjmo+wVcEA1k7wYL/4YTA6SXQrCe+EMkqV3dd6ACpj5uhjwdOopTy4Dw
M8p+S7DL8BFUrYxRpUpcgzJYufnCEIv3LAt4dO1TjY4QLZ3+rNsDx52GS0FS2WyXgvhfQtBZUCFa
qs7MlH1bIrzsZS3wO3uzrVeK2Sj59QE2clf5ADuLF0kfUipZ3n5A+WMyChxL7/5DI9BQqzFM3O+E
xNdOgqJv6NKDtEhHLvrAlrs3nK+8ElzeAc8Dpd73MVuHTEcto1zaUOrhw2ZtLlp7bHkxD/oOfjuK
PhyYJAFpg5RodXcHjDfL/V0T10K33lBaS4pByqnpmVUxZC7fY8BPuS/FlVsCguqzbAD5RXu+P+AV
ejnJ3k6cnBElCJ6EertVApg3kViidugijcfYbFuVA6DRLasXEXMKopp1hhXg943IQLJnL3D5e+Z/
s1yFZszlLBD0EhIMbWAHa5cRru1ZEI22tHddIWToPHK5e9dGCXViZ3pXW8zXjDmJRjT7Ep5/eZVE
WnpD8BmINzXJ8n8a3V6oZ2KzBuzbzm8YtDB2Cu88WoDR84ww9q20xiCeV+rbIeydtLk3VNwR2jTj
UAZtp+ABbunpDLaKikSVeKNi4MVox++3rTzHM76HfyxJP3RjrJVKujh8BKTQanHBO6L7A4tG9nSk
ap3YUjOnn4lzEktnjDSR9jIkjvL7XyVJNyJGUS+8+1eKC4dF8BNijHW9lffgyCPyvHtLjca7xqZu
cGzXSA8yZkZa+s20l+1kNvzBYPuZEBJTy63vb0bNAg392CfIgCluCRUghY4T5proY/wB9BgVU1xs
l+Qwp0nhsB5lUp9uqrfHG0ONuFOevQT2fTtCobvcadKaC/Gd0/5QTpq6O6TwgymDf73xE7Qkug2I
XPZ34OrMxM0PKlLWGDodV2G9snQepGCR0VpgbVtrryFCdSUNXRn8GPCOA3lnCLRwMp7TwADe4pDt
45SxEf8Vad3OhYPutrGbOIZfKxvhjyuJJ8sYHYukdwRkqAXQQFApH2I5frE9MwSJkcTzPwaQML8c
X/hPji8fyFmmzLSsBCGgLSVCbJc3cL4VyhOtNuzeb2DcgROqHfLwvyDVDBFD26QHz785NcyB/G61
LnOVH5PX1/vX3FuChN8k0dzw//lO8sgDyKr1BCYWCPP/AoUa2moCO+H72K0TZUNAYBKCVHkZTddw
E2OVOge99d8TMzmiL6SuASgyDeJVx6aKnm3IH2kNjJ2eqRqRS3j0/d+PUr0fnO/Wq0DzCAyP7c/V
gJH6AwMH69+yMXKijQ9w3sC5dwLrZBrdFvAR29uouA9pyZE/k8TRIgErIRAOIufRCu5XC35Sj9nX
gJBy8/WjLxRVvQd7QbpNbBu3WAcKkSNqQItZIVDLm9rfz2ACYx+u2SDVbroRpLDiR2jxe8k+ZF8Y
gfYn9VjjCd2eXyEotDX+MTYuXJQq8oXlhTBu5ri8II8dNp5lANJ6JGfGL8DnLd+S7Ws98U1diLLE
u7CP/C0LJo7uQgJnvrOGe0syG1tWnggZ37z73ImIBTQYlPd+PJGrsRyWUklE9ChtZQrJZZvt1c5W
ZrDScEVkh4dRPNPy1JP3RzNXXXgfdKG3ThOoaT2wctNXDUKRNx5FE6cJoO7sHmaYMo3gCD3n5Zzt
Zx6wiN5q083DZWNqvIBH2diOFu76iZT+PXwUf/ILM+/VkC2iwOmUQdGB3A7lAvrqZ937RpDHEYvl
Ch8t0TuE2B9eHxAYF+Z2vDUZ1NbdZs8NtEPEfPfHxulZQT1mnV/zeX7Qw1Ewvu1W3vi2m3OSTtjB
kFVQdBQoLKIOAfWKzixAWpX/lyBkN37srzsY7YTdKqHKxGbjQaunGUX9D18z2m4w29+0OBOsI6uM
RukmSG/lkwTUubC2SNI7GroGtlr9TvCOvPbb3EK6hWBi/THLXTri93Jhr4i90Yvuu7xsPZ2tpZ7X
eWV2XXCLgZHk2FRBSpOXMwEaLmO2c9iRp25jsEwdhpYYG/mC2RP9m8bW6NKmy+UxDwf4j3FKX9XP
pSJEAe0bhVRGiS3yo0IjjGJ68NMrmjHotFIVnWWoadkMgnFjRlehT0fmdfj2Q6IWP6zM2KbHU7Wz
dP3CJDyEKzxMZ9frRt6NR92jGa4tNmvw+c/Nr/G1WPxlytZNbCxC5h2vFoE8w8G1/fBMQJHbSV35
qjwXQRP6S1bv6kDqrpZWxe44b4cQkbUftGvJuBT8y+GVZ4gH0y/ixVKYw47sOXe+VXRJmbX919WA
8FeUC2e2+dbR7Dq3CICPL+hX9aD+NoreL92FgyBVtHc5kT0IVdb9fBNpkOJihwFMDhOzXUPkY34O
YUH9cV23DN/DwMGYR0iK8gL8G09MZpb9VlzPRzb426RSwnZUdRMbzpjB5t/a3Gq5bsOQKpmRkOh7
cnaz29c5AaLr7AkYLtclp7Zmri7HKvfC6H/id2DVwDho8B8ZaTmf1ijeuPnnmZ5uBjmBY2WgEWb4
HrYJtzbsA7NpRJ+x47LYgonHy9B+dHyHvmWdPE9C11GYeQZ1sSQYjXhpjbdAh5ea4tfcEOIO3Q8U
kLbFHxf8e0UfkPBYPFbGYFjLCGV/NRxUVKlHOtxBNQwtrjFGbAQo9O80xfv/CpyquPEqsQi7U0th
8qj8ObUZvPzDJHtoJ3kqVpYjYCK6ugnJR3o0yb+cYvDwGC5TNkOrxxoIDDDbnwMSJCz8IkRK3D09
ED/uu4pZFlm24qeOj4pjbb5pVV1vTh9IcKO1iRCnlFRC+dbFH8Fsr+U8S/cmqPHEC49diNLt0L34
osisujgVRJVr10gzeEsmmtBMsn8Kz9AColIQM/7r+DYRzkfzpThT3C4Y2XlqFAaNmftAq+1ap/gx
1h/wus3TfginHNcmdKylHH/6zcZEvI71rzQr5t0RKzpjHWmwprjCv00sTs9iaQBxdZ4BBq90laRd
Rbot1uSwvNYG1WDYg5k7acOXjTT0Mg9K3kFmq+0DpkI0IkfeR7r0CK4W9agXzEGGIeDszWQvJfYz
Z3aXEAYl3XEw/hOqh3hs9wMiFmvQOKVSO0fjHNWnHWKuraiAD7MMV7hiTuUONCzBizHcHx4Lp3KX
z5vd6zoTwzgfYS8hD8x+LQI/MT8NS1RrFVjFZDj0cXEC/+WP4XbsKztHjmiVxnwpxWWUzq5tfjr3
0DA4lO62JNG4AvXOeB3iq3CUrDiYRVzp83gb44f+wQTpK3JlgVb9z22vPXyYelAs/r/v/udTk6do
kPm+bkn9naifLhyw2+46oKPT0gHhttpUUy/fedwg+RF3ulWoM3CEtWXtBKZXn4Cy4VO0jR01jXZt
Pnw30BWjpBomsftSKn0Wh8JariLGdFsXaIz9+A+e5PBHRHoJssS1JBjBiiKLjl1MfJIsqUWJEAZ8
V0lua0lzQpIU0YBKktNBvZTX4xk1W1Z5cBWDJFyCI7rJ/rBTyzaVQizu7y4mLNSj2tWYqHuZbiXI
K+ZhTunG4DWVKKOtvi65fd2qFhWAuF8dYJGQGcnZkEvSU9xx3AahTTeXxAjxJnRM+C5o5dP8Hq+x
Y5meT5hs23v1kLHJaWbth1F2zF1T11H2RZwvxukoRNZMA7DVTl2PM8ilpoYE+N0IyNvQSgeD1U5H
g9JXDO4QWXbzYrp++vgi+frhFRpfDDgdLqSKy5b4EGFGKGe3MDZXwBMfZoY18GZTA5iIXEH000er
Y+1kpicwEbdRtoxQHMf8SHNNy5NqAvDFpgkG006tgViAD2OdxNcKomQizfkv9l+oa3uUTqDRWTfc
uGAy9m7TEQWmtGb58EoiWlBg6VFVVCC/gDxVSqa1cx0L0AygwFbDUKwBLd5CeDlzMNe73u/gItYq
g1UAci90eKSoy6MhB9pIdOyvd7uncYXLZ9B5m4uAqNKjw301ysKv8aWM4KjPODEeawyrcbSTqNsw
+cLkoqQ2T3p21mkp/5zz1gQlJQhu9nfz79HGvxSZTn9Y2Vi729xzGKZ4vw/YfSkvHLLwj+AULIIY
irw+pjvYKpePBLurJI6X+3XETjmbK6eh3uGbE75YjZL2wj6Wkf3qTci6uTYy7BM/W+Te7rdmBAHn
rU1+hvyAhLmZhFiQSh4iROb0AoBKpGjrTpC4v1JdhHzwp2bo7Za+tJxDNxkKhmXKMLL8wpOBfwf0
kC1S/a9omwc7GvC4yu3dr/q7qMOOMXQ9pbOanTnp2U9ugObVYDMmaTu0CTTMdXCmLvg6P3ylt55N
8nstn87D1VuqTBj5WWnjDSiHg17PYAc/A8cRv17ULqFRcIzWOlNPCai5AY6MDJK2b3RT7aLqfmst
hKqi76W/TmPTsqiRxeEv6sJuM+D0KtR7SlUPEd6LoQ9ue+93AvLe5AIw7//4DOEFAM3grQw9g31T
TLQl+XCPEWiH1Oeupfhe/ZQ3yT/UWrWsse5JgdrCDOBe/pEQl9KARU8PgxHyjf6KFomM604q7QR6
62WmSOL2XbUD/PzY7OBEbyCtZN5GiG4fuvGgJelqiKXSBj9nvpbX+A7B506AZ6EggoPq1sLc4D1Q
zKpz/S8RlUVTZ8fIhHTcsZXL9ioTgtrBb9vyzgEPlQjQvtybKDrvewAZvIVSGq8YG71ggCUwRbL9
Z46cdHm9t8WnpzCmhMlPS31mltdQrGZuatBXQNs6KG++B8mn755FqIOaQ7xQnUNNJ2TXhheFyfgX
mDdXfLORPoNU8amzS1qaxawl+dROUQNdLSbDhW2EWZ2cFkdsvIHz9IsRDBYGZCyGjszoCN40M/wB
LG6eWPdHZJlKh5PQIjpS1FaMk+zL4LqzCglNCdBtDo+swJQsP4ycKvrY8LRA2v1BcOr2FgOrJdzh
xdMczVmcC3SIOZRz8uyAxXuv768MYM3oIMjM4LOUZWHnUn6nYCvP2EYfxtS+oW/7WUOVRFxEj17z
/nItHMMvgvuljXC9RdrBWHzaPMECk92ZYzWJjv42NVuNFOo5Sb7zX5jIvY0el67wHXdlM6Qolxog
UumpgSjnIangCe+4LPmtQf1PIOURk6/oVQRuxjlLXrQgS5ob6o2yhTjEwZUBUljt7KeshwaKWqyI
yRVyanEr5TAYqMjZ6Xs4iFd9eIYoMfRmRUzrlMS6kj6KAKv/ibaTDvgA8mC832+YvO84+9UKKaDQ
R4FaugPz9b2DMOo7/smFIPSJM/p3IQzJpEX0MkRwTR+Xccc2UeB6CZVZOA5eX4PlAuOxlq4mFK+H
Per9lx1NpbTqjmTxDqEev1EkdIhch1gtsGkMeNmHvl+EqXESh3HJY2xA0FpYpc88TEmOI+bIL0uN
UuBlT38PGB6sAV8NiTDiQWbmxThxGeekjB27rqMUgOVER6WxxGVts/FpKOM4OmJpLHwUURL5fykf
7SwCoLUyp3Blt7cz8nOGSKiSrykrXrYWWW72T2ZZUBfpkazalhd0Uxc0xAdp4jBaEmNcGtUVene/
UP0qVch4apYMzIt6iyw+G8NrbZtYv5jXhs/Izmy6qaNGW11wf+VHyymmkoslC/RZ2/2/DYrWPklg
3hHFyP9DnG2J0OBNwWl+Kkghb/+gBZnSv5zCG7NrSKYPmvG10lyPY9JAzANOsIhEYCszcLUH0COP
EUYoPPe9myBPxiDmwcyRpbSNl3V5M9Z90r6oT9VQB6nTsrMLbtNouhiQdusK234yNQue7kauAbhw
rftCQ59MB+qwdPugKkouZgVh4Ut8bykV3QtAxT+TI5E53ylxs8Fbk2z90zXQJMB1TSEBiFzj7kZN
rzxUEN/4HBtmnmwEIkxtzSbXKPMQjNXLytXV4jQog11nEVF34jHw1NMjuahvbN+pdR0/jmlbgPRs
9Q1R69TYNh0h8o3vVb+P+CsHxfOI7XZXazTakP9Mvl4f89jCtrQDv+8x0reCPOyMRxmnTt9EbMTj
IVTM/zoRMhGU20t3wC8oClpHLLuffB6sZx/P8Zp6dEbUtCc6H04iReTd2g7j8XJAJMCC0kThyShC
8X8AYl5y0QzuCn6cvvj6Q/hNcu72UxmJ6j/nCMfqr7WhUZZwJCAXwLlaYLBVXArBE48+2bPb3rNd
ATjh1BYjl2+4GFBJFtmGY7AwgKW8WfFO3P9DUiRjZa5KROs117HWlfaCA38Bq3HfXOGJwSCSixdf
FCSHdn5GmtXAh3s7s2Y22MuV+unxaYRI30STqs0tFtNRb25DSknjvZZYRHMRlZZuurFBnDFHLfq8
Ve1zM4pjhP+MPbzS7XZK+FRWgldxJoHvj+mv1IML2t+plnGNp5NLWx2ht7ieWDP6tCcjkQ0JqRIt
BXPT1XehnxYGtsUSQJOZWreJZIUNQpk75hKww/meZ15UYwcYo5xk2wLuRLtYysqxHiXBmOlWgnLm
OFFkA/6IwLCeCfD+zM9hjEhcTAw+d0wvIt2PvR8tXET68w+3qAdK1Ntc2rZy13WkwBBYfKEq0l+s
B9Cf1btqc8gbSwwesB1/DBJVGXUgxliqS4JCVANMxv/7mboqp/ROyx50C+J6vG9OiY3j/DHbn5od
uNMUpD4B1h9mwUNzqA3sg3DljNKHPaSNCbpG+Q1gmQ3FChOt8R94+K+TKd/bHXjiJXw82gLvQDjx
+XpBv+T9wepwFAT//VEbGsXc9MJpl6wLrB9TrkLDlgtk7f1CB8QbbQnzEsDpHky1PlQ84hHn7I8Y
m7pRymgb1LFU0xx2JnSH7mth27v7qU4cPiBix6rJF63I2vH2ZI/wrbwwewiJnktHpDlA6lfnDj6I
z3qLU7eBM19p026TUZWNbyXeXdzE8/bA0MrWjCp9aedvOq7xgFsLsFB7/KJUzAH/bshb6LAHkzxN
pOYmtle2tBtFVJeT6OzF2s0niPaXR0iZxUOdbNtUUlBk5xXnm9wW5nYLuX3gJTaxdJlus99ROtAx
iI6iG8rSqytxGpVaZkQZgXqiKiN74RUItx0/7Hlet9iJmrVE1+pDvF2V2wK5k7G5dPU8qTW7v6xS
fIIci60bDS77aovgKOoghvecIqzTsd1cz57C6UokAtP1rI/9JL20p1XHj8cUz50Ulbpen1XxUuc1
f55WLbb8WiB0Kwld1ugBqtXYWRgS0sy4455TJAVSSs3P88nq5ocWIL4osC3CuPSdVU773jZSMOe4
SivgCM1zWiIdeZevSVJMIHBaQdgL3hKWYrMgMF0zRehAKqXPJ1jtGDUsefUB+X6OGxBF9+n9DX1H
HA1FJNLu3D8SrrWOSrXiS7YxI629KlWIqe7brIpn4o1XcXCX/Tmro/nKjRs1R7Nyc62qLALN8kLO
RoH8iwoI6oemJiBV8tYSFkYaVd/1PZ7jchCx/VHj0W0TYuOV7fCk0EDonopKP8Ixttg4HfkBe2FW
Si1F4HrEmWevpL99bXqwqH7jBWUFdwckOTI4Azri5/ftss/09jzn4k2oUB+hpL8Iz1nb20PiPsYF
AVZaUWWuQAgGF378WMv6hrUYftY7DajZcnD+bKPXubr3tL/BFYeFe5yems0GaSo7vp6BlOOl2PYL
QczCs0Wy/Sn+TtDMGL2Qrkktn7duhkhoh0QIrz1c8K3FcgbC2ICfFV5qHP/x3oB6oR+11qNlqb9N
FrhDyOaeKtxpbIsSvekvs0budPD6TbOo5jrLzvavfuVfFqM9PfOn9jNO1yG94t6seX+S5lY3np6A
8jNA/VHB9JEVwdiPSCaj6E2kxD2hPW6SnLzNvpCKoqobuOvddT81212JMhoVn607V8ZDGMK/0Kn1
2wbX0WUHo3wdSdoTAqF4Df8i43VnqV6olyl5X4HaVutfQEc1lQ3WoEIxPB/LNkRI5Ry1ZiCWzmcT
WOBBgYNeavMw1yOQ126IbfQN/1z1xHrI0t5WgvlrFsmOWDKsDty5iPhYHDiMkJ58TwfA9f390hTY
5xo1FhOWOW0oczhp7aCQ87U/1VT4DaGJ7Z6a8D0wj5FuHrBPw+Wbz8YtIzinOAutHCsKENWv9HYj
M0zKmkw2++63d76HkHmxWHDH0GMjK+vjjXw2XqBes8iqOU3PnnvUxP2oaodT7EiP44IQm99tbAk7
w/hnK8o+8W1HgUVdAaTN77d1xlcL8ja+JNWbWWNOttSjN+n7Fn9g0g0auW/V2/zj00V9rBVFW1V+
H/ONxkGTwdyxFvQY/w6lWwpoYXPx5toXzMKNNINuaNlRsMgfM/wa7f9Dis/TebuXglnHZ1Rb4X8a
vFOsd8vXKQt6I2d7VobP7lVLU+gK0kvfdpXnpfV1AZkZCONvdHLtQsjQ45ijdSe8SeJYkRGdZyvN
KFKyyTCcQVG3kgDqG12QcCMnMUGQCjmt+GS/qrKMJzs+kdDWKEJb/D7UaSljgko2KkPDo+f5I7bQ
FOKBdVjdrPgOuW+z2uzzP1cuaTdWRk+rV6JBKP6S3Y5Af2pfG4V30TiQLpixwJp4+amGMC1uF41z
ZaADILfGqrMCYvmXNfgLaYFZ/KNvJruXbZ/xs4MXvyxveMhdjj3nM0iQhpLSbEnVzKKxw0f4TFdc
QmsBzbyk8WxYFiGT2yrUR1KKTj18C/6LuHxXkoZ0fWuhCZ8ox728z3Sw/HZoKlC1KA+fE3lVSjB0
25wuvxMABua4h8OLC5laqz26l9Q+6yu+cBZNLCWVgdE2wrGGEDq0XXqXSFXnAXyMYahSg4TIqQjo
X0dQkJNc7TERUANvDGfQzEIeejKIGxBWg35YqfbvHLeMCOaBseWgmHIx3I1jZZWCNFKfXU8yD/CG
3Pi/6cJcCuWxO9ZnUgc/PTjQlbm18O0mQ4CCwTM/qQUU4DrLnxc77z6IfjrdgBa6DJiEu1cc1+td
zceBn+Qo2M/YnwKvRPA4GNRd7BpBNmLwKVhnCiKP9OmOL27yMbUSsoADIqF6KgS8WI8gH5Z8rRHT
nc44Q02MgdI6ki6YsIK+KXLvuQhsnfO5dqMSQGRhq71bpaa00fQ2r5M8xNgug/GP9TuLMWJZCD4+
ohSVfCtJaTJRyt/3nvYj1+z7DLeh2b5QVlxWIRUzHfNAEqJgWqAPNnH/CvkSwH0QMLexWFNzmdNf
w7SY+9P17o6PLtSG06LweqP3otc0GlLAQZhd9+1Yu0ha5VkyTSCxeVdBO/oEqwfng0DKw+nOOt2K
IJgk9UiNjKXg0EJUwfRE+KKDdQxnZ3UBXAwHaAstcc9RL9LLYvcOuALBt7uVWq/G1/4Hu+cQWxuB
qrSFB/1WKKCpUgVE5pnUmHRbvVrr+8KvYbzAaz+aDnBOsuzEtxwUWVYU3etrKwQlEyr7IWpS1WcE
grteKE3Wh3y8r8YpkpCFGWeJvFTE8dzoBkQ054/ZUau2rFymoktuU5MpfsNKlfnUB70d1X724zye
9U6lefoWKXyMXIIMwEK6DM5k+YIkreeDs2KBS+I28gqlNttenJ/OcUk+X7MuWt9Rp4h33Kg/wUJ8
7HZHd/Xch4SQsRbcwcxOhZgPuzLtctGWUAJtPaaAiPRRSIZcNn/oHe41xCmkDFZksDcaBFmNKIbp
9WIBhWR9LWI4wWoS4odpuF7BNGo4L7RsfiZBzspI5vMijU2ExHOEAcnG2Uio5IBKaMPzRb7eQXso
xXxJ4pvT7Ur4Z2VBA+F/BNIKqVuqKa9W0mnHpfaWhVODo+H0li/2JWpGJFFiWZNxb8ci+sj3cHiw
KaiyNnKje3FdI/PY5paf/SRSXkGMoLP3d8G+LA9vz/AvmW1kW9qHa+40Im0P4h3y5N8yPu7bkvKm
3uDtJHyvicHz5B3EWRyGYr5OU3UdzWOJ1PMsxrzMOD1U6CUvyONp3Gq5r70S/CU+qTnQRXEdQJK9
0df+JjEmTLYpJtb1d9GGAkyYJr3HUx7cK59t89UHT7bkGfC32/S9YGh0nLAYxMSL69C3/eQDOyMU
y3KmugUCZSi/hejdhRq3V2ZxZryiFaSg9g5+kSIRsuSUFXuy0ljIjeD2/9ZZJneDbgGtpKmNwlPK
9dOKaxJm+5/fltx0fMyt2hR6+ITx1naeq2Bh8J+pzfZNCDEQ0xxdcWRIksrr6f7bSI1AbTr2gzPS
wlzBLKFeCJjDMhlH30DwwZmTXZentSfa1cQTgEQ6XU4Iryf6SMcM63E2kWhKPGKKsjoAsdzMDc2w
ZdroYgSK2GVAesVpU5QixCR04S3xhJ4YUle4y7OJcqPTC0fwlmRahQ2q8SY0hZJBzGKwd5OTfUQm
k9Srp+gNTzHXemL18mUAeIb/8VT8b/mcbKPjfqyoyin5r6VSzKipUZWm8VnkNrW7sUQQF/Fc0Y3/
KD/3ImaHO37VAucqccS/wGuoqtbTq+KT7LXW6esP2eDhIsWLFwsxuSz47/TsDKQ1+NFseMNOglhv
Qck7mo3zkrtk4aMz95OMLvIizWQ+CgBVOfZuULYJ7M8IqhaTcnmUKIK+dPPMbRHo88LVI0bFoljH
NwFgPjo8CteweF+JrkrGaSslX+0phDRz4TcyyMl82s09BkKIPqpOghG45K/B9zQgtMuSYlU0sR4m
bxcDwnCEMXgxaKsqMbBY9bnMkOePejZVRynBEni6K2CCfNNqwvPdRlDZ6H8LgtnATI4TQrIatMZD
lhoFpN568bqBR/NR528uOwRGzegkf+OG+UCg74lTCM0eV0EqQUHskpOyosZYpKfwZCslvwDr+Hc7
WHZFBvpg4Btf0H5jXhF+b+ItdJzeYQgQyE6GfnuJcyNXeelYd7MtbP6t9NL64Vf2XXjVFs7BZ/to
gVQQTq0/mYlL0+E2vGFSCNG3f5/kS6wejcrd6JCdt6Gq0ccgETgdjXWYUoz3BBAqKZSiYfPGJoFU
piCv+46gD8VTTdl91/sZ6Kr2aYX+RiO9kvsSlhB3vPHXnHHGvtAi6pMxzM2oyFL1sUiZi3bYZAmS
0FIIcNomYUoSqyg0mazGB6vxjao85aWNObk4jhwf5Lw73K2ICS1pOu1N+jdI4frgkLc4kz0r2Eo+
GujVcyfycqhue5C7S7sVN0Jp5CBsXIXq7pbzng0svFEpEjr8e47tI2UNZYO0f+Hb+CRPgaE8KioR
pR1ipxLvDQBmDLE/g+C+FEd9Qnbbbp+0VV3TDSs8q6ke4Nd0uy99eeNDEAQhpob7s0InnNAucZhA
rrBLH2bwY2jkPOaeLzPVg5MniMrSN3SJ+jRYaDhrg9V2DhlkkkFV9u8hc2vvQNPfXkPUXQ/7vLRu
XMTSF6q1ggAxCbsI+jVsk6uRG+IC5itErHnpjGj9+XQNdShLoqFoh3IPfP/Ck7DDhLHGPRkBNEMb
Cq7DUTfcfNxkrEurLBUBgM/TE2TzeKKSZUOXQowGAatD63tYYZNcY9oZ+T9knzNc8hCtvJfEqLAG
PWf7E/0PNFJve/N+JwkxyPT09AZeXhCw7rnkWBq34aYYhNpZXkwRO04Wq+xcaaBYpOXV2JvvUNcz
Imh8widwIBq3BBZ0SWb3whqvr+01TqZDQosylP0u+EjBPIBpzlWlSn1fBavZzUCE1OyoIVwTZpDj
qMqD8o/sZs0M2/pEHaoj4lkcNgztyIUo+iIEuB+c+XKKUNuuu0AROIvOCH8VUL2qdc75CbHCx9DT
DsVomQ0Trktwem6U2J8YrSWEmJaQjwrPegHORkXmpkRfi8Bi5nc1E/kGG90JMMyP8ioeyc0yPSaC
M+LWkkprDILIqSNQZBPEHx5DFeOKX6tRvPZMBVGKNRYCX02DreDOWa72yFtlWmran2miXdke+y45
TXuTqNzJVIea/GeIfKD2FXk1bfTsOUA3ChVp9HyIp2dBpelWWdY2lwUvccxJY0llNw3xPqfaFjey
hVpvVcPdww2MuewdQcoprQoB/LEp5pVblGDD1x7B5QEy9AABI+dVsZycJ0YV687bEwcjWDY7PZ3l
G4CVyLOFssSRy7ri76nCI8BPpCBH2AfmgT/K6h/1AMmyaQOdOpyew2TOGq3TSNYVlQLQVLjKoF+F
S8q9/a9QMaqdX+e1CF7MKwZY+d36GZqbyV6AmnqRj/eyy4sf1FdriGMFgRuN4eJ3SqMy4PKGEfzw
7/04Im6LzkAX/n6+9CWC4YdFf+OGKOYVdmBQ5vrhRM8QzWFNN+eYoX1Up9jnPGSuDfhrGdhIq5Xn
PYJq0maXtoaYuecwiiEJhY4JPpnQbXP4ACMU24bgBkHaTTdQBNoRnw4oUlnyJOn60V9fe7blGyUF
Q7Y8SV8Qs3QrwSSfRzlAoqP1IsAVvH22Tx6R/TlzDpxqHlmJC4OGOiRZyd9Xkyd4WtUl1ILnaNND
Nsu5JZDgplGJYlf6Ubf+eiJX34lYOJvEGFApItjLn7ViPyXTPcC8HYhl5Kyf/tOahjKGZkg4pMQi
wKElG+2QAN3Y3KurJ+/GOdLYP1gPcISQj2mw6LUddsOkEgEpX2oVZ2281WKcSiNRGxslZLdJxlRb
8LOOGt/3YTdA51HaZJfuLxARgvBqwdS4X5HXSs0EXagsKnPUnunqVk55oTqzsRlyKjzM2mIBUUUF
1eVCLqRUxQFwfiYFf3ElrZLPId6k55IaNGoOZ6GbmKAAnGtUsHRhR4689SF/uwAqTgRnJ+iN6cGJ
o92ZHj1YhMJ8KNhdPv6JRCkYa9aa9lRP/tlAwcAqYZsBu1Lb4v4xIlWceetiahhnONop7Qv5pqdM
Intuz7GWvjt7lAIjS7/soqpBizz1u131IJgoi8pcJxmvEI402oouhZZDZg6dRt+xWrLh2g5CGseq
uLvM85HoCWjzCyfbLs53ZB6a1it62HlcU457qdHgswm2gwArtZcsDYZPw2wDC+WYq42ocIC1672p
77vb+TU3TBNICaEFOa+hmG4TI6hRJThN0na8K+bV0cUDny3PQlGyk1/rATlspcHx50vn0zaiQs1n
jnssDrUgrB8AApO1TZTJHD9Ew9wu4qhEg2fVxmj0GRQujQFArjdxwQM4cjWPwza926X73x23dEj9
5eUgjGvAjz0oyAvgsoY9Dr3rrm3YYMWn8HRDCdN6+0mwL09Qpp0ID4taNOssFGmV9PuxlzL5M/xr
qRO++ivwjYin6yi3tcmpPKbz1YqGVyOJaxwYO7c5iBtdagt+QOREavshDfffZWKZXINm4pqFpsVm
wbf2QHcVZC+hOsTzkWwjX2g37M/3BBtZToLxw0Lmyrcmrmg4/GenfBUWAOjeD0vk3Vc3JSH5BEf4
H0r/Xr3Zu/gatuZ1ZL7a7S1l5qRvDZUq8JuKJ0xw2PQbBBkERJWhgZ6jvHkYTQWf50f9/EbHXnvk
81YHLtcY41BciEEMBZTCm7eHUFfIYKZkPuZZim+FpTYPI+79Vwvr5v6/7komoVCLgnrlCTzaWQEZ
dRm7klucfL0x4o6oA3SjJtbqZFh6KT5RZgooMRTjt0OZw3EFCdthWJoufJM1xSqBhnIpH2yRO/U6
qeAqVAJqokHU26dF7ismUxrsijnJCaJvuCOwrt604dO8ZL/YjfuHuVgJrbC8AHUWYvnEQEhOxq8d
2txzGC/2VFmHqcrHMuRhVSGGW8+o4xur6Y5ia5Y8t3piEyigpXoR8MUVhXJtjAdeT/9LN1TVCnZe
ofna7wnJqp6LX+mXqRreNV8LGziq+HP3FaejVEouX6dGrM35/6+dJYILwhKUT6n9FDU5CsH+bFDS
zWrSuVWLQFCM90GDbycEyGuuxWd8GpUG9ixRoObDwZ0bS+CEI5OvfRwcVB6re7lb6NcOQpFvyAmh
z5U9GrziH1B+rn2J4SsasI0Z1ZwHBBSa7GamPDaPO5M6G0u/Bn6Q51v76t2+C3qcD6/DuXpGRM07
v9JEKmG8+Co1yQQOiqQHDrbAYkQAPznhBAqRd+GZTtH7Zz2t+QbGQDXcel4Gi8N+UJGGAJ2ZAmsa
P9Gs7X7w9nBcYzbGdvZyTEBjB0ayV3XJOy0fhDdn7xexaGuZ9KC/R4m5HxD231uAEgvuBunq2zL6
C+X2+PrRv1P765OxW/toqdgGPFCB+sMbiVHnhfsuMat7SI0PdZBevnZ6zCEkzGuUK0fo1S3kS5Fm
oguaPg6OedUPUurTNteuzcf+eynQoG1R+iIDa7Qap7xC9GrwEp/MLXxRKhUZBy/as4b9nfDyqGrW
uS5ogxCKu6kSubK5vDN0Zztbo3IzrWZakTnsEbSjOlh1Hcbi0r52zawwZ03N6ZBaS0QPi4d3/Oaw
QAnXBaa7gSZG7ycD/lL9L7g6gv6axizrwMYz8xZFUCKca0PXk8dFdMqwuDY9hBjBa7h1anzPrPLx
Hcea9ihQ1EcIe1jPFwUwJdLjWiCO5nnSokOfPyZwYrRj6d+zT4ZydwhVaORTwWEhN9G3n7O5zWN+
x3ReQRhaIOm9N2E7MldHJ4p76qSAVPqWX2EK6qFDnQdoqTqFf/9xlBNtpPj8QhgpTN3kJO33tJH1
9588Q3TulPy01jZClkMAPqNYaeosIZ2T1ykAJaIy+j+pm7HFI2sfN/3VvXekTB+N60trNxI7TFtJ
D4sBDIHUYq52+aKLnP3ajtERz+VxsOCB5r4l7zvg9Lmcd7UH6svhJtmJeGoju4sSyoFI7IogDAbP
xFJTQccUVFjmTcG+t2Pi85r28VcnN9/Sv5U8b4jMELAOollVOeNE2kQWybgjZFu2e9ixt46TntwW
hNejzzz0bsYEhoz4x21aP6eE9cI1CT/WEW28f/N1YHrI5HzEalyx6qswUeQoMpvHESwcpAHzoEio
skxkhaZ1mLXJutsqEXOie7BfmrG22OJV9vKBrb1dZh2iYQjOPDcm59P7TOBpGpQ8drvN/cFoMz3f
SuVJOWtyAmr8yj0/KfFgZhJLH6mARBrFNaelVETlPu4OHJbS6yaOHEVKI6cy4LWf4exAr4ohxYJL
CMWUGMY5u2hQirftYgTmOS9dLHi7Pxjx7eTRVo85pkySisZSjXDta7Vm7JgqHpGxXZ1VxuXW+Hx6
K2zKeLbBAJsZOU/I4Q0Iya3P84jqkb4WN2PVLszb8JnHXkux6YD6gb2AnV5s98n3diYwzVrf+yh0
lNQ+05DXFljSLHd2SCB2rO8kfl4WDvi7Q8NxsdMnsoRe8DtGTjJAg8MCJKEnZJj9/HlGa3Bf1+Tx
GUmfEerlY6DXrb4ywMnZwcgZ4K6nAyE2/yB0YeLKCB1Us0wbi8ROCj7wWtR0mkWE6YOTC9rNxGVi
3wZKrII+yh70e54jUZEFxGMUAk+yCobPb7AqlqkZrZBBYMZ/UoiLO7dINeTqMBtM5yG6lmA2+4lR
fAwKomUjHp6GA18mIeZBVlCFNl6HPFxgh/LwMHTF+1GxyywaBbGo6Ecph5fypobnWsrAAb0D+YBD
Gc5kgNzBP1yM/guo2hQRUChUoOYBW4Y9/5pkDcsf+95QABox1vzaTNX9Z8jyXQD6vcqFS2RF+hIl
M7fr6GLtEQ2YtWFyPn61KiIjNtGmnCxGJmP6WzBQDLjLjtysJ9QGxmBfG+Z/50oMtE9ues27eVl1
qdVlCZoDUOWNwIrQwo6ma4eZCb4UORqu3JJBFCXQLOb4lyYRdDw6YklRmtmH2cLithoX0c1ToyA+
11tT8JIzJrOzah9g9MxWIk4IcK3fDCaK9VCKUda63LippZUT/AT3PY6PuXtqCgCRhjYQHa/Vs+e+
ACmDFlDsae8laKh7iLp3/EHXYu3vvkOEZ4oDKRbsJLuQh82RCpG0tn729JIv2c8ZVImi5J5P7HU5
1jmuVujAjGbgryKYTElYEPzTRtpQ8ggS9Ap11/SkVQwVZGzWgsIkoVeyfP6cULDGrqO5MQjf9dNZ
9G8i0uaXL0X4JdxwYgV7nsOJlZ2x2ZyyIlZIpsNHA5lr38XW7m1Yer/0CI3TcVyRliJpan8evPwN
Qk3MGAIvum6U5l+Xl2yz1GXVy3dn3W2v36yrj8DXn3nBpLhpLIJBvb6GxCHC9vogFqTJrxb9SBUw
cZlUC/solnuiWwbc0OdIqA87YD7ro49ADweeMpDs2GjzFKYkKktyqN1/D7ctHkTgkx4P6Y2ryTTa
lA+PUtjmcPOxTbpdmDz0mw5srupBHshoF7KCJ35mEpvcXda5MxkxRx50Ckn1v3riOve6ejUVR+D5
SS3u4GixpgascSyllTWfvfYKrRr8kNeOzDZHTfeeWuMa0fCJ02d5D+T1sTuCzwyfYMOK0eAHBkWR
cOWA7QhjLSUXOxdsZtNCwKFSAsXdrOGm3+zLNihyHk8h1xrPBW00BHXqrO/X3ks/B8eZi1aWWW06
V1LAWn0iyDrZ8UkhyO3kbfI+fXWy+2gLuXi1QbxJPANJOlCNizK3iApxf+IJ9NLccUH9V/tKjAle
JGh4vb6OTVFFwvDXz05GybKTsQuCE5ac0XAMOJa6wkyRe3XYzewTty0awViFDryWz5UkZTr6sIK7
MpQ1rwQCaEIn189M9WihzbKG/4iFApV6bHtCXGvaBeum8QcdM5XP72xroPu5m4jBDGwyXQke4wlv
GgirEnmakQgygfTVmEbOHXRwjBewoFIUnXwRZkPmGstljfvs+96w5mrtOHP57WIg0CKnsqrWpUe4
TkHcSLeZC6HdERVy9x24qknRmYLNqg8ntcqcZCY+Wx6brzzmyukkuWyGmUzkfpZaz+yohwCjs2iw
sCGldW7K9oPJFextF7bGCIeJeCAU24fa0FDu+MH62gM13zVb5Vcp4P95Jtg0ARtThGyCtjcJMbEQ
/JoozoBpJH88e32O+RpOl6M6/qbQGW/YiC0Ux0ctQZnFdQvWH3tn/EjJhWNUhEyG3Sivaye3DG9Y
e0wfMv8ksBZJsQlF7tQMc5PcYiX1NRrKx3ConU38cDCLq4j4TKGnUB6eSVAuFLhC03I9FnS0l8Gx
tWwuOhkDg7VXMizFyBKG5ZCRiKkOr1dHEk9E2KqG5BjJJrpkj1Eatk4xH1svoMRPAH9DqpyN4Qzh
FHmddYLDaB5og5nUUHuXYApRuaVd7x28Ff5sbEdHsORrDpw0LN19UIIBiguWE77zACLYd4l6Bj/3
4j9oqpY09IfBchri/vQj5nf2wAPoqLqrUcY8eQLTTtVGpsP1L/4BTgPQPL2oRa65ynsImI4UplVS
8vPWD3EBRm1CXmr327qep6xpzrZJ0vwlf6SH4o+8y/eA5unFQLnuFFR7AEqvpN5WOdWhCo3rJEch
JootAHqzbTFSGqVUClvitJnPLNy87FxHu8mjJ/TGsFjZ68V6LWXOdVTa7PxjbtB05vJkO0Y/SGoT
7JLPq1ZHVdLRG9ifQNj5uHdW6OxL29PRPcQWF3wbXoIpt5y9n2tTKudc3bF2F9eZwaPJ+AgvH7TI
ZREza7wgo/5GS5+O0KYNjKCS4IXqcG9aoS7j4TwgKKu6Of4UE+GAOVclqIbDNjdZYN+fLvGnoOLo
oTWpSTMvXGda7dwund6GRld42108CLnm+mJbQU3PJpL/DHIRo2Ma3EUX3GUTQsqJ8+L/y91uPYEw
S2Oxm8SX+bFmz3+jco84s299kVzd4GGtODqOpiC3uESymkA7ouKbZXbd1l1td2Uk9IIvlicNc8Lr
qrAaeVDl6GlZd3lYNOg+7R2Qi9JArCUmCVmLmmAG+pVl9rte9XPhPuiW9fTee/qx6XQkWVEk7WpQ
R7xdQphLQ5I+br7culk/j2SYXnKHpGOHrGAE8gqCdl2S/coZRMGtONNIHwOXPVMo4xz1/a8egeKE
8hEEhlntYjczF4DnH7rJQ5mchj94zTFmmpM3zXjucL2CAkVfwvvo/FZ7i9Kwsb+ifvTZkK46xkhg
+YOF3eo6OAoqTzh7i3AG8/ZHGTYsqZOvYbPM5uRettL/OwYlhUvZmD8GT9/t2JK+7ruNf/9BAIEa
CFi8c1ZYW7rKoK+w0YBI2vMuxtfU+81VoIVVRI5v3GeoMG1PSjIGNwW5j393Eicc6U3Z1/hLNa5D
wQMvPFRbGBkqNY/iDbkLzFc71Rdeav/KdKW90Hju43eO1l8D1lVeH5WE7d6rXOtEVbUjOBpmp+m8
20z5inFLVamfT4XxeZ7oXrmrltDMMFP+M9EMgHPZbLlOQbN9aMNVfN9h9Fa0GIxrflX+HUTihIBp
5JWcW8+IlV/J4erxX3oOd6PGHcUSFB48xnduLN8CG7pxo1uby3L+Ee9dPmJyFzWzuObCXNmvFG6z
spd3TKb7p7q1wKl+GrIcVcWiQAuSxsRWYzZmwLJBResTMgTKPouOHGjwz8G/hGJ+Su1N5F7Ll3ME
UAszmo1FWVcej9luZLbauylSy/atXcVXEmL36lg5SkUi7zjtZZKPEP0Sxsx2VOESdR/Q4MLFD+IQ
oYIyIIbKvjDKAnoyX8z04PGJBbjlb49ywT82g/EUKS4e7MccqVa/Y6WMQICGRZM6IudGZSoyBrd0
Ld7To38DDLkGTBE79F/5Yy87mWPt7v9KhQfzu9CmMijANJd/gRpytLZ2V/ZqQ+W+GAdxnwrJxMG6
bbuHUv44SFR1PND8a7DMyhRlWjbkChmYyUH8ZHGb1+5QWO2Bcr+DzRQez5W25BQBXRaQrm9kZO+a
kI5wP7/c5x2PA7V5c3B220n/aP3BKC/8qXfnD9jiwA42vV5ze7lysAPZd4VaHAuwlseT+oM2zDOP
YbU9hE5QnCrm9Nm1xWNSpiuzwqBGVPf5ehTC+XMLR6dxtyXTEC1Xj++fgptRIgUoFMOOkOeHheD8
RX6ivyPGLWDPtUlpZnbhQ24ZwdTYjVOe8DTILa87BfXBvagbUlKWZm9tY++ciS9FKdodXVTsNnXH
P1uwXqsbMBaF0COQ6tTmIuKBCA0T6gtgt5/O0hBzGz4Sy7tdw4OXwrBRrgr4lfqAdVwcWU/TVOSe
+63sV+7HGVe6vKatepBkbt5at2Sqkudmq1a5FFHU0zghkc/sT8yzkCR+aci+MTqd/Ux0SovPvU7F
ME7kUISZR//1PDpbRSje76wobp+naSAkMtatOuEn4FQ9tbpaKJApKSxj6n3mXtKNVMNRmIsqoKyY
7jldkUP5scWemdF7YMa7zptFGhytVZk6r3+1nZdRe4w9toGdrCSRmJ7RU6Id9GEkLAqY5iNFgw4A
fp37htMmFJTJrtvidS7MkuXT3eyldwLgO9d/zOcRJWFdtrg0ysugzMljb+xPqfCadLToZb76E1Gh
YHCahZ08sNP8WhvCVQxH88iPhVq1MTFen3l7PMAz/5OaCNSdF2/zEO6mN8cK6MAecVDnVroblDe7
ShcCqfO86tzM0m5fBMfei+tj93uWQJeBiFGrN0kzPhRRFVS4269BRQITcynmHm4llKp373qmaGb4
ttRuxcNduCWqeBxygivJEn8cJRunwZZ65G4vHd7sP/LNzp6eeys2pzyNdrVZj8Tmk6qdkeMBnmGj
s7bG8Ew4EVVChSuOjiYLKUwHA0MxDYTQgANkjhF1sNit6zTsf5jZ7Si8NxSjb3pI2eKEmPYpe0JI
N108SEapq82UrTVjWHuTKKC7jYy3V0B0CNwNhbDYDew7iXxKz1NbRwlN1Y3KRbSben+PMzCMWFwx
tGn390jfAbPPLKUBzYptzELQaSAg93vtOeFdhnQ9s356DCbqHYYje7K/gXg+GioCrLgPoIktkcc5
khTZSeCO9UU8f3bqpJDwDY5ped57u5KpgRQrYQ8EAOrU4seYRZfiCFHKP745KmayJzzE5rLZtEh8
A1pJGoSfBXeFaz1y3S9WoJvtUQzF6S5eu6aHn+4H0sSuGO13qAYjHxC21L2mlIZQcboEcnMVbzNQ
c9i/do7mFpWFWX1ciNonEfL2ccWpvox66XFvLx+xO7ok7/CZwiWDSyXmmtmPIeHefEu8N0Z+Lbr/
wnX/iud79UUfs7Ejlvv9jSbcclGVC0NIDqa7dwSBbj7g7rN4/YpWuHfMsmjYqWjO/31nT/9FZZGJ
luLwaqaU23Om5OFtjvobxBGsShCsJ1SJH4h9XqCSKA5axReecwVuV9e92Sw9cVoajqYOOGboD2Ua
A5bZUNjK2RXm0UNMFpIkTlJ4zDPLAqsg6EPvmnvDCm1BkGpOm8dVsvBqAGNWuz/vzNZYBQVBjaGc
lKQVr/4H8F9m4y8AiSKV60keJwHV72sYpLv6uTQfz/ZnftjvjjVbFCAWKR9gCgxHNFiMgUgg/Ri/
YX2etuc1WTqS3/uso29UvHJy0bhofcjHUQtWSiuFca1zVDQATu21/mAaErO8ooVpGupsrXzc3+or
U0MhBlPxPZtpTe2/vT4YkTmj5clCuBprL+TtGFn7mVog3y/LcgV2g++R5Tmkz9gvtJS5fMNMeIqi
bjZUTGvPDf39Q37nxzNMaLPyHDXJtCVeHDIjutHWvE8HLiNxl94v9yfAUVjp24GYM5uHj0Zdsyte
mQIzsi5GxMHb5zFmEwKG/B5PfijV9mNTq2C4tWnifN+yxkj0AIpwcg/5+dpq8rcCsskHtwT9WMam
7cYyk/pG6XAOZ9r5rftOLW8JXOytaY45WA4bnIIMp2SoXpov+si3IRfvJXovYJruYr1QQ/bYdrHU
MooW9+JPXO9Ln43WbpDT7yeRJ6JOcqANyDBgE9qOfgI99ckmMHM5Nd/+vTbQs53Jjh2GpPK/Q23l
nTk6lhuufc8jFWqsi2qQfSbSOVy9TB8LTk9XXH4wxTbSmgjSQJ9WsXbl8r9sjYeqFYBbGZch+JEB
AoYvarWaFZAVm53F/nmKh5+SFtHXA+RnJGKpRgbPn0f2gMJjxv37ryjohVTEoJJD5r0k6SJl8z+e
/zINXTpqSTPT4MvSwVGj5NdD5in/HeB2Dv8N365l8fIN9WNHwJShkhjajLhcuN6x3G1aCK8uIMa0
adROuNstJaQ/xTWy5Csza6nFt2LtGgklCYAv/LlHZc39PFvErMDAtJkWSoMbAlsUxGmnR1S09igi
LY8yOCKmhTpm5EQMkanvRvjGj/TZ5rck9i52NY2BQPYdFuLX2jtrYjauwC+qlPk4D4p/2UpfeZHt
Txlusqq9I4KjSKzV0MWGp3GwZkyMwjh8e1aFg+mspGYr60du6kdgN0bepZ6YtLLZ6t6qJH0eRJwy
b5ZgY7s4dfzA1HlpMA6w8TXZBqQYnsA9R7mfJrNkdTlQkNX13ZytWJ0iWXOzTBWaiz5sz23vjvrZ
0NxhX9Cak+rx0U1PZBeurz8kQjBl4p3a0EphKBeQqBATs8MQGKghrHmgGmze+B5WuHEi9T8TfWLR
89PgHl8nT+tzuWysg7gpK98fFoqDLYcUlbVEK9BvnwM6kw7UXlcP4rgXO3iEp4oExOqt0UfOt8sX
RwyTemwXebFwacWd+6JO6LwXRfJAbdqgwHUa/hHJzfZqxeFzM/LenjVSncmyKfw1lzYDANvvruzv
NRQy6h3b8XwBlPMLQvBwtHWMfVuS75GBJtCsttoUNfkc252SgB478kO5A5FSxohu7vBVR+JakAjL
ptHILxRIgdwEfD8fLDZ47euqHkbL9F/TYMwVe95uN6PHAplYoRGrfiY0uszdEwJgO6pQNZyDy3me
pPc2oLK9lTDUy2TiJEwXsbSEHEbQgjHwlgSG+3RXXGsP02QQ8CiwmoNoXsn+3pJYQyi7ykulASsa
3tKBkIOdSaL59NvgHIfZvEqrLKRbIsFQHO9+vIg5Pu0xAS1cStnT/Hqgp9TnCyP8fXCv6mTPBafj
nATFSNWAdOmUbgLGBhYA9CDp3OxV8UiYByiCl84TfExU903tMyNc2w0QU+LTDr6K2MRXeD+RdMXR
ZqnFpfm7JK7u5uwxRpUTuawh04h8qf6pOk3CWMF55YIHztPXzk1I1U3IpwvUnRep/jN+oRIVnmAd
m38dqs1BlqIkTYDJOPyitex1Satau6mTapB/7Vw2LJt2STjWPFpWxXpn6QWnySCU2IWtvzCCkuD6
Hi6QY7ca4KV0lsj+9Q4ySUp6JvENXfX2Zu3IQxz56KAwrYHNQTqfAgM9hq/B1Mf8eru4xdHV+1am
RnCT8IVoRuliGqErcMIiEcEepxQhOJ3vc1MqwPCyEMoYmGhd5+h+d+MRH7EwADHMGMYu0ysUTUBi
dIahvEtYMNnjyMmjeebHwhTok6PG3C+TYtlpzdjJEOMIFJb0amyvmXR3t0WjLFuADndoG/sc4Hp3
6MmgkhH3XlsEXJS2+ZodaEoYGncZt9z6/nr0HR/WXPemARNXuZTLYtTFkFJeAXe7mQPYpPtR+wtg
itA70jEulL+w6nMme5ve+bgNGE7FRtkZxivEwtfE7qXTZFK/dEHtNcGHfhbFHbAEQiv1La/7c6Yd
xexjU3ZnVez4N/MSjgy7X40ZQNXIYv5Z3+J79sySJIdjF5AXpwSo9mkgIJLB8rPJXl1JezVBawh/
HAFdmfnpcwe3kBCf4oDb4+l8/bVAoYZMUdtQY4GBn5HY8vdc+ktYn9JjBxhzunSs+/OQtv3MGY+I
NBCEJjlu7GRLOGYzm3Zq9t+r4YVg+xneNlysiL8WMKl23N+OSTELDJyjklgN1gBHl2Om0lqeCXO0
fBBMpi4XFkeiC8W2Aquh3cLfqbUgSlljL0gMuBvAgRbx/Ok+pBwBGIwD/GMmKqtTDczSRoekXSkG
eZ6HDf6/DjtAcGWHZ3XZ7OL4fW5Uycpfk2Hh0G2OZk/09gYwLdJjSBNardR8XVITBH5oJg9YXevC
nAA0XWWRRwfHAECDKb+tuGgMWJBmAU3C/fr5ppoqv9JDMXW78fn0CebVwVRpgWEZnJbbv1fxTIdP
h7rK1QricdgfLqPwBevsXqPNMRXJX4bnorfSux/MxyPSmwHFbd488g2g1P8+DAgPr7918dLcveSU
mrSx7I3oASI2DrYWG/ytxeVk3Kb8MBYhov/6ChVNWYW+y2bu8J4WS86EylqwnReUE5eCYes5mkdh
YWjzi8jkO6Y66SYjBF9TWaD13e3VuOMHl7t2kskYDL/W9MWXqtPeT2gH966GPhhWoA4zGgmkgtXr
eQ3QEo1wpUL04dulqFOCQvfAfByreW71XuMXJzTKKXf1WB6aejQoX0yuW3i1aYYk+xBY+h/YlvJI
N5969v30EEq2bz2dzTLxZTzVcRPQJl+tsVSzVY6OCzc85Sk4Q7/dpLAHcl+Jm2Gc2ixPPgyW/Szb
4I/B9Xg0EIp0Kl6PXeJFBm5IZ25SUG0KfoY7BkqoIu2H0XQYMYlsAp3iDlVLVWSg+/OPKnlj0Pj5
7t89jtGv3ED7UX/i+PRQXXHWttpF72bPnQohzHEemfGZsmbig8x2KPB67lWgehTR6r2orUMMUMo6
8Em/7xHFLW88bVrhD4qEgqYTgyxsGMtjDs4f5I0fzjY1L1urFZyHezJfKHRUxLwjfM8dtKPsNxm2
aTZpkMqgFZ9xG+Qn5yFs3l6esuMKqlEtjNhxmKq4mel0aBvidBO0g5Z3swP57g10+caSxcxpXyBF
R1OmBJHmJw7aliDjYqdP0z4pOg9kFp5nHOotscvb5SZZKQ3s8fpR9cjz0aiqqoJZVzxZdQoHePwu
RGR6JKRKQATIokTDM6ZeXfjtkuA22ziaCiQTbpCd3dBKj7k5r1uZUssyMd1jl9rDY8ibNe2HCeRh
gKXyEa6/6BU+DTkM1X3y99DxqmVccU/emAC2WcyPRigWcT+ltMAEOozuZgy80IQUBtzYQ61HueWJ
NHsagllIVLXfEhYlmSfjwo76v7tpKJcxC6eEQEnG7kvJhtMXDy1vlgq5RRpo9rhPIQi81H6EyEa6
naiuGQpZLEwZmb9wQhHLPCc+aQwsbEFQodEFTEpmlwhzkuVwapmiFkuiulsvkyvUaM/p2iJWZnyk
g1QHnpFXqbBbnLBYcIRI+0U1gR/baeYM+OJwBHm97su0cErFHAjjbM/PRO2tH2dWPuJQX2sPgC6m
WpCuX3s/hEm3Eg52ZpoT5BvWNqtvzM5vROmZDqcJ0q2b9tlYSEwMJXlYdC97dV1vFIhe+7+JXLXq
TnOdhKqNRk/Hffvghn0HUASyPV7EkOso4zhAIIxpkKA4hltku9+9dyNiAgtNXlLuyfVCMD0WcxmG
0TGeCEzwKL8vFbEqvl2lZIWNJRHvPcFHD7L1gxUuyEZ0ZRMXiREIPXb0Gr4gfNaUQmNdCfCBZFjj
w74vPfKJyg53Z4ibwa0c3wqhc7WNHReBguOvhi06Mj1QnPI735UhqYwC6yVPMkNEAmZkRhxfi7fs
D81Tnjrt4FI13TBICyn8eM1kXM81r9xXdIX79VurDcJKgrlWs9YnuInePxKjz7BC1fsjg72KAhbL
gqAhbyodupCvZmg+PHq88hj/m1TJllwxW3083Xczqpqax/LKfJqc2JTIvMxl4+MPNApP20DnzWHd
ftzt2dQ1T5902XUp1gLspagQP5GK6QFDnfGjQh8a8vxjfhsGGd/5HdX4Nz1mekYmJG8wnQkVXB5s
a65PC0V2edpTY+Gm/GVnMQoLaZJjV7hqm44JDZjAXd/ALnQk2FZdEDGjpPhktRfJqQMMjyqDpbXa
ZQeP1p8ftY7q3n9s0M3uw1Aw/yaHYKkGau743y+aJWN18WbEsxarKU3ZkaBSP5xB6g8uPlTebU09
k/k9D6QhkFJ1wFoZa5M3yE7oZwysh6CVaAG9LR99A9IXb658mpnI8/3fVkn1cdrGesw6+1szZGFx
uDDKW728NhEv7U+u6RDtnm0F9HE5W1bp4ROLdP/58lcPlBB7UnwwOQCPwCb7KSo8dF3FZE2g2GIj
XQfMevherztJLLpvnuU5XtUCVT1+3QSyNqI8BwpO4bPA+VWacZy9leyXk3caFrJJPPy0WDcvYocw
R6n6ZdN8SqfkvZ6C/fO2t8VKzBllh2evY5oaqfy+SKA5EJfew1vWTXx3a6IiYN3KW02SN6EfRtSZ
W558/0rKy4tjVcXPGOBQHTEt9VmAvj+fPdrcvv1yuu4Np8XWhexmHsnAmwDwkbi6QKOjFmC9ErY1
IS7uZRUTLe1L9o+dnz0pgo4rrPWTUr1vno3U/C42bCYu55A26Wf74YJjeB+tSTxeqbYNbN3h4WZv
0kp9qBBkG/vsevdj06LGbQ4PHyMo0BMCUq8kvVlAiPXsx2tNe9JhhhuRxrnUs5gTTGeipID3VVnn
/RttBVO/1w9M8WX9WCdtrZVcPHmPu1ypn7xB2YaKgpbRYkh89udl1y5kLGto/sM0z3TC+Hnlaas4
pEO8/aJRXnlWMhhRDQknbhOLe7bk3VUzCDIeM8bY9BUvkuTp+XDmqAmecsx3J49b/eSgzxGqHXof
kLidVrCTEqQThVDc01gWwTSFWLpgyGuIQnPX3o7jYqPOZqIdcI9IfI+h45uDkD2EWyJviIjyJT8a
BE4xb5JDsyDsUYST1m1q5v+IhA1fI3jFwBM0z7RSpYLesebQDc/CqLErYSfoj78l539ndySdl5km
kc+JTUVA4kVo7DY+4YjtEhn3Nt0ULklh2VOhqZT6hAdmB0r4iBOyZXtFrfakqAeo1eqOrft+uZBo
07u7dE3oo8YsvQxbB4WzBRq/zIFTI9S8JDMEmjvUPE9ALKTQM2yMyyJ2Eq1aRM1LmDfDA16jeQF3
+npAlGey525hHu3iPMVKXiOb6huMLaG15NoF6wJTUHh9B2mTSTfgomAzrkxa1tzC55EQtCNwNtxV
a2/tOMexsi51V6JZwfX4lhmp56GKfjm/V9l/VcIUyMfFLDvflK74882+5z/fedYpQnfkhgeAuD69
Hiuq/8wl3Gp6apKj6vuNREytxsFcRHS+tGeTsQH3vdOCyu5gqPXxF+/B9grAlq9t8vbDs4g3U9Rz
/H5KLBEcdNyk+BjmJS3bAZ9tS6hmbVmIsogBdkEZ92HRx90Ra4+3q6p6LrRLdSqUY9TEay96dVBY
ZbG/S3YqLW7/i9GndKueH5BwnP86ZmzQL/6nHyrDqYkfmM1xGqidg1XQSAaN7FONmr0+hVNTE9i1
gMB8j8zTQTk9YFtAAdiw/5xD5GYcq41yNY7Fx6qMtvreZLK6R1R6+AmRcTdM/W+I2qzz48t4aQTQ
m/6jqHiZbkOiCRil1mjkRHX7HzP6hfKRS7urk3Z6rk4wz/mKfHSGOMe8YN6VzPVxyPhOX7OS8Y34
bVpElBbP1yJBnrAzYQOKSle4PsxUBQChdUqbw55/OxPhNzRlAZg9JRzAdrUOb/kiVwmaDeDoZmdY
8Iajc2TCts/SQcHdg3imtytsHv3t71H66odLbTuTR0Btj4mMV/MGhII5nnT3BcpY1GM9nmAat3GB
C0D2N2ZtFJVUw82GalbXraGuQxrTvm43WxED8UJSByzDwMmtv2r+eUNovZxbzTKtFzTZHfJpCTWe
qEt0tDKe4tr4kzMi9VFd/dPOTkbI/tCsfvOLyA0nksOz/wNKCzh0b0PRQXovwG9WpsOWhVzLdEw+
02X4aOfDyxf7IgxS1RgRVKDRVb08Pp5I0A5foXCpH8e9RtHezqoZfv4FYEatFNxLnx4p7ZRta2ZF
px5SFORVWIjzS1yCcxfAOgw5uxarYkw4SAvnSkTibBBbSeICPxgeMP/LdNd2M9MdU5Qnt+zULZhE
wPMv/9cHi6oIX98C89HVR0SzBmuybQVPVPSGafisHXFVIK/7ZI7wcVvmIKH9XJVbdRqGIoGHHibr
aAptqWHS0ZvOEekg+CYk4qDajvGlQtsq91QKB+wk5DRFiT5zFR/RP5qHucPRQcl/32RLktHZuoHk
znYyLUssVSow/mljQmNnQ13KaOH/5sBzMIUU3u0u4qKy1WS3yNtO8+g/t8L2aR1OtKFJOh4vS32J
a1aRK+bo2PaYS6LXA1LvBZ9wk99a6p66piqcpxrFRvF5anDO2y6g3ScYCmFL4lo4zI8Ou8k1wYGY
XSlz/N29ko0RuIx9zDknJ+4+7FVvFXLFfbT2tbiR72uQbZxqvlaNLsREyIc/YTMbyGrVQeXaepja
PVQ/bhihjQuDbCKwcFZC7OB6q5GqJOH1YCtOwLiOxWd2XTd2bIMM8JfmcGtdIBfNQUxyZfcVBocV
QpPIZFLaiKP2iykjMmBhmZkBAAtJTlP8sC/U0USwwrfIQbms0dpt6DyRUGhiJ2u14KsiEGk97vK4
wCvQ7fEYFeQC9mtO0uOd8h6mUgic2ATA0AtAjJgS2m4MFDP96CR1dkR1kgo6FJ3Qz17sT+nsL/c9
HK413WW7MkNYxZL3HD+qhVeQlzWMxfJCG9L4aS2v1hHNPE41DasZj07B1bqXsUPQGATnjsUC7WLI
ph1DG1lEYl4Ht7R87z+pNni5Z7Y4fRuP7JK5yvEL4vdbmwCpWhJv/Yy+IM6VjKtARzhrp2UWYXZp
J24Y8nz+4L7FqYvZTjAsQAtBu+gNwaRaqqPHteMXafz6bKioOT6ODTNZDUObYwE1B4CWOxH2M81W
A1Tyiywl9TW4WCSsTEgUsTdE68v/8SCqosrxtD9w6ttYkZvnixkuSEIXmLahrFbvXjbLFL6rF5xf
VADEXURUdxwaf/DMZzflO52tW2L8Z5B3qBsRSNK8/QzWUJAeyAcbaonrXGZKHteSvS3FiRM8oPEr
6ELLtT3K40mF6LSF8mW3GEpwQdcisqH97PzupoVm+2ImQbUi3rPOQtqxh82qu3WA8kNoDVM4ewEp
vqPK7nAiYgAQhpv+LiLUNLmpr8FQkFo+7oFOIhH7TyCumrqhsC461EiFm489dCzh7UcADmUPtYfn
3qi6eaVjn0xFNkvoyy6YIsONFGXNkMm2KcKxbvmd55HnsyM1CQAunEn1RXlQFcuBPKf6MO0rg5QR
PpX133Xjs160m2gO6SEqtnSAR+djj1ST4yCoHFJiMGVcvGRYmM+WCsRzZjEdqihQF3aCqwzSPE56
iMN2PBpe4gH1xmwIAXH1689HtgPRPNNdZ+TZS+LDrUdyz8+OqJPQFHSuxTfiVhnzHwxIsM14nIO2
7ATxx0hNqUL6o9JbNXc/+hNWBKJn7GDhr/fwUdcAMbTL/mJajiqWBmYyv+s9ppY+JFupZef0iYz8
s0KvGaWQvh9d90OPia5BoOVBw3gqGKPoCfcrfiJpjtwVx476oUlgbTUMTRREDgOTPmF0aSVkDMVn
E1eYQEVrngYDPnlyPRblUGS4c9kdK0nbQRdS4hXO9GV8gyMdwkxjCpFjDjCKrAScNToqXIztYq6f
CAiMGcols+qaI9ZuXj97g4J8/wmPojF4rqmHz4azd1gQVg4nkoJ/hBo93KPdr2ut+4JeNhPrRnb7
ZD6STrE6+MNCFfrlzSQvFoEiUWNmdB7GMX+Aru2GnS+fAuAa5B50JJS2yLDxlekNl4YJrEvzH+bZ
WecafiF2AKFfLWVoTU7nzJwS7WXUxJRssHmhiZ7plXXamA01ZurUrkNZxJzmYTlqxUAIepzi1zxz
CXwSU2S/kj8RkBZK62zqY9lWCGkHZsw33cKN1Pnvy1pNtaRtVs4SfHdV4TYnka1eRJfRdofXMeWL
DkTnhvaKaIXPa4vSAZRwRAD/P8WPpSdvinQ5LyiwwwQiH51sW9s14QMUponN+WTY4kIy8KVlJL6r
SjG1SKQ4DKPU8+H0UDt1hdJ7Q0uS8UlaitoNUUkkjVmXQ7FpfqkV+63LkLLocvqfjUBxa9+OQR/B
VPVK00j9pJqCG/lfb9cncrqxiCAnIZz2bu98KtBEVKzzoaXJ5pCqMlRr2yC7DkMU++Rbki4EUZo3
174qNA2GEnRlmTij36ccCgYioptEwpdV0HDeyOeqNAi8dEPoBtG/1ti3bRGN/5u3K2Y6rkivBHTz
RqgXoEMgTi1RKghYl/wxiI4PRrGCPjEMTfKMX1XlSLFFNyQLS7hKEVcHvr4aQf9Zf0/jVKaMpzTT
cTPATLmn/Op+dy/P20dZd8+D70OnQ51gimSfeYzMOrqu5TCj10N53fmkzmYZveuOYGu++/X92qfE
GU4bdqBVteNSclXwyO8kXIGgCQIxJMvGptoIYXaV932q9QxBNuifvkB/GE1CQvbmLrYUrIQrfYxY
Fw3SkWDbLS5a0jrmcZCEDa3AyCKENfQKsNDDrap3Aw8w/fjQ2nHvWInqOqmMo1YuzIvGqoDvbrud
XEbzKKlleYJcYg7DIRjh/UMCtN6Wo/VxbAFJ5HDGl6ENSN5PzDhRcV5j0O51MdkXoXzN3wJpob8h
+lnc9fDgWhDgi9hwnIfy7wEX3G1sAGWWSndMgqigCtEWw1Y26ye/bKXcQGqICiJdEuLOQGc4Qttk
6P+xbZXAZ+ohNO7kE7mCtfDaaE19dfLU1G9qdr0gCcIxcUvYvNwhd6sWRGab5krK13XYGWfuTtX9
qkDZYYc97cQ73fen86xSzOv1UVQjdG65s85/PODqfsl2Br3OPS0OJ+HZaNM2uvqDL+FZShlZDcEE
ZCM9Wlaxa26vnT3dUUJyd4njLQRNJ0D0GRsflULNK+dxyELCgnh3I/fIWlO1OvIQJvdYHdFOku3m
7r7qhgdW9dPMpWLHQ/+/gDSqso5KmRq5W7BLqfyxbBJZeo/PKDb3Fc6KTZs65i/+LxFiPRcV12Jm
2l9vVruQCRxTFBKhVZRwbjeTdwPDHC1mdc7HZvbv+hXq285fDC4kuzxOvQfRzqIGUE6y7QEoSETo
+ui35kv5GBqHI4oDIwljVyK6EIQmZLlRWQeYGLsQvGYzhEo8WAvACGaye55UnUhk5IiyDkNn76r8
gtJK9jKTuwFbiGPRZpSuh7Qrocs3ngGdQNqTf5L1ghKfmF8TEOafnjTCCB2OcAW9F4PgiAGtD/xU
l5qjO83AVTpEPKexq85nItmEAqLNOS5VuqTAq2slMgjHDB67j2WzuCNzLiN+Koar3Luz8CNvfbwG
XmguZ4mkKxAKzVTTvupyJ8LURulE61jHrUGSYJpkEO8yKsHJRSMLcmuN105MOxGGT0XuMoYKtv9B
4rJkALFhvG5uu/VWc/GTJLE4mZ0ORYfhiXPflWNDAadw9AR4iI1v0Pu27LkrWKmukmbr0vZMo2E3
atikOOlbi5de1wWz8syTyzGEuhXzdQb8C0QGyV+NuW907LUAY0cNQSGIBgA1IbG5zatvg0p0ZvQK
4m7p6XCQYYZcHrfloEQwQ/UFJ67jqWYOAabmySIEfQbsp7PSygqtSZIL+QJXJ2wHsUu100OT7olO
NiC0KUb9kuaHBY4S/qREKA74HTRiezJlfwfOZXMTotI0+KGlD1ZBFMpyqo9yUReOlUOBl7Md6h+E
aISx20VbuHHMF7ApbVY6GL7cZQ24Y5ebqfS4LPQitqNH01VbrIpxU37D9AVBhCam/CYIZImyjZgV
uZu3wU0HELRxz6Z6v6es2n6JCUYrinYNuWN6kisb54F5YEATmGHSBXcrmSl9YGcW1VV17KZ2Xxhd
uJtrwcMLS4DOFWY6XYxKIcjvV50jMVkaXD1oRdPEH8LLYxCmKuI3UT/a8Wx9om9XYFljgNqjdD3z
W/mQQpIhPMzBcn5eKBGB1sQa7m5hmUmsfMZPl1DeSkHorBC8LnD/KqDOo2q/Bw9HmnjxtpaK6+Hb
obXB/rCrkb4R7jhY0A20jq79Ngn6t1w4fi5QVN5F5XlVP54bqDYGYIJqoRg+xo4zySc+FVSfToC6
iwuMZ+/jQHoithcHwRPKD9n0YxzP9jEEmd1DgYSFmMRrt7MjsT6Sc2E3y+iWVvWXphBloh4v77hk
iOQO5iFHgsMTTLCztN8khm8JO/AhfdO5rW7tGbNGcwllJr55jaRgisbjsfVnQF/WzHUjPsE+qlso
9dPdHWRiLZwq6t/vRa7cXKradMTnYQhMcRc6//rZN6nrQnzBk+qwdKkhY+ILHjqUyVZrAShJMJ/N
kYvhXuSWBG+QW4i7pCPvkZesRlcmkiYuPxrRYuZzGHGKyb7XdmKxPXORXMqnWCBVqSpSVmNxy/L2
T0d3PCsCtCcsiy5KgHHksKGbLipdpYENksgM1N9ivQLOi3h5Dn4fYkv02iepddFDoht56jfPdF02
98BVxzqPb2Oq5y0yTDYb37hXr9SZiVENLZJ08iXOBNtl72i1aIfNug8+SUcHASJxKqOjGBVi1UHl
+MGBBKyE4TXvmGuqDHG9Gh24gWyJH2Hojyq9IWso0ByD+rVIggkAOyuJF0Nbnoi/gds59ZeKysHV
jOmBBNKuOhxH82AWTYT4y61M3+ljwrY2lZCgZQlWSQeNoW0GJkXYFpgppQoFUNZP35DDHi+Ds3NZ
SpGkLmVjy/lxuGBhebausI8qnoCBM9bqds6X9c1CWWTl7zO/7l06FISoEgyTEsFoLeVZtNULhSgO
4YO1rRV87Oe74++hSzTthxRSz+3Mdgsdiace9rNTg8+ttEup1ErvzbjmbX1m/RsOFaMFYdPBWS+p
AwqgmpVGOBF6yxOcPhbOUkPwVYeup+jAqM7j36t82unZGf5E7DtfDfrXyqr1VXAKNyY2q2ARbmSh
OhSXB3odg+u2UFbj07RsKPyzFt8aJqiRZILUpmRX6BQFEm6CJKsNQgBvHX+7A5eU/ocit6shBc/B
kFJ/EbShOu3S5DFzJZ8BiAFUtB7bwrgP0ji616SJFy9jlvCuiH8RyS7zK6o/1Mf727MdJKx63f5A
sJFlvye+ugJzkqsqzYjtBIZVFjc2QNrLfSdTSz5fD2tZFf4zEoSBf1b4C6gwHFL/lZ946h1sqm1Q
wAO+G3R5rp95XcDOurAJcZBVB6IMSUYPu5KIwvEbNyu4LJlAYbnjfRdESh67Yz/1NqoGvk6t3IgG
NadfgoeIm8RTN1GTzWaxCqYyfR87hE10XmWSiu3Wt+8Wye1G67/j5ogeHi57h67eRQcISdRvIjL7
dNt91AzIPXwvvDny9G6hwgOQqMz1lIQr70H5vgMjaAJEYQUQngsZC8/HnSfGGLJH28NR1954QIC6
HSxIrYHz2XS7glzdpy3R329St0BWC2Yk8ZdhqK0bhgSDB67KUP4lbj9NQWZjW9pQLu1R9O32QMDG
IoCAXi9PuuSGXT09sfYUvKkFyBGzWX4GgWqMQLwflQ+ncgsUBKz/Z5ydbBMb2uly6VkxKSjYC2xu
9W0CSquuGE1PgMq4pur2WMGAaboW/XGeIPe27DePaMxjhU8wygtgzdLS7m8KIuQKvr4/3RBAJjf2
WJgFxZFoIs3WqCbdgPXiuKtSDXfFmiek3KYPYwjyLItxf1V0CO2ZJpsc3e/hwZ/FFiwDdsuPCKQc
NArH28As1LLvv3WN0qGPrM6paLUIm1LVlwBmcd6q7IzGfY7FA8S2OSvZzv4yON6eWGxF7xtrVo3j
eN/Yhx93xgPdvmEcGBCCqTeo7DWAWf8YnjzzkKhqzglWIqwrUNZ59Y8upK/pjzoHP1PNSRlHgikL
Ff+YsUhdT1DAgPO20oH8UgcvNpIdRRHWrQmfhuSyvIsYDYtYvLWVA3NPPZ2tzzvhcaSDsjiM2aes
tW4t9Kvt3Te+F4HYX1/BiSD1si91H1ChLm8NlQfK1hWp5YBwYU4Fq3GGa6ic6Z87jFmYX6RUDCEd
UlBzK/UHOPP4pw3u9SQkXDq7Je6PE+ccwOxZuM3iB48paq3VcEiDwr8ugLmKMjU9SkhxPSkdNAw7
KVovLNLzjcVW3Gng1V/8eNho8m82/scTbP1WvQFG2XORVa5tHluTZA0yUAvMEM0GgE7v4Ja77Xi8
IXavXqIfQTBr8wiI3Lj5GyhNXVzAY4kBR+XfK6uF+q0jkdF+cWfzdJ1AJ+OVtQj1Kqbxg1O75R2r
fCtiIcUTa74LrtPvlnMUsSJbgBO8g3Du3K6dixFs2LrdU6rBXeqe8QugiATB7g6b+Cy25j5pK+b2
0OiHkf5aXZLkx4VRIG3jgwqTqL4ioiGUM8SiOJumQel0HcjUmkWawnurjQMjH3o9J7/jkwKBqoeL
Ugs5V09q9YP7A1CS0H/0Ln1Bz9fYV3PTy9AKPGiyWes43EliF2m/Fw7g/0CM4KE1dYw8CscQ1qgO
60V35XYZvX1wd12lb9TtKsxQsYK0u+UfCOX1DUOBIrpG4Q6s9DH5oerp7LZRmmlzOm04Yp4+HGr4
SZfFG70TGRdYi3OPIfdFehthVA40NKwYeiacFf+QTMiTsIdFVRd0S9w+BZGSjRpTa63yfuhGWyTj
UTxPMUJKXSwU+NsZJRPtlHzR6Ld17CtKeVZwSeHs9fJAN4WTAEChJ9i/ZLj7/rQrT5xpGrtpMkPV
Zj8OOzzUsq+7ibjx9N88dCRVomMkegxq4vQW2INKm+6pK9hx4vnM0K0g9BAILGO2QOjw7byKwepI
Q2FyPilPZ6Hlja27mlDCzU+tC3vh4vBT4LQCal5RdPdI1LAlf7Ae94/wEUYDusy2QkWpMqFfAQ0K
xRIL51oFU4JHeT3l6wMjFM7uIAni+3lkbMxmq+tfatlZa1kksOBnpOFLiyMU9Tif4qjpVNy9sbk+
Jp2cCTINQNBkrlhvLQ99vQx7H6rF/VdFVEUwhrEqFTTrDB8fr8OHTtTOrSspA0rSXMMPYctLr/vS
e5hBIZlmMFXrNssjW8l9KIIPm9H3bgf3qYPho0um/MUSjKfVOijlfWXM0qAgsG7ho847oIPy0JvU
cOakgBojSrxxOPL7Rzv4HMJK37vWfVUaLDUQykr1t4aKeip5xx2o+ZWk48mbJ8Z8u+GZBoAat+7N
0bUq7qzrm+Z2dMli1d0p0gDoTdo+1ZXv8oyqFXJ+LATgByKOJiss2z/8rp8Z+3/SlL5gYKd6r4Zq
fgbiw7V0U8DXYiSZbEsIfRrfL9Oau664VqZQ67F6CsIHNJGBGWvtrM1tJC5nije+1nfVdQnTXSue
SN6HVnfiQIC8Re0a2Q81LdBnWfN9/pAQ+KJT1rruZQiju6SVVLVPtzyk145Hu6CZC6vevw9n1vFh
ZbPiNzaIUrRv7TxcnW1we2wYvXj0ApdDv/gynn8yzm2iClyGKl3uJlm+z9ZX+NZUfoFMaUfd8UUt
0BoEYYTKvh8yDwPYbm5lZYqMO2Ir3owIoI67Jj8NAQQlDytflE01bQtImybS5RLZScACeGb1Y3Mt
TdPOAUTRtyRE8y99s3CSdsQUv4vsZokSfzkScshZVJFz9l6KzCV9ibKHgI2GX+vzl0SWpu6tb5+F
XP85PudF5fUz592N/uLtoonP6eQLt10ez0QUxNCSdbr8P/6aVABa+lf5htbtS4Kg38q3y+1NihYj
oKfb5kKbjdFYPOLUx3pyci9ivSsqzSjSC5NPidha2W4xBZO5N4zotn0OeZmaHKn6hU5M0fQrLiHY
9cf9NYfCfHJH1R4ZGnQ79+ZVmUHOyZQOHCFDKY6hMa2tlFxxqH1xOtUiiOwMoKAxr9FIinid0U65
M88jQtozbJqiZUNdoKOXVD0xQrTgXrJc5CaH2ugevdrsq2XSYn9Qe11p2BcuPusl0mekmnAHUnWW
6//hWzfvKPFEZJrVeR/biD5YxCegsT13kAI+Uloi5nCVXrPiIRb9xqCyWccUBCw2cebZFaXDAgAE
0y7r0f1lfcd9jdc+fdqkK21r69CBMERuknBOQEdMjkpHaPum2I86FO9Ms/heIXpWJxBa/3FHbBLE
+yYkKvACpiXhDKInk0MBQG2O5agER5bRZlUPNjIzfBlLIy492bUkg8X1TYpHL0lTlWbDUcLkamKi
U++zYN2GD5WeX9QP3LGZObrSxmoYfgh0Wtq9TCqdyCrPFHYjjOtSGzy6tBPdhdd0B1GtPupO0CMT
LD6jcdWT48ETS6IxVKhG1sDxGRbdQTP5o/eN+/fL8ZPvpIHnULlcl1Xbg5T6b7VUtCr1rxuwMfY2
0MOckyt9xwPCMNxcPBcrQQNI5ezQlypASxkudNcpLep9GVkVSobdUHcOGxV+GzPHtCVXQ9N14L/7
8hTNFx7f69qntsbVICS2UVSBbYjCH2jO5SAK4sYaLdee6YZBS0cgcDuu4jLbE6/zYdxyF0hdaljI
/edPwhc9WAXK9ovqTxOmCWFnvWMV6p6vmqZfuzpu2zZZ4J3F1qvstN44Jsgr6sQWTf88R56sDJjk
JcQK8iqCUY0wvHoaDQoUJRCRgsawiVN81uru0Rt0Hri+DCKlk/2eWGE3aI/+hBi54epBiOChIy65
+yLUlY9ZNF5x5YFIc6sADNMVJTy3XG0m+0fHEBXc/LGe+lalAdZBbNgaRTI4nWdO8rf5p0l62dB+
EHF1LsUEtW+5LuuBVvdz/5kvFiqcG8lMA4R6qNRuSqPzVyLWY0YcR5WAVeB5yEOg9eK5hRWCczoG
sNE9cLQDZlVfYlONHz2FEK5gYvaTKqssK74ro04yOLf/3qV8JqmLewdB+KBVTC95BMkamaY0+y4d
VEq8cKEe/TDr8VHlfEvub/5oyI54wYlxWGE+1l29zuB53JHti32msQWbQjZq4qLKQdFjRJJUW/+L
Q45D/JOti3aACDI0xo3+SXAl4WCcNSMW5Pe6kvvwSvLr6Ss+mz3t9iX3gd0feqyA5lZTGoZ58/db
/ZdsfFtTAmuFjOCgoO9xORYe2n8aSYZ9MT33yAR0tNP/YwpcyYOKCmKHu0K+QBCtbzDY2xpxEJ5L
qSsDGXRrB+ogWuWqfG1nqwLXDWm2gBTzT7lFtkLVOLcM/bdjcC7OV02mAWtjB1MVz/Gh6s/Dk5r2
UjpIDYXvVWWFTthWKoq1fqkyUq9cAi7LjVoc2AL6ba3ieVRb8dQKZ4v9PNjFJ036tGW7nZCEIK6t
yx/d6ClsTS2xhRptUFu3mSWlO3rkwtjn8B33uzirkIxBHQiOtw3FWeYwjFVmLaEnuntmfyyaLS+f
9h+XhVPvLS13ZCW+MvkVqAHmrV5ey8w7HQ5c6sPg7K28IiHdWz9jvSH1w/K/LGbmcfLEuZTqQKAM
ye5s7eNprrtTJzU8GQcdd5YI26WdhgrImeb3Lm+eFW/PUTCP0xKQl+kzsG4J1k2rxjtOtGDVSRUs
cIPoZSl8AiQtU8Vi+BQOAziBHMY+rnklcwC/A2aKE1e3dLn35AFzZifV5Z82+/EtBBfM8AcaiHpn
eCIiSUzw9GK8NfC4ImSHRoshJYGPfR2Pknk+WLRO3kcrRpxqz4g3Bab8MDrGXX1UmVCZ5aWvQYIz
IWhInJgc6we1b4Dul8MJl2c4TuX7uKsUmgGaWKqytZ7Hlp8O50QUuV/KmfmEDDkZlA7EadpkZ+Xm
8Tk/Pb6315Q8ou3RApwnzj/4BRJhiFSK5ZmVvUhWCa3MrzVphlLXBmdbe2l2AdyL44+evIOeckxI
WGM/dQxBoVLpepf5xCYZtd4YJIZxK+V+MgPcQf3oFR44kna7FuwC6bjkKVM15gNGFtGy1wiOI2E+
C/jiGvgYb6dImoHhVBNPeqmmYqPTwdcoTz21jBXN0bLeYg+qiEwkDYn4EGNyWUPWnFRyNriMNBhf
ULXT9XPRbgqntyounS+OowQucN64RF/QosXmaywACZ51atvnsj1LZdemilcynC1K2fU28U1RTiGV
+bUSn/AYY9RaMXBNwOce6vqwE8YjlCnlDJ+1qgWX2Fu3xWEDsg4YzeuaFsd37B9oyF7s4DqnCNGz
aQRcAyiNYMf5ZQ8l/gmn7IZ/901QPfq2A6FcXESExbRrEz3lYC89h2n7ZAUT5NV5nyNq/BU/qluJ
PHYwuGhZevpNBg7o/RDysO5NlNUku7Khczb3EGXbDJb06FXOu0h82tXKOPRfbQKT9yHskwUNoWIH
5O2Tk5bksz3lgU0oi+AkAYPmzQeCVHh5FAtYkuHkN/da+yVmy5QufdBKUvjslkE9ozmVY+4+n8+q
OeuJlu6bBCIyCIHj65WQ4HVzcXDV4nsqt4HJhsQAqtJwP7WtNhA247xHTa8lTMpPjjr82tiBrDBt
Ly9iPfkLKu5nHJho0SPBR7479qoMf79nFWIdsv8KAmknOPN8wokcM5UF+kpVTjSkNk/VUoPPlSVW
9kklUJmhwZg9JyCO05bJiR8rTErPtx67Uwqo0EuO0f8Oncur1cTbtVodIe9OlvoAY/T52KfNX6aM
dJRaM+i+TmE8CNCaoxj+BIoSALFBBVdo0qGBASxZRU/PLrcF4fDmXuhTa6047FdA9GmZEOc4kN/F
shhROThgTLhn2ZANXEQMl7zu+RpClJ0SoaABC3M0ibQMwSfRaevC85nukIk73RH/1ouixr2qblwn
y8CBZ4vFahDCI7bZup7W9vkLUJlTHHt/lwiWkP0sHwjbrS3Cx8cLbPcWPZTXxTFytBzjrf3IY7nQ
JJPz1WbzCrcTZZjTx8xMGjyRef4NGVlRV/Y3+hZpRV9lmq0fnRUuWTcGJ64uxiNTnNv4KNAANbJo
G/sHQNWEWz2Dkb+G8wPRUS2Dq646Of4MNUVs1GebVOEdINF/zx3id91F3FMhNffztGeR4D8mg7Ec
sLlPud4hQZrWK2poa/UqXXLl1PR7YMDY0WldnpY70QWDE3F35kAnHxegeLkQuPsxH64s/sK8V42b
xSAJu0eDALgBzUlcLPgU0OWQ23x9qcFGsXYWsFmctdmxgDrXwLC2xnt6J225qDU9aWjdEBGwYGQd
hr5SWVsCkCiVSeknQ141/QhYYt4H4vgeLyDNd5ZwJ9wbvCu3hlZwB+7PQTTPgY2NWTp4BgZck7+D
cuNt5rVl56FViGYUy1035VgezSX9kI/r93FxBHPtJOR6d5XA49O/t/HIehdNF0glJqajF2p2BwfU
lYpS6F9DrLXs3pN2xpMOYNILCrTPmtf15Oedcj8L1OY7xZrtfTX9WjV4ou2663E1W77s7P1zLwtE
DPqPAdBjgbSMgPPgHDSARg3t0HF+bRuAZb8p3w+aVM3YyXsflUYaEuIkFLgL7cGObf8/Dq6Z06/D
GgYhyQ8YEt+YaTFumKrAyYwIt58ZcRHeKEtxdE9dJOILFQkMeQVPg1wdeSFimndeSQ3Gh//RKY5l
Cvyso/tqgkXvrxmCBmMcZcgitKASBcorFtgRl5OVNq7ZLD8fNKWJHbb3kQVXZlqMzJFAxJaehCbn
DknfJrDkKd+s7xsCqFrKmM9iCguR3meVIW27KNycfu0HzxwhDjUY7cMCNn96Rvts9FRO6qkaXqKa
2Gi2QGiW41yNPo+2ry8jmyvHhIHAt3kWH+xcy2C2gJBTne6ngell50jgieXFPIQT90t8NMXFUMjC
tNHzT6XSh4LAh68qNhmI6VvcftTRb3myfwLz09lZb41+3CBgdah+hNCDclw+RLU30dciFxTRXsLF
j8Q6TVP+4pmPPTAU+yAqA3JMzlGHRMcgdsJn2l3K/7tNfJgBGTUweLIbpj+/M5pPLg2uharXCPWn
JFX1/dtEgsCOYAFTalvdc+oTQW5o7OiqMcmib0fCPEOBrmfmYmZgPWzmIIQiYkVcj92XEFcCtWC9
JnLiwBCM0OJd9zRiOyo9lLaFq72peKKhu1g2SVOpTRXbfwWTIe3GtoMOWda+M3hv5YYZwzkQdKlZ
xn1YLapR+xUO6ISHnOnlwV1FoNX4cYI9NimMBlvH9UAHmpTcq3jBvXGleMHxuezYsqwQtLE4+MxR
mhaeh5kwjcls1nLHB9MzMhg2JsIGkcoH1zGZCtGzS62Sd2kO4cj5BaGerCzFOLYraFSSw6W5eNS7
WI8HT5sRGRnORFK6awN5z/Idl1d0OkDK3rygvzu8j345XOUzeBtc3mJUjg56jme40ik7Ua2hJ9ev
SJAB1DojWI5dA7T8W2wgqlrAiSGojsDQl5ariKE6y436s59pjzmKjtPCj2RVCIp3Yc0smHc9G1VB
gcYcuSH3yEzyUQwJcgl8Bs4abeP7s+SssFAb2DKCZgm9BBcVFlcRANEfoxKqX2DRCuVTgQDk9m9h
wRYSpXVqFcRCrIzzmAA3O0I7UHav4dwvdRoJjnKwbpV8pwRYlvxgJEn18iW3DrWfJxifMYORZ/Em
pYYlgXiHYHRr1JU2H6ciN0lWOrr2FRGdMdnR5nnglaErcSGbSa8i2Z8vJUSC0e6V725Mraauccrg
gE1EEQy7pOrYvHvLS41niQBtArrq3684Kg7VDnfo6Jc0139uHl11+/BZ4YegfA21IvUAdF4P4TY+
UzK2Isq0A6lrdA+NZRFDCqcpNFLeh4Z+2zPQzv5BFfU/m36YC2+XURkpqrJ1pxoGd6AI+lib+XNd
ThGFU3yUF/ZhUuwD7hCAhDmy50yWYskzjij4ICrw7ejB1JQ2qLokUSGWXj5ZSQIKz31N91xVDrAN
Gs6NiNdY5pOs6+aec7WDDOtalgfQtj1uO3GSbkUBdovBy7A8pAAn1Nyydp404vFxDGLfb8LjgQYF
z5irXJK4y7IIevwIOCQEGLj6eCGQa3GjKOmGRUTYHqTmSXOjYjNLRpqslDuusHXegJJL3lc1l3y8
k/5H3u5IwJ4+WOS7weKBEYWkal/AJY/iN8xkdagueFkeS/QzuTWdMT4o0XGVljkwj4BjBC89dFMi
6P7E9jehP/xpPY6PX1yuK4flq6AdzdL2sERmdLNozEWKGXp+Of2nFE71uUkV4uj01PYkZPC9j3J9
yvf2EqGvLHyGcsEiiMe931uUGNSE7Nm4Dlp4C8ymPszU48JAjWPa3Kgo2dbBmueIBb6VXKNT1nJg
aGt4Q+Ljk8a13/k9YTMKpZFmogqhFG4MVxzBetWLPTayK6W9UoqtrntHFc+uGS2tJE07vopBaV27
Q+sQW5TXOe47Tnt+Z6wnf/R/racc276Y64nJojidZ3GsmwX93lQIfTkalRCmwq70QZjUQNILnHMr
FqWXK7JOpPuqaXhsJrdEx9J7rAndEpdIOSA54Ed5kdKBqNy5439ZDSjCTGSuvYCcXY2BYNAKyaWa
47RgKK+ZfYVfVkxEG5uJUSGzKur9S4/rRc87zb5jOA/ewcT2xl98sT9jMgYxnNjR9Hsj5LEUtBfE
6FZLnp1RyhSXfuLkhmtFA4L/jBtV02GqFWQez0K+lDRFYk2TvSJ+ZptMGl0sdkvii/GSyk6Gmnws
L0jtX49EPlRkJ/kxX6Og/BfdH5Ib+xXi5mHmbAMnb0vhAQp2sk4uvhgQR3XA/FwUVXCctfaqQEEF
M+Cm/ChheKH194aRxrb2vnVP4pjADbOktZJDV4vrxIpqBqAOekgiSaGZoV4kDW0gf1WrKABfM7E3
H6Je3HKW+5op7l3CWwqGVFZ0sqsKSBVhNxWyNspB2mMS+LCYCfahflSbCYU79TE/tPpPFzQvuPz3
m/swPuYwt3waNDXSBPugYc7ANFgnJzHYOMP6F0CCO8fNzjzKS6OId7c24far1a5B/vBDxoujGDCz
zxvo4HLnewC1/k0JVk2g5gai+xcPX2X4BE2XmOIthlAxzr/Y3tbJ2YgUe7xi3rTZHNMru/7XB6yU
Htlk/E1Gfiomz3DZRiH3bD+uv5UcnIMBQlProbZMzbFucDpbFRS1dBc1KlPa9nAUghdjHZEmS5Yk
Jmx7yknl+NoP9s5HHS4cx3GdHqJ6XShEmbLrsUld8M35Tt347lkD2in+yrW5P+3aXkHXKZxO38oF
shwdqbhLCN0vJEMjCV3/D50SsiV551dh2lxKeF2TJkL2KTsATWE5zZk2ehZY9SZ121BSPoFGx0+v
xOQvoVfSpBNItvI7Jq7T2UYM8TS4VVR6wn4UBWMq19SxItDrGGple5Psslbv5b6b6cjnz+048LhS
fzzj/wD3qGJt2pb6pEKSbB1jlvP8GF/MHdfzu5W+KJa+jn7bx8ghXbEPxoTC3ZhmwqODX3FAPjgo
bAqNGq1k2tBI4es+MQuV8frNARtk2W73t75+m5LLSXvcaUdCM9udo1xKDX+2tSMwrSSL3JecbLB/
ixpLObL0+xTyjQeUo6SZL/VuBKndldtx5BGDpH2OP9u3RsU7cPwWSEV0/j7ZpxFDsp9WXA7FYDaz
1jZrHxT4HAVRgTfKRJJoyUbLX/UdicPGJeXxg42Ij/jBTU+aZhNrmH11gHGvALjvAco9kz9+LA/z
hpeIOtKSOJm+QXXavvPWC/XY7UOfE6j2EKOdj+sAuepWg6Ab/T29RoRjatqZu9C/8/4FacSwPSIr
+q6QnqUVNfkRcxIsNQqgm/T0NDaEMU6CSXmfYRV+ZklhxUqP39kfTwFildStNT80lqIbxy49nbwF
D52JXv6prNeLgZyUCnN1EdRZm9N+OiAKC5Q2LsnODWCqF6hyNrI5fsQEjMXz8fseX9UqOUYLA/dE
rZhlRNcscDe4/UIwFuqDspQ9TwrnJzFlFqXolgxiH+R1DlgL+eOeBBcUKuluFJhtyV1ZSClizV3o
LH5WJqjTlp8DNXDJi41AsWpprdSP36BfOvSaGA/Iqd1loLp3quD1lpv9M5c8N0My90Fl6R9LrMaz
w+hKPsR+w8erENeBe4y3U/FWA4NaU05PObIRwgAqIYZMknWom+v71qV3+GjUg1tf0Uw9G6ACDeRz
znx7ZJaPF8zpZLliDMysipMmxILYgU37CmizDRQ2UA9Xi1vGFn6p+HCVP3gg2MnuE0xRUb/5lM1q
pcX1cW6iMyek0T+VN4cXMVE/6bEYpSrImXyFVnJuQY3J0LBN8hYqm3+oO9Sp6mmd1A1LOXhSV/Iq
+mHYnrztOOVc5qvrKXS3lGMRLVCxI+l/pe0QHfdWpG6x1CXcliV8yzGqAsrbGuQSSMn/FrAzBJdA
uirzRkrvdfoddrkHhQRdeI0b/buCE7hMTQisS5qULc+IEGctGeCNAgTcO0NiPOH9rbmqLMlj7uiI
prtihPwbzYigYnIPBs/otBVVTYs7XLHWl/6as4AUBEIadt9Kx3MzA6TaCu9NJKl8RCFYmRvl0qtf
TjUJDsuojFTHdmv0sPbDE1nBZ2k9Ug+al+gli5urQT0AJD4OXgi66k/Ltdh7c1M9lP46K8Wt7RFI
tM1cPtF1JrI1OSDPQrQSg9lKrF6+SC4tCmkbH2bzfTDWcfp+kMFzgxxteCv8Qb1e6cb6byLHq9v7
KW6pFSZm49Dsk4YCn67dC/UCmNb6oO+dZqpv9dB5refxVcZ5d0KIyStsybqolBGc3Ll298zlgZwO
KHxZ1JiNdg0k1225PS/57N6xdb59KKMWFHKfmTZ2htJI89uLuuBtdAQV8H6q8WkPUm1Yl4QuvnCV
n+6UVmx7YY6tNWFC3L4BWyTD/wT7R/YDkvSerYqlvjK3ULzLhnmoKZatgb9st35mWo3mYXP/bK5A
4L/aeU/jhRwP2xdwa2af3uIOvtT6Dbgatyb5s695fU3EbuS1QXgR2smZjZboN2UdvSJXmrnkntfb
DAclpAD4SktzOOZPuswE08XvYQg0nnW2cy3cTerqMbBai7l936Qmw8USY65+4G3r9aTYOEtxB7hJ
0fLAea0KSeJdGlLu4hJRSnnZZJnJ1+TJfv8g7S418GSajmxigP2TOlytoLfjZAu+j8v1ulCA8Rbp
148beFKdnTLUTbfAFTOTBQMXSbFE1X2i+S+SugbHmj81Fhx1p9hNKBoq8rCC8XSv5j5/IBdSLeVu
1e5N0lO3zSm1PwxlG706Mqt+P4ScjpZqKb4JK8nfdeseShK3p6fI37TsFFTou2PepSUgS6eDGlw6
8qPwLGnuXCkgd9h+fDfhHbgvNrgCI1ehvrE4mQR4hdZIsl70pD7bPXiJf2gwaVK2fsfovxUy87L2
U2l5a8wRxJXnad0nHVNxV8toQGYSnjNJVl5xOVKRVFaVq4gntqiwL7q7hDCKlKUMVbQWDcwZIlIO
q64KnJkmNODqfibKJB9D/C7Urh7YHcR/eRGf4MYXk8ZK0MYmLJxSyhyDWEo3JCe4Ef8JBj4CTufO
G5Z6kw+xwZPo5xAYYAoIIfU1DRwdGIWbPbPl3rt01oZvAbiTsbMhpFI9NvJ6AOYDrHB210hqU4FD
/MPmxV0DlzxnHhGVS6gcluKmydBA59JQC0pHOoNmG1yw/uI+G3Eg9KdwWDOgE53Wyf7j0tO9f4eI
koUi/MI428OQOS2ViBJWXebxpXQe9pTmOhPi0hpKuJkzGDPkxHJqDPkJ4LngWLwl0JKnDecAzbe5
OreE4PGRvfLe59YubiNNkF6e3LfNJg7dabCarkrY8nW9ns85PW2ad47sxp2jCV0EpJ5Y1np5/PDW
fQJtZstRU0T3BllYiqAm/TEZmCaaYssJ2hQN7pD6tDr3VshvshC45Q5QnM8v+CyyftQUcZDXBSzH
xFG5j3cc9z4fKgo7T1xne44pB0sS3FWEhqFpfg+xvCSA0j8m9aFKwCdK6LzmcQyYgnRbc3Kg+hZ/
bGZf2LQ+LSVj2DL7U7VxFWa3KXEwYXDJDEI5BzaCojV/W+ppOFieaDnGFGwV5J8kitQ9cB/foKJu
PovMC0MxycwuZZRL5IyjoZQhPWSjbu/XlgjwNHxPa+owVdhKMlyxIgxPJ6WjWpyKa+Yu2YpquuD0
zVAS3stbc6HVr0PdgmhkJWKdVvW31b7d+d5FyCBb4AHtpKWfAyCcrOnF8AuZZAW2iP5LiqciKYUl
sHcr2cba/RDs0TFC3b/5dXcvOFrb7Ge5yhVWz+UCOMkbyFhv0yKavhGH4htzBNX6JqkCEU5+szvB
NC0du+BAlfI8EwTH/aGPB3PiF4PbvnPZwSc0OOQBM4ipEdO3PodB4UPrc5qgRUQR8IpQLkrk+/j8
ax/GiETQ8IzNH3KOR1F/idP+b9pkHOVJqlKoShFyl6NVrcds5jFJJJ3M507++bOI24PneJrfu+uk
DDuVV6KFVE9UVFYYY3maBjnDZPzVYuEBlcT2pIFLa8VD3IBAWCJYEK9A+IYzt3sgw5YrydtpRSWx
KoYzLAvSH7zTNZqpjZaf6rI4XVBPlWnZvC9sOcEfOhqEDPflCvwW5oxSYsA4zhS9kawNORQw8HaI
sM4KV8YgqzU9I/xwNf3jFZH2kmVmLJN1JSR0KaQW1S1lq/zgoPok5vCKQRFil4ks+BnKFYT31r0f
iFhSvPfA43Wyh1zaxtPqG4xgZxU5kuAWlrBOBQsqmOcYGhQ5tEs2d5nhArADnNtfv0vE2X5CGvwe
J1bDPtVR1Npk6SZw3jR2PLJj8B3dWRvGX8ujvPDyHYN7DZtKgU2zAwfcQKjYv92WGnCq7JmW+Gmm
Sr5XxbuhyiDczqlUWRzApDu/U0XvqWGw/QbIs8pxquSCTEk5mur3PFtLZzMaGF4Dbk44EbnVRaSR
AAzX76FhyzX+5Gqq5fWASHs0oQHFVnmGwU83a6jblNkO5FAVFBvQnV0qXnaZE6PUUuDXvasjHUq0
C4pXO+uFtN3/72lQp2ZtsR6uyBA9CMelMBUjlL3/Ar7RqHSaheh4nCcsbw8zwCeyyoOXgd3cuqRY
eR7Txl8dKPGltMpqM9nnn8dmhqLeadxYRW1A5qJHcq6VcFIXjsZhYPh/2SY6ib8ouW+g+4lNVI4h
RZo9RmznLBSiIFDiNloeq6y83TL+kJw/Hgfmrf0rMXSMFylFULTbjHYOsk70W67gPpk9+Iz6Hx0S
uWTBnvb/REAcu3+7YNhWRDTRXEgyfQiVNNbxNU2gR4pBPIBqIPCPWRaDTOAQmp5DU5MgTFENr3Ne
i5gSPNn9C7NBU1qHhImAStV1o8L0yLfzqnXrvSe/r+1w69T03OXzH31VerrzUNsI4AhUcYm8XW6L
0gtg60gJmsd1TqxMCKx3wU6u4+z2Hg5nNM6ZoQ/h+jjxrO3G8uFJQp8jkWJCvL5HXwtGtV4B44ya
D+Q8WLzpdHHbcFWEOnlsITdKQaZHurk3GlaAgRDXxjAbKFLSZ5HLO8q+/2TVVc5FEIRO0nd0BwUL
62F9CMkSZUtzQrIRfHWQg8YsRDFA/hb7RmYNc7EJy8yqA/OpRBQEQG12yZ6gt6UqyNWISf/JH69M
ATvdm9LUVC0aPU/uAfjTZ7xKoIeglJ6LkCjzrW0HQJK+wNzAZpaWcQhCHviiLzJnvPg1bor+vhmP
foUro0VJ8PhYB99eZygg4pLgYUOu2eXFtnKkmVUK2u2W2WpS6Zft8mVrJ7F9OO50FxLvGbQYavKU
iVWuLsNFU5AQa8BCLVw0RvknvY3msSFB9Dti5nuwwh8alz82xi9SkJ0Jrr1xC4iUx/6tU6Jiq/Ep
liJ0OJPgeNbobVNP39TjXjrY+sax4Z6fD/Xqi0XdbuZb/PqU1uSGdQiAKMXXdHXT4h6Z2+8hQaLd
qf+uMZGFJrtmurwUdDjxuA3Qh0viwFfXT4v2hSeCISVpU8s8u6tBd24+cOdxLF3gfSEpoPXNqb6h
6vdUQfv8lfumw6DrP/VjwaEmrp7fBgTB8rY8olwKnNVBd9VifMDMBy8H0ctLHKKAF/ySxdf1/k+F
m4NuJZaNXORun94+q+uNrPaC+hL7MAMAtINvS2t+T21BER+URrsRI3FqaVK3xRX5QF27rLBxkxRN
j9f5goohZe/zs9WYNrOy9pp/QbqNdhHxiscFVIat63RNHR50w15wHNKaBJrOntawQ7R846l/UK0p
8THGZ66Ze8PJF4H6zfGpSXs2W1bOcNB3PwhzYhOedrIHriW8+2dsipSoXU1K90Denx1IW07sac+V
WK6Qhw4Df5GCJyiAYX+9cC+aoWqEZfR/UfXBNubwguH98IptodIdh64Zu5PZOgDIBvZ9ibZhBsQm
u+Rh/PxJg5kPq1DNvVc8J6/A7ou6varkNE0U8pk03uLma4bTap6vWmJWnewJjgf9OO0EopM1rDKl
/b2DyaPuZaMlxhbXVIgt2SF5gs7IR3dgPOAZwIdnjA65akwHQygiKHRIw+2p/n7cilQ2ABHPMGyx
9Mj7Z34cckqB+/WjE6F2ByAjPIkQcTNqnU/cOiSREgWjtbBmbly0AVpdxUDlpq98uVVKnXFvN+GO
Gx2zpVonmsKaiexPPPgHZeF8nLok9ltnLDcIN7JWYh33vlkPAOumZr2ZxqM08OSGRcrSQVcPw8Ql
yZA1kwSH5D+oUmWDj/HPE1iX447Qv+5Jdc03JoCPzlJaC1lWdezfy8azcj0iolVm4G7JotNLv9tW
JMEYkYaf25rgJZuCME1G09ThpOCP/cJ0XZWPVV1tlHRCbYaIqgXbGvnV9z2DefqtTBq6too4WFIE
rpxlR/ogoOEIBFGu+9OYgjSwSlUM3JaMxdQ9tUid72CflXG3S0of7V11JmH1FY2C/DKOP85dApFc
Xzw8DzuVyZI0Bo7nT/RZCHuzyixB0gJ121c/iJ0ea0uSge4lpGUZgc9TZ3FN6leIhNHualeTl+6P
Ilqjdgy1JuWJGxHTPVFisXhJ+wLgcv29k18l1UKxtQMLMCbvgt07LlK50+IsqL8BCw4wu74Asy8l
7V1IxH79C69LmH94fDjHZCHqwpXkqASRZeG4nfPebLKymqF7f4NlBx2VaMLtkR6nKrOrfMLdle1W
VhxUq7Pm/taiBESacy0IV20j4E3auwtlbb7EPh2QwG2ftxxUzLF2j3RGzP+hH1BRI7X9quQvLbZe
JBiIdN6gMmIpDwDjYX7La4FNDofxtUPaajHsmndNbG1DnMQ39CGBjts973XKJ9MKtv5XLelRQQ96
p/FeUKbmjh6bRbOfT5vc5wHjDd8vM6q5bpeqyvLPrOOSn2ztkhWUnM1bLlMvflYW/w+dU/2xEPGG
LiHKY22y9nvv1v9jvLEHsMS0ANk0jS7ogZjafwAAhuzFYVbNeKbr+gjqj/GEBT3x0xVtkxAlfXIh
ah/cR+RFSIZu/+i193Mwv09+ffTC32foMN651MeSATooAl/UQp1ZCtZkruu+cP1RYwB0TEVD3T8S
jMelzfeXCN0gkMP9L1S6DbdzlNp/ZLEgHda/GueYW+5KRfnpyhVV+NvrBAxfm+kWuaKENFARWSZo
EviODXypIZvfiuTfHcaCiycRNJias4rcVknj9rM4i7MBKynpjV0FVqsWaX08mc5+CI5Q+JOTAe+e
VSH/c4oqyMSwLt6I6vRx5gIbBuiO1BhlaImKX3b41FOZ6IEemK/10CYurIK6F3SoTC/54Rh3zRXs
UKzv+3F5DMnp6NroeIBJVdd3CPBTmSUMEQv/Cp4Wqeb+b3ge8XnpkE2avEGQDFC8UsnWKe82J5ux
OTgqgjK5eTm/pVW0HUp3U/RgighcGmFw3EaQ1HMzEjmg5A/UIPjHdk8tE9NQVVIfoJdx0URIZi/n
sMj9rTHMLPUZmbYpW9B2obF2+q/5M5dqYTWKLSEVUHj1PjV1oQmdUumf7huVtm0MJF5r1lXpeRBp
plXm0HnVqQhVoFv0Ym9T0/OL9va2DbMVaFOZqt/7TRtsH3BX85bY0/yx0K/oMOYTwo5UTUNN94K8
Q3VH2RNPNt/qT5mQtRvsJxUBQe9yHi21pHI2ZimfOIkLNCDQNpOn/LT7kLfpzzy0T/TFz9eYgBeC
DM4qg3tdmEBBc7LUFavulHPjM8ZPh3u2NqbVpPmKn8L5eAlltUOlT76qTJ6hxWJrXp2LFvFlMuQF
G1LZMvxxtXfM4wNXst5RyWKygJ/2Kky2k3vMzuwPloH4efEtLmhvvIMlsCS7ue49CJTvshHuXdo2
NdGaISe9kx+izlmdnp+4F4V9bkI2gXlK58+g/RbNSge/wiJHqScJBtMYSjcsT8aP2fHUbEHNhqa3
NpxrWR8iOAyYVCH/QGGy7lTkDZzT/LLpOr3W/KAgUgi03cRfPYzWXkaX8hzZPxfqDtV1oVJJooap
Wi7+afI4J497s6yW1JRChRmIc3yy9Ga1PA7zjjcdsBLUvGz+WzOe/dmO2Z337UR9ZlhReu8KxUwz
a0tPoBgw2v4lcYKZZSp7cYZ2puK/pwDTMmIuttG8Z14ULn4Yr2vrP+4vwr3eaN2f91Y8taazQNb2
xqI0q2QXo2U7jqJ3ZoNCyAQAECxpP78qxltf2T8x4bB/iF8TloTdj7b3w6E3liEvLztRL/iuM3Td
OrqsTKP9ILDluXK9TtZvwNZO0Z491gNalAgJ9FMmPEKDDFB+fshcXozvvfEBDHvG9b370hsBx59y
TiEbEK/9PklMH4U4+0Ku9LBE8H5pPQMTEqkTPC3Sn2utKJbM7nwv9tuknNJtc28WaDxCEePSE1w4
uxLzQs/b2XFIJ3poExvNbOHJGnfSbc0zMVilB6lUI6rzfr2eqATKnC2s0XGuKXibU9js8Q0b21Gy
CtmENpyBb/HN+uFbeMRCeLn0i8yS5i5UBNuW/SLgZblug1YDwawujDF2+WUOuaFnC/vj1YlJs4Ve
CPIPB8GUva9oopKn83Jq2bRX/Deyq07Fn3W3v/v5tV2BU8PwDbjxPktRlRY6PlF/SB9rBvmuvKYa
qTxbetgQOsMeFbZMyExvZbSFzFqHqWPEsoIw7+Zt8vTE8gHyJnaEX//oaJiAedyM4e/jiMGUY4UK
1i/NnL8sio8L3jrGyeukitlaRZ37ULST1gDvUCQOVhGtGJb/mkgOns2Vl639yT4eUPGdjjbTAnOi
ms+4w81o6gpg3Zkwsc2zjsVWjqYjKuj8yqBfCQe0+k4KZIa1NFBLnexLDcsxFxp76ReZpUfJmM7b
Qz3ImxST9Ygr+HCug9bUFSpK/woJ/FuCNi7Lnt1cyEtZ5pADL/d9zcp6V+TBLKkgirFfKt8hWxf0
sNlTpgUAX6TNHG4arqxdBq/6sZInVaOlEAc8vKdf/tqW2SHrnuP/3Ejwq0OsGhcLkGvBr3fkK+vS
Liuv2lw0LuKj81ctzDiFLMW/qpRPcwyVv8A4DAzTlp+DgdKRnrtoqBtLxN6oKpeOpvDsxMsxrN/C
4/PiUdlx/DuXxj/fCSnud4G63piABZyEmCmN1j79b9R3FOUVW602K2XzbV/WbvrPMnIICC7I2OFc
QL3f+mYNrikvF3FxuzZuI1fZttV8g+BPayRmJlDB8qvsS6GEPmkQCMoWqu9p/5HOqDYcfJHQarPd
Et+4jxhsjVME58Pw0wsUpTJFWnJKodveoWhK6kzC/P1ZVSiimAcxK2pvTOn7E/l1df0P4i1pR67h
LmkP02REh1ltcnnZbtMfhMRQxAbxs1i4qRE8ZeNcJpyNMMCc5jCKzcx4A2bXWxmio9MyPjXYr2P6
BoT2+7qNognul/gfnJthrGZNlr72+gXAWtqPUnK9sSuTa/X9iYJ23EzDiob3xDYUmzkB3NzQQ/DV
/me0kJ2FJCnCuQ5iuA3sHTdANrdPDlnJ+UPTdLBGMBPbzOVj1Y2KmRTtRzTPb9KmRxYsPtlYJ5dt
LJ/t0VIi0L7A8OWHpKNYBM6ReijwXNqkFk7WM1+DFUaePBDGjkaFNGoHGJVHshGG5wifbsaS59xh
zvTh6ljgD9iv7R7kXnjizC+w15B5Fbls3FQlb6Iu0pABsFPm7QOjoDy4NwC0gxh/xNUG1AwyRdJl
k28QINOV4V4MuOrYzRGX0yLMy2zVu6he5k12QYxKN2u+0eCy7ZjD0/Vw25rGzNPUGDclAgrEiWEB
l8YO54vwDrcdnj4yeqX7GtKxtU1YjElpGvBUxMuPmFyOHK2yLnSnSkzmBZHbdlgbZ0znlVhw6GOc
McVi1lHmJ7hVy8XWOLa0Cy2Cnn4fmHiCeVqiQsRrpmX9dMmvonl2544lA0fCECBu8FflnEbJUAHx
eB3XKu3WIfYH9yltA2eXHcr772mv29sByZJX6IQL72aHp+y8PZ+gnBGYLKEZHv+BoocIzBiI57Wo
Uqjin8UxlcE7fN7LpbKI+EZyuak71eNHQQ8ZOY5DrnoTY9St6bVBAKInclvo4c9B0/iLfX7+A1tX
aaCrJ28+La/neIClZg9hBKTAKVEOBIuEyGvS41filvSqVZCQJMJd3T04Sy/j0CTGrEKgzgn7m18V
813WWcW0WyNUSqtCoQffNUyiuYanJNhNrtdsWlJN5n/tgmicXJwKI/jLjZe+6UNInAObCNnn1fD+
4bHcvVA6My12y5ryEXVThiGvG0orYNIdCk3i1pb/hBTPKt6THlGBQFRFX37GRT95UHOruR5yrdCl
vG86UbPMng2UnRkvyrzQVKe8eMfBnCUtSTjuLoDxb5Yh5rkVrdo6wci2wzvGLYg4t2bDyR1fijtv
Dql8EZpyB/NjfY1IxeI/8CpctdiS3of+zykswhwDkmcVDf1F1HSnWNz4Rs9wPlEi2/dJT6HqTJ6F
v7H50pc7BTh7GgFYnYi5i9ZWUBa0+CdkiZtEnkgiD9CzuNdn9e+B0MsFEc3NFJMqtzy2s8aK9Rlw
8B35x5Wj2ZJwAhElx32ahQA5cUT+C0v8Fwe/md36vxUqsj+C8211XkB5kqL4Lu20aTVTJC42D0aN
4niZU43DjMVoqn+aHtIVWgWSw58zDyHhEFndI8w68pIMzjkP3z41iTVzdOPfL1Az8ArxPDWKQMij
Mjle43tU87dZ0qBf3sPgKuQHg0mwNQpLRpMp6UdfxTlB71PIV29jwh1Zx8Z+/IfUDPTffv3DeMV7
HBtRlbvZR7RMY9HsJMnu3ZRfL6JKzBJjc192bAeIAr7/ByuTbnZc48fdCFZZQ8ji9xG+yPS80/UR
3DuVfTk5rY8tq7V5hkWvCTVUkR/Likbn0LhrUf7xbw96sOt6V8vvOdbIdMj/1IDPkYY6oAbPW+gD
u0cgUCajJK4Z9ub9gG00JpFxpJ+aCKRfgB4djKeFIuKfRba1N957etG0lv/mFCGktvdjGpoNK4su
FgPbzJjStZq8XPZMd/cWhjIRPgINLAnVujWITdbkhOBa11RtH6Y2wLOx2CcvGWloKOuqOgpryzJX
kGKAK1WA8xJpAgLqIlEB2hUSu5fkfFEV5GDfDRyjY8hfydLGJ4IdPu4RuiJG9FnHUXN2OnGfukFq
SjsbbqojCVZyTvjFWJTvWk9rcfY9FI5DmWu0q3+TyB2cih9QkZxCrzwIRWVv0IF9GW/PFCfEMyix
3GlJPYYYhg/Y32IK4oK0aoGz/pbeaIY6fapxuomG0pH/LtK7Y/tqFmpnTcbhhyNaViHlaIkf4zK2
5Gdd1j+4EwKKm6ooZfho0Msh/doqUMvmurvDkHT0Ng8d15yDHUNz+2YHIuXzQmRFjtnCDFC7EXiw
ABBbQNfl26zpTgzORksmXXdfqnaLqxnAwvWauF8DIkzTvH73ZgxN2dHhgUg7XvXYPWMYSdRK25+Z
2jN/4BHktW/kJHQZOIxlD3QbyHEF4+prdA/a4T0YVyZyM+ubGSNRw/NZfryLt12PQYDHyl3UZxd0
ADU7Emv2zQ2LU8yh4BRPfYOJ+9vU1G5ZEjoUzbdLcFTh5/tkEyYd4VFS9qQYADGLgygtcPuZqw0P
PeiglUdeR6upHp0JsAY9UgUdxY6Kw6HdlBBI0VRznI8yNgfFzcSgzJlTEyhMUvxmbU7leyM501rX
UxF9YIr/AmZ6+UsOOdopNRaQTiItXx4EFvHCfyDs7a7LvO0gzBPorFQTInTbmiZ/UejmqPfIB+QK
mCrrTHFVShGk4VxXS0c/l/rRtFjcyVAxD8Yk6jL5m0k9oe8nYXqCWCEDIdq8LMLPaU92a6tS9D83
FbsVY5AS+ltte6yJcrnk/x9/GlqfpYJko/xCdlY9Urfn0TXx7Qv9sNzoe8tO3H8sRDIUNKHQSlj4
S7NMUhZOyVCz6cIVJZ+888+WFO975657x0rVoYAY+LS3HCxHp0R/gvcOMdPUKBNN4kIPf/rfYDCu
t4mcLjgigc39KJGLG7I8ef/M+ykBw5YGjZdEMIEm2ee46DuxkYgKjS2DKdqIZLLu6vd4lhlnkkEE
5KPdshXGn/J0hWesPQnKNX6BhaSJSyNX+FzVOAbxQUInO+Rmmb6at0xzp7KtEDX8MXHODopn38Ni
/8SOFnVmxk+SRDNH20bfc63XFn03dbnh8nkQ8vzNiUaj4TTlo11KLKr8qMVxIUsC7EHNlCb5B92I
dhPYeDUDcvzKAmj0eWAA/2kfg69o7JYWk516Nw39MVoWCZYhPc6sqr6HA34vhJUFivFreJZzT15m
cEc3EDBxFDQBkR+JejmZ8ZBtGqA/d6tRqAmLiv6PU8ccMPyAjMd11bCaLz3hU7LaRygzdSfCGb8z
pGLYlSHYAE1nNltzitlYti4PEkXHF7Uy7Wo3G/JCel9rXHkdkWGmHYQF9hPRKoUWvzWNKVzg9Yjr
TO282Evut0yTbdVmbsQkAKY8dk4Dai9OhhEpdYTiv+0jxa4gaJKRSqqzXUwAzkiqZ61KsNgQcAtO
RcQ9hSkpR4GyVx2A/1B8tXqAo/buWjxFxuNrKlT6J/c4rTRkKbZYfvMcOKjF470Eg72hKqo36zZf
Tr7WB5YRllqKocrja0/DM4kYUr5ntdaPmdmDXpBcY2IlwRajCG9/4uOVidMZ5F12INbVStZjLhCV
5XoR/Emk2vCg/Q3vwCpMOBHQSHHxUs0sWcAhs2JvPnVGy01ShtLlADTPdgwhGk9lffJm+JvSq0KL
EzWrjVkWk5kxRhAw82uLce9xFQmAydWPy+ve7AMMcPRs
`protect end_protected
