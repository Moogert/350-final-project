��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h���F�f��!1�+�0�,��?�>��1	���6-�$���.IH)���}^���p!�Z�S�'��8�7Tq��qT�d�f�����d�q�y�� ��Wz��6��b%} lt�'��IÒ�x��S4�ѓ��@�}zP���kf���(���§?,Wנ���AD&���ce�����m��l���av���wq 8q��淏�oL!����E�ˡ�S�;,�T<
����+h�8��Ѿ�:d�<B�DZ����1�eF{+O��;������Y:U�#�l�i�t}��V봋��#n�>��6��)���рȞ8�j��1]_�o�R�/�ߝ�Ӝv��F���	���7g�|��fcJ���j���jF��X�$��%���U8�$
w�{X��헺2\П�\;ܘ^|.Q��ʍ�3J@�4>����P)�*ګB�v}Ь��oNƲ7(����bxy�v2��ϖ��j6K��+�j�p�xb����瓃A���H��5�L�zPo��*�@����e�/����R?VQ��\�kb�S�Z�To����>�YkD�;r��sC��F�Ě�RG��/��eG����������?���#��9s\�N(�&�L��%_\��ѓ�����-�����6zr��B.Zȑ����a������� � 9��!?���rYsHA�k���򶱟�$V��J�8{�����4�D.�t���Q�nTBJ�\dh-���)c�RC.p�j5��`QhDM��l���+y��O�|��i'uqc+�(n��ݻ�/Y��U�U�
R�C�H�{_Q'�u�i�I�c�H��G������ĥP؇�Nk������.��r��qhꥥ�T֩����M��Y�ӟ�����W���I�e���R�F��*������`�|�y-����U�(�v"�>�ĭ���)"E�n5B�_s����<� �2�objc�$�x���y���,�DA���he�%�9��_�B/]����"����Ϻ�
��)5=e,�W�?x-Ƅf/���8f�(��߄n^_�.�u�Z��Ϯk�m�%�t���n�_���a�8�s�ty\L8�㬪�roa���^�?��Š2]�7̥�۝�VX�=(/W#�S���98�Bĝ��E�I_Ri���q�'ש �C�h*u�3�ϑ���7��h`3���+���F�t�$���8��-ݪ,�W��g<�;�.�)�;..�4��<��1/r�.��c���c	����>Y:;����L�X�����3a�j/<O�в���X �CK����`�����M��X��nd�Fʓ�M�	&��1�/bN�E�	�b��uKL���p(�N6��'qp�a�$�A4����Ʈ���:����;���0���n��5�B?�o�&�X�q�m�g��L��{����-!�!Aw-�7U�X�;I�F�1����g�nj�<P��[j�d��&��' S�f�L�v:Q�B�;���)ǧ<BJ�ut��C�Y�_�P��f/�f5.D9ɦLA:�cpYD������k�,����1;�S�ڼ6W�I����kŘ0�-��Xɑ6�����{�y�8�&F�7��-�9"�����5��Ϗh��0� �Qsքs1U�Q�*-�0M�Z.��C��1ӞT�۠*��f��.�n\�Xp��KH�@5ş3pn_|D�wG$��!�O�T�f6f%�z���p_n�I�,>�L�������(�UfF9{��ȉ���	q�>`A9o�u�Z�9թEsU[����f��6v�8u��a1�Ғ[�fi<�,�?S����%R��?T�R��a<��JW,W�eC=7�ίq��G`W��M0����Z��c�����F�^�m)n���	��5ǖ�#mO?g��|�b�0�Qs��S/�5���<4n�y�WRh�T��^���������O��~w^n�*�ʊ����θ� .��h*T��t�쯘��u.[�W����$r���y���A��翐HsyP_CR�Jra�/k�?���6�p���)�=��=?r��U��n�1Bc��X���F67ݑ�y�?�^v�lg'OT���O�4�bMk����FBorj�|�7j�R����U/��[�mC@����҆��<����DKN���^�yӷ�i~�^7h��$�ט|AI��]��0��woW�>�MN��݌;a*���p��x{�\���w]}@@��i�L�|�ko��'�:�)k�[2�f ����a&q��v�E
��w� M��e���!��4�쐿�W>L�����ed'�o�Nhx>�5��e#M]��r��*3�R�Z��V��̓����O,�I;rG��>�Z�����"��
�*�$(��]�J�H,`��V]'6�g��^����<��j{�F��htM�W�p�e��R�8Syu����y�	?a���a_J U��Xt��̴��7)ߴ`=�x*���W�r2�^�JA򠡩},���?됈����G�P�tg?p�g�/��a�M�A����+r��.ܯ;�!nh��W�Cv6��#��������9��a�~�M~�@p2��a0@�%}R-�^���\��P�]�&���-�@tJ����i	��g=�Η�K����� ���2}I�����V���^4zs�O\��Dud��1�EH;F���-��}g|���k�#$;����. �%�7[�/�4�[˖�����[U�z6���dT�o7�H�U�IΜIˋ>׼`�6#��g�+�����E��θ���+�z�(���1A�Ǘ��dɤ�f(�y�K���VZ�p�Ll�+	�+��e Ht�_s� ���0Qk f���e"_�8��0��p�1��V�h�pC� �#�+̣KR��ȶ�vT������$�}�b-XR�)�yg��(��wERͩ*������+�D�:2(�Пa�?�ar������	e�c�Cq��i��K+43o̥w��F4��ۅ��)�$����/c�u��];��1�Akb[����҆ۤ�1,n�S��?j<�6����Mo#�[R>��pK_�&v}u�+�T>G����aϒ��Z��6JsCv��8�ep���A��Q��֜���&z��y����,պ�,���roR+z���i���G�yo"����~���`Rm3�FGnP�=D8A�(��f0X��7ϕ��R�h{qL���jT��.T�TmY���}��U��� ��I�ZUj5��H�Zp�]�	�ڨ!��N���i�g JLR8H:���CTC��M(&0?w����gXn|�H_ʶ�W�z�լ�8���$�N��Sګ=Z�t�����(��ľ?��ѻY/�?��D:���ZI���~�*���G�3t{\|�-��z璝����w
FU����ć��U.3O1�Sht0�kg��eG���86��5�8��-ֽ��oB��AO�w���Č����W啼�ݤ^ղ}���kઇp<�E;$�ye8]��D�l>�iJ���0�jK��_[�B��������>/�p����P�ޑ��>�U((�TZ����:�kʒ=qA[)203Eeޠ "����>������+��9���6��j4���y�9�J��XL�Y�mZ��ޜ��h_-%>#dJ�e&��5���a����<�X��@�&Zn�W�`Cnc�TN�����2I[����
��T��Ɵ~���z��s3`$۞%N!��vɧ �����쯺i�\z�	���|"ffݾ|K�x�V� X�<�Lk��Am�^ q�ӹ0��^)ʀ�UL��N�8��ϿV�R�z�o�ʢ�VI�g�0��]ϛ" Q�#jՄ�``D���9i�3�&�QV�D��v9���`M�h���bW�G)��2�Y���W�&i�&*w�U`�1�������B�f�J!��ؗ�xvV��}�D�Ѕf�5]�v��r������w�i����k4�7��=��9�3hHH�8�Vut��⌬㛧28t,���-����W�69�pE��Th���T4�,s��D�7.:,��L����,=s7��H�J�:o��>��?�L���#�U�F�R7�e�-�t�h����d�x 7�P	}�ወ�H�P�^ڂ%
��%ǹv�T����6�7P�4�qk��F"��5鞘Q�@��seb���"�U52K�ȇ!���g�ծ�b�5.5���w(�9�J%FE����|=!���*�����&�L�}�-�?��o�$�X����8Xb��@�H\R��k��n*e�*�i�X��_�7�[��
���bς�K�݉�!��ÔO����`��>ܙ���E���߫sЗo,8��2'�SqrB\b�۬*��5�|�ܞ��*��ԣ+x�gi�U������}�v��
�����e-_{�xX�Zj����$lh�<�"ח�#ѳQ䗧���k�d�����9�Q�[�,/⴯X�- =��q�3?r��k������}��o�����-�~��kuN�3��sk]�w��w�(`�
��X~��ȵ# �o�r�ޖcS֯=[��D�2��w�o�n��ٰ\��i��*��n���q^T���}X(�	���S>V�!�t �ed
Ή�s}��ϳ��E�Eo�x��wEY��0�-�Z���*�Ⱁ�V��^��h�MP��kGyO��Za��D*�Y�4sR�R�3ʑ
��CS����v"
�l�ߌ�S]�%R��E�Y���\.�(¬����[�W�>���	�-�߼�R_�v�8�>�����3q=�V�O�z0�� ��5���c��l����ǒd@ދ�*�<Q����ɨ�����6�C7�3	��4������C���'��МLs��cO����.s����+	H��Lu�`:&ܝOz#�����؛7�K5�\5<�^�%��d6�`n=��+R�*`7����D5�>���Ͻ���qjE:������e��`ٍ��tFU5���e��O�5��vd�ݾ��Z��&��Cw���v��L��n����K�%-C��+@�#��?�m�s�� xF�Np�S����+�2	�!�g��jV�<H��������Fnx9�A������\��9�����Nh؀���@��C���e�R;�m�@�0�Q�(�Y�!Fe��&�5�|Rz��L����f��/	1\T_�a`������MC0��aBF-u�~v}�����Ӟ,��ύ{�����WR�Gz��o�t�<V���9��b?Uݗ�8.a���}-�c�uu�P}7{�������ӝ�jo��V^�G�Γ_
��Nę�V���@�<�z��	2"�K���J(�"r������]��E~���z���2v8TD��	o�"���']�P�	4o���� �b�Z�LxJ�d�c��#�c��S;e�-�5&��i�?-.}׌��z�}������w��7��S{*k�R�1�c���گ2D���0�g�J~Q���D7^�_P-�7�u�Z�������39}B��"���!&�r=U&H00���2@q���	�p
�O"Ef��>w�L`�3��h͎��nym�ulEL�{�&+AcG��>�Sh��}=�Nm����]E{$�K[�� %/�-�Wپ�xM���;�+�ͬ�%������=f�F���`Vh�e� ��i��D�5c���/kO�?��
��Y��@�6�{}��\�ε�h]؛܏F�ţT35���d|G���@Wٖ���;)��c�\JJ/�x�P����� ��*�B׫?7��(�ƛm.v��'��֌i�֊�õ�ā�-s����� 6	���
��GՁ����ƂE�=k��үA]0�uc�(�s@Զ�Ê���֛�_h�ᙷ�.��[����`�p�ais{4�vԾw9{օQ���1�:kU��3���H���u��<��a�ۣ�1�}��#Ѿ��Z�e2��C��= �����n`�)�WL�f ��8��+f���zxF��\��W���ٖb�]��Mx~���zZ���u��7�S!���}�NFM��xt��k]5x{���C"x��D����1��G�ͨP�?�1��L �ʝ0���+�wR��&�=�C��ᷲ�6�R�qgc��n]vZx{-OX[��K�^ߧfL����.9�����b���%�,-��#�8�X�R�i_һ�tV=ǁ�1�6�zą���^l/���������o������uֹ�IG�0�!�x;�������%�=���Z��o@e��YUUo6���؁���κ�dg����6���>�C�.��{ͧST��
���|6hv�.~Oy���t��f9�	�9�Đ�EK�D3�g�*
8cԐ���gA@C1�l,~�r̓��q�I*T�wYie��(Bn׉���	��á+k+4�gG�j��9��!�P1��H���x�2��R_��-rVL]��Wh	�����be�)���U7ۜU�_��>���g�;-����d �6Ze7���]x�F�`2�6�FUأK"qC�܃|�-r��r��l�GFo�OwN�5D���ԓU1 1p���Ë-��\�¶�o�w��C�����
_H�y��hǂ��"h��iPL8P	~-�ć�Q�G�sBS���.���{I�=�� ��^}	��W�AT��fv?�q)mQɘ�jMZgM��`�Db�8���~���d��e�Gqh�8Y��Ψ��y3hL���9n��ˢ�:n~�{��o�<�%�v�M
�A|��&A�Py�/fzXN�6*�%��q��ŷ&�p'����L���̰U��W`����:\��]hx�C������Îd2�����ޖo�(@�x��D�����D���	j~(��{�X�X���'lbX�Φ�jxG�c��"����jJE�z�֥z��\�+0�2�`F�C��~]�P�nӒ�ek����8y[D��|��0���%?[�n;��'4��m>>@mb�\���F+�j:L]_��}[%7����^�TP���>@�L𪲔@	Î`�J7�zڈ	m1HI�~a��K|.Đ!�3rB�)t�	v��K!� �jq����E��7T�p�v�*½�V�%{��לm�eM�v�W��)v-t��W��w��P�7��šZ�6^�Q���8ݜ��e'@ĤF\�7��-�)�J��R$k��%r��3S�}�'}j�/1�x���2Gw�n�5�P���DG'�&FrOT��.&�Ba�J�&Q�+?u���8]�H���k�ufWe��b붢!�K��@��8�QЛ���kN��3�)>3�(!(Jo�}��<��1ƘѶ#�����p�r��T�o�3ƨ������B4��b���dD����3�����	��aVߞ���<j���EI-otIm0�l��=��@��Y�榈�b\L�q�����Y��X)?q�^*<��m���� ���2��Su5I���\�(��ͣ$�I&$�+,��h8�:B
�+e�(���z+�2�q�{9�:E�AF~��b�O����G���&}��
n� Ԭ��V~i�b��ц�L�4�ي��?���B0��"���w,%.�ʂL����
�{2	Iք��F��c*.{��lZ*��KMm��"=H���3LW�䶴������WZ.�7��rP��F��.� ��-��W�V�U&�+��UD����Y��F�sY�j/���7�8PV@�u�g󆭎6�S���P�o{��B��a��/��'��ZY3(�(8_��*��P�����I�[�C�
�+vl�6t���($Ҙ��(i�|�LwX���F�uiw���/<m9�)�]�����}�S�@��j��-}P��G�K�O)ce��Og>U����\���A��&�O�c>�hv1O��l_��)v�8J�t82|�L��K��J㡍�CX�Gw,ԡ�ܵC��R\����� z]ޙ`�E���'[��؊�?0�uhKq|�?X�v��fC>R����?��ɦ;I�+���vt#����̠�3�4Ѧid0��痭��7����gY]!�f&�75P�~��}a����0g
͎��B#T)"�l�~��b	�Hk]�;�h���J�X��T6�g�����LU�m�}2ؑ�ɇ6�ڒ7Vg�a���x=�M�s������5s�z��;y]�c�j�IaM�,9?��'05"�eo3F�м9l'�d�(�љ���ރ?�ɟx	��R�\�fٓ2�D ?	��Ňb6�-�j���?��,��Y��0i�N�%���*uT��o�!�Q;�)ĉy(ޗ.[����*%/F#ȭݿY�L��>x,C�M�KZ�l!�����_ʼs�ԁF��{���E�0}V�q�~e]���?�b'�C��D�[yB��'�4X� A�?�n�s.��3���F'#|�P���Zg���KAb� 2%�u'�H	��F���1�a��~�b���ܹ�o�	�'#��#A��u�(&o%�� K�w ^���V�4+��%�-/�g$\�����eٶ���y0EӤ�w V�%㛯��ƟD��~��䔘��h�8?&mV�G&�.9ȕ&	��c�N�߅��&��W�i�m�������b
��~�l�$��m=���L ]RNy."��o�! �ݨ���H�Q������Bi�7��P��y��?�!K�"�IЙDdO����w2�'��YpL`�tM�t?X	�r�����eﵔ���I�r+ �G�,�P%�=�K��{�Cߗ�A��E�)�P\X��`�[u�R��i�$��ܟUP�m=�������y@��YyS�FC��J�q4��N�v2��˫w�t�0ԜK�&2��Ң�c�^��1�P��x��l��=�^B��|k��&4�� r3N��5d���Y�6&�J�E�έ���a�e|�M~��e��kX1�E���Mp��C[r*'�pm۲N疩���%3����ń�*�o�p��퉂�ҩ败6ls�Ͻ}n�Og�{:S�u5<S���NJ���-5X9�J�a$s��X�:���m�`�����((Df�Gf�Al!����5��b_��+��КP������v;_�{^&�������sz����D�ϲ���u-�(�3��S�!"�����M��'s><-����hl�A��<`O�+��W�l���w��$�.o�dϸ�:m�Iӊ������dt&#���4_F B��}Ȇ������xY|}�eL"�4�';D�o�li"���E�M!e<(�$.wn��Dݻe� v���ph���Fq�EA�
��V��A� :X��8K��Po�xnxT���q�a��e3j&�~9�c�<��Gԛr�)q&+�_�I5��k痬BnJx��`CT����O�X5ǡ�MKc�����B/b�_�6�{�zp]�E�yk�v2?R��k�kjR�S�-{(�0~�aD�[���r�*��e�Vh絸���n�y,�Bwx��E���m��&(�����z%�hp~�,���~�G��5�IZS>)t�ojcXZ�s\���'|��1~��d��֜�%f<������������0,R�T�!b��-���e���D l{�fn�}V���$u�0:/U׿��u��Fp?nX��z�Ǆ��$G��zf߸Q����3�䔅R�5s�?[\���~�g�{���̧�6`��K�r�EH�}�j�d��j��PG� -zP�-9T���ޖ��Ѯ��xn�#��3���r������@�����2!��?�	�g�.���d��;���Vu��^�f����S���O�T�.�Ժ9Xpaz����C��N���&���QjO���q�t`�%��/N���mH,��XI9��7@�r�4# H���j'�g/�&mH����ȯ���Hf���=�u�_�i>Y�Y�w��H����ӛ�!*x� �f�/	���	*7����6J6�s��������:��#�犊�;v��l�H�#�3�V\�/���Qf��C�=�c�#lOJ��rо���0�g���*�%%��"����;3��;6}�Y�[�>��/����X2����,���9�9q��PNT�]l��q�|�j_�S�0�'�x�����;���D�7[�U��T�����$���'<��5q�����}��~��h�B0�{/��l�y�`�ʾ�$��#�����/�w܋�0���U4$������l�8g��91�*HZg�}�2g�3�� j!�Q�U�%��R�+&z��W���z8(-����'�j���`@�q�����P�*:����	+g��UH����-H���$�;��Ӄ+^������S��1c��İ��Ғ���A�@t�A�Ѹu�X�o�6&�������ğ<Dj3)�
"�����!��*�8�~��Uf�R�{1� ��ٍ[>?�ZڵwǟJ[jyZ��۹�Zj�<Y��>?Jr���f�)�܏�J>���߬�B�Ҥ�k�k.r�,xs�U�Uk�ol�N�A�ˍ���O=���������2���fM���ｓ���J<jp�-��Æ3D�uG'�&����B�?U�I#�IO�E�e5�]]�b��Q����?�W�3%���~�Rӭ��@{��
��$�ѼD�>ᶻ�o��ɸ��~�3���}��3��*.:�{��Zs�CD��j����6��4»��c�0�P��c�Wj1��󋹭L�܊g�끏��*ȃ@(#D�T�P^�&2lQ�.���ج��;桡�v��x?A���?�G�#}Q�!�؂�����Rn��	���a�z�"����Nq\뢞� ^Ғ�٨��OL=U?a�M��S#��&�:�{��+}.���'Xb!�-�� �c�S�y�o�ϊ�%�l�"���_05��pĬ�+ �ɜ��e�2�p�z�s�p�^�D�g�A�Lϟ�����.�[����e\��Ɗ�GD��"�aV ���[HFߔ�rMئ�ʙ�z��x��6�4_�Z��1s���E�ZvX��|�z�'u�L�x<$��&8M�O	� x�$��:�\~�f\K2��#��uL�~J)W
��fQ좷�����1̖{W�IH)9�>5F>m��w����DH=�� �KQ����]��5�j�Nv޸�6�$������=�џ�H/�+��Y��ufO P_�YM\�^�L)�'a-	�ܴ��w_�2�Z@V�oP,_5�[��P�ݺ�|�=X�H	_5p=� m��;(f�|i\��!�q��Ƴ #~��5��n��nu�\D`f1�.�Uz�!���^�����I��0>glb}WTD -���B�7�k�~�f�����\~=_(/B����N&�����I�L����6���޲ft�fM<�hH]�� ����HcЙI�TF>��F�;H^݅+����r��:uA�%-&$3DԙK�H{m8D�陈K��y�T���Fo��`�R�(3��}�XS�iG'�ޯI���p���B_�>J.u�[>�.�D���z&�8�'���ÿ��62/���F];zq�!d�D�jA��[Wsop��;�(�>[���H3�忙	|P�xE���+��:�U�W�V�"͟'6Y ��xյ'��I�q&��uJ�������}5~�0n�Ӷ�[�-,s%c�8��� !w��"�fk�k��?�4��B2> Z밀P��p��H�K��9)����I<��~lUo���s�r,Oqё���V5����}`>���s � #.�MK^���&�]L�{� z��HT<���� a��Y�����
A1X�n���h�������N��W
ȑ_�s�"���* Ywt�����p�X�/���;��������V���-��&������"�=k����d���� ��7�/;9��Q�� /��jDcU?�|�s�4!�}��>�������΁� ��5
��B�U�cS'li�κ_�N�&bh�Y�����S�$8���˛�_hU-������^��h!B��P�%�]�f�2 � (󪲨 ]�D(n�77�fS��Lа�.�*Xоl�`/{W	��YJ��T|�JYR��riz˂~:���0�v�m�7�P�~y٭(v�g/��|�����DP/|�\�${���Yd���\"7!�8�Ė��3VX�F�y ��n��]-&�U\孮�&&qX�*�`�lY*�7v΅o�����)a|ﳍ���<��"��������]����`ר���_�[�k�����`1U������̽����QCѠ;Y�URS>ۚn�}��N��WrWW�(I���q�'-�;z�BE��3�%�A��">4L�R?���;~����0Q�����k�k��� �^v5����]��	��:����}��̠�~��\Q���&�Z�A�� SA����i���0�u��f��VOO�i�1?�H�p7_Ĕf��J��j8�K��=�����;N�?�^]Q({���?���勒�`�}��$H�|2c���j ��v���:�
d[�;��Is���M
���!SWn>�� �r�t��t�����g��BR&���11N� ��*�l1����NCՙ5:�&z/W���m*yj�����0n|['8��t	�ei�t^�P1�-hF�!�����p5U��^�xz���m�V��nu����O��@�0=�K)�l��D;D�t�8Ԉ���22I���0c=2�\D$�d.��Ț۳{0�K�A̈́|�$�%ɩ���k��|A�!|�ߩI����0��*��Ş���Em Ö���4`(q�T>Ң|c�My�U��w4�a��k�Kf;�8��m}�%t����\#���y��m�ҁ�
 ��_��m��ًW
&�Ã����ŭws�*�o�����Mv'G'��&@U�m�K���A/�#�#�]�"1m[��~�P���UߍX���՛�W�@	S�$8�X'���x�����6p͙7��LP��Tܣ��<�K�*�V�7r��Bt�HK��O��W>nM�l��l�����a҈$%��OaZm;Cd����W���s%������繮��
:�G�E"B����&FӨY�#_)M������b�aH�Y�v��<����h�8��%�1�p�Z88���N*u@�e�@��x���ը���Ng�p�mP��oD:u�kݺ�2o����)�|V'�^gq�g���S�(XP�yӴ�X�ު�.�+����
!W���W$]�4j�K�j'v׾񭢧�o�h�MoJ�;!Rݎy��E2���C����o�ocp����c�OU�j>Y\�M��^���qUI{jL1q����	���m-1��������J��i�Q�~�C��~M��3$�L�[��.��ƕ;N
�㻿���,ɡD	�rz喇�>No@B�2"7<�҈X���c�umVƃ���G$o:��I���M�4��]Γr��laO��#S6�Hn.^���l~o��"m�a�.�ft^�2U���/Ap_6�a!���H����Kʀ-�8�u�?���[[,خ�tئv$���<��	���9\b'T��E��!p��xD
m��N��~iB��+M��M�ow��o��WJ����<fw�gE�\�7�P��k�����˺�S|\"��d�!#��J������u�f�ц��ʧ��m�pF@��Y��^d�kr�*�HaE��]�n�F�C�mp�T@%[��1zﬕ��'F�:5>�x�V�e�Ѝ ���jw��1LƄ�p�����D��k}D�)/C�,�_ ژ��xv����I�5�m�88�Y�Q0o&_&���c�qn
����M!�	�l�Љl�*����.+���1_��O�=��3�a���T��q���V�xL��J���`]?�SU#$_~��P#A%FR���������n�Tm�W�-ob`��]��@�Jr՟�ÅI�$mzݵG�?:EJ ��07�RM��@�������N��/u�Hg�hߘ�1�O����t�2�,O��2姘��U0&����%�/s���q�a=���_O�����R����KO�J�>R�����_r�Ꝣj͚�/�d��N9-օ���,�dO� �2NĪ��	1Cq��D�m��)�&8E�Ա������&�G��H/���V��ОbW��Ǹ:$/}��\%�e'�8y��+�Z�חdMa.��Uc$�Y/���R�kYD�ꏊ���CWhJ�I�
FM���~;El�0��I����kw'�ߟϢ9����;3���0��b�����2YRQʹW6Z�.��� �0�,olG�ڏ,VJ�]�����V��f"�?,��P���fA���F��ۭ�t���V�NoN�3;��R�L9����[�E�м9Vtc�ƢW.tS��+��9�q���1�[[x�g?1���3�"a� �����dR��p�T�5�4�Ʌ'T)`�FL�G��R	A�̹�XvW�+�iz�7��?1�@���+�����I��6g������|ݣy��`b��)�S|&_���6��G�Ӝdb�=#!Q�,;a��?�8C��tAG��&.Uc��)$vy�I���9��*��]z����8[�Њ�dp�So���Sۢ��"�xUW*�
�<��HR��(<��^��c��gz{�˞�,F�ў�b�^��I���P a��]����g�<��4Y�(�
䄩	U�Ɵ�ܿ4g��y���'�Y�ㅰ	U�'�2F�q��,*q#�/Y�[Rf>����1Z�$~=�N.>�K|$���K6���U��g����t��V)�l�4^�vi0�S���!�:���vК��0�u�Z���W�7���܎k�kؑ(�����9��G�JS��k��iO�5�X,q:>h	�b{�#8o�$��O�O�K�މ�%�D-4�����b����'�n�C\��Y\��&9E�{D!&���#-A�8��i��E4{�S:�{]._�����L,�Ƒ�����0#�T;,љwj��.�pD�-إ4�b�5�u=s_l�j�~���s� ��%17j|>�m�O�:�Q����xJn��j�ꅯgr �k��������9F�`��\xٹB�G.��X#;���#��7���r���I�¶|H���@w"�ɧc�϶�:����3�w�1�yk�q~�FV-á�l[=!�,.s��\�{X+&?��N@�g������
���`��zcu�E���l45|-���T�V�(�z0%jr	(D?],������ؽ�P���W��w��"׀�v�Y�搿f�|��Em�~<%�	����s¼��{����t����42^�������3V�>�/�9���sǐ
8q��8T�G#�B���R����Jn��ה���'m��&1�3ٵ8{�^7V�2Ĵ9h�K��P�4[|0H���!�������M��4��*On�N�)��B��^��`��إ5\�&NQ��^�.�
-�����b�JƊ$���V��E�'���/�9���=`�`��-��I[as�>YPs�i6���βѩ��%�+[��^t-d9ڨ'b��+���t��L������ ԝ�B���ʘϱ��nj���V)Pm�䪺?���H�I�i sɞ�������7��:O�AK����y��(�^�p�}����IIX��?4,�ϲd@�*�4.��c������`E�����b��9 h�N1�U�n5�\z��R�=�666���M���ն��w�jTqY��~��$C�`d�5�t;���tq�,`�Q�o���y�;�' �&���G��	��U�{�X��0k�m�g�7�*VLm��KɇT�kj�n����9m,
��'�'�m�Õ���&s���z	�4<&t���l�	|x�h��!���!kE�ˉ�tSNM ��P������%m�L�~�d�4G��zbr��D��0��Ŵ��	����5�1��>��/@���T:�D�$��d6�	���I�r�XS_�URUc��L�­k������8��$��	J�J"$�2� ;�����F^���¹�uodo�X�ot��k� ���N˂��$�ɣ��ƍ��/~��)k�'',o"g�*O]x���Gcn�ʐ�2�K�.��qU�+����bv_�e*�1��d�Wu[�A��1;���ۻU�w�j��#s��W}�@��ꅌ̩>��K?�b��xQ��|�l�t�����e����'���F�h(������:��J��� �Y��{���v	�X�Zd�=�SH��P�Cp�-v�)T��ߴ��z�J>��C�g>�BR	K�!NS��7L
?=���H�*���M��ݖ__(�_-�b��O*u-�K,�Bz[���l�,��5�L�����_�O��P�%��/���v���tojva�&@��G�A�yU���R	ժ�ye񟿴%s�F;��2{�N�Wn���T�vZĤཎP���֬�&�Qh��~���U,��?��T�T1�Э�Ӊg�i�!�ٓ<�#����7�yB*��HXr�⒓�P����:�8����]�5#A\{5�N_�����w�"T�r�O�����,4Hr�A����ϡ���947��6>3��zG�����;S�?���8ѻY��
�&�-��U��'��:���v*��f&�?�l吊��)r�9l,)F�x&JI�5�V)Jb�XX,��e?��4m����F��d&~�]����jZ�R�	3�4vm�YV��S�wa��\��H����5����z=�t�����Tw�g��`���vH����9�����n���>:��P�����gg�;'Ȧ-���h(4KN�A����ٯ�!���Q��y��wr�MP�6&����Yᨳ���Uį2��jc�Y��wzjy{�h�[=��� ��m)�f�#R [��.Ay"�ظ�,�<d��R�\����H�~n��5a��>�і�*Z��]��ǭZ��5���̽JiU� Z��/6��A�����Z�rV(zԭ�>3���,��HB�,�X����q��	��#W]?�|�/C�e��a��\!����?\�f'/}|c)���1��/Pw-�5�T��@��nmg#�|������z�@n�(��R�┅`�%�S^$�tl��$vR�Gd�CO?C�	䓄��C��K�|[�ɽ+8�ӹc�mJ���g6g>^����pa ��@��ytB�/��""�z���Q�'��������ׂ����p�-L&��܎��gY�?[f�+i��a�Rh�b����z%9ޓ�c,T�}�C2L��?K�8��'��z�����<~C-�ܻu2�8nZ�Q*	�ya=|�B�J�ԫ�{�^��I6��BT	��:����.��w�U��j^� �&5��%
�;>ӏ[
��gTҖ�d�X�x`�_��ح�m�\U0����Q?yB��p�9@�Th�j��J�c�-ά!�mɜJ�d���3Tl�a|��Č+D$5��	�t�Ѩ����-Ӝ1�>���@yG�����(+�έ�x(�=�L�h�Yy��̓�O9z&U��lF��
NS]��{�ے �`��?m�7�􏀲K"r�l4 
{,�ڵ�����9A�%��v�py��[��2�,������?C�KLrVᨶ !���d�K���π|
z�
 ��^eicE�z5H=#cZ��>i|���nVR�W`��q���m��"G�|�lb)f�U���@]m���$��O����5	q�����5���Q�2$7�dT�섮��mG��Z��3���K�:ChY�	����|�ZHю�8��C �3��B��~ǹ����.d��Lm���]�J�J�D��@C��S4��y}�E��t�)x�(��i�%m�=���I�{���0�+>V|CZK�}'� �g�w����f���0ISy����j<RB�O6�j�>��Oos���)P(7�y���Nw\Ij�Z�Op�������"o�|_�7B�zt�?����D���x����td+9�s����&>�_!nCt�sH�1��^Ћk�ⷐx�P1������e2.w��iG{�S����;ѽI2�+�H�;_�$c3�ڇ��\�y�37O2᫭8�)��7=x��Jq���L��]6� �~c|0��FU!�;�Q�,Z�Ң��N�������#������D{r#�]r�.�.P1Fz���%��N�j7��Yμ��&m��}��yR5y�fE����5��~��A!ֶ����K�$��u�y^Ø�>�J���|� ��S{
�����&��k��/�{>�`��
���GU�%������Y��O���0�i���	�=T��Q��Pu�=�T�A�dk��0�-�2�w\���"[P��x}� �UdhH�*}A�W��.ؓ�p���{��)�KH�k�����wȸsٲW�P��F�hCKP�.���Υ�%ܘ�"�;l�}��_R�Ϯ���N��*�t~�� ҷʐ��Oe���qܹV���K[Ώ��JB�\OJ��:&�"\��bmkG��[���o���AQ���n��s4�T����������X�����Ѥd=[uV�JW5V}DjF�U�!_fA@+p	j�^���N	`���#�kF�f�%5YE)�\�D֍r����ѐM!�$��� ��Q ���wD'(W�糰�݉�������X�7�R��_'ɀ�a�<@bϵ��`l:
/'�r�>�e��=ľ��ZSY��A�~4;*�h~�����>�?bb�)H	�
��Z(��@L�^��P�Q��%YrOs~ǐ?���m�k���uA]�-0Q�{��h%�xu!*�߼�ZM^0��yCj�l�O��^�[����8�h�v>�XS�ǺI8=��K!h�,��M�Z7��)���h�0���Ӄwg�T�]�J��0Rr����Ed}�M����t>R�[���#�w�Հ��㥣]�g����z�PHg�q؏��3�I[VƄ㄂�X����m<a�1q�IF���Δ,N[q�@�X��@\��['b�FWq�fE&���S�M8�hv|�/+K�2m+%�NO��1�g���;f$h�0��tX%�yu@kb1y�]r۩&�f����w�=`?10��ׄ*�H�T������#�������`?ZP����f��t�"�&]��/E�2�x����$w�Q󾘤F��#�_zC��1:�s�Q�&�Ň�>"T�z�C3�.[�0��X��4�� �b��J��ٿ��ɢݎ� ���I�!�c�%�y�g�t星10y�A9��e�� ÿ�⹷����}� 	�����/f󴿛_U�l��!�J�n�� \G��NNt1�Y�c�Ez�C����'lMK��@%3n�%�yH�l��e��DE�i	0�{L4�S�5x�|�7�گ��U�����,ǥ���G`
�rG�ު~]�V��ЏKi�.�7ļ���p%�7�>�1��UB�Sp��>���t����Н����Pڹ���@�6JP�k\�����!r&IH%r��Y�J�]���
�N
�~��/�����B��vw/�/�ꊶ�a�'0fI�MFؾ
:|��w-��֐<�s!�ꑯI���U��m�A���Jn�揭x�V�yE%�?�.���*�/m��A�6�te^*�g �=ݤrb[��O�2� �+�m�3�e����#���ͷ| 6p�� �����R�*�{D�Ai���r�g���0M�Q�_��&���:Mek�"�#�J�:�����L��j\u	������nI%�l�.e�8�uc���^���|^�EͼR�n���VFg:�
ѯ�M��a�� ��ԥӉ`f����p�����呅� �0S����Ä.E�".�5��?V�K�Y�ġ�VC�b��_�����+d�52l]^*�x�dhe1 �ζw~C��o٥�P_06x��zrq�E`?^C�oRV��4���$�qS�A��Ss�ER6՛��zJ���|��t�b���@��$c����Ѩ��%�:�����j{�CN�9}5����:��V'f�'I�����@�sQz�����]b�a;�۴Ln'[�;Ў�1���*a4��ڧ���ՂT��?9JW��mTŶԧF	+i>	ZKk���9[�8��4��q`���f�� ���.f�,����/,�@�$ �N=TP۴ܿ�l��'�{���]����(�hXNg,n�Xn�S��
�B���y��>��f:�s������P"M�*�W+OV?�)
���Vv�P��	e���%�j�D<�;���y�pD�"ğ���SۨH�Po���v�;etrױ����U�11�q����k_��_-��a &Wm��d��'�X�*T.��
oH�q�D��+�M8�P86��)�pEXa�+8���tb�NC{���r�/(��(e�y���5
����"�|_9��1\k/\�I����
UoF6>s���))^��c�h�  ��P?9��LIg��c���ÿ'��Ck~�ޓV�u���Q{+-]���X�3e��Nnj�~�C�6i�.�N����Ә����IY��@jF[���0�6[֩6hJ[ ;&�$l�Â23o�B�֯����	�s&����V��Ǻ�hڲ���%�@�#�j����34�4mӹv��!�M ������c�N(v�'jb�[��-�ڞ	�:��"���O�:N�L���s1s,���w1�{MJ�Ke�n����Ԩel���[�(�o8�o� ���mF��"�#.�|L��;�$>����`����@�t�K��s�������}�.���:�;�n�¤h�(�(CnRX+�+銶�H�a�O����|�!�ws�����bcC"�f�@��>�ѱ'yg8`�:��e6���}��g���O� ��Q���e���v!i|���0T����G��+F�D�QH�)~���g�?z�H���c�0�ѧ�&�j��ۛ܏����F��� ���n�=�7��_߹P�J+�k(d����~!ay�������̍�q�hl��f��9�9��Ps�.�H3
ԫ�)��ic��N2t����st2,nLOF�?��u�Ι&��z�_u���GI�i4��O�ݴ��{��^��H8>#1�e�����fM��A�Y���L8������U%���|j���]~��˜�^�ݛg�	s0��6 ��/�H�h���g/O[��J�S��XJ9��v)~R��E�#��P�)
%FA�z�����'���>��O@>��i���D����c���|%"�V5��R�fg��7[-Is�R��$׍\��
��s��.��2!�e��}=�Џ����+���{�gL,�yRq��+ڑ�-$4�o�$bMa1e�����t�9��U����0�U
|ˑg[Aw�e�V�ల��Hw��;96s���|ŗ�i4�2l�pσ�i�ܺ�=(�n=�a��Z6��!m�gWI�(;�WYw��v(�A2wa0�,ק�!hJ4	
�	�����Ɵ��v��U#P�&rЭ��E�{��j3yp���=��ǟ��6)�n.������[p��{����_�Pl�2�9"����ݜ�]�G�p�����l�IVb�����rA-F8)���O��<�CG��aXl 􁂀%*��\�� %4x!�pJ�a���w�G��j�!��:�1�|AXwJ]d���sj���G��{�8��8�C���0�_��e9]ҥ�n�fX��R����Uk���%�r�l�����$k�5ӷ��)�8Ju~��5�[w5�/����<&'�� ׻U6��A$G	���ot��;D�"UضS�+����I<v��}�Ծ�@��@p��b�Y���N�cA�m�����s���9�:ʌ��!�Zr�N�����G�$��DN��D��;J�ViL9m$���}��1���N���a鮌��6&	MC����,-���]ImAĎ�k�m�Z���萫:8�)	90B��W=���I)7�NFo�Sv`
�߄��:@L]���� ��"�*�Ќ�II�-a#�`œ��7��]]uܑ��L �)����{�yU�P�>�WRVݳ���~�o����9_���	*�>��X�C�~�<ݱпG}�u�/�I�ђ�l�!�'��X�|��.!H#5/��L��cc�%����xl72k�z�8ʪ{�G�&�Mo��
��q����QC1�l�m#
/w�Q�ĉ,y��d�Z�w]<sX�j��7�PK����$���FG�
���������~?E&�㉦�=3N����զ�'m���3uZ��rI��D�����W�-ݶ��}�0 ��B\ך+��
6�����i��F,����V =MX�}|2�$��*�L�e�)ܽH'��π/k�m��1Qٮd��C������6��\�������\��?s���  `4�w���P�,�K�p���h_O悺ǥl��z�C��Q�:&\$��f8a�g�J��1p���t�0�5 ���$b�/X�LY��϶(���Ą�6)lJ�ʪ�E�Xh.�hjvu��Ba!�}?&c��I�h�$y$�?�����U�-+��I�e��FB508C=����{17hO��=hF��p�)����ʄh7��
M�#"]Fa�R�����E�8��	��~�G� ��� ^�3X�� Ij�g���23��M��fC����i�ӭ6]�Z+m�}4\��]���łL���3x�w��3ZT�����?�y�G��W�Ln�C���c�L&�l�N��Q����+��*�k��*��)gω{����Ȗ�嶨�@M�_�"A+x<ǆ�(�E�P�l/�<|������ �
�6_���!.*��Ǹ�%�H�o�Y�K,������Qv�`�0�)fzx�(��a���g�z�����g���H�����S�a���͠��c��Y@;:��ӟ\�̮��C��\��x=��*� ΐ�5Ā������.p�&���,�YD<p�֨�ݗ$��K�vYQ��:KJ���sҙ��w�@�"��O�Vyu����s�/��+�i���*�/�������?bR'+T tJ0ܑ	t�����������O����E(�(�G��:HPvfì������J�J���,�R����<�V�LF��F5�����o�����A��TD�h{����V�b�C�~M'n���ol�2�FG9���3`�\�K�!���T��M�Ze�%A�;��U�]����g3��uńu.��*T�*�1��(X�)G��8�w�"��� ��ݤm

� S��0o����z4O��hN<Ȝ��gj��)�½K��Q'�G���� ����6�pe���(�n-�Ci2��o�z�3:�Tц��r������NR�������)j���,�y(�z��훌ak���u2dx�a���ܨ򭾡!�>�;���W�o��н��!Ĕ�Řm���n�t��8�u[�U�|@ĺ9�Gq�1?�Hȯ�Kt
a"�H����H�F��Q����'y�.��~�*�(s;�@lҾ��k-;b�^q�?�����Eo�8����g�f>� �2	v��1�A�ظ|&q�MF�8������B�h�7���L_%�����}����=V/�*���82��(6�c}��Gj<�Y�f�呣x�(9/�i�k�L�>'�R�E�j�҃Q1�:Lk���<��$�	`^-�D(n��(�g��/��������?��'<kGO@��e��0�҇t�]�w����>Me4���fQH�'!��!r3e�|��nL�._%���pDa�ֺ
u듔I��{�������s�{d�]XQ�:IP[)\U&�R`3*tɏ	�n��/w��&��ε��� �
[�Bnr�5�;n�����_��rO�s��Xz������@� ���뮁A�j)�	���g0N\���	���x��C/��͋?8��j���~�R�b�jBo�Z�K8�c��k��y��`!�,%�H��s�ע*�7�s��\�^�����������{�䰙 մ4c�r���s�۩w�L�4�Qt.{ ��<H9�I�${��FP�N��f0��4kw}�(�iR�4���t 	�M$�k� O�;1���w`6!��˾��ђ�k���ص��oU�+(B��P��E>��t���3kT�{N��y���X���ㅚ(� +��*��HP��քTL"���]�Y�wrR�q*"e�%�RV���JY��Pyg��.vn
>k�l��y��[z��6��������#�F::���� ��P��z/Y��tv	O��Z쵘Z�I�M�(}���c0���8��|��r-����Zp%U��ܪT6�yY(p|d#BJ�:T�3e�9�Q Y�{�Ƹ+X`�8'��0o��I~��������V<�{%�F� �u`��l�S헻��=��J���Ia�&c��E������9��������ۈ�{��[��nD`H;�\o$��9�t�	wx�L1��QQ��L���͓cHBTJ����m�$X�N������8I{� �Қ���O$i�r��"]yfz�����BFJ�\� /r�xq���pO(Wx�x"լtv1K,��_&˗��P��:��U`�-~H����KI�@7���%x�}���+@�EJ�Pr�-�E{���S�y$ �I�Q����m�`_��-_�)Cz{3��ٟ|�@�?�Z̽|>9�dz����ęNf+��ml�8M��$"�2��5�iD�wۺ\����%�d|�|p��ۀ~p�kPMT��4[N_nn�q+u���'[�0qB��ƐV�y�XĦ��Y���b[�w�e08�߬�2Z��DZ-��B�����-L9�\�F�\Cl�f�K�ѣ1Y���z��U7H=-�\u,s+�D��ɽ�Ƹ'TDC�|]�s�9��u@�?��r� VX7��S��纊���%��n�xds�;.�ٶI?
��\h�cU�jeY�����7���K^��舩x���P<^��9E��!���.�悳UzP��#t��bl\����u8����+\ˑL��<�ϲ�~��te�۔ʊ�E��q�5��9�����bj=8{��З�I=���U��X]C��s�`���i^�;�lŇmU�[��.xKlG��h�JP	L✥ ���,)9���Y��>��*T�)�G<�7�Py�T�v��qm&�}&�$�O'������C��U��¹2�!V�o�����ݗ���,��#.5cH�Û%����w��p��UQy�L%	GO?��|�a;��a�����W�fш�A�W�	��;��c�Ɍk��Ŕ֋*���M�gXۤU@!�#�F����X��qߞ��M�ɢ��Zt"����33�Lg�8�U�b�m�A���[HI��0�0���f8�j�
l���<
/o�(l%�z��'�2�8�A���*���1N&�-Ǝ(nL���vtwʕ<�� �s
y�~�.K���,�p�k�M��-�� uwerϋꫧ��n��BhP�6+U�\Q,@����i��~~�V�p%���j<��Ңk:�Z��$�r0ֶ�,|6:���
i�)tЂ
ΩCX<F�9�x���a�&r��+��fNP�v����-�L���P?	 �2w��l u��qqI)�QX4�*G���h�A��k�&�Hvmk�����Z�!�=(��'C�=�N%[)(�Oc�-�S5���h�E����?J��fO���
f���S��Ic2G�J����U��VS��
���h��͒}f�;
��5 �Zz�JSY��m\9R��� 5\U
Ls�W�LLt��P�cHcD�9���}߱shdܸ]�g7��ƴ*��=�?;��h���_�f�K���D�VƿP���/�U�"�<E��yu!g��#�Q�&�1�8>I�b��AhnyI�b]���V�Ǹ
�I0F1����VP	x�;�|� N�c�m�n����g_�/�e ԅ�Ͼ�#u�8I�9�鵷WÁ0r���C��۝�j͖$�W�O�˧�V]����A�'�@[ǝT"�����G���PDzk�r@�1�a[z�l=$İ*��e�K�>"h����D����oQ�V�??9t�c^B�ԩ�b�������ں��`��?v�{?���������*_ǻ����Nd�ow�B����ɭ<��ڙP%�'����~jt@	�xDfUQ0����Q��4e�+Ԕy^Ld�.�of$!D�KU���j_7�pr}��!�f�ˆ��H����V�Oowf,-�U~I
N>&vB�O�@P�zX�K��V���_����vP����~���&pܑf^�Ee����L�"5�@�I駎��M
A������pF��VF׷ܣ��U�Ľ�ƹ�,ڶ'��C:e}�!n����b�r����2�m�2Q�*���o)3������6��#VA��~c� n�[F{�)؆={0֯ߏT�Gٔ��'Cz�^�y��`�`�͵�����7��_���`��m��~Ї�|g#�|�>q�IF�h�zk�����A��~��ˬ,��q�<!��e7rQ+4B��%��R�tO�M��_�/Cv ,$N�I�b(Ӝ\�p����2��)��2�JBF6��PE������RO�$S`����a�2d�_��O.���~{� ����l���6�t�jVx;U����f��H��{ɴw�u��e��˅hG��=�A[5�N�����hM'�������\�(�Zo�"e@�?{�4���T~z��SO-I�=�����),�������j�����iuk��"�C��ܭv�ma4�n��a.��ۻ��,�rٻZ��t��cP(W��-2��zWpd��O$�8zv���.��ǘv�\ԡ�L��"��X�>8���2d�y�YC��Y�y.C�v�u���A����r�O�q�L2�VG���_S$�2t��lì�\��µd�J���Avd@]��TG;:R�!˽k�PUf��e���=3�Hv�jiL�,��M�.'���S�:8�J�A����~�1�}y�N3C�]�~�l�/�j�t�S��OG�AC:���W�<<*��AR��Vۃ�O
�ӟٱ��/��J섟��/*�a�6Ël|��e���?�^�@����%v1
����}����^�u6�ڀ<,���6�D���b�?A+�6y�5}L|�r�9sti��F���M�W�lz$	�������5���ͻ:�ϑ��XfݯRF'_u���/�/��g?����]#�/d��>���,��+�g�d������fu� r���qo?F�Ӭ��ii��d�m������	{SXC�h���HM�UZ���R)%�%�x35[矕�k�wF�%|UsE,����6?1&v�ɕ�$�^�ñB����'�"Ϩ'rݷ'�"��Y�ȡ���|���0�~.�yR|�$G�	w�O;�{a���x{]��<�fr�7Z�-����!.�ouL�*w>�Ԣc��s����<;'��>�в���E�>�%n�1�?v�E��O�n���q��J�B�r����0��l�M��Ť���?���+F���2�����$b��h��ǽ����~XauA��
�#%s=�SN�%g�:-���&�B��|ZPA2���B��4�8V�����9�� O��(;S��LZ���/C�\�9�0(+��m�v������a�D�U��k�_ص?�"[������,�Fi�ˬ�.�Q9���Z+�ds��)�3�_�`�֙f�0�N����W���$��r�5i:�I�m_�.`~���R�6��	'��������-�?�"�D�Kp�A�En�7rX�y��ö�-��E*9f3L�C��vģQ;c���g�[����YaiT�c�`�q%k:�w4)�a��i˘�����]��,z��_%:�L�#TU���_�g��,��G����<�a��	:!ǉ˱�d�g�W��qH��%d*qt�'=�}�$�=4N2N��ǸVw��?� B�����+d]�N7b���j�a�ݪ��\��k[��o���tih9���T�&\&��7	q�f�^����o9�_�%��g.��\��?l:�s�
]���\0�c9R{�J?m��ު�%�,�9���DQS&�D�+h��pj��%)�ꄦ�%�T]�	U��I��(VĜ�@$��b��Z �-�!�I��pغ��8T����l���lP�m} Me�02����6����z����J��BL#�|�uf�� ��b����W��qb{	��Cj�b^�]�[�i��0��	r��<�5)�dV�����U��إ��~#���	_���<�����ϳf�zc��v4�����#�|��??�m%���股�WmLƚ��5�G�.�5��nNhx*b���+�k�f��w�v,!�I�"�x9g�Y��~�>������W�o8�ͼ������F�/rNRwN���s �wI���&!��� �a ,_
��^����4R@M]��ənIr*ח�0!�I?�TH��	�1�W5&�[��L�ʕ%�fS5��6~��,����bI��ִ7j�#�ͰPSq������1N� �ŝ6qʀ�Ǹ�Q��}{*U��c>��K��#ξ1�3�~hP�e5y"����*^�q�3�t�,����-'�� Jۀ3�Ǡ/���Bz"=�v���n+�{B�aj��:9֖0�8+���	zc�i�z6��"�ӳ�B8oV�x�qEsՊ�g�����J�Nu`�����ə	\��*̓A�XcRf�����ۮo�G��.���!�F�h�.��� '\_��*�-���7�T�G3Aq���D�w��.��ÍD�+$�Q��r:k��ρk[?�&�*����'����8�a/� n��Y43��t�
�CI����� O��l�ĵUg5��.r����ԯ�^�{!�T(�0iB^.C�Q��G�L���Cw_�߈���|�ў�.'��5>mLr�G���`��=T$��
"A��\S���0���XHC0H��2�݇$��8t��Tc�/�L]�ÎOo
|�������*|�ȃ���B�t[�)Z��� �㦻֎Z��H�Vc&�K=�WR�|+�O8<�S#�$�KF�i�����P��#9�a6����*��^��S3,��Ր��[t�K��8�4�@�bN�Qq�0�m�����/�
�eKj����P��2>��>1}�ubB��V���G��m�5L@�w�)k��%�e3#	~���#������0��>o�<t�b;+������/�8hW$���"]��s�����L��F'|W�F��W�F����.G�c��z���3��C�1��d�}�`��ŉ�����78������Δ.�sT�{@R�bq�ɨ�[)��߻K��Ƅ}S�� S�0��7������*Ğ��5��]Dm���pw=l?�L�����w���M�ȟ�=��C�<KL��R����,�h�T]�RЅ��t6u���>Myؗ�a����̻X���"[��è}6����TȖ�;ؽ��A�Q�	���9���Q6I�)8����p�:�}�s�M��p�]�/l9d���2��I2��7���5�@��d���j/�JLu!��sW��p8�/�?^��K8�L��DJ5E��
��S���b?k�oXꩡ~vr����Μ_�L@7�Z�ߘнl&��z[�i�	��q�'�.�/Fgs��Ӟ��Ň4�#����dIZK
{mbH�'���UM�86�KE���&�dX��Y��XS���:Y�����7�3c�@x���r��(-�8�qqd�V.�9^g`����Q#��@P���\�~D� �vsሹ�9��b:��*X�`�֏�k�����%��goù�� ��q@<��N���K���L��|�c��o]�{�j`��?d��B`^LP2�!N���w{��Q�Ж�/Ŵ8I�Q�w�A�]<m��7��َ=.������J>�\��_�L�䘝������O@�/��P�\~)��f�2�yz��q��)y����@�j�xȡ���E���K.O��*�떣ȕ]r�9}���772'���|���V��{�&�o_2�)b��S�+tzjN�㏺�-l�Jig�M����Ն�@oz��4$#��b�z$�X ��� �Y����-A�a#�����:vf͉��ըS�G%y+���Z_n񃞛⋱Y@�ľW�N�4C0c`P�%.�g�:vL��uوc�z^e�6P"٠G��o:�����V�%�rW��ZfO�LYTi膢�1G����Jk��b��ͪ��zO�N�/�����rD��f�]�chL��x8w���%y����۹�Lb�y��ع1�GH��z����Sw���0Xh����`C̣K�AR�y;=T7<�{�ۿ�k�D�O�kt��Ir̔n�'78n�Z~�F��}u��kH B���L2�c.a�^�z�82���LTǟ�q<S�<��u�C�.[���9����E�&�ͷO1�m�Mm9 ��f<7h�%Pluij��\�v�`j�	Q�e�bי�b���᤟��l� Cc�\�|��r&؅�j�N�\��t������6����-f��2F������& �pN�X�?Dt�1B�u���Ŏ�Q3[�W���c��h�;�q �r��L�pt�������è��G]-���h��	!� �u]Z�商�$	X(>	�.c<�ϔk�Q
�殫����xDg�N�-ٻ"L���g(w�:�!�Ȋ�$���5�"h�v����Y>� �uFg(� Ǆ���O%=��*6�Ea)�)X:�J��zۈE4Yp��+����L*ۙ�v��R��$��sS!1��B"�����M�f����E$O�żgoQʞc�(�(�`�Owvqd�M.n����v����_�_dn����r�Sc(ò��.��+I�'n�z�����:q����_����/�=��"l�~HY'���7?k���e�7ԉ�#@ �sg/�"�<xy1z!D1�(?n�i��`�L�Z�T�Vp��h��F�T^R�0Yݲ��3���Vp��#�6ژ�߯T���x`)qo �`6�*�@�����9��<�*V�u��Zk���sĹ�~z����W%ǅ���gmy���?Sa��� �����`�d�
^h
P���Y�ټ���IiV�C�!��9��e��TNWE ���~�(;U��mY�� �w�U0�yՑ�t�M|d�5��<22���Rr��-f:`G�ԧg�&"�"���'=�̒���&��d�V�_���vV?�tu�=�����(�z�G�˗��I��=�/��0"���l�7X C-�f#\��ڡ�i��0}�tF�ψ(J.e�*��x�'�*����Q��@������J*��"Yg2������k�\vKl�]����.������o���Y�w'��C�f�QAC&t��$��iլ��) +���Pq�z�jB��������gd�x"�&S�"���C��VɈR�3�j+kS�CO�*[���,�ޏ�P��<y��ēܟnm��Z"�IA�̍9]S4<'(���l���=z3��D�-��_��!`>0�NP�P/�C����{)U̾g y�4�< �����!?���Toxcfe�B��e��!�y�Ĭ�,
RZ'�MMl�� ��U&t�<�([���]MP#)�ˡ��o��f�Ȉn�!��xѲ*����$+���p��~�L�(���̎�����̋��hK�f���;���99T��p�|\�Y��O�"<�
�`��$�EB�'; ��:Y:��޸ E�tD"c����}<���:`��-�$%' �����霡U|��Qu�|2dc����	�w�h�hM�b-�NI{�����>4��I)eRl؉D�A��m�/X潌���ߕ�y���{�A��8VNM����-�w����b@��K��P�F��2��q=!����6����_����ZQ{��n�6�~-���0�d��e�v���oK�_W�Μ�B�u�č�謁E�j�ѳq
���܅I����p`�9��RGTz��q���JX���Ʊ�������,p�D;8�u�n&ٹ�|�4�J�&b�l��� Q�:	STϻ����3�}�r	���	���/xc�0�O�'�G�������//�W*���Iֆ��z�RU
�s�X*�_I}�DܜJd�x��Y���s���ם���,S&�۪�v�!�2�"�PU��rs�����ݸi���X����֒k�u�"� �[#�*��ܴu�rn���0Zv*�i���!	���Yqީ�R�;E6���o�K�$�!C[eu.1�^�?z5�Z���Q�n�~�̠qV��C���z�.p�%X�ڌɎ%@��etS�H�-�Pr�
#��AۢY�M�r��~y�0~yw��q��QJ/8#M� RU�W	E��X E;lt'ε�r�W�s�J�>�ڤ�<K�[�3�y>bԞӃc5p�Ib���ߖ&���]}�L)�|�� ��Β��Җ�s���u0�0�E_�\�Q�	1���
�օ�O	�<�ǍA���Ӆ^j�����0��ʣ�lY����8�tKb��vE��]"�C�tyLEk�H(G����?T�0�����U>�=i1B�@Z�,�q�!;@&���ao��
U�EZb��0ϰ��xM�y��QO��<űx��9�����ӯ��es�R/�Rv��JU� � ���b�q�?��{�#Q�#Uy�h���1��_{[��v�e�|��ڡ7��%���,�<ZV��H�V�Y?=��<[����_�p{~�é��2�{V�l�aN-j���|o��W�H�e�J��7<Rh�k��RR��|6�� �c;l�M�Ay���Yh?���z�L�u��%'�ݖ�� u8��-��7������m����=g��r�ϯ�}yeL��Չ���M�J�U4�x�g��:OI�ͱm�d`�-KVl%���4�y��T�=vh�<��j��¨�����|ތ�@����XD�:{��[�6�^����xܚ��o9G�����7�U��=���I�C�@�����V���/

d3|;���������c_ͽ�$Q" �;�c���Q��D|%�8��Y,��s��C�� <}MF4Ő�[|�^��6��S6�{5�]��ۛZ�%���wL��Zi�\���EH-�:FtQ`�@"�	�d�DK��b���[�̱�"��� �3I�]70`�{��MB�e?�����g
��WLs�u<��E��~�7%�ɥj%f��w}4�֞�酙�y���?�9���j|���m�L$�#>މ�R/��ÊSlQ ����Az��Z�+��y2DW�af��!�،d"�Y7mK[��ß���r�pJ�!�O�խ!u�	N���h"�*��<44����U��&�q�&[�O������Zt�ܰ;=D��&Fw���C���ڔ�q�O�i<-\��<j���j	��pG|�g��0\��/�8>�R,����~ego�/�l�������e��	�"���đP6��X���G�s�Wx�;���*�;�U������N�"�֑�"\-���蕝&��lC"�D�}t�=c��E��O2EϪ�MJ0t/�i�������^A;P����7Tt	�U
?�ש���7���@��&8w��/K/���g��o��Z�& �@-��zQ
�n6����.*D�l�Ú
��y�ٮr	;�X$3ŖQ�P�z�㰖>컣)�������z(,���k߷2���c��
�"�=�e��*^GbcH�/����=}E��O�1Q������b��%9�W �<�ꮫq>E���1��G�@k��{#&�k�Qs�p���2�#s�����i�ᶷ\G�j�`Ne�v;	o-�I�?��[������8���j  [� mc��=�t�掅��_�s��V乴v:�~&�����������3.4�\����C�ҁV��6��P2�~� 'e?����
�3=Rcb� �Ȭ��M��I���>%� �~�y���%�}��	�@{�UR�7�W��E'�|�C�I>Uu�?Ɏ�1NW�KG\�ۼ:M�h�W�ٴd��hut��+jE��iyJ��_ܾ:6d^fvm!N�9�y��Z6�(#�1�r-�	�Z�ZYV�P29dݟ���H�[����Ͳ����$��j��s帻��>�HY9��	���H�z��H{�-5�> K����Xg�EVs/�[̿�1���P0t�:�1K��/��왊 
�f|�����ؔ�#�Auyp�r��u���"A���G���]�S�;(���|���G�Tζ渂��	��T���:��}�0�	�y�	@EBO����|3RKԵb݃��)%�ᄥ�R��L@��g���O{��ܠ�"�� �͆�A9	�J�u<���dq���zF8|�'j�;w�`,��=���;�C]Ք�]���Tд,y���	b�Z�� ���<R���3�=��ċ?��4���o�8�P�r��*�lkX<J^����;�x�ٽ�k�U5qf!�)���X��e� �R)�j�w�o�@C�s����d|�H�.��ءj���!����*�W4�|��K��m��0l�r�8�q��<�]��Ob�R�eo���ռ��J1~��5��c�f����n=Ч����NisoK�	����0Z5�?7|t�hE����1r�ͧ��|@Msԭs��ʒ��1v1I(���bB���|�eo��{F�r���tR��$ˏ��J��C�υף��E7!���~��>��av]Zݱ�_�rZ!|��_t ��ݺ�&hb��,^�,�j"�}��Mޏ�&�P�n�U���앸G��@G�A��({vǡi�!L�0d�
�MM�v<����9�D/J3��Q�]�
c~��i�@�7�j=�Z}�(]:�&�����:��,�d7����e�L�'3�D�Κ��DuleD��w��>U�<�F�fT��|�٦�8�-�F-w("��H�ǆ�q�J�W��e�B3u��zix�2��í���"o�*v���xL���xI��M�p�e�!�Z�<(nJ���"j�R��n΂=ؿ�Ʊ�� 0��OnU��
�#��z-�I�U=�G�OK�E�m>$�i���$_Ge�}m�Ǚ��	T'��-z4J�e�<�g6���+�**�Q.4������c�+J�8E"�gӆ��N��Kc�TA_�Q!���^�t0kv�V��T����&2a�'Ͷ����x��Í_�H�#�Lh�҈�ji5�g{�0�<0���"������}�m5L�,j��n ��$���߉��-_�0싪�-�쮥r۹r�>:�A4���2���.3Gȴ��M���`�����U�e����	�_j�W�lG��D-F�<��)�_�MR��,�#wL�X��d�z?w�e�M�ND�+��?D�՜�0x��C�[����\�����b��=�w�S�`���S��gk���Ҡ]Q�D��1�����?�O��շ��|���ϜZ�?�Thط���P3{fk�r�QC��@�OѢ��g��;�] Kk��F�J	�����w��ė�_���O�>apW�VCJ_�J����>F��V���-L�{�tk	+��ՉZ;�M��ܒ[��=m���DfD�D�A���]�q�M���E�&��R���/�Pn�`���u=V�~��ܕ��pV���� 7��8KP��誟,�2i�M�ϫ#�����z��Jl��H�U���~A�{���x�*<�%�5���+�Ż�:��h13��Щ��t0V"���@���18,�Ƣ��z�����b>*��|��FJ#���<������O�8�Q�d5���8�Ҹ	�/�=>�d�p�pe�6�xT۔B_Uz�H7~�q�.�(��֝�یnhN*��U��3�2����}h�N,�)0|��˟���c�g�F>�ƠR?B�
�f�E���Ԟ/�wpi��6/]���G�rT`�R^�N7�6_�.�Q�j�g3p�"n����r��������H����d��~�'u��/0pZ�F�+������/Yu�Z���V���.�&<[ՂbQ�X�ș��0l �o��m�P���i������әq������"�ò��S(?�ag�m�E�:\�-��Smb�v�5Q*��~��`!�$�LZq+���{"���C�H<spԦ~o�s�E�^y���U�neߠMLRv�/Fn��$��ސ �����E�f�	�V�g^�|�䁋{�`��.����̪�������F�L���_p�*f���:I۩������E��c�^���vkTۗ�䴣���Tud��U�γ�Bn�0�gW����l����V%�$�B��V�x �"=����7�Jׇ�-x���)�놘h2	�%�கk���)3�yBI>�@+���:6�/���R�D%�@����~7���L�3\`�� �[�ַX���Gc)��q�?\n^�	,�g�6�K�G��f�Jl�k�P��<4�������#�.cY���Ec4i��3��ro�z��K40�X�,�̴H��b�7�	h��T�D�fPp���	�|U�6Ls�����k�x A��h��Uv^j� �]��kr.�ǺR[�\hK!��Rv{����po�7���S�kw�d=�C5�Q�	��T����:�s�إ�M�������O>�U�:�@�x=���Rȁ�a�He�B�2���@����yh�z����"������fO�ZCt
Q8�C�Z�iй�L+�B`d�/;�N͂o;�]2{��SI�fhfX���8�3w]t���Z�ը])Q�_F�����RɊ���{�8�qȮ>D�"NPٌ��,_�WQ%h�a�����7ư�D�� ǎ�p��54&+�>�dG������%���%�k9�h���ЃW��cH'�����#P�C���Y�&��x����}Idi�Ynx
hc6�o����P��NW��{���ߙDΐ+����QX:Q�6�V�,g@�q������F�/��A�7��s��V3�8ʱۇ��S��1�W"���z� �� ���'�a�H��獷��i��|���E�\.{WmL{����x�J�T���t��f�x3�s���<ȱ�DA�E��£���D���ർ�4�TU�;�]8=����&B�,�D(�_?'��,!�M$����� F
����󀄦�L�y9���#C>�a+>��ʒ�U��]ڒZ�bX������5�-c�|�����k��� ]�n���r1�9&E/����b�wu������cU�@�jD�<Lxkq�~�h�$fk9�?.{Z�?���7O0O�J�Α����-��`$���}��b��m�͢���Gؤ��̑G���$Y�i�l��۶�S�d;!���V�B;=IͶDl$��x$Ɂ�p�$S�T16gaaI�0��hfU��t�o����/�%�����S�ۃ������1�o��^;��_Wj<Z��(r G�%j��ĵ���V��W�u1Ӧ�m�����}�t�lŷ_�7��^��jjX���D@"Y,��T�il�r�.  �D�R'�d�ױ	�4�k4����k�2$ޱçvN���F'�e|�|��,�u��ͳ	��9��*;�9�� �	����w``p���h���4��!��`���q����՚w�ָ�6^;rl�#Iz��s�)���|ڊ;�Q-8�س��fs(ך-)(��L�4�3�o��]C�C��g���L P3������g�ӽ��',�3�9 |M��4;�>��Vk���?�`�F=�:�5�iU^���C ���ޒ $�U��헾)6`sY�s:6A����D�����%\��H��SUdn����	�k�ռ,|lç��a=��/��1�����&5	l�ξ9}��c�k������|�33O���ͤ1G�d�z<�&_��)���0�ݝ2Vc�
`p�`��V<�R^o�/n}�,\�oӍ���u�+]$b���n��G�U���p�����.�(�v�E'�5q+B(%7}���*)�}a٣�hc�"�B�U&��BM/���Ƃ�����`�1��m_�ݵ	J]Md�<��z��1��Nu��	ccwlB�!yŅ�mF��G�h�e�y@IL�ݩ���ΘϔFR��Ig�%E�
��u�� F��
��6�>��)�J ���O�^�<�۰=�o�X��W�~L�QX0]�o6���Lu��Jã�h~�r�+!���I�ׄ6ڱĈk�����O��SN�IS6΁z�
$����$�0He�^��9��Ҩ���j'�/ښ�cYT��@��-}�țG�8�8P����"!m�u���3!n�������썗nv��j�;}C{ތ�k���+��km%�,}����H�*Y��{��u�c�ouē	I/$�߶ߍ��֘�E�"�Re���#G!�<��i�=K���&�jR	a��Y+��}�U��i�Y�r��	v�EӼ!g `�1���P�os�)���qd鳮����-�_B�w����N9�]�����h�sh6�.�'�i��1?�|�l�,�b�DC|�o�M�d�@!}�䪅��%��`�^H��r���F�8�N	D��N����̊=�M�A���99�qd�~>d�r��c�x�ޙod�l�B��\톴��:�0Ġ.�����������7��@�@~~���Ǌ���Ny���5e���CT���F�� 7�l!8G;�%H�݄lfM��T��Ȫ�S���w���1��G/p8޳F
�~��YI[q��%)%W]��,PB/5��통�[K����(���x�_�'\��I���,��)\�;(�&��6����	�#��*���!�(@��v����W�;��Y ���V�WA��5��߂7�_O}�Qs�&x� VH\©��y�'~���G������6��׼�n��x�b�<�C��J��%$���#��w/�/2j�%�h�c{�J+<�'���tk�ڐ"#���h��w���T�P�ԆYO��?u�L�kV�"�=/rfp����'/y�pA���_u�O9�K�KuA;�Kɪ�t�Qĵ���S�J�΂Hz͋uf�f��M�"#w��:����_��������X/P`>��.������i�Vb���!�F$h���J���o5���^����x����ȍ���G�7�m�J^HE�x~�X�1t�:�;ص?�`X>�qg�.Xԉ	L����O�6��*���H��$�:�=0�T�񁸛+��Y�"����C�5z|�+Ƙ�XQ������a=�4���Y�ޙ��d����XH����p�J�s��B������My�!�U�:9m0G�b}�s(RJnv/���[�r9���9{ұ�������Cs��^���w�<�T��r@��jRW�èzS��YB��Dh><�z�%i,	c����HGDq�x#�gꆳ4=�>�r��Ճ7�����opm�EZWlVr��]��!��n(¬,�
Yl����W��`�>�v[]����êeعS�;4J���h0E8I�9D�:e8O��֒|6�/�C����Q�&�v��Z�  zX|`]b�37��d"t�F1g�}ʛC���٬�����(�I�#ϽO�ң}�"$J�׷��w8!O���Vc�m~�s�gD7!E��O`CA�9��!@�5D��O̕}�R�1]�$�����y;�Ee~@��x���m�'&��>��Sp �9暞򘃋~.��ш2ó��E'��씈�Wg�W2P�����Nkڙ�Y�`��a�l��vp���堡�L
�LWXIF�L�4�f�*ݭ<��*޼bր��m��~��(z����
�Ҵ�ci�J.���ϰ��'��϶���3G�֗���n�K�gH�孲Q�D�Y�WVZ�Fq������<�1�999�R��V��Ħ�u4T����xg�#��+�XW��u���$rk��h;A<��^�\!ǅ���K���c��������u��ZX6�5?�Nr+�w�g1��_.�]3��Y�ujV��%�����Zߒ��.����/N#1�xz	xVK���|m��nvB����p^�oL��^�c5O��Zn�7���@���T͜8�'�?��HQ�^���`��8°�%V\CS	��Ur���:D~���ĥҢ�r�\��ovmb�L*YtS��"G6U���8����!�Yl�ꐠ#�>��?��T�0s9�08~Q��rC>��{�E�pRN7t�<E*Sw��A�[�]ê�d�����TW�l���VC�5���K�_W&1���T�ЪQ���5�E��g2%������]�� P�I�uW|��9�N��f�^���΄�p����j�4�֠�M��/�8��O�tm�N��W�3D�N��]�����w�*n�2Yg-��❈���%���8p
H6���Pn����X�~��('�kVJ�¼�KMj���4%<���5�b4H"���P������؄^�E5Yq�_Zi\�P|��"��b+����;�^�l��o�)�O�&��>���⼸�`7O{[���)_c�F�����S`���@����& �
� n!СЇ΃�.�$�Ȑ�]5Fy-Vr!���'�(� �'��a��!iJ��'QՒ����{���{	��,4��Ls���d�Rn�爌Ã��ć�k��QD���0@(��*i�ZC�"$oE�I㉳��|˫�@�R�i2�2��A^� ւ<��
W���Ϙ���P �~�W��e6��<{np+�3����ͭ���BTRt��/�8�ߖ]~��ucSiG�t}v.��s/=E�ҵB.�
>w:�iZf��ɹ�Z�ܔyj+oQ�'��X���Ӱ��ڤ[�;�a�Jʃ�5Px��"w��0^��ʹú�o�>�a�p��T�\'mc/,���`Ӧ���[��]$���9Hie[	~gڲ��O��P��uc�TW!]O�8��d{�3��{s3k�����)�?��ȚE�8��K�s9�Jq��e;g�_����uй��P^���������&@ֹW�������tI��K� ]���H��I� :�n�-G%S�i�b���[�����
~�� �}���>U���j�J��쪖U�B���7���������^ pA���Z/��zg�:�?��@�0���ׇ�'X�%���.5��SnL�@���TLX�a@�{Bp����z�L�cH�(Ulw��~0�ʹ�RXh�1�BI�#ţ��߹w�}�$�e�c�A��yf�X���2Bՠ��$��9U3=�|D;y�+ '̫ZD�䮀m�o�=5(FvЉR�ty#m�,c7��&�=�8)�������"j/����C׎�\�l�e����`pE}���{�ICѥ�+�:�����&��)�}j�X_+�-0�S�E���7��PK�B]����@�c��ђ����)W�����|4qG�k�'��v�p��]��m�o�O�c�9H�FD,���cꅡ�~_�-����AS0��>?Z(,�^�%���X2Q��c<�Q���ǖz��Ee�$�d���֋Tύ }\�uI���?�i��Fg��gY}L�s�E9��釱��Km�yW?�d����8J;Fs�A��G�L�i���b>{���[U'�Dy�m���Jl����JxU |"�ǐjBw��|�^{	�H�4p����^���M���7���@���y5�"R=p^��
xU��o�t��0��)l��"���ףm!�'�/�yv��H�ߚ��߬��E�#���xF '7�O$6��Q���k���#���C:�.��`��;&�L�^8�|=�pH��\��`%}�����i�6��J����i4��ٲH&���wL����=^o��^�(���1:��x�e����Z
Y~Pn`�.�s�~\}�`*I�˺������t��I��. ��wE`�04��?u]%IV������1η�:��㉜s����*�2Q�|jb =)ɩ)�4 �H����h��I�E��g̟z!Z���p��BE�l�>�<>)�1&�K�7P�{n��g�UԶ�g�Hۯa0s�4e��\���i�ʭu˷�6�_Б��^���Kz�i��C�ȅ��e1�����o������׎��5�$���mľ�t�G����*���S-T�3�9dW�ݔ:��&��ř�ʂV��'i*s~�r��a�a��$���~�h�$ioR����4R���7� {�	@��h�Y�.��f������&W�1z��b1�'�!�rD�r�q�u���ۉ/�2B���4��#�?H^�}�a=�����ۘ@S֑�<X. �.#��D�Y6�L���6�[1$F�v���O+=րJ�Hs�u!%��{�l[ ��];��N���Tr�+��C�͟�.�%qJb��ռ=�aB�L!���CUcD5���Y�j�kE��6a��"�xT&���H)�-��t��Ds� ��	@��ժ	O������U,C
���$�5Fq�v��
`ua�B������_��뉛�]���ц�:l��7�s��trTg���pVE���NٯiQ4\��snJ���h}�Ғ�4U�Q0<zy��ǁ�p3|� �|��[��;�o�|b���{ ��^����x
tܵر�����"��I��i�u��ex��|?�DO�c�k\Ӗ�h���щ�����&��y�:���nt�V�MW7:U
~�zf�G��|���>�?�x�kT�JGzdQ��\��Z���_1��o�8Y�Q�Z�=�]���`DyPt/���'uhv��ǃ �D �}r�Xe8ǩ�Z9�n�"��j|E�<��û�&�w�K�o���ߞ -��,�[
��AV��hME�c��CS���攗1��I>T�݈$_b���v]tn0p���E�uIޜ3sw���Ak�Y���UB�������+��,��&e	������#�}���܆#6��)��Y�Lk��K������o�Z%�9�	�Q�G����L{����jj��(nh�c�h���F�T�f��飦=oJ��f&��a-:���55JB��I(�N2��T�>�m�����g�����f��܋T��K]���J����7xD�X�>��Y1��T���N\���J�k=��������k�HP�z.��ڏo�B����K�˗�M�����D��d̈HY }=� xOQ6���xl�;�m%��� ��u�k��-�8���d�F��	�'��C�`L�f���� ��K	Ä�����B�t5��U	��5�J�Vv)���B�[�)��1:�5!��.%�h;����:�����x/���	��Y�	h���RSo�Z5ûժ4h��	�̝,��K��ޑ�UrW�T��Q`Y}
�X�/���#(?k˾|��V�=76�x�M�¾	�űl���셡X;��z�Go������]�����0t���ҁZA\��G�Z�E&ȳK*��N�ҙ��'����Z�zb �O�n�CR�Ho��{Ų!�-�8�z�m��l�w�"����I�"�!�������h�iU[�H�J���S�ݼ nD��S��p�5�є-<Zn���Jǰ�Zh��*���cP˱e�:�	�УWv��J����f�����(��Dj�v�3%��lΑ 76�w!�/�n7�A��S����?���.����Ah'��w��Vn�V�j}�?��K�p��
����7�K`�_��
��hثP��2{�[�a��l;����Bv�XiH�Oyg�Z��8	˟����{��A�IH��B���Z�V�۷.K>���e<`p�iԴ����H( �D?5���P0E$x���\(�V����J^���j�?l�em��nn̹RI��&7{.�D*,�����5٘ӳ�����p22g7�����ψ	�%��^���H�=
�p�_?���EB2Kƚ(��Fa-u�;2C����}^�ԅl��ɩq���{��U�Sws��j�}p��B��v�k{O��4U�6���l�Pg��Y`�^%h<���r~)�4�X�5eB���VĂkD��EI
��\�h�[��몆pg�
ڶ��ﺉ�z{� $B��3X�`Qv��[��'�>����NO*�(���2Yxh���$c�٥�\�:�5�A}�����!�$�R�L��8�Y`�zRi�%�g�@P�^�,�� j��<b�,�<��5�L��^oz��}��v�l^���!CI}1�֐x-KF7��b� `�Q�D�˨؄Q��Rs��	���z~���r!i�(��CVh�<e���h�GlP�<�|A�����f�Y��_G��7Ց�}�=�WDO����a��@%.�D���*��|Z�����$a�|1w9�TҶ���u��乇�p
Bf�ġ;Vl�J��\M�O�7����Dw[�Tcp����^ ����UW�����~e�o�D,`�4��d�1�ނ�Ī�g��\����D)k�7�"�U�=�9��4���=V���i��n��J�Ҡ�?�`"�D���%��͞\i�R����p@�{8Ka��*_Ġ��!����Β_�^��+����� �B� ��Ყ��8e�֒"2C����a�k�m��.i�/�s���U;)*(�j�LW<x3�C��'�F-*�4� ܝ8agį�l�,�ir��]d�Z���]N���r����\����f�9���`�Z��]y�0�/1��/���VK-*���0�y�T�\ [0�0O
�u����u�oC��`��M��.���ǩ��4�=�x�7�׌�Gg"��},�o��ds�ۯ�C�ʡ�Ƣa��o�N:��6(8I�ia�G5����ɸޠ^���dA���pJ�J��)�}Z�-G�͕n�������zVGi���X\*h��-��'e0�Y 2yʣ�� i-�tu5sIO�ww�u1�U��Xk�\5ݽ(�:s���W�8�B4����󽣙�N��+{a��Sͨ��b�����_�
.��@��nt��
���연a��S#���z��մ���a��)���ziLN�A�z�����%�2ԯI͊"ןC>Ѳ����<? �
[��?�s���p�Mʚ\�9h�P⨐��u���A"nY!L�g�S"��a�F6����~��u��
�ʑ[hRJ�$&�<Y�����~�t�P2���wE���s���6z��|E�n�K�ځ��5����V�U+�N'�����*xr|���d���p�	q��x�*���`��n�#T��
�hW�|��	��zE��[ٺ��	��H翟�m(94��T�p�;}y��)��b�"M���v���b���.����2�6b�B~>З�H�c�x.��&k��X�l�\O�~��
��x��h9ﶬ�i��b.u@J�BN�J|whx5��H_e��~���	o��9D����r�i|���X:;4O�N��G��[M`!Y�-������L��x�K��ǗH��<�V�^��
��a�y����tŌC�n���%Z���@􈒂7Ȁ	�O��a�9k-2��6�����c%����ٌw`�ۍ$���D=	j���Ir�
�z�Tr���.�y��J ��|q^d�/HY���F�x $� ����'��-n�+*'[�J��F<��m*LC�MNa¨@�NB
x�Ľ?�#�o�ܥ��M��rhEU&�\͌v����?Xua$���2��T���]�Lʎ���0�H��2)K��e��ˆ�c��,U0��8�bq�֔�$�9��+1��?c��1F�[�\�v=���?3�N�����*a=:�%B�9�CKFI��P�x�`]vMD�tW�Mwء����U>jrF��������.�k9����8?/�{��=�ສj��ܒ-~(��:CM�"�-A9	<�qH�����M�YE�D�z̻��Ѥ<0*������N��|I��zXҩ����	�z���C@���V�@�:K��A���e�6���ֳ�:���;�Rq��{+����ge����x�y4�Sz|l���a �k}�-K���� �Y%�O_���z.vB�����X2gb�ne�p<�P��lz6ĆW���*������������8��T^Rߔ�վ����/��I�q�'���q�B8�����q�Wh����%>_�P�&Wd2���r����WX+,Ai^�d����Q���3��^'}�>��^߼��Ԡ�O� ;�%��"�m%M�I/�]��뺖�ղ�g� g�M��s���rh��
��gA�SlL3�i���e���6��Hk�b��ej4y�'�r
B<��sf?L_nlo\4�H]�G~;L�7�ߜO�&'ٜ��Z}�U)���t�R\C#Ef5��t��d2��QO�~�=!Bd*���?�լ��v�#�m�\O^%�8��NT}��� �֓4z|���۳�:P�d����sN�6�S�(���R>":  C
�	���r:���:8�&�\|����(&	I�#h��3��2������R�\���f)���z6'�'��Z/���8��2	ݒL�8�Sh��尷�-���oo��e�'����չN�J���N0�y_��8��E]��|��L��� f���Y���'~DXFيOI�Ud�|A&a�e&_��!lμ����T������0�x� �
�w'A:�q��&u����vL�I����E���}�[jn�OvL� �^8�]�]$�i%�.���஥M���)�>U��ѡ��$3�oc���Ϻ�Q\�zZ�״5҅⢺���z��q�k�/�<D^���I�{<<f���W/��Ņ^�g�@�L,?��8p2�t���Ck�.��X�:ԅ��)`�Y����u����C�ַ2 rϋ��������~˗iDȊٸ��F?y�=�׈�@�-��O�ǔ�|�I��=�
��&_!��'�$�`�v-�-B\�j����i������z�%+���KN|4��#��*�%T��u�E��(\2
��ϛ>MZ/M�n�O(���ݪ��#��k��!ȴHݣ��4�Y�8��F%���7��Q��=,Y�f�DT^���@����Q����آ�2��,����<|�m��Ͷ3<1}l͵QN-������$(�Y �>J��9[�����sb��Q�Rᓇ-t|�����K�#�}$�&�F��0��r:�,�/����$�=.
T���t(�M�	���}���?�|����� �⻛:B�I"F*��ڻv�"`���N�,�e��.*�>:׵���kqi�S�dt
��7����̌0�ƭ+!�\�PK�O�ݭ��܋o�_��I�
_��2���`��2I��s�u*��"���}�-L�0+ӧy�>dQ�t���#Ɂx2V<q��`�������4yp�4�����Q�R�����`3/��1�׭�yT�pr��KoM�9�$X��¥�4ְ{5$/�oK����:����*�c{��zG���	Л�!��������M�012r:���P���J��{Z�DNmnu�3�U�O��)d�6�h{(���V���"����73��Y(Sc!�a����"9Xx�������J�A�#�Y��Qn��X9�Ҵ;zLXàQ��\{�o��w�d���Zz�8��)�τ��Ihs&*��羭���M��4Y�Qf���U�����>��)�,���g
�a�KzV�m$��"Lq/~i�!��8ح�	m��y<�w�\.%A�O��F�䝪���ఴy���L$"��,@�@���}���5��-R�N1�����.Ҩ�����vO��@��c���5ī;x+�������nU�E6J�9ޗ|@XNk�����~ع�eDR!�v����[B�1�K|o�Շ7w�H��nxd�<-ҤSۑtɩ�T�-U�� O�d��E�R%:��̚;AAU�]qگU�~��"�nx, <�o<y�~*��K�e�;��_h�Njsb��B�y��⁝t�K���c�O(����m����^>�xP�?��a��F0w�L;�o�庡���f
��m�	��o�#D>�!�q\˥��WHI�1�<m��n0.���V� ����FM��f5I�C����O:��[��v	�s�Ӻh�k��	 L�R�+D��8�Z��(Z�V����u�]�d�}�1��=M(�K��}���A<�`
�F�ڽ@�r7��G��2����:�8��T��l��E��QI=LeZ��z����_���|�����N�q�'�N��s�U�[���v��g"+ߦQN��6�lr�JDP>����bO2��#��e���9����6#x�;#� Bc�$5�H�=�:��/����9I��c�Ŷ��������qH�A�6�x��/A������V5b�>lwD���'d�{�P5�ou&��ޅS�B����'w�9�Է���1�ǉq;��؁�}��*n�<��'B�ԟH�'�j���g�L;��ORXlA'���Cg�N���Ԟ��k��p�{9e�a3��  ,s�m�i��!�W���
��媽�#V��U���D틘#�ŤY�1R� ����
��t%�2*f�rI!V�d>�31��s�4�L��P�_X���R��6.�Qm�2Ͼ�[B�+� ��FV�j���HQ8�9�\���[�X|J�p�%�Ϸ�����&4��,��t�{�?��i���5�4�����ɒ�2A͐Rs�6�y�R�ϸ��ʃ�+�쐢~K�v�vPai,���7��S�U�ѿ��׸̩��՞��8龉DT,j�4�Bzs�+�6���5{�}��j}�+�-��0j$��k:�D�N�-�����K��_Bh&�h�~�^����<Q[_͕3k:(��?���M���W��5��xY��c°��%�Α���n���Z��Ak�v�8�R�<���`[�`�̛�DJC<	�0ѧ�:�����H}�3+Z����G`3��҈�1;�܃ �m�.p���>`blܣ^�X;�Sg��~T��r����l�$�[!`� IJ~�]�x��=���D�h��i�R�q.��Yŋ"!�m?Z���Z�� �$u�"C:��;��3��8��P���U,�Cۄ��_�tJ�&ò%���*G!��61
����p�㾏�<0{�&�&�d�x��c0�����O�K�c9�KSz\z���+,G�5IrF�k�9�����3���J�U���-���v����C����1k���������i<#�.&3x�x؜�Y��SE֐�7��k��U��j�7l(p��+��#�G�1k
�2���+�@��=⮮�˒�?�J�u�g���'�N1'X��_4NK��Pg�8���;:X|r���;!�Z��z=�ь��`��&tM�����k�Suѷ�� �pT��n��(� �E��fFS��2�*s�ډ�k�_�vН��[��I�-⣝�B{uY�ne���@0V�=@иԟ�Y��Â z��%�Gy�!d��Sw;R�ќϊ���ݦS�'\>�q��/@Y=�R����<������(\�ݛl���m��
�Z�ݬ�
�ҡ2��QI/��o����u�е�z?++�~��6���m,3P�2�0��o��~��~i��\-z��*�WSF9G���y�m���|ah�9Q�Օ��k�\��2�j�èYi�U0��\z��r <E���q<d �R4$XWUf��&zm�&�B���"����iQ�8�X�RG����:���L����?=+�'`������r�-���}�*Nq���W=c6��5!*��!&������s��-��TH��k�%pl�m������ Oq}f�10(�E�/���_�XuRW]�����F��ǘ�0,�}�,����!��ܴo��s�ދ
��<��,����������<1�+6U�_��/L���L@xu�����ýS`���`~c�`�.��U?��	���b�<iyA�לN�������	��ʖ�(
@�K�fڤ-�D&&�:Ѱ�xw�be�~���.s�Mc` C|4IG�� �L����[�V���U�D�5ؔ����������X��������͍t���k��$�	{Y=ұrD���-�tN`#��Eg/��5�!��t�i��T	�U���P����Sl+�3X8�)ۦ��'��u,u/1�g�>?��d�O�1��8?����ydB�n�2�[X��w�;O.�	/�f���n�p`ko5��i�ݕ�Η��ur����uwN���P�D���t0��HK���,����XW$��eU�Z���̿���U whH��6�*�y��]�n��]Ż��$R�����o���;�v��P)�����t77�ߓ6�Rk¦a|I ,z��I^�K"�/q�R;!�S�R)�
�)��.�m�o%���C\1��d�y�I}� 2�`G��s���0��������8G$�.��7�wN���D�~��}vq�i c�`z��=�Q=��ՠCi��m����A�%��?�ގ;�	����b7Ii�����������݈!�>���3�d�-
ϻ�P�ֆ���N���:_��m��	� ��:,�/��B� p�'/S�����O��;��~���DƼ����)��?1����avN�×��������DH4� [������ț-��E��qa�OD��f��'�BXS��X�6��*����w
SJ�J���c�*�Iz ��+�N�g"���Z���#4�0����#-S�\,Q�m����LY�"��Qr^��躠�j�ˢ���X�Y���
\�^;y�^y�2.�͂�־�;:�����\�Q>�"=��1��	���c할Xq�@�\��x��֝�l�^�|�����V�{m���0����Ed3S$c�ħ�Ծh�������� ;�M'B7	C���,lc})���~���	�G[�`�!"��C|Ɯ��:��9�f
Yp�o��WmxS�{!��p$��=��؁)r}�Wl��O����T�g�&��J�˭5�Wp�Ӽ��k��K�@��-�&����'S��l�)�b�Y�g#�v)zs?���V��\T�y����9��
�q�5r��;w&���>׏P���-yп��9a�Z�w1�����!}t���H�d��:{�9�C����A)7 d�����Z�?X���9���^s*�8���J��T����PE�y�~�|ʫ��/�^��!گF�Uwb�L���n�Ai�*Q?",u�*u������cL�y=��,^�$T�N��&����fڂ|����9Ѫ?h�$��\�%\5���)(�mi��Y��\2����Hڗ^��0 ����I*�x1�9���@�i��LpG��_��[�<=|��&�m%��n��2�Ϫ��]�R����}�?؇I��X'���)��e�c�b���I���`�Z=ňk��d��υ��c�h���3�El��̴�"�����kC���>8x�%����Vc�f����8^�:]��n���;�ŏ �1��'�e\?���J�ѻ*��X0�|X���A!��tD�.��H����"���zh�� =��U���r�hÓYau��'b(��M���c>��I`#�jHY�	@�BS�j���|i䬦����
$Ng^|��{4�?,['����a3Ϲr�����a=2v<gɄ/�=��F��rJ�}�;�s5��-G�Pw���*JI]t6�F�"?4�C��Vl���������uHl��
�Ё^��w�u��mv�CmؕJ��O��*{"I�^bQ;��Y+t2�*�Uf텰ڼ},r�C(��`9�cX�&�����mw�j�ֹ�b�_V 8��x�2�5��vo����c!A�#T�&�5�	j.l�<�}!Kr��."��ga����_��v�/�)��C��7Pi�ed��-��j��>su���Bf��e��.m��37��t�g%�p��29���DT�m���M�ʚ8T���<�(Kd��}-"U��F�Y"�od��ƞ��s/2�;�A7f*Np�8�ƞ�es�D��M��;U^��ME��"IC�\1	Wp0���f�K�oB��7�2�$�mC�[�|�u`jT�X*T�����f�y��t�\��M�Uf]Խ�'y3��8����_1V�ß~�>r!-�	�+�[�\-���=�Fj��okL5w���O�8D�	���V���[S�dt�]=#2Qs�'�0�4)��D��ٲ�Y~S˪�tnm��'WIl���� hYU���Fi���*���OА��p80��������M�Jb��l9/�����k�o���iC=�v�B�����/��| K@w[�X�4:QE��Q��w��:&(�a1���G�`H�{����e�R5��;+{�ӰC��i,$\�F�?ޤa_�� 3�q���-�%[�4����K3����d~�I8Z���N<,��i�|e7��nb<bo��iQ� �����#�܁�X�<�N��-E���]��U˗��+,���^nO�yNu��2'��;��6��]BGQ��H�*!f����7kô��j]�4�m��͂�	���V4GY0���P�4%�]��+­�b"���I�3���LDO�m�y�,��[�D��{Aۦfo�=�N���t-�U����ú�,��4�F��-Y]��Љ]��UX��=&/��YĲ���S����e���Y2�ut[�V؛U�'��
:v*�u<&�z��N��+�>�o�	��	GRͥU=$���L����Fd�-M��h0sz&�>H\2�ٕ=�|y��jq���gڕa�YT��On���~e��5�����d�Y#B5���@��%h�5oK�����NKK�&�F����קYw�>L<i�A��QbJ&7���
�|�����a�t^���!g�k^���g_M�R�Ȝ3�|7����$��6�wRӣz�%��_)E��,[��#�hܥ��v�br��8�,�3��
]|�qO�����zeE����C���E|���M��Tُ�ՉGLid���u�.t������4q�1�ӏM)t���YM�tߚRB�n�\�)�qA��Uֺw"��*�H�e���m\5�)x�+��;!���ʥ

�Ndp�
��1i�� �;I~y���S�>X>���ETބh.+F�EL�M{>�
�	����J\_̈́�s�g�a�I�C[4g-�f�u@�ƈ�X�opT:������a9�(h[�
^�x!I0�5��sq�@�x6��i!ν�I���o�`�q�*MB���$���KC�b� Ȃ�
Gx���ܳ�q��A�mj�ޒG�Tlwp�l�����`�&YF($V�W
_�m�|Ǉz��a$� m�h-H�iM�a�N��{��m<Q+�j���i�@V�:B��е��D���I$��s-ڲOJ���	ă�
���+DS��>�zP�v%S��ua��2����nVx¬���؀���#=��t8��Z��,Ĕn��S�*�����5���|�H�������z~s�WA���%.4��puP4_.c�D��R+�8^3/��b�D7��+[���&��]h2�B6� ��8沅��Z�1��F���՘:�f�Ưg��:�d&����~������d;�-,Vl �r���+��Dn�#)aM(|2�enE 娟�kӟ.Ũ
��J��Cfih�ؚ�*�?x|�E�! ��jט�c�t{�aЮ���h�)�>7�����U��L�I{�4�@,��j��z5��RI�Icr�l���<-����W�����Ҡ����V�9�>A7(�W���9����]�q���}�b�,��㼸(�h.9��mI��y�c�U��D��>	r���;:��35�M�C'v�ߋ* ��Nn��K[�.Rp&/q���7��ި��5�V}������%* ��B2y�r�DHP�L��Fz��9R�����셙����vs�=+�;��g������=��=>�Oi���Rt��C��`��Ƴk�p�ʹ�E��H�I�Y+\x�,�ܥSp�I��C��o
��q�ɐ�(Ab
K�5����$�M�~Տ�/�R�LooRI+AcX�:�	�O{����[�\����k�\��y�=c���c��ūtV0@��)
��)���_,c�F/���k���O�L֚P��H3�~���T������+d�!�Iz���RG��$�-�	W19w�#�!���Pa8h� VB��S�;9,�#��o�5��Q��'�Շzb��C\*����)*� �*��P(��,YOמ����Q5��nipCq�F�y�lM,q������n*׌{Y��t�D��X}�>x�$�|e*v��Q����J��������
���-#{v�P�K�]k\�bx.G��p8�$��c� �/�?����lyѺٜ`�����F0qZ���P�>+=Y�&o��G4���H݈��-�6j>1Ĕ܍��&�=i��сՏ��ruR'�q�T"O��sf���7���� V�5�Da��2=��Sٸ�h� �c�|1~/Z�~�"��J���4ǧI���� ��3{��N{=j�zm.0����I	�'�Klwļ��K�M����=ǣ�}�f��Sd���R�0CJ[J���y�R��6�?|o�#(���HW���U�r�&���,�&�1X�S�#Sg옪U &_xj��h+@�}��*E� �
�jN�>|r
o�B<Y
�|���cRk�h ��!�my`�S!"�.��N0�ܹ��!��f���m��\[E2���ټ���� �ѧ~��f�I@#��,W���{�Η�1�\F�Omҋ��~�Y� �g>�N��~�߁[��$CM��K*�V�E�3ce:$)�L/%�qn#ʮyHX(��W4Ha��Kb��x�:��|�?�u�� +�o�k�̨��\�e��vל�E��b�Wˋ�٥�"��?;S�R��:�
Ս�����֜�������WmF?��sb��듒�����<�4�?�O�r���>-
���::�}�F��	�̿���ݾTCX�~�`o��=c��V�`�ԝ6K�9���P�����-���Q+İX��
j�l~r�B ?�K��e�V�L~�������u����4PM	4ք�l'�II�-������XϬ��.�F�i���>�����k"�kq��P��]��_��+H�#,Vގc*xK_K��5�j���ne��;��ۓC81nƥ��0S�.|���GA]�!�ʹYRd0�	:�ś��D�4��,�jx�J��w��_ӱQ1�ݵ3�M���=�a�N�w��{��3�O;�o�E�^�B��)�(�E��_k���ӄ��۹�� G��IM�&�4%���+w(9�y�"�.��P���a���M�7ǋ�q+3���LzEU9���9���%%�n�l<Y��/�j��%��Y����<�[����j�yH&��د��3y���b3j�?���*�Qز�<݌����A���T���$������ҏ�L\0p�����ќK��h�� ��	᫿_� � 3nW����)B��	=bI�,�Ւ>{�Լt��t^�E��U�7����o�RH�e 0�l��L�LP����1��H'�5m�{cgA��pZ��dd4��Xn,��c��)��U��8 ^�5R)�z�W2����N�����O��-�7�R��5{�<7v��`U����Ms���.0��[�&�Y�^D����������p8�|��X{dF�\쭨����Qb��B2H$V�pmMݩ������$�|״�h0�8�5����Co�F��J�$�*�F1�r�$A��u�'a��u={Y|6B�j�1TtIx'�����:���pM�郭�yI}k��_0����J4����a1�B>�lVa�ck�剥��Xp˰�n(�U
wn[^�TD�u��/^������������������N1z�q��dKtS۱���nL�����d��s��eQ�B�x�`�})f����"6��;�-���Sf��H
�5�9�OH.��g�'��	�
Ak�Z��N�Xל�N�LN��۵_脄/i�:p��"�w�'/ ��W�^���,�W��W�6BWul�L��9l�x���td�����G�~?m`�͙&<`�@��A��o�z'GSd�t/���xC�U`=�� �;��R*�j0�Yp"�再����y�� 	|�g�n���K�Ȑ�B�oB����/�WA�S� 	.�-�|�+������j!m�Ј���  L�"�	�(|��H���no���Dj;�C�*+6aޡ�D?��:\���˾��g���}%}Eus���Oם�t߿=�`YT�a�C�ۙ�>�z�p��R:Ȗ���wR"��C�������=�����{�u�8�K�N|[S2���yg\e:1�A'�����90z$^�*\�V��2P�Քg�����fĠMC$Gػ�?�6$�(���x�1Ƅl̂OfЅ�<�w�"�T�9w� k~��AP�p`�øĳfu�^,��;{�J��Uٴ��uĦn��&M��VS��`{!G��HOt�۸h�5�z�~/�Ɏ}����yZh��������?���At@��<���$�I�������o�Sn�/�� �E�wS�+�*u 4΁�U>L��RrD5לH��,++|>l�I�s �`�Oԫ,����ĝ5vg���jT�/6�~b=�rh­�UUI�a�N����^R B���ţPv�5O�0��;�g���o����v˂�y��������e#���))|�Cւ��o9�N�-4��[ِ�J���{�d�l�А��L�O����w#�K]�fVtK�[y����b�d��t��1���N��{�V;�}��{��ֈU6֟h�#�~ʵ��]c_�t���D ���]��+tW��+=P&]�v�a��.>1fK�����f�J��ivTc����`=.Co_��0[����,�|���^'2���#ѣR;9Pk�;��^>�z�]��{�\�P7y��+q�Q,��Pʩ�D�L�"�:W��L�������EX�G4x�F[������@��nc��X�y��w���ސ��eCA��X���Lj�mgJN&��@�j�X px��%�����H�i|��0�݀��v�FTA�3��t8�9A�R]E]1��Amb���t��.2��E6�O��?�\�M~��h�̌�	&ӑ��c^ȌVs&Fj#ل��*!��Xt7��s����8�%&)�?p"a�1(J�����7OA  �E�**T��Z�<���W��o(E�A��������	8�*��)XS� ���]VV������P8cJ
w�ԁ��Am�:�_�Z�Գ~�_Y�SV�����*��0��0ն����Z��#ՔU������	����jl��U9w��_�����ğ��J[C3\\;�:���#ȷ�bgh�����sM�Y2�ޘ�TZwb��G���P]`eQ��#�����B�T�u�.3ЍZ��- 0(>~��_Y_iG0W��&�8�G.��5����oA|F�N����Ԃ�M�g�?B_����]�
�l[%D2��pk:���u�
��Ɍ���!Q�:l�e(�4�/WޯG��d�T��L��o,s-���G^ӹފ���ΌF���>'���~���2�������j�;�!x�ؔs���Z`���&w�5�!XK�������������Ga��3�����Tߍ{����_�E==�ŤuK��RY�/N&��&'2��Θ��-�L>wy�1E�E>���@ŕ�t���Z��3趏q�-(D����+��&�T7����`Xwږ�t��;�Wŋyj��q��?�Kh��b�N0:E�4�}ݑ�T}�S�ۑ�
�q8�I���	��Tq�?��kLgʪ0��%slj6g�"o�+꿼p1����fH���bz}d��Y�9��?�%� 4,c�����R ~Ni�X��"U����SP�DKй�	�����eD�q�j�ۋ�UZPi� ��;�ٟ
TS¶<�`e���u�VĽ)��	Y��R�_-���9�}�Gp`4$��G��L�������b�F�Z�8�fZ6b�0���8H���VT����\�R�l3�I0%m�P\����:�<�����]*&�ǆ��r�co�y-������F��Ü���Z����n��O��{��y�uY�W��x��/��9��zO����Z�3��v��3���=�qrĵs~�p�tc5T�@o�D��=������k�#'�΃�"	����6P�G�Mf:�"~-.�o�)��|)���E�=7\�����o�����1�h��_�������cQbl�R5���4�T#������ �˳��̠ħ�<)G��	�2� J���i���J9������[|�,Q"�u/�u;5�g�ث�����0%8ɟ-���i#n�֏M=u�P��=���[��&�s~Sy�S��WmTuq�O���	N�y�|���������0MXT��F�mֈg�͋B��x�+�,N>-V� ����O����T%��p���hdt��9#g?ʴ��ʫw�z�����8$S0��_������h.R��0ՋC�x
S��f�➵l%n�7MT��Gp��i�5���y����c�6�_�Ǩ~Dk�U讜:/�a~vUH�����6�Z`��0h؎{�l8��,b�X�DVj]�:���K��f<��\�؋5^�̒�S��y�BpG��c�Ye*�������w����i-_I�4R�*�{�6}:�vY���DR5�	3�ل��E�<�R#�	�=�j8ժ�KhǨs���aR��r����k��/(ն��Z�����R3�ڇh�Ê�8`��ߪޫ�R��5�.��Ai�y\f�(��1�N����� iJ��C3�o����������Ʌ�t�/*lMI�`�/����w,L���AA�"l|�ڼ(�U��7}Υ�5djj�tp#Ƙ�)����)���������>��\l�Z����*L��N^�y�_�d�o�����+M��%�S�g�ɘ4�fj�h��+Λ�L���/t	�gc
!����UW���Y c!~ă�P2�]�1nUb�,�s�h�J�h�v�w���^�Qe�ɸMA ����`�i@�bY�]��?Grn����$�h��� `�qE0������7����hi�P�6�+^�cԒ�Cw!�0�K�㵛�~�L�����%�N�^�[u!�
�<b��/Q�|ܴ��j�9�A���3�-*���$��OO~?�5J�a2���<�T��ߪ�2/Crv���ѕ�!�O�7��Ă9�<�KLR	��U~�[��Oos���9ݻr̹$^�%l::�����F5:D�o3PK�{E�(Bg��e���E/gV@*=�(�L�هi�C�M΃̗y��`lv8v��C�LRّ����lP�4Ͱ���+�����5ṗ�
�(�j���J��rQ����*�d��p�x
�Z�t���Z|�	"D����/ֵ?��NR�uuB�W����>X>�������<OP�|ټ�^#�&�l(�^䉇��+�qΆ���M��e��B�۪�>.+!a�ˠ��*��D�d���t_�[�+�_��~����wDb��;p�������tՐ�����H�e�����'#{ͼ�_�&gDfs��{<y�P�u.k^���R��zy�r�8�o�-G,�T	���k�2��w��ٿ�p�=|7�&Q��~��d/�{w�Oܠ!�7��%�-p4~����V�~'�2��LC�/�Sg?�]�����b�HE96{�s���c��5��C)w/��c�h��w6�z��O�f��Rəks�@u��ۧ��'?���lO����r:{�d�ēr$u�~Qܜ��~@��o�����=�=2hG[�߈��`��Ά�27]�0�H5t���8�S�>�7�cZ�}�WNh�^1]ҷZO�����7�ϟ���p��B�@+��8�ʱ���ĩx�H�,��`Q��[e���mu|��;<&"t�ym�z�
�hi
������':�}����Ϙ:.��CޭE�(���~�mXJ=3~�m�Jw-Qtn����$����D��4����K��aoN~��J���QH�i}�Xe��(^�2^����bY�	�Г��a�c.������(nt������,.̉{Zy+��.��
���������@��w��Z�y���������а���(@Ċȗ�����``�ы�P��vn�g?��u��l�Q O�vG l��fa�1-{%��x@�O���;���_�n�Xɿ��g��;�� ��p�Y���Hk�I�_���"�At�#P�c������˔��~ۆ�*�'e;ʲ�#��Ɂ�V��l�7A.C 㝣Og��)~<]�}ݻ���o��غ!�`R[��^��A���I�坷n��u��Qy(�}g�'t��%�3H|���t��Y~r ����|?�+q��1��#j����L��d2�Ͷ6��ڵA��ƻ��sǂ}L���冪+ف�`R"b+ʞ�i��zh?���5�$�koz:^]��v��X���f4�J�`)��$!���[8=f��[P{��@`~�������3+�a��R�����&O:�R:�%�O���b=N��y�����)��f	I"�*|��+�����8t��*�&�u�5S)p�Ң�@0iHa} �t��
f����W�r�~��n����I��Np��]�h<���O#�arj���=�9j#����̛^A��@���UZW�5ܖ��%��Ss�`{V���s|���7yohO>�^<�I�]E��-��K�G����:�$|
�:��T����@���s>st@;f�{��<W��I[�~J��������U|N;Y�+E��s%2❒)s�B�����E�_�xK@T�˄��WB��	����+<֢\��&�Ԧ$?Bp��\q��H��fG
,�_3�Ol$AjHP��˻��b���.=����i�������_n���m���tc$��-�뎖�.}p�Tf��ZA��D�0	"9�������� 9�6�x�FD��ft�1�	�ћEĬ�M�@Z�^E({r���VY8ݩ�zp��m̔�A W�����Sh����b�:��꺗�d�^�
�O�E�hk��'��̒&��ct����]��6st�4ufҙ�PulFg�_Sre�i��xB��u��J��h������W+��|����I ɞ�:�y�@'�Z������@]�!�ɱȨ-��hZ�S��<r�~w���|�6��jHx������gp�� ��&�[<�@T*��]�g��j������?��<xu��*[Mh\76�85n(v�d
��{>�lSqL�a� [q�@+R7hЭn��2��(?��*����3�5�����0%m��2���.jl�wCYV���ycT�c������I���*A��yD�\İ�P^�W���D���Zx�(3�f����>%�wK��&�$�lj�u�D-#ݷ��M1_�Rk�.4d�{{��`;����p�+��ԏ�箽s�b��A�c�#���[՗�g׏xd{>č�I�IQ�%�"�.��w�a���\r1��n�b[��F7��������?@a��E� ����Br.;�A2IX�͢�GH�m�T�i��vK�R�Q�ʗ��҉��^�`�.�⽖�!C}rhL���e�J%��軛�_�.�΅N�o�9�X���,��i�_~�#��Q�*�9�� ���?<f{:R�W"lJZ[ �c�ٚ(��J���܃�pMnAu:������1SH���j3)55�Έǟ�L�QݥBp�6�UC���]w��G�GI~�d#n*�hWqW)�ߧ��'lĮ�΋˄��[h�ɿ�Y��3,�F��[KAé����쫃g�����^$�% �4<]+��9�tr\ ��+�sJ3B�@�z&@�.ם�"����"���~��9O$��(Z����k'�T����O�'�}����h\�n�/M.�*|�/��f)�78)�Ё��rJ��U����� �u��������}h �!	� G���~���r��76��Q�-�o�tl��I�I�ɤb���~�ޟ$�s�\�L���������KW��f��Û��oϥ��Ca���}T4h�T�\݁S6ū�؅[\t��K������p��n�z��2)8��%������k#oC(�K��M`Ͻ]�侵����)mT���	W}�0��qY_C����;��WX>�2*�WT��n16�P �AFMHQq`�����!�#�|���-hS즟��|��^����E�]:� ����5H���ne@$�3]ĥ��֞��E�Z�B�ܡ�]�P��f��=�>�fK��%��sq=��)��x���J��1I(�,we3�R�>_��yK-�j��L����#�U�Ƞ�hgNo`7��(�������e�j����.RTb�L��?BB۩g�R;�9�)J@�(�(
j@.�]��Ȁ��T������8�\���]⮇�ި��b�R�ӯŠR��=yˣz��Nx��@������-pR֊7�{95[CdW���MB\�/�=
���`M�t�i0�<ڧD���'��"�*r(�Z��ة0�g��6'���uV���p[pf�P�qӽ?wU~$�$�9��'FLC�����lXqk�8�� L�Չ�h�']��g �*m���	%�1�d�J�J�(��S�%��U�A�I%�i���Ё��o$�e��~�veܺgSO<k�YǦ�5Rˬ+����D׍(d� ����A�+��scR��cFZ�tD8�v�]��?[Hޯ%W�6�9cR]�Th�Pc���l��a���ב������&J��W�y�']��+�V���36/����L���y�ܩ'��O��"�CvY�mh�5bl�������6� �gb�Xґ<ؚ�A}�Z�#�kl�K��Ṙ���K�?�QKC�*�����;�͌���5�%.O�7����nFR��K͎�^�(&&&$+9?Q�/��0��Dn��_U�>h2v��2�ۀa��X��c���e����
��5g ��s�Ѿ���#j��Gf$h��v�Q@	"���� �����I�EΈ��K�FO�*�m6��/����.9�����LL��ޥ��I��q����U墺�x{�J�G�t��S����bi�4y�Skg����'��b�؂�N}�����4��1���?!�m;|��S�1��1�K�'��7���2e���c�t�W{�>��/w��k�����܃��:���V�Nx���._�����Hp�6��N���H�>Ȃ;�6$�J6He4�k�%ׂl���/��I}4s�AO��O�m�����v�jF���).<w����o�����[NM<Ś��nޚ����?�K-�b�+����:z����@��U����
��Τ+�{3h&cb��K�?MrbN�V8���q�Ct� ��h�*V���*$����W�oKb��%�y�(����D0N 0����g� >���&"�t����3	A�b��0 QQ�)�@�Nt1�o?ѻ���B� �m�����K=�)�A�����C�^�n����r�����]Ю�0p��[$�����MҮ`#�_j�瀏�-����m�T���! �g�`
�QL� �H��XIM�*à���/_�۞�l���Q�K7p_xb���ͮ$�	V��N(�d�y��q8�5��\���S�fy�ܤ3OT��$�M8�~eE���roV8P�!Ri��&͟���������3�0��²ۯPU�0��eܾ���Еe D(N؄��8u1Y�Q1
|�{¹���F�xln5�w���b�	�T�k��N��}׀S����v�9�e_'�;R���4�t}�����}f�����q&:0E�ɔ��#��.�Mt�uAo׶��LB���\�HM9�������� F�|���8Ɓ$vkF�@�߁�e}��tX���"�.��F��nA-����-��q4��iNC�n�xB(o8����ãG����n�F��9Q�Μ�.�����T�O6��t#����{~+�d���m��ʙ��v��Ѵr)� #��V^眜g���-c�tcт���e���4���7-O��~T��z�����;:5]�MO7�_���}˭[�ɸq�TA�*Y9�T���b���t����
)�;�u�����v!8�U<��b��Ћ�D��Iv�؉��nx���/{�
gMq�\����V������[��"O*��H�a!}�f˹$)���Sd�}���-nL�����Rl����_�\ܮp�|�	K��Crx'������swZ�xo�L�I�?M^x� �+��H�*⃯������J�&��G�[A�H��oe8;�<[`�2>Dl�8�&l�4N��i��wUO�j �<\�+g��JgM?�v2=�&�����B��|���WgQ��Ì���f�f��􈉱/db
Rf�EI�S���F��⎤X���$�K�f�OGۦ�&��#���MN�3������ v�ϴ{B�3?�˃p�(����������c#��q��E����TpG��T�ُّ�j߅t��Сҵt�w�8l[*S@6�È��lꟷ��B�����QSP��_J縐�`4P(Ē�q�8��	hC�a�i+�uf2$����<�Gn��^J�:���	P-2C#��e���O���/=�6Џ\�D�<Q��cɭ��a�;t��*��n��O6�Cb�t����7�����|�w���`�	�,���z����SGc����6��q�!�I����`YF:0��.U�@%�p�a��Mo�K���P����s`o�m-1��a�ߍ�J��	z�#��xެ�Ƽs1D�䊀�&\K���hp�BU�	�(�I���v:sb�A� L:�˜�������l����
� B�t�F��l;��%�(q���wo��q�2M֭��j��I����KN�+�;GS����̩��0#U�ۿ����(�����#�*���W$D���
P)���p�4B ��gL���۽��k�DN0��2�19yfzI�P�F��$ƶ���Ѵ�P���KF�fH�nP�5/l�
���J�����z�טyv��Ǎ���U� �y��9j�U�f�g�A��`��榈;������z�0�h��#������~�[�N�7&�m`/�r�p1L�1R]d�];}�����Je?�;_�Nb���}�����ީ�����B�c=�mg�p�7"���-}Q�۫5�S�׽y�Nj�fT��H��x�L�����E��2�j'RN�����N�p��R�ϣ����'��b���!h�3%��Ic�����Xq���v�L��H<��5�q}�����8h�ƺkT��"�S�� Ә�@?�7��X � C��ǫ�eX�L%�}#k�Qב�;]�_/�0���W��o�Z�\�(s�M�\�'��g�1�N�%+�:��?��`�$�ߋ&I�����B��/���<�ci(� �H��S"����$�䀩�4�-M��[�Qs�vM�̞�bo��kx��l��`�R�_@+�k7��<�����'!r�S�Hݻ��!�W�^`��²�ľ�,[��B{���|�)���H#c����ǈ��̦�����$�Z�tǫ��MT����l��P�k�ы�Җe���AQ@r#�Q$�����$9��,�P��N���#�fNш����wھg���տ�{?�g��f;ST5C�^d{+�߳�u#��@�	��d�x�m5�a��>�e;�)��,�Pоl�s��c]^���0@�����S��;Np�-Ȱ�6'�ݲ润�:�`�j���!����G�~.�M�;��۬��$q`Y��ϯ�90xߨD	��׋�LsE�(�����2�$�K^��q]�C#�1�os���u?���TĉhU����[���7{7:y��tu�)^,@�ͯ�MU��JP3?(� 	���.B����htN��������ZG�	ώ��@�>n/�?����~��F;!L��aZN^ڌ�B����*V�BO��x�0^^�lDЙ� ?I�Y�b��yNvܭ~��B�V�co{OG�:�;M���1\2.��5Bb����g�h��Ȭ��o�e�L�&�Y�u�S(f�M�()�(I���5F�b���;���NB�Ou��`V-q�˧>t���q�ƭ'�Q0F7.,F��	F�[��;.�ɺO%M%����(�;�?�1pq��p?�J�UG73�f*B2`�L˱oSc��kq��W8���,g�M����4�HBw�����x�d�k�J�O�����-��^W������dT��gǚZ��O:O����6w��j����>��t��LS�_�v�U��M%B�^�%��Jy�k���X��q�Z�ne�'��n��?��(� �b�t�<�p$��,���'$��3k������4�b:��M�ӗF{�\����=������6<�����|+�V�Q_|�e���pn�\-�nѧ���T���Dz����Rք��":`t��z�%A�,Ի����$w���O����.%5�,��X:�gI5�����L2=��h�3��'���=��`@��M$��йq8��D��A�$�d�����_Z�o����Q}r��a�$qv9.��a;7�M\�֞�a�i���og3;<���`��X� �5�p�w���4U�~��K$��[�"��(��>���P�/�����}�x��)����YE`�ߓ��j��a,	�i�*v���L�shj��E)ɾ ���Q�_X�!�yCN=��)),E�dyd�k����gkQ���@��UTVT<��6d���n�%hB'�qxT�h�����D���h�y��CQ�����@b��J��7�;���(t�j��$������b�&sj^��IQx�PLU�x�Q����/�*��w��|}�%�