��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g������*���Li�ĉ�3���R�\��0}��N��i�b�QO3s��N��㐝p�W ��Kl]���BI숹�(�a$����=ZA��Z��<e�TrRd���t�o#��K7�QX3��O���� eT�2j�Ŝ�5�| ҭ��\���I$��Ng��^�i�cۣ
,�P\��B:�CN� z���� ��hc��GB	:b�[�5Rf���il��.Q��</4X <�Z*�Zv[Sr�w�P�����˘��C��\&�η��zR��bA�AE�Y�w��\�7¿ȣ���p�A
 I�!�C�^�@��r�>��9�UJ\�r�Ԟ��n�c�ޣR��[A��?��"��_�(3��n�(r�K��ĺ�vhV�L:-�M����
1��l!"#�v��"���@'�,�;��z]�pѵ5�Nf0`������ s���Mތ��h�F|�=K�zm%�!tY`0�ߗ��wߥ�Q����n�PuQ0z\x`��>��x�m��}�(Ʈ̳�5z�N�t���2�\$�Ec�#���O�vޱ� 0�E^o��P]8"	�hX��@�W�s��Y19X�H�$o5k��l��UuK�� 3'���h�-0~�1����1���+m��`E~t�>60֯� VD�I�Jhs��hbQ�.w�ǫ��1ņ�f�=��7%b�8������V����o��%ߥˀ�$I�+'�ibK�ӂ��N�Z��G)+)%�3�	��O�U��k�5���һ�����@/�����I_��M�*+�*��,�/����S�J������� �'E�18M�1�
<�B{qq

�����:�|�S&����Ű�o��J痻���ivdR��ڈ<����t��cQ��n��+�C��TV2�s愱f*�18���ӈ��T� ��K�lP�IsC�gC���_��;Dj��	�**�0Sa���Hic�˶@�+��t��xF+a�&�=���EqS��j+�/����W��a��;�`ϫZAM�
�qM� ��c���mW�A����^Bd�[�s��f���O�9{�P���iI��^�׺�&<7��H��Gy㱺�"�]^n����V�U�^�a	\����׹x���������{u$|��	b�T�O�����8t�b�U>Z{^�]��Y�{�+V�a%�� �2G��瞡�.b|?:.�p��$8�SQ*s	�]�Cf��]���Y�|�W��J����/#�7�9�E�E��(��}3Ӽ�x�#1�Eo�n��#"���|���@�i�eĽ��)ұo�J^A�/���,�C������z�<���%J����.��U�=�\8X��ƪ�6~��]L<nꓜ�ץH���eɎA~#bg����f�-��Z�+��	>K�n���f�/H`�8�	/;|U�
sÐ�`c�ihk.�&E�(qeg�_��z�:�p�� d�� w@����5�b���T;I8���}2"�Y��ţV`4����2��~��mu���D�u5�;�ȣ0h/��׎P������R�����6<zjm ��c ����v���0�n��:�δ�]�$���S��yS�'_�\�)IB]u�y��`9
*9kB�f��,�&�6bF; F!���rG���.�QA�	1��W���z]�{�CЁc�6�ER2~m>q�({�w��D��c�s뜎�'���茇�ϕ"�Y{��_ <�)��q-���`�d����V�A�xQ�_���7gA���1vm�y+�����5 c�H�퍹����0��M�Z=���/�����b8�;�X��fd��IO��6�]v�ٞƪά7�;���{�MQ���F�Y(iY��{K ?Myb�IP!u|��Z�:���"Xb�]���(�����m��3�k�>�+�;[� c�����DX\��ݑ��}�q��-T��H�6>-��,7��l5��ZC�U��������~d~ׇQ�r��z��]>d����Mv:k�JR`�dE%&�(��q�p���z����!�~�]�&v_�}M0�i��3���yb�H���w�h�}�]��>up��B]�(O�GѦtپB�daz��[��&~��=��c5q����rɉ�T�{bU�}v:p@obRh�@2{A��)/���,��O���T�1R���+�;�t�	��~��?u�3�?YV�a����p�,�|����V��_Mi�PH���m��·�zAv���Kڳu���-s�!���_��ըr}(Zg�H�Y���Q?!&z�D����藉�#Ed��Q�v��bj�]mKJ]NXx_ � �q��8f�8�p$��e�O�J���gMx	��iBn��&�K�6�(���c�T<�c��ő�&�ی�M6B��t7h�6�s��Ukia2� ���(/����e�n�@���Է&�ĝ3�g�w����F �&�<;��Q�ye~�ԙx
��7���R*��|9�;H�$V޷inp+���>%ƟB���c	��$F��N1w5gC]��u�pi�s�s�'2N��I�	f����tr�ܒ/L; G<��
D�Hm���0ڒt�H3�z�I�X�<�nDNa L"t��U���1��"�Ze��r���*K���k��z1�иf�uK���q�~ϊ��O���0��FP5J�����E��̪� O!�è�㴔�aʿ�IAHIW�* �@���X���A*�ǼMY��[׎�d�4Rȥ��e�`߬�5T]��������P��)��/�Q�O�b���d9�*j���ge�+Wq���7q8��R�A� �wY�����M$ٖ�]z
O)�b��ۀ,>>@�/Y	�*��kb� o'��Tz�Ǐ;&��ȧ��������AŴ�C�O�2Y�42��mU���������,D9p]�D
�o�Yh�ˮ�:��$��	�v��[H9�Xs���%���|�b��*�.[�Jcl�G�8&@;�T�k`qtQ@#���$��J���d���7�j�g6OaJpj��$�h@�!��?Q�p��ѵ)���45;����'�:�%�UxުD���G���Tn	�e���at�`,�I��zx,~�h�w��Ub��"�?`����╖��ܔ�71��ٲO:ңÐ���N�ú��Q bv|�KĪ�y�3;h�H��Bk@vV�X��/�{NH�����]��x9c��B������:�A�P��E�5��@����>lK>��@��H�ߩ�`���Dc�5C��g���� d�����!���'}j�M=.i�6v�YI��C��/f��Dm&��(�pf��g��0�d�f'��P��-�g��r
�	�uQc�ތ�L�2��|�u 9q��9}�\s��r����YyAl۞>����W�Ĺ������%͞H\�6��K��ou���bLl�qo�� ���K��BV<�c�Z�Ƶ��0�����zo�#S!��9ǁj���h
;�9�\�+�O)��An��ф�����6/x@z �J��Aop�|�����W�A�A'[���j���ꄥ� �Tx�R��9Dl��dw��uk�/����֐!fY#/�ȩ��˘�k1�ٓS�߀�Ǡi�s[����Ȝ�۔����ϧz9���5К��'?d6��Vd��19�����C�@�T�T�,$;�	���-�uȦ;�'9���團����ؓM����#G<X�yk!��,��Ь�G���O�@�w�d����JM~�"��<h��m�PA'��JK�5b� F�B�v��0K��=�&�uKCRP�҇��i�ۢq 6�<��T��v���˒9��0:}����`F�d�(�ۓ<k(t����cc���=a����c�����P�d2��*s
Z����kҧĹdikΟL�OC��N��^FW��nl� y�|3��[��aL��y�a���rPɈ 	��;�8�7{���m�ɛKV�9=(�"m0�
����D�X�E��N�ϳz���@�j�\8ބ�4\ܟ��Q����{�7�/��>y_�G�_�U�&hg�3h��-a,��g:����s���� �9�*x�N*hV�]Z�GS��j�N87�j���4<i��N[W��%��F篜I���&a�Ra�`E�#;�7���7e�����'��O�w#5�p�{nL q�ԃO����#?����B��ݳ&�����`	q��N�9��1ۉ/���;��X!4nP��UV)�Nh��>4H��X$s9�c#�e��n��t���F]���B��P<� �#~b1� �{�!��"��_��8F� �t��i��*�Aؕ�����V7�7=87��������v	�!L�3������6�����U���nW��ԚC;�����j��r�a(8��a�G[��_`�ƃ2)�:��Ķ1������������/a���w��;�x�U~�ʩ���t��)�xS>���(+�v�`�hx�c��Ad��2VG���:v�?��`�v�v�S'�m�G�,�`X�>�IV�a�m�ƥ,%/�n�`��+��[�x��t���x*����bCl���:8C��(X��iE����a�G8"�*���b�0�+	��w�j�'���I �'v~l�$`K�'���/�F@��P�~���� �l��.��)�+�J���)�V���e���`�J��V��5!5�%�h� �QN����"�b1��>�������Z��^^� ��}�k���;RCX)���2�7x}���^��7�UT���&�F��d#=����>~�H뿮�Y~�7d7Eք���^qBD-S��õ�{;��F���u�|�M4��c�WП2��,6���w�`�g���<�Aa+o�p`�&T�o�ZP����xoWR�3�͊�����(B	;b��ә͏L*h=Pn��p���Y� ���Z��<�AfEW����]}8Ȇ@���AERVD%�����ϙW�nhe���sMH�7�����I0�>�{Z���������K�}0�mx���_y�k(�gJL��$3�<�Z�@1j�tey�ڐ�E9B�KsYƫ�[-Yl��,圖4Ȋ��Gl�E;6W���^�c�h�����U���~v�����ݷ�!����A�Tl1j�Ե��.V>��;����Śwq�i�n���5Ji�b�9���S�l���� �Q]g{��w|Z���̐GO�>u�N�Dg(h�AȻ����Jaa�r��U�H��z������j�D�):���]̇A�wB�!sǒ��3IU)��8E�Џ#���b�׻2�d^v7�*��/��$�j嵃��[�/�f�����޴:���9����e�3K-�������JܔY��YG�ڴ1���4�"n�[Jq����r�b'/�m��3yb�=A?0ŀ"���D����Q�9=w�f(|}Ъ��ZQ�[ ����n0��ǻ�IFo�K�ʦg7�9s]_M�'��V�7!��X��y��\���6!�H��,)��~kE��n����JeEV��CG#$i��{~Ý��B_y���K2���x�K_K0�7�S�	��BYt行��L�z���k���C�����`�)�	��V�%�G��_�M�Hw����C��DHv��k���|Ů=M�j�<���B�D�"V��mwj�r(�K˪��U@��Vl!�rp��[�#-�zj�Y��ܤ��o�Q7�G��#h�?LV�9@(��NU\О������N0��vW���v߬V��}2��wp]�2f���}/w�t3l}��&i��YX�<vy�9^��A�ZZ�0���g����z�y��!$I��7X�H�ȼ���n{#�������'q�Gu]�ϴA;p�_�����_. �5��>�.\��+�6,3ԥ3؉�S�)^n��E(��Z6	_mW�B�Q���=SH/[fC�''/�'k}�1�2�0�\ǣdޝ�tZCG5��ഺO�x��Z���2a~gL��1K����k�S�U�Ӻ�$�<4�A@��&1.\@YG��%�Н��q��K鰉��mgP�频!�cvѴ����>0��Y4G�+��jݶ�d���&�'	��.�C*�n:l��!!�$�sg�	�j/�v+֢��$Ih�Tssש��r����,�v���&��N���ft�aR���I+0�c;Έ���k-D�6Tp�!x�N�yDHc�GzJ��[,��J�Aў��J�&?	�$�� ��Đ)Rw`���%��ۜ��}.��IH�z�	�;_���%����ߑ�gFp�@e0����#���g�$~��Ā���B^��`S�B!��6���8M[����G�T54����z��q	4��$�R���*'g	{+Df�vP�JܟT˨XT�8u��e���(��d���Y��e�*���9~��eN>5_.��K�Ǯ��0�B�iC��E�E�T��"��t��d&����&���1��l�P�8bͺ~��� ��rĉ����\���	�Ѹ��9�'6��Idꇰ�7��_��M��F���@�>������I�{-�?KP��I�L��Z`�� �X@R�J.�`�: M���	�r��5��:�j�E�;`����G4<��/����U����s.��U`���bΊ n�1�j1x���6n��`�6�`�ϵ���w�nX��D}m���Z<���lK�՚�r���뀱lU�++��5[l�Z�|5�()�~��4�����մU�� ({�%�يO�I�m���z��>��J>݆�or_�Q7D�q�	?�
�zFЅ�W��ٞ���}n�+��1�2f�@�&�Ňa�C�V�Q��H�y��;�m"��;���}��=V�ʣ�6�ҫ���PT+	���$,
ۥC9�E�ZÀYp��|�Σ�>���@U2`�a���V����(#����ۡ���^�!�k�
�ѣ@�c�5�O*��tt|'�Jա�C�����`T�; ?�:C���l��5y9�+az[;�ێR�?�RLR�ʊ�Mi�EBq�]�a�6F�0m��T��V����B߫s�@�Fc~D�7��?et�80�����,��Lږ�O5�>;��9�ɉ���Bֻ��2<��P*e���M�f�|
L���38�{M�ˋ0_��$�������c��L�;��o������f A���i�1f�9J!�������*�<�?�8����X�dh:/�b��Dݑ�[�TIa�Fxe��V�Ϊ�F��I���^[M�d3s�ΟE�K+��/�s����*�D����GI���^�|6ƭ���%dk��"_ L���%[v�E�q�q��:��
8U���Z��C�mLI!>z�=�Y�F d6$����u�<�/�O�{6�� ��]O�4��~�a/΁�D莲��H��cMG*���}!n�x��-���!Vc��)x��xt8_������%��DL5.�8$8<]�bs�G�TL��kJ�O}�v����
61��TK.��Ӛ�q�p�9q����x��C^ok����9�A�'�^��L������<t�#�i'8�l�G��LC�ە�����|��Rk\�D�HrV�1�M^-��<�o߃N?^iT�B����y��"�z�x!);1d�Y�ׁ7���dŃ�/[�L���ȩw��M�t�x�Zň���%�:{�pw!cܬ�&<&�_����;��hw:��1>`4�i��lDS�E��� �!�,�m��=q׉�85�&�_�9;��-P���h�v�=�é���k7�X��h�)@�
X�>�ε��qa��1 7UP����S�B�VE��o��,�9��WQO�����[1nvp�|i�_S�����#Ƌ��u8`vUK��z@�7x���t}le�R��(q�����N���S~O#���c
��zuL��}?���i���Ms?�|'p���-B��Zrln���}���nX'�=��f��ԃK��7W����3E����cv�c��3�s�H����=�)�UmU\!��?�\�G
���ā�f���
s�qZ���^0���c��)��>��S��t����'��:�N��d�Ԉء~R=��D�����.��t��O��ܧ>�a�Y�L,��-.:���hH�V�z,�u
����$l �U5�m��?9�DzN���2_��*�<��J��rUN�D6,Z�#d>p]�]zJ�3r?G뻸UNp��uU��+82xi��*��f���܅�)c��|My]%���P�e`�Eq{�6N-�W��*�I;?Vӫ3��nm8���D1��9��k�$���%Da�GgKA�IL!�bh��.��q�W�$6�E���5z�dGx���$�� [tǫ��k�u�E?�F��K=�5�m�F�z��m!*�| V����M��硜1�Hg��S��o |d���̜ �6�PQ8:�*�*]������C4����@�sp*�&Tl����V��i2��	kr�Z�E�C�=���+x6��;�d;� ��� v�fX�[9�!���"�b��_�ȿ�����WS98uRܑ��fd���oѭ?3�	������tf�O�7r��]Ta!N4�g�$s�E.�8͚۠�za��g�WW ;u�3@�]�sFѧ�E��,�3j�κ{\�W䯫�}q�n�X^C�7�Kv�W�{~�jJ�ؐ]:R'��	5<��ဗ%���"Q��<;���$s�N@aé����U��R�7�X�46���;��%��~�Q,w
���N��_[
&���a�,^����D�2�]m��4�9��r.S������.꒑��r`_m'T����\�J��"¡�1�N�J~椦�yT4�E�-_���^����۞���B�(28�"u�J;��1������""0����(b��"z��|s�;$D�
Q	�G��Fl�q�֕+I�PD�M%�֧�5~.�w�䏸��$��:҄>��By�Co3����㷻�,wF-�Ԝ�-Ҁ�O��mo�UA!Yޚ	n���d�ŭc��/}*��R3kI�ѭ��|Bk�v��P��eE���6%�P}�x���4bӭ<j��U��8�*�(��d���D��:)aД�����PQ�*&-a���kߊ��Shd�wt��3 ������B+T�y��	��bP��p�5���r�Z�_�OG��ThR{Z+0�y�n��ޜ��}���+�~$��|C��S�簔Aq]�yH��/#4�[^�́���H��� /:��whU@��"q�X�!׶���Ck�l_<NN�d�o��x[�%p*�T��hvv�%e��UZ�g>#��|<���P��4�2��H!.CL���e�M����ƿk?�F>�d,Q6�Jcpo	ݲ�����O]*��v�. u*,|��F�K��%<o"�Hk�f ���ti��� ,�ctRMFc����̀څ�2�Q����na\G��C��6����"5�&�+E�GН;s"��eK9�ç<�%׭~})���ݞq�<|$�и#�T��⧓U�N�ᘔ�"V�����NR�����~lg��<�evޜ�`C����L��A�
Ypi���$� ngl]���nY�h&�!���so�u�Yg�V5���d�H\Kiԥ�-v~vl5� D~��ͱ��औS���F�R��vzF*s��"�ÁUQ&׏߆����J�%�]r�+���BoV����m��G2���K���wdX�ey��� ���W���A3���W�
BX�
7�[~�{<w�|��P�
"L�8�d)����u�<�@�$h�鲕c=�BҮ�+
L�P��zsds0u�K7�(�)�uU���v'C�.\K��R�|���������]���^]�c5�{�L& @PA�O1�*�G��}[��75 Đwq����NI��p��B���p��^�}�}-�ʘ�GL���Υ���ye�Ί�.
���S�w�[E*���>MhC��ߟ�k�r��^�=���&���^v��n'��mD���p
D��t��6
6g���gG�&�ts�����aC�� �~��>�ql'�qK�ҽЋ��<�� ��!0��}��5>m�σ�fB&S�j�5x�?�%��e�T70M���&�=0��S���!C���"�^��8���d����*��������zXn�OqX��pF��K��w�/�1��3�\ĶfD��!��zg,�X6]��74�偓��W��'�/�BAj^	�땶�� ��&�(<fMy��V���~Z��D�;7�Xl�m��w�3��ã��u^�����f�=�TD/���{3^�]�:��s��t���$��@�M��2�`�<,�I�i��Ύ{�������5�4��w1"b�$�'`�����O.���袋#t)�$�'�tp��Zӕc��GKt&l�m
�H��%�$�#��a�Cp3P0��*��j��b����-@�����t!�ґ���j�f�������gf�SԖ8���*���V�5kH�Ҕ��Mi�/*]��7���E�Dè���0ЁZ�����i�E�*�K��Tu���v�N����@+u�	�n 
�#l���&֋k�f�S~�5G����l���VO��P�c�=�����^�#rì[��t��Oy٣�*���8"�%S2���T�������j����L�z��YiE��wr8�~I4��~���jU�4`GcqR4�Jo)ɬ��&}����Fؗ
>��?A�ż��c��Rj�**,(o���(b_��sd|�cj��
�u= ����#v tJ���W�I�"��t
KޯЕ��w򲞧��ܰbMڎ������������ ��-�w=*���)���S����Ը637S�牸r~����Ɉ�Ǟ��};�Ptp3��o*x����^��!\��H���y�
��ւ��f����6�r��LX���K���<���:!.��[]�[��`��_��M�G;�%3��^�1{�.�Ӧ�m�{UA�ak���;��"��h�D��Ŝ2��H��N,P��o_������~F� G,�Ui�
.�����l>������^ʃR��uI���<���VB����:����� �� Bq/|�Vߺ��]�@�O]��[�'?�i�L��sE,��AH�������gazt�TmMk�t�.�lXp&��d*zjpB�{�ޅz�J�?��K}��������8����b������	Xq�Ë?��_��Pl���.�=�|�~�2�q�-qQ��GM��R����,B�"�6¦�S)d
vNI�}uDgVBCy��t���3��)*I�GИ���F�����jH�f�ut/��L�e�v��A��6}��w���^�x�py6e���B�x}
%����=j��~���1��@����!(���i!Tb����n:(A5^Og�Տ�Pi0���Ky��%�<#����W�= ���8��>�'�-n�����[}E+I���F�{����߲��a�'���w��_�+Q}���]G�{B�	իƋpF'�|&�������Z�m͐Z�B���H0Q�
 �(r�`����e�v�$o�#��Y�U�Є�~X���a��[��_�Y�wc�|�)bT:M8l��$�O(��BΓ�-�&����ߖ���|�sZF 3>�����y�X���,��Z�X!2�*2W=/w1}B�:����E��KJ�����l��}��!�:�3�6�r8�eXK�c��^����L3H�ۇQ�l!��(��F:���k�l������.�n!s���;��a��r9����NY�:�� �j��;�$�a(���ʥ�^;w_�(����yB�*S�V����R�.i���T�{��ʃ&��yR^{z=B��xIj՞����pZr��p�ge`��Tɗ[��A�Q�̝�On����p��\����k��a(�A��E/�M��%`�vVT�Ɇ�/3����Z�ݱ(��`ԀJ�V��a6��!,/}��N=;��>�ǔ%�$D|)W:�|�Z�3�E]�3&��,�;��wT�JǛ��Y]%�"����s|!�ż{�*$>�畓ߔ+9�U%4ҸkW�n�}��m(m� �n��S!^S�w�,#]=�?FJ6x�/�0����{2�8Y2��Ϥ\��x��E�N�J�:kn~1�c�ሻ���NT-8��T�s���;&28���.D�F���t�h��3�쟗)%-PN���eܚ@{�j�2�f��!,H��UB��m�^�"�c�p���<lQrP��q��J{�rc�Q�0,#�PW���MF(ȉ]����������n��P��7FL��8������p��$E�I��8��Ͽj�	�G��6�)e�̃
��.��hh��3��9�H�#��x��E`��Ώ����޳:.1L��(�(��¹L�9x*5j<��>C��m��>��P�LƵ��B�
�lW�se8k�$aƕP?�
��t�BA*��̉=�~:P����T ��lt���4�a5Y
�x���~��o<�*�F@,XQ��UԣKD׍5X024�eYo��ŷ��r�~�1�;�����a��\�uwKB��Q�iw>�t�s�2'L�R�"e� ; r�@���,��qa����pm�����Q.�1����JW�$00ξoHQ���B�r:����-"����H����o���XN�"���Е�Uy0j��K&��dS_֣�zK�.b�p�TG[C�fh������tx�p.?e;�^f�5����F)�;�����T��*y�YH���?�{sσd6;�Pd\�/,ie�'s����d�Z9�Ng�rd�����)�GH���çS���F�����t��G^���$}t�����k�{���<�JoB���F�:6�
1f����Q�N���w����h�?Z��,k3-�
�����g�T�g���a�Ey����=�x�_RcK�46�G���ZϢH>����=)�o��=��nTO�%7�0�R�k�3��Յ�ˎU�lY���z2�љ����ۨ���	��Ci0N��pY�9F�W�$!j�����X���8ȸ���'��c�(�Vf�{G���H��������j�y� �U.�,��H�Gh]���e��+�I�EڧBU�qv"t�9%ǔ	��f���+���"�tYGgڸݨ7��s���W�JT��R����_��
���@,�|N�;����p��(c�·��1�vnT4K� *��}�Q��t�����(B�Wۉ�G�w�>G����w�H#145ҏ�KXB�%h�����Ȕ���<�$����3��L��4�j9
@������&ce��#�lQ_��I�w>Q^�����G����5��0�����B�F�_�j۞?��j����2,.�r
i̡F�rM�4����K;z��&6&�W���v�<�>QJn��K�~+H�Dr��w�"�[Y�d���[��P�3~�+���k'VJ-	�>�q,a-3��I*��є*'�Qh����".��.f���­1oO��89
��#�3���3m�6�۷�� >�uw�p5���"��ʨN�
o��w�(7�.��.0��#�p�j�CM�# -���z���%t������(ůs�L�E�r6{ �<r|.��1�J^��r�%�X��=�!������D�Ω`H}�J	��.�%�N�4 ��}��������1���qWAX�Y��
@�N&��~��}c���Z��˲C���G����±�,�&����G��QWp^)�
*pC?���h�d��~j�$RM���{�fvN�<�ӻF���"q&���X9T��gׯ��*�c��0.]P�_�b�y���=�ԉ�K�.E��;P�]/��L,f����MW<1eG�m��V>S%�i�b�xd��!B`������2��G�.7A*]Yx�M�op;�O���ݺP�R�p �\��o�;p�`Q�}`@BL$�=�q͜�kǊ�j1��F��p�xe�e�^ñ�0A�nG�*��M�k��6X�g���8��1�bM֌WyW�=�� ����Ў�e=b$>���:A#�H��4���e v����]�lYL�1'%a��hIn$*v%:?����%Ϭ8"�w������[��:3��!��N�>�~Y$9!�o��fv�Քd�i`ı|�����V�z��|Ulşk �&`y��l[�b��0�Õi����h	��F�)��; u0��sR#�[Z�h��1���wZ�j)��?�L"��hl|.˘�~G�eIx<���M�pl�Y�~��?5��܌�����-B䌓�H�Ve�8i��L�����-�R����#q�f�#������Y��9^�<+(��ɨ�C{�Ͻ�/�UĴ�X'��q����]�K�r���u�R�}5c&'���֗}ux.���!�e�T.<b�W�w�1��|g-kc�nѲ6y"�Wj"���n~|�����m���Z��w f�m������<�oĨ��C����)��>�j�c<g��D �xRe���P!�D���9�dL������m{/�����]��*�O�6�a��@[�f䗽�^���f��-tB��&0@���aD�%���
)E�"b	���4�]��&����Fl"�7����Ms���w���:��\�`h�I�&�ъ"�~����׼��#������4���Ra)�=/��f2D���t���0������! HҸi9a��fX5�#��X��'ϟ5i��o�:1�n6E�*20�,r�h*	NO~;A��,��u�&��9� tƜ%����R��=���g&b�Kb�$˂=��:�ǃO���~!�EDF�w��at�;�G���!��%Ro���z������t|����S���1�"<j�׃������E/�[�MZg~��?#����5�Y?H��fC��ѿ�
E�2[���-�I�ڗx>�`t^�J��mk��������e�7_���(�nUq!������Q��.�L>F�����ol�n�uK��V�Ni��G:�Ӗ3!x���M�܍��2�k���3�k�ܦUu82�g�
���M�@����r630���N/9��|�<	{����-p�Ok�B��*��/�"y�%�ݫ� wQ�P�YA�D~���ƴb�a��r�2��f}
��y��PI��nzzE|�sc���Ie��Y�u��UTi1Ĕ�K}�1�s���]f�E+��
F�ғ���sl�J�#6wX|�x��:�"����36��cd�D�qbAd����'4|�ZK��0!qS�K�3T�Ov�vH/�)ʲ@"kw�^��������7kv���d^Ѷ�,U9ou'�md�s-����G��RC:�h �?A�2���/ ċ�_)�1iU>�f�ܜ�P
�8�D���KS�U��%n�)��c �� �ﺕ�:)
:F�.1^�F���fS���3��S�|�rF��Q(*qF���m.���~�)���M�9�<�O�����{�7HIP"�y)3�p��b��!>oU�R���� �0|����\$t�{E�8���7��S��q�o	�X$V�����t��M�{�I̖�8Qq��GY�K ���R��Cof�M��\�w攘��� H3ZM/�hu7�k��nZGɭ4#6��w�F�0�/�u�����Jȷ�~����x$2M-�̞�l}ٺ7.|��>�5��"%X��zv}�J$"���D`�/6�|"���>>��9q�.O|=�9��nrE���s�'i�Z�>i/^�	E�x��l[U�d�U��0���z>j�w��_ྚ� 4;�Q�Le��@��j(����Dt��@�dJ�`�	�#�!����2O�6�E�3�_?_L��N��Wđ�('�0K��{K�(�QZ�
D�Pp��rz�6�}
 ��\�:BJ�%�g#�ڧ��7ޣ+7٢��ܶ�w�6�P���;�ď�������W�V�T=�?��T���xp�6��^"A�aƱ^�3�S�[J�����H�k��Ou��Vw���:!N�fi17��,��ߌ,�d�}�"3g8QG��y`���}��%���D]xi~�0�����{DꟄ9}�=���d@�#����w����,!��X׷)q�@��^�Ez�����~<T��x�� �Y̬�
c�lG�*����E�oֱ��
G);R�`��c�p6I;7`G`|5��7���J�Wfq. �G��4�C>]y����׏tS�����#�������v�P���?�uf��ƫ�b�_�]������VuY�'����":?�#��(j+֓��E"5�N�1�^�2nd{�����urѠ>_�5�{H$*#0�H����A
v�/Z8�t3������m:�r����
)�߉?��}ԇ�ܿ�`K�ւ�������}]���A�GϫǢ�Kv�b	�ɷ����e�կ*� 
iJG�����e4������\�ԅ$��������"����үJ�#t��DTg|)�(_U��!U�2�vz��>`A�~�@jq)T�t~�|�u���W��3��&��H]�H��Ey�nOuE_F�ݠ��ږٰ���<iLi�e8Т'�|�D�ٗa��`��a�$��\�cu��վx�K��E'�~��_���G��'�9���6]�`/�z.@����(+�i<u����'�B'ӛ�Z30+0$���6�RU����w�Eg�W�l�\x�\N	&�xo܂b1�Y��CĔS�|~Ӷ�RF_aBT9����rU�����BL�ߪ��x��oC�Y�q~
$F��{5���J�	�����HW�&Q�Y�]�Q�R�!%�����7}��s\�"��#�ۖ��~*�I�a��3�]��F�k!r�5]𧱹"��?d��T�wrϚ�aw�	j�1��D�x|���,ٷ�{p5�*��či�	?]~���s���'/&����iŌ�� �-e���6Z�������~t�j�뻢��X@�ӅvO�j�3ꏙ�����cNG8�
2W�6b�1h)OÎ�;�)��� �}.�U4.�0���K]�$[�eZ��7���u��+E9d�x��l�(���G�a�xp��3�����l'tfx�B�������Ek�m�(L�W��S-XC��ļC8�� �)��P�܄��O��yo�����:���zD��d��&�o6C$+�!�w��i�%��`�zd��MoӿQ��ʍv��+�S�U��n�ięM���|�9rGX��7�o�xS}����x�ԲNr`Ua�(���yٺ��J\�A��@],�/�B��߻?�C&b��%W3̩�ݭ9��\IF������
(���D�*܅1⑻�̧ܹ�Lj`���)���Lr�LӚ�g}%m��x�!ܴ�-l�,�Y��F�?N�5�2�_虤On�v���i�.6E>j.�������M��ډj�@���X��Մ^�]�M�*ih������j~X��Xۢ�I*i9�O�z��Y��p�D�ƹ�ֶW�Ҳ�=tN����!;?T
ZD=e�\�}-1Ϧմ�ׯQq�p�O�E����S��?��LK�`�������%p"���u���J�:Y>�x�Dk��kFW�ߕ�x�έ��߽d`�&�fHѨTۖ�2��y98��.��L԰�p/�TG�lm��Y�@����Ld�G֕��tۭ�K��i"�?���Kb�%6t��
��/}{c�����O�:ػ}�ao�#���,k���`_�R��B�m�+i�0�f�f(g�!��M�4�Y�k�os�;��S�sV�ϲ"j������ Ga㜧�u���2��`�/�M��k������ȡ�Y+vgŕ�AS/��������s��zFW䍂�U<&%�6wY&0������=�3+���i�nŋdj�#鍇�8��H�'�n��j�a`y"���G�,E�s��oLa�����W�?������,�vOY(��>�3�������1+Έ 0�	�;���,����w2�R���F�L��Y~��䀓�F���H�Z�E ,�{H���0��7���9�L
`)Di� �<��`���y�7_/�����@���"ǽ�эXF"�5(���<�a~v�/R
���B��1�u�?��ܨI32���7&�U�4.S��q����J'?�}� �ͽ�&���&g�G���� �IO�i�@N6���P^��L3��<�p�((�;�u�c�5qL�_ZR����T��2�:c���k~�����c[��<��.͐�'���8��5����/�-����éE�8��B�&I��*��Q�����.y���үc4�9iǢ'��=�8���x�k)��������:+I��MD�����iJ
{��O��퓋��8��ѭ9t?",R�xL�u��Y:�;��ͩ@[�E񐾧p(��x���*�q.�����>�-<2�2l�$p�����C��p�����]<^�<��L@� �\AmyĘ!�%�]1(0�Yk���\�#b�U����`�<o�~�';�Ҡt\"mf�@T`���|�;��=�Y����}�t�&�%��w[B���z�m��p�j8��9�ϗ̺��N-fF�r5ISEXE��,a��Ad>P��FP��2��?����S[��=�/�@I]@5��Os�t�������g����	�����/)�X&)����eqAN�LX�6	������E�#U��ew��K�.�l�Mְ�N0�����LZ�gbXB� e��YV��G�̕T|1�׋z�;'YzO���
i����)�&1�_c�%%��R�������	��1��^|t�k!;��x��
m+%9�̩s��i�hX�RI�Y/ŗiP0�#�r�B���i��Db2�#ONZ��d>�g�dn���LW�����`TK�N}�pd]�� $��[���W�Ig-]IN�J&F.�)D>��k��P!�H��_�|�G��D$�8�#�Vdlh���fl.I�d��/B�8o������$Dp;��ԙM.����o���f<bѐd�(!�4��	�{����02�c��K�4=�ǧ=G�phs���<��:���$��ǯ.A᠖��7�/x��sg��^<�=�?��^�;�.�U�`�ycY>dN���K�H�'ꏞ6Lk�&ߗ�:F-�=�_�ą[�_�+{��^O��V���aw�E�c� ��WT�h^C�k���m��S�c��:l}�k
 ?G�� (	3g[CLk�2D��ֶ���$��rw���=�\[�r˟~~v�-:�����(�?�E��lz�k9�ӼjU��,��LG�@� 2n#W����p�zk,�}�~-��qn�������@u���%o�LJ¯XY��w��l���'���31M���z��7_XImms��Xb�9,(�Qpia�J@����W��j��c���f��>4��)���ɓ`���v�#�N?v;JE!Ws��T50n�l�d�J�w���l�3�>�T_��1�P�9[��;�B�F���H�f��GW�Wf&xhl1��|�:|�R��Dڔ�=��@���V)��1q��QH�dɭr�b�~F�L�����C*�.#���+@��p���� 6�"3�j�jX��a����'�EI1��5�X�*�&Nd 
�d�4�@�S�(���՚fEqEi8v�W���2�.���+�TR���m;{��޷{\�eB6H�A�v��������J}����nE9��b�R��9��/-Ay��;�Y)�c���!�2��U�ӓܐ_+i"M0Vl`x�߈i���Z�C�(��Ǘ}X�σjw�(lC�j������Ƣ��0��. v�e4ۡ\�?_9A��F��ص���mY�o��9��W����$�l7k�\��{B�\��I_^��_�%¶��� 	"�g?�*�SE��X�MaO�ra�~�\�	xὀ_PN
�8*ho�)�S�9L7�'���0M����]�Oz��$�I����	�k����'�澜�2'�xV�~���A%�K�e|�(7���kncyπF�Ӹz635 �R~���Wa���`����}G����e�c��|�����)O�n�z�<���> ���� ��~䗵�8�"`�'S�i����0�����_B�e�(/��>���@:�B�u�u�'��nQ�AB6�bgި�Fgj�A�A#��S>�2P��������9��Q�h.�U ���a�U:ҵ�-��1�.bX�?�|�a�o�pnQ�*u,p�7��2����DB���w�.���f4+���l�$ؙ�)w�J�x?L�"��]`���Z9��^��Գ=�B���AbϺ�uL�ۅ�-��qAp�زʫ�ո"Ӄ��[#�[ҽ9Ř)���J/=�t̓ɿu��,/,4���o�Y]&�)	;Y�}!��k'Y�ٷ�� dǣR>{���:�m��H�B��vD:FTx�Z!�v��`e{r���ǀ7p|�?l����T'��P^g��Ob?�rK9��M��wN������@Jh~��'�|m�+�f9di��;X�O�K�k���g@*.{3�Y��
��r�� >U��&M�n���rR �
�oi��].7W�A���j�!�co��`���y���i��ԛ�լvm���{�C~�%٤[�0���?G��C�ه+�ud5v�.9ܔ���O5LZ	%ݺ��[ �,LC���9�%�>�>-}�(]Q���FƯ�r'xI:�6T��*7E��퇖"��!����,�u�WIְ�����ǿމb�0p��[7#[c�BW���r��M�{4��\���C�0�T1֥�u�(�qǽد,� '.[��C��1%eѕo�.A �-Ϯ
��qhT��>��A����n�ߦ��M&n��!	^��2��C�=�H�o��ZM���R�������bE����e:H�v�+Z�c�Y3��e�P��� 4iid��[9�Y�8B?٠[��@)�>g}���Dp�#���D��|blPo4���18�:L��톫��~�xD���#�1�ĵ��h��q��?���pC�Za�2�.�P3��z��+K��l)����+�>� �G��K=�hlB�k���S�,��s�ӛ�&�^L�I�.^3�nx���1�o�:/nn
��@C@����[_؃�g���T&���T2C (�WQi�
�IUW1dU/E�f6�s�\��d�<�WW7g'��O���1����|E��+���*��9�JY�^���ｾ�[`z������w��@�+�y���m��ʔX���@|��XȐ�:���w��]I�'D��c���<��ڶ�鴻o@x����4i%�U����F�e ����r�O���� 9�￶i�R�.�4Z�o�eb�M#?E�a؄/U�q�!F,MR��c�_��qh�t�\�}u,O�4�r�.k� ���z�V���Ѿ��cG��D�&�#0�ϐKej��i�e��V�l�Q�񚡿�:d��0�at)d��qv.;���q��\�`��Q��Ze�Jg�@�t��Q�a.�������t�-���P*����)�͛���yy��+��T���c�u�b�����SQ:{�S��Cw}�T.���-�S�Σ�Í��Vn�8�9��ǥΜx��ϴ�!���uiY�
��xJ��c�!�eUl�p����j$���;������V�d)|'i���@�	�@�C��'i�2R �\�O��L�i����4C�*��qWݜ;w����?5�,�-���w&V��U��wzR�����*t:����AGХ�?K
S��Y���_]�*-�{�3O�r�|n�x�ru����7�	2�𺿋��,�p���u�G:���3@�DH� ��K(�BAr�g�R1����$N�@�K�},/����-��2Xk�;4��`�ןr�����|������8+�]$������[�P�&A*����ŕ!S��Lcqo�OB�Y�"�GJ��(3&�?RTS=�w�0r�mDL���Ĕ�z�>�O�����OC�:CXӡK\&��4��/�>ger����e������m�B�֞%J,�^�8�7�^ّ?�J��0{��Z������a�%O�x�bt�ʟmX��=>��
g��PH[HK���zQ�)�hBE�G1��rw��65�us�m.�_�� �I�B�b�d�&���-J>)Gcz�C� .]ZYxU���+����+���ܶn��(v�q:�(װBOo��OC���ba���}�f�nHL�վ��අ�V1�ə�Z�>V���~r�I!d�2)������f��F�3����}�l�,�8��3���n��~�/]˓t�o]�-���R
�aQg�L�#	�<�'�����Xy��f�E���H��鮰�z���C��r���fw��O
��� ���p.��޸�^�w2�7W�-�����Ҵ�2a~e���eu��?��Lk�XwXQ`^tS�v�<ה�[�F"�f�&��D6伪�2�1Շ��veKS��G���"�X򄥖|1�Î��q��Ї�j&!�q�e�F�CօC��=��=�Hy�·Ŋ5���S�aJN�wr�Bh}��G���ď�:�\����d���J��� *ݗ�y��L<W�?�J4�#yBvZ���w�8Cܷ�rd��:}����m*���?��p�7>�KR�q+J�}Ͷ7 �{`wX�� G�!x���C�+��Z�e�k��dia�Ţ�kC���l�a@���AG�)�%��a0�\v�3�#kvOZ�� ���>⏱��S1��4��i���Y.Z������2W�U�^�y�3�Jf��ҡ1��z��-��N�X?r�P�˂m9:|����Q��O�,j����W�9��E ���l���(�L�"ؔ^��ŭ��-%K�Xl�����̀���� l1F�D�������(Ŷ�W���>����@w'� �,�(��r��v�,h|��D�֢��dfua�yI�	aSf�o�M%�D�x#�9ږ��3�_�N\��wƓ��@�3ol����a��ŀ�'c�=t�sk��u��_$7t
�Q �x��O��<'����PD8�0�D�O��&���N��=C��@��߷tX�*�5��xj��ax�����@ѯ%�{�˂߀��}3�X@O�?3�t1��@́3eN���b�x�z�.���'vؓ��.���27�M��Nx�iA��YpIE��0N���`��۰l7���Y�у�W�,���
i�ګ:���ـo��5�d4Ё��\��(ɤ⊆iA�C��_���44�U "��.-�uB��� �I�|�%��5@�MA�r��f�r*���\t��<��������	�	�	�)���qs�,�ե��m����!H)����?Wn6�[� �lԃ��"R����d���
���1\�Y��t��O����*��^[�� xJ��\8�^;JX�י
S���~0��n��_�S73��w�E��b\�N�8W�����	c��������JK(�OW(2���9o 7�o��Y��&���9 ��9w�?x�-�����/���HƜF���61E�#����ɧ��kp�/ހ"\�d>�x�kO�xz�o7,�ejʑH:@E�⭲���PD�?ʎ࿍�`�g�m����s�ّ�Sk���`�pD[�G�=S�2ໜa�ے8���X[�<��ڰ�v�m��+ϰ-zCEH��q���r+���޷�u<V�E��*&�K�C e^�TS�ki�!���%C���SX��ZU�\����]�hyሌ���ў�f�
ш'�����j�|
�2�lk���2�:�i
rI;;&���=��� �	q\e����5|�WJV'�2�/�j��M~5^[0$��W ���c�C
#�zd�*'�ܜ`�g�.�^q����RU}�8�x�zF�>��}5�`����E(��LI|���)�#OA��K�2u_�4��b^��<0X���:fk��P"����Zg�W+|�׻�C4b�9+���iLf��=�\��x���ջ�������s��� �:�z�Pp=p��i�����WK�G�w2������G|�����d���t끜3����,���`[�Y�J�-/L3+�q� /d���
�$�FSz�5�n8e���*�2�hgp����j>��h}�t��:0��5��>�5���T_(Y��&�J̓��J�A�
Ye��GsŶV���҈fݭ�閦(n��L QlS��9��@%��B��
�=���,���Hj�9�e��
��@a�͔��-�W����w�y�Q$���5[�
�&�-��5���6	n��~�N���oh���w:��%�������5t�U�d[M�.T�����R���{���ksk��!y5��h�Z�
�3B�`��6��Y�L�
��l�Ul���F�4�a��>���W&F��Ĺ�<�r�]� n��Ʀb�%����bɸd��	�|���$�o�K��(� �4Mpy'f�R�3x�M�Benp��L�}K�;o�8g}TrO�V�sgV�a wP<i�x�|S	^�p [W�P`��7�w�v�J�<<�GeD����Ͳ�ȳ�ۥ���`����ξJ+~y�o�=b�t=���u}I���LXa�y^�}����#�h�V�IAF�y9�kO_��� �����. �U��]�O�6�\o"��v�����-���.�S���k�8�:!|�߱wm7��Ҍ=���u�:���P��{�p6�F��k�N�Fy|�����㵌�r.�=��b8��[@�#-e|䭲��%�-[�/԰�۽����թr;�/�M=���:�68sۿ\�=�BT�,�H��I�� I"F��Pd����R9{	{Q��l�K�m.�7�ܳt�����*� �l�x�]A@6u������W��N��W_O^_�
J]l�泐U��V�7**�G  ��nD�P�Ӄ�}X�|�m�㝵$k�Gx�Z�+��zKW��z�`��P�w�����!=TXV۞�C��=1�1�?Uw��F�pL���ݒm%�	!��Յ��}�9A��9K��?���ˆq'sÈV= �z������jѫ�@K������Fh�o�-5�����L#����Qn�J�\�$}.�J�,�;�e7n�_������eAZ=B]9���� lkN8T��`�DepX�,�D��6�H\֬�]�_)�2Gʑ ��! �SóYnl�-��6�s-lSm< JE���?�+������谭�����z�$��Fæ��b2�=r��&NY�w캃d*^|�=XS�tfcMxaO�gբ/8��tr�G�<4�G�^�:��Yq$z_�3WiL=����Z/w�׳��u{hg��{y��H������t���~i���FLyȮ��\PP���T'{���id�i���G�&�D,PU��zK��0l���ۈ��n}���;&I7�~D�������<@"/���"
���ktް�u�0��~Y,��2�-�Ռ�!Y ���n\�Z�^N��k2�pJC�iB%R�,J���J��wC�Ʒ)��ώ.,��	K1I;�A�e\R���pxZh�E�K@j;���Ω�3��HR=�yjhLsk��Zsn_���B� ���k����:]�ܰ��.�cIj�����cF0;Γ�]���&ؾ[F%c��Q������d���?����LpQe���W��^y���]D����
q���`7U�ާ�g�.���0K&-Q���6B�*����A3x>�`���X�O�GX��������k��]���dۣ`&_��}c�D�y��l{�z�<!F�r憧 $d���N�[�%�8�p�Pd��롒T��5��Ba?ܣ� ���r<����&�����~�����l�tb��e�ʲ�,v�!���4�F�hO��~kѿ����h��x���a~,x���b)��������-P�z�P-�b^>IS���̚�r�:�1|�Hs9ڂ$�=^v�frOT��)��熔�Eu��d?z����k���=E�%����
i#-#��}B���˿9����w���s��;|�U��� +�X�׌#3U��1Ll=�C���cZU?Z{�PH_�O|Iu�R�3;y�$�(�z���(�	̐�Y�;��`�ޅ�S�p��I�E���62��!X���)!�)B��)�"����.�f�|1�O%�c��$��;�&Ȥ0ʟL	@�T/���4*��9����숰�{3��%�$�� ��g��	�c.��� y9r�b�>so,Ugj�%��W<w�3�z�"$�]2�?��
+-�-����O<&��۶�Eѷ�rZ|q��7��ۃBB���!�����eJA,>�{7�ڮ�p"r�Y�A�Y��[���'vC��OH� V���c ��`0'��m�9|��3r�5���Zє%ܔE�:�d�wY��j�,	Lxh��i?M\t�G�d>�N��]���|�<(g��R� �f�tIň=�vM~���i��{T�������00R�ۛA9���t8��w��<PnH`~�L�&����uv����#�8-�ך�c��:�Zx���"5<�c�:����B:K΃7�_�z�3�V��X�?"��`CY������jKݔ����^��>�DJS��JS��U�	��2v��g�z���Q�?,c�{�F�OQ��Ò0ؔp��ɴ�HXSOM�}�S�y�#�<]P�hB������������	PyJ�I?�)΢ӣ�/ȍ�<�mcQ��z���[���cyJ���i��|�M9M�U�e`����
`�{�'.�r|�~ ש���̗I="�d_��&#Y.���=��d������o�`�3�sUb�2��V�+�0t2*k$�ٗ����3-Ř}��/�8�ޖ�M�P�'�Ŗs���=�#R8Q鍧^�vv���1(H��=[""��h^K�!����G}We6����0/�F5��+q�
�Rd&��$��y���� �X#�G�@��UJ�l���;�1Rx��?@��4t�k����|Sٳ��Zf�w������&��!	��"5I�v}[�ucƸ��<���2ت�c�6���N�f�h��]����`B�[���'��C��KU=���Q��B__ka�O,L&J#��kV<#}�boc��8�y��=F�r���Af��G��t�pA�@��Y�7оH4�h��ʁ�)��|�p6D(ߍ!����"3�3�%�5.N�|�0%#e����)�3��_���W5 l��Vf�q|���@�׃��@���`�����p��oH�\7� �ꖺ�{�������~���`����n�T�7w����SQ����iz[��ky�Ԏ	
t��P�n������&�W5��i�uId3<l�&.[����4��\�
ၢ��H��lQ��*=�]��I�=-���`�H�gdϛ�D�z��o|;	�O�E�ḅ������}f�.��������f60`���i�ԽqW1e� ��봘}�L1{kp'�����b��S6��{�h��3�e"Y��m�W��4���M Ca��z4Z����H�]��R��8�^O�������0ʠm8偃|��e�����1���$�C��$�ֺ9c�ˬ��cviy`-r�	�Y��ٓ.��L�E�F��[��k��	.�,�l9��܋�����zRദ�"g3������p���Ƣ	Huƚ�W�;�F��YfE���ʿL4��)�596�%��SW�ʌxۛN5k�5TF8�7+I��ݞ�hR+ˁ �,}��=���K.�u����D<oe�.��"�2�H[���^�{�ï���(�jX#�GMac 7>�?�}� �T��(@P?��@�cyi���Hp�`�# ��.�o�w������ꘈ��n%�/�9x)+��|���� :���%�,v��?��2a�M_��?=`+����o7���(@�4ƈ{_Y�D��q��Pi���K�Y*b���q�aB����o�9�QFn���z��h� �Lh�b<�xx���,,��ŭ�+e�T��f�v��B�)H���z��ɛ���"�y��4��=�{��d� ��R��P�e��h@�Q�@��/���o����t�y�`��7�j���{!�դg.��:�6~z�S��6)�5QE���qn�̀�J�O���B|ъ�D��;��ڱ;�/]F���;��"��߫T��sr�g*?�׍W���<8�p_�$��F� �f/S..Wم-ԇ�*��^��Њ#�۳Q��8j���G9r����D0�.¥���A����*�Y��Oq��U����3ɍ��Ք���r+Z�@Ł �jH�v��@�5-�i���tb(���Ve����z�$"��� X�����b(8��&���N��V��{�I������ެI.�f_�52NC��pv�����G���Y9������C7�ȁjۈ]���J���+GA=s�.�iI�eKa��r{i��0�7�>C��X�}ݏ��F��v߬�8p�h���X�g��#�(-�buŊ��].�T��z������=E�>����/��zi�!s�� Ҋ�B�2��0ԙ�Q,Ր����˳)��ɓ��	��C�J������+M�Fl�jo��Xd7(��ě7�N/	�v�eXڏ�[fl�'E+�QL������.�t�IOiIJ��{X�)a�w��#m�%EufB�
b�Ua��<r��t���$T���	��:o:�}7#�x Y�ŗ�{�3�'�*+m�Z#��!���$�Lٝ;�5�����/�>�Q���E�lJ6���>� qC:#+Յ�J�wA���2���Ss��`K��>j)ң���2���l�n�m'`������®�V�?��S<���'E����W��lȃ}(� x�+�"ٳq��+y18�x��m�*���.���9���D*�GO	"��.H3��S�6@r<	AYm1�8®�H�K�*>TO<P2��w�ӘJ�	�O�mĎĪ�:�G�frX�A��X�9}G~~��Z�@���y�t?����w�k2��o G&Ay6��g��._KZ,���GZ�~o�F20_�KM&�2�$�5Q�uy�-([��]G\^n��i5�+�r���U/�*���iak"�a^(���ь`��e����;��h^�Vi�Wl!���s�*��u���a���r6	�S���Q��L`f�C�L��q�U(�ٸ���]�5%�e����1h&���o�k�,S�>t�
F��/��0ڦv8��R����Qr ��0À?�,hw-͊�b3�\�)�P��M�E��[j8�A�j,�j�U��&T塼�,u��?f$ʪ��'�r>&c�0~��]c��͟��S��"��tBÍ��UI� ��MP�J&�Mn�[�]^�-�����	��e���M ���=�Yuʊ�����ê���Z�U�^�!���ۇެ���	�����{:����V�IӠF��0�����>�@�J��R �sv9+h��T�p�TL�~��I�92[��y�zv����p�K��+k��� ����*�?̈��������֕]����辻!c�7�hP���X��L��X�Cq��HS�XoGY��q��Ym!K�`�O��iA�pH�������7/��^cy���d[L�~�Ĭ�?p�^)b�\g�z0w�R�ڡ���ڊX�C��T�X ֡2'�w����Ą��`��M��oCwc��K�E���'\G�z���1:V�о�C_�&&'v������pD�͔��G��Ɇ����W�Y��4�|�}�5��s���f�KY.�,�߇��MY�mw�r�(GA�c�/�ȑX�3UFt�n����� ܒ�m����46��s9�?Vs81��-<�7C��v�������'
i��g�v��[7	�e�Ę!���|����Ng�ܟ�s$�����섆��%>!#��\Rb�5�KE*Wu�M�r�q?����/O5@�S�W�$p$�J��Zj�D�f�z�+�j9�ܱwak|K�i���l�E�
�H�u&��k#���_���>k���3��{���W8;Г;g�J ��Z�S��݁�O<%��E�{-qk:vȽ����n�Ģ ��=s�f�)_^x��y�e/3�lK���&d'!T�+��f/q2��y��!4��,�{AjN��A�,E��/��yr��G�*�w⋸Dq`T�'7�Q�����БK�I�Q�%@N�$G�Qb�_�P�]~�]F7:@p�M�S���	���>/����P��G�7��%X�n�C���ZB���	[�����ʃ��y�J��ۿ�<E	��IRH��T9������)��R�>:\��j�J��G�&�7W���긥��I�c�Q~���f����X�xm�H�M�4V*:�kS:�c�\�F���,Zm0�j��~i�����\�BO��Xɫ�^7���>Ϊn������.J_#�F%�R嬹�][��{F=U�t9m����M����P��{S;�qb=Hk�Đ�R�I�a+��@Q�J�щ�J4�t��������:�������ib��o�xd�i���<�i�¦�L�e��-�}w�kC"CF���	�����i�H��ih���<7Ho*�u��S�;D������,>	�د�
�y<�"�����~�,KV=�#����:��/������=�O�~Ϣ���jڱ���9H?F���V����tY4�p�R�m�z$����������4k��Ij�5��Q�-�1��T~��H��J��C���uh�<������3e&nS������E�L�V�c�����)۴B�Zl(n���ha'2Y���:QO�t.�E3��4[�6C\Lg�vjC�������y�;�,�"�˨���t��c:o.��E�h3ki���-[r�[�z�i ��"��q�0��Р�\��Tlp=%�e�w���cī%
�.���T�`a�5!
��:�F�T<��ȦG���(�x�A�&{�{���?���n���vk�X8
NX��-B3��Y��/�6�m+'�w:�A�2��ӾQ
��ڮ%�PVh�@I̹?��s�3<�����(E�F�Z�h���M�������)B�Z�@��5�����S���.�[QN=��x�q[l��'��B������4頋��8z��;�*$���m�(�k߉�U��d��	
���1��$.�{��3�n��z��<�)z���[�R���x�^����� ���pߤ{2=X��W�D�a�q��
DU�	a�Fu�4
~1H��
����E�!�@o���T��Ѓ�#�w�~oĔ����r��k�=���:�ɖ;o,�8Wi
���H����w��h��B�ۻ���C�%��8��KrK�)��j8��S�>�La��&thA��n�R���Q�o���ZW�g/x�vr׿�ݔu3�b>6�Zu!C�}�ZtE`#��	�w/�r_@��:O�����1�Jͣpz��깕#��9�>��㒐k57Y���f�J�|�U�MHj���7������*W9��L�of�e��2E�D�7�0
�N���~?9��I�t�&H9.hJ#߈"O`���	�e�=|�2c��(/	��[D�����V��S>�[�D�)_�uF����S��~�U�EX*�ei�o�y�D��΂��0! �H��x2L��`6H�.��bD���V��`�W�^cZ#�/���ͻBF��:1(��)B�&�㞜�p�~9�@Cj=���(��R�7-�7����#�'����/�M�W+���9n�N��<~v/By�֦h��U�M�M�K�U�|��޳W��N�¡�W2k�<����1&�VK���0�ԝD���_LQ]j|(�%˒]���jqP� ����?*��E������>ɮ��ޒ�۩������,�F�V�G3>��{��SߤM�[ُtoN𼩎�v�!s,�.N�*|���kxV�����l����I0����wYg4�*�� ��3q��&����g
~.Mʉ��ݮΦ���v������ծ`]�U��q���望��$�+yy�t[�
���e���	;�sp�_���e���������L��B��?V�fRk�H�z�l��UyT����$&��	TY�J�dsB(�:ŗ��x�2{�	J=sw�S�-��`�!�QC��N"#dݡ��������2p��ޢ�ǚ�
�ױY�����g^X�$�Ƚ��_2���hA
��Ɵ��:f�~�]���u���vэ˘Aa=��zs���&��=������f�Fh��Ю���M���~n,Mt�4]R����]�+����Yx�7���ɳi	[�μ���<�u~��# ��7� i �����)F�U��KJ/����y�^n��Ǩ,�*mg�6�n3?�ۂ���^K"[��f����O�W��"�=�֫(��ܫ���k�G�ܫ��;���*�I�����}��&����i��4��GM�w~& ��Y��t<l��L�'�M;���c�^��U.'���5��)���-�u�o�xvD��N淧�bg"�	.��	�k�3kĂ��:��њ�`��tQ%�!��u�~̆Y��"��O���������j����g�7֦Rꄫ�N=fR��ǅ\�Mb$^Ưoq�m�3���	ӧZ�o��U��ن�4^�P�X�a��ᡇu�^œ��4Y���*�����]� '�%Ĉ���D�-'aUW�Za�
ED��@�g�D��~�O�Ϻ+�^T���J���(���/[_M���FP��zq�JU��2�j� ���k˵)iP2]c���$\�i��Q�v�'C,�$I��r��a맃�F�Ve(>�s!�lmkM��DC�