��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h\a䖇 �;M�l9;Q`l��-"yݫu1.P�L����ip�ƛ��[�n��)?����]��
�}b�ø�@��$R�
��`^��N�t����x�b��o�L(8�?��%N4=��&�D)���=���[5֊���G�s���M����
cÏ�_�	Imܑ�������P�i�o�:��iI������Y�u�Í�z�:,c��
5\��nbD��<��As��Y{H��&�F(8�Ck�����z���	)��. ��~;��#�(��,a�=��s����l(m[�`��*=�:R�O\�D��� X��a)��#��AI"��
0ˠȩ������<hkc�:~vGp^<[c�L�Ļ?�l��s���9`/@kw]z�f��3����w�D��P��L��O,��(�V���q#�WH�yh�9���֜'S�;�C�jĲ$V�S����2�qī,�SK�T�ԥ�k�J�sqz�E�?6�6U���(����d���𲍦w��N'��=.�)/3ֻ5��R�o�`������зb�>Gs�e<��̵�f�!~� TU��f��qt7���悴��N�M���-8�`�G[�+��X�П'�>P�Z9?:��^�2e]%t�U�U_f�!�͜p��	� uY*��y&B�.����4�j�Ő�߅�������X���
�X��^�N)?���DS�̳d"�z�� �� ��M-.�Xvԕj�;y)K}�}Jw>���49)�w�FwSV/�P�|o���p̈́3OS@$������)CY��ꦓ���ҫ������?̚�$O3�<�!���ۑF�,Ս��I�7�RE9>|%�����Z�_�a^-����.���Z��䱣;?��mJm3��WbU'$��N��6����|�ˎ��_�Fz���y�\ja�E�R̥�ۺ�D��m�E˴�%rM�5�0�Qc��D�ݸUϣ�Q1�w��)�k�>��G�����K���>�����>���,2�#ZpB�ir$ʁJ9��&�G�2V �Ъ+��/�
&��U|���k[��kԘ���w������q�zI_��T�5��BD߁=~��oSE�g7��վR�aB��ECr�+E|����PPE %�ps��?I��1��X���8�J��q�b	cX��0�6�3�o�?חh;2���{.�b{0�)�PC���2�*�I�&���4 ��|T!����wQ(�������8��%��:!�Ǒdʄ���~t}�a*W��-j�����
g>@�IR��?��g�$���eg`�Qq�J�ܒ�!Z-�}��w,�4��1Ί�����Y�7��T1<Y�>�R9�����X�]�5U"*���V��4�Yhi�XuM|_
^��jR�&Ƕ��@��f-&�/��*�T������TE5�_���s�=,�2�
�mH�� HyE>�W9`��ȼ_���	�<6��n|��~O+4�����Dvl�>�bp�K��T�����c���(G'ɂ��]�:��nj<�=��9;!�y�]o�NY�NJ�}{�pj�n�ǃ~����@hd�$}%�(ͦ� L��jq��>�&�����Ti�)�2,�nB�]���㴕[�Õa�om%���O$4�A��
#Et�	 R�F������%�|�=���lW݂Z�N1�����i�^w���c��wI����	�uQ9�3��_LV�a+�(��`F�~3�ݹ-�h�<8�̏x�3,M��?S�Q3e���	}l|u�¶�x��uz9���4R�R,"^J�Ɣ3{�,�R�K�%Hϛ41��A����`~�gQ�(nH�LE�=������?K�(pA�l�8	ї9V�	��J�U��S˜�N3���x���j�'���)`��c�~R$UR)v�g7���K��I7��l��8-1����T48�t�5��7���t�O��(��zO���4n69J��4Y��\�8��/���|�Og��ʑ�!)��o��F���mې1ݼq޸�k{6U��E�-�td}Z�J�[Q�¶6%i)�ω�U�	#�z��Ns���Z`2�
8[҄�:������	-�k���m��o�]Δ�W����3_g�m���ylF:%j`S<ăFO�];ʾp�gm�g��_�G�
�	���O�3�)����~���UA��_�`.������4��eMQ�/�.㿝(��	Wh�哗�"�y�r�'*B�P����[��)'V������-C��=H�P�TP	���wk��͘;��XF=@;d � �<��o��'}g>V���(4 Yj�o�d�^^Ӂ12/������E�E��&ۋT��X@}e�^nP��# g4�m�{��GhE}�h4#p:�{�_�7�r�' �4�_�������5���*F ��[[?B֒߈��<����)�r;++�C'0����p�'1�v"����䅌�w��C��{N��oI�6���:�|�\�;څ*�6G�&���Ze�� �ր�-b� H�(.��wd`������.�}�\���ä&�	�g	�*�8N�5�?���y��!�4�,_�	�>|�p��o�#�2'��}
��.z8l��7�(�3�n_�@�q+�Xo�p�_Q_YMۄ"����������5Ax<�UDTfl����ƷӪ�vB96���l�����	�|V-��v�o
����k��Z���ut1r��6����t����l&7D�h0���	����w����g��n%�y�h{L�G�<fχ��6���� ٙI7e�e/,�Oׁ ��w���C��qz"pm�Pⵍ%�Ow����Jr�=IQى�m��w4׼R�l��,Er�����u�X�:�j#݀G���	����[Sq|�𠏬ڳ�)��S�hrZ�&�ؠ��n$4O�!4�7Emn2՛�����X�{�܅��<`/��H������VB*8�i�ÿ�.H��=�Ƕ@�N�|۪��]k<Y��st��2����:��3i�E��i��gp�&%��ފ��/?�8��:�p�;�ro�.&������́�y���jә��$x�J�����9�Z��b�х�;�iS;�xN��*��-�ℋ�2�ح� �����L褧4۟��@�{�@�ٓ`����-�.g$C��KZ�K�v�O:f��aU'7/��K�T��l
jr�#3�$�u�oƎ ^���~���	8�g�'`$�b֤�VIju}o23�j4li��/g]�O�Ug���WE�0�}Ou��i���~�!;��YG����w�Y����a�SnFJ�q|q�<��=/AsU��Ȭ�w�6\����T��WM�g����1'�A��o!��?�a���U�G��<�|�,Y�\�B����`�p�Y���%����UJJ��{�
Cf�Bi�up��&v���W�A�G:���@���7���b�><@��I@0[��̩Y綺Bm�[@|���H����;(��g�м�T1ܫpi:W�T��t��8���븈�V������ta�v�ꕮ#����!B�CGv�P��~�.��t0n���z<s�� ��߰�4y`qG�(E@,g3r���ޠ��#�3*!��B�W$��D��A=�h��9&	r�t�{lmyIz�,H����v���on��ES�JT���MG�!id:��}��=�b~vCL���-G>��2���up��{s���
^A]F�Mc+�Ee��Ś&���6x�T���}�%S<���v�J��.��������du���GZ\B�~�v�5����G���9��'��% Ϻ�#��i�
�3J�1j��T�s%��Ł����Z�`D���.Y: �*q��wG�1��OÉ~���"C+�8,�+v�qP�����q�#�	A�y'$,�i(&�ޚ�{�:ex|�}��!��ޱ#�.o���M��%�Cŀ�k�@SE���x�tV ���πa�J��B�E>P�,��� B%0��-�.3TSU��s���2h2�rV��c�9}Ոʣb��k�4f�SU��q�
�H�'���c�˿�ͬaU�U��Q�!_y�v��[T��_)�������/$�.�&��-�tX���k�Ç��Z2��M�K�I�q�b���d��e�_M�*�g�e�f�X"���R0�������Yf��F�73����}^U�0>̀7�
�;w�������p.6��7�q(�t�����*�^���<Z*����ͅk�Q�Pu�\l�d.ڇ�ęq�*F�uL~�� ��5�lO��H5�`��`�:F�&2@���iu&�P)��ˤ�!�sT�s�V8'J����U��LZ��r;��Q����킧
�����׫����1f��>X��)��iƀ=p&1F�I%��-�,�'�b}dΙ^�hѣ�����~�j�������~f���٦e�ܗ�Dݦ�_��Ę�z%ۨ�R��tv�E*'��Y��e�a��3��c)��+��m�>��(����*T�ˍQ��(k�k���|����9�a�H�K#�T��~0Q꥙NAM��X����es~�H��uZVSɤrą�:�T��;U�G���|(r�%Pp� {�������K+��>�^�I��Ѥ�YA���w��K�	7Nd��$2�]I�}Ϩ����k��R��Iac��|;��#/��B�\i�7��h���i����8� T��a���!fU��_H��Os��y���{#�� ^B`w���u+:1*��Α������p��5������b�Rth��/p)��ʠ ���͐�]�O�8��β�����Oe$ �Pn�~ʔ0j�h�MXY����"|9E�� gK	��6л/(S��'�)"���E�z�b�0�e`��~�h�t�%��m�*��t �:Ow[��o�ه.�倒I�� M��A�:O$�Y�k�?O?���9�t�7��u����k����Q�j�t���V�Zn*���W�"t2��r��G9-Hʈ�;!�0Y�y�sd������N��[�ٜ������ �y��}��ݿ��}TK�,�khE�W: g��jm��#\q4�_�X����7- ?yO[�
����R�hjݎ�Wy"?yr4�:�[�\�K�Byc���t/>#�o�p`��Zp��4�LMJ'Xj!Ӊ����h�M��3y.-��e���b.=��&�N�;J}�q�"e��]�;A,�b��X4J��q��aKx{��(fI��!�hw�3)��*�b�O�lk�2�l�/LT��%�C����Nܯ��ur3��1�Sf@x#E�ɚ����M�>�}2�#��3�:��Lr�-v��#�>�����Q��Q%�R��d!=���#Z�߷��,����O&}J:L�?m�����h�I���)Ҡl;�@��
J{p����X��J<�v��ie�Z���!�ґ�`<
��W��iN�C��7��������E_���>(|�n8*Q��:@��nҵK�"������x���ao�+J:�?�����:Ik����!E�{n;
�,v����o��m�5�c
��i���UPz�R�Ů���H��<�w�+ckG�J����x][=;<�k(�WH7��W4?
�v�&:	F�3/��#jj�����ǅ�W�)����cQ�&�VKΉ#��Ԁ]��ˬ
�RZ�&��P��8�����ב�]��:r�۬�q:�׵�by,�|8��ӝ�8���6��GQn#"°�3��y����K�!^��bMon���ҙU�k��gGɏ�Jj���̵S�X�$Z�1`�ZV,�����n�'������=�!���	�bz��|Ј���X�]���N�傂w���[�1��9��.����d�o�c�������ߢ,�ʩ�#�nFm�]ܓL��'�Y7E%�h�	���
J�k���������Ǹ��D�P�}��)��:���A��U9�?ޜ��].(;QҞ$aW��Q�An�v#��t�B���C��	��+�3~���$�0�R�w���x�g��Z�!}v�2*�G�HH��~P���kP�V7��=%f����+Zͽ�E7����r'7;�|I�T��9��hif�,�s�7h[Ӭʐ��H�ε$�#(g��Ֆ`�hHW컊���Rj$����T1$�̃�-�0���k�]�]�꣣��	�V�7B�*R��W�4��
�&�.���ߴPj��D>�0@�=]nT�n]Φ�o'KD����`��4�O�����N0 w_��}��s �~q�}XZ�D{C.E1�J���aRq��cQ��=={�jP�w�S����̕\acRu�XP�4�)�+�B�xA���U+h�OX����B����4�D�8�!��rt[���H+�	�#��e�X������}bq���mdeӐ%�*aБ�5�	���i�֨�B�,+��$b�OC� ZIC�;Gw�5�N�q��f�v9�}���}�;�D,����8J��bf����~�ZJ�A����C����6Jm�Ϻ�]�=������ʜ���ٿm3��U[m��꿼!V���Lk�u�d?aet������>��,2)�4���6�}2��w����&$j%�3�\�=�����:˫��,�;�ud������b�\�\f�T�.��<�?Ȳ��
���QA��:��lF|��%i��a��A>�4��`�_����zb��樋N��wB17m�)�Sw����~x���v'��+�!�`��w;M�i7��|4�e��0w��5ܟ��7K.W1 xz���0Y�<���x���ih��I��T-���AB&`�F��tyʨUH$�t���Fq�ac�1���Y%l5��rh|X��X:�E�>�#J�L��ݥt��u�X/��
,��k�s[ʄ�_7�:����$�S(~��m� gk�q.ÎE��	ٜ��l��Z����V�wVU�bM���|e�l����/]�ᩙ�N	�	�:�@�O)�{uz�\���r��8|)���$\�%Yr&Tb|@PX��a��P�B��l�����ޖ�>��:s(���S�"�wt��aL"v���l5?�kwB�n��㸲~�ªz|(��&��| ��9x�HE@@e<
]A�s�j��3һCK�F\z';q�g�Rg����=K���` �G�E��j��@B��mv�y̩~ݓ�lL�� ����8�3�
�y����F�R��7��M��+�%�룍a�e}xqT��\�� �e0lʅ���!��OvY�I�Zo��8�+L6��u��l.�*���T�Z����+��P)��3��퐃�|�v-t�z�)�Y%SC ���p,Ӕ0���f�Jn����S��5�:-l�KhQx�C�"��d$Zϴ=��9�Ӷ�����Ӽ\���[��jD���
.�ײ,���:ܜ<R��"Ӂ�ip%�e=��T�ۓM�����٘���|�&w�h�O��er)��O׮��E?�H��z�5���I�q�54��r��l��z�Dm����,B��h��������l��`(6s�5s� ���	y�\�;s;��Dx�s��` }�4E��#/����ү���8�e�bd��9]�u�ajs/6��ɱ[M�F���7�1L�ȸG��H�#K:��Z/���g�$�f,$wԶ:�b 6wǠ���jY�ܯ��K)ؑ1��Z�g���}�ny��xؐ������9���"rV�A��S��H}�N����4���N�U�j>t5w!9H�cJ��ɦ��8���Af؅=������H/ط��qx��-�D����dF��J�2�$�Xx�-p$��v�
C~#��"-�kj���C5��7�xRl��$�D��@sT��[ S��[pX��e��
d��
�ᚿ<l����ap.0��h�A�2͐Jg��'��S���O�S*����5q� Qzةe�S[d�]���Q���S�T;(���!Q�0�t�k��f���qUܺ���Ղ�L�J5<��Px=�4�6�}�4ϟW6SɏDT�c�͕
���ŞY�3���
��j���ğ��� w�+�LO���כ������F���;9�ڏ�=%\s��J���@BQj�x9rIt^�Yy�&���y>�.ҡ9�nó��!���8:Ep@"��j�����G%yB�)
��݌�\ >��&�^�Qx���3�<D���F�7�D�dl9�nv��톗����i'����,��C�]l��w����/0��!>w1o}�ɮ�O>rR��(� ·`������XN�@H�Dj>��W�M\3}^��V�}�-y��Q�mv������.�8�͝WH�fc�q�bs�b�$(�t��b�&�`w���(��-�1῟��r_�Ή;8�t�nЉ�����Je����2�69�8�����C{�����t�RX�����!��KY֔�Źbi���ɧ��,�-�����{��.�jk_����^��d)Ǯ[N����d���٪�GnS��I:D����ԋd�Y���^²1��t�'�<�nF]�G�%3?�;���k���8��5"�oq֦���Qhc���"�|�6�m��?B�=�8�V��	%����E��q�OsŪ?���Y\��dYt4)x��F��dD�����z3e�zn��̼g�Y�?j�����P ��Xk��g�a�xʽ��`�mD�y�D
�z���+��R>�ے�>���/�����
�(��P���R$?k�W��S� t�I<�TL��;�|{�t�c���Ǜ~���+OH�d�G�m���B V1��4�$��gʑ�#��b�C�_߉P��`>�8����I��vu������ۏr�Z�G���e��*��F2����y1�LCO��ڬ�W~Nщ�mb��"j��U�;�E9��.6�m��_��9�e������q&����P�4�\�y{�Vl��4^4��)hVA�LİUR��ρ��P�����/�1J�ӷ�u2����"�3�ɜ�*�F��N�v��S%�2։����1������g�C	���z1 �>^�(Yw|��:d�
x9�oT�q���'��[o�K �� +�ȇ!;���oT��5�ẗ́�a���+��}��鹭�'Ͼ�.a[Z?!-�ɳ��qηw�lFg��<NI��u'l&��@�(��GDs�̷IZ��q
MjHjŮ�K���f�R�;��m*g�ۓn�FT�V����߀%e���Aٯs��������{����-�qd��%����#f�6W�Zi�F���;�$ 8�jx��61��0�$���+��q�o�c�J��x�z/��H�����+�>�Q�O����m��5 P�£Z�G�w�$5&��tg����5���sIMϗlv�ED������Pű���B8�toZ��F���G�_Z�R+�F�"VL���7]x]*ò�I�e�����`����G��I�����0�)HΑg"��QO/W2J?c�t�*XwV�̴H���B��5����K)
���~�U)c( [����;Jo�>rV׳����ށ|Q6^l��ѠXU?���.M� d��$&�M��ki��j,8߆���,}M��GXe\����&�:h�s.)m���Nwb�r'd�@O��I?��`�
�oVD�h�]�g��'�}�{R�3�!w2p�b�:A���9���\��{ J��ڒ��'I�5��%���]�xMM�$������$_��eRB� x%��w�'�t�+'�Fܰd�3�4I�[v�twl����[��|�.�f��~�ѱ%���\.㗑!�f �^w+TM�I���B��,Ѵ�I�h��~t	�!�Wp����~S8�?�Z<�}<L�tBU'f\���hĈÙ��M(���6��@��N��,���nܘi�
�;-tk�B�`f�d�(�.��s�p���D�s .���)�"�>�;��\��~6���s-F���V�92��/��:]Z����K����Jcъ�?{:��ͪ�/x�BN�yZ�������%W��� xh��Y�4\^������a�%+z�6���_d=�z��ѵD����8��U+��Pn�2�"���K��T��{�*�8�x,��X�Q}�R�o��I6��_�X���GgQ��*���
���ť&#�`����i&ڷ�>b�.�H�8��Р͙S�����:n��4Ϣ<�*�enZ��Zc/M�­��v�"� �lU $`��@��F��x�� Ru*-I+��1�����rZ>�Q?����֍8�6�	h�MeD���Ϙ	z_g㿋�B�EB[&qTC�:h�!!M��q���62�i�����#0#5�}���2��x��5��4�>c`�1N�펅��J7'����X#���5�ؖe���ڕ����s�g-�����8A
����9��
�����[8~�C1�;r��=�5h7I\Y���u5��Iz��uɃH�-8���܅*�،�j��-��躡VX1���=;:���8�JA�����[i]3�k�JP�KV���A�T/G��CŐ����:Ү�V��2���p�O���
5Ǘ4�U_�>��&y�y����`T@-��
�����I�-���Ҭ^\��LG�}̍��Ώ�n�(V�]o��$��vϲu��T@lWdjC��Q�/�	����8(-��I��5��\�C����z׭�x&4m��/QGI�_l���,V�ŚU�!�n�0��s@�"�|n�+(�Ӱ+��ٺxS���m����=�E��Ҧ�s��d\1�Ov�=����� �+�V� ɾ�������M�x �RR^�&�����	2�U�#�*��y�D^<F�L���I��ª?]t�\~�g%��5&�B�e��6����`�pH�Hkg���i�H��*�y����Y��k\��ȣN��ד���®��奚~{�(?��j���E!�Ħ�j��p1ْ��;.ga��q<��B�%��u�I���_��W�:{�m��|��eHzC�P��]
RS|҈l�Z%�#�m�h��Fcv�훾�m���c�aVL[I�.���8 0��eq�T))���F��Q�=�"�x��U���6B���{!3>�L&J/��qQKB��y�)����3@�5�ڙU��i�� Q*��}����u�\���K܏{�x�$fp8�~�����%�:�>o7�\�eM]�S7�2��U���MU���Y�m�����a\�/��7ȶ���k������i:7ۚf�c�J����6�9#�<iF��$K�*W��@Q%F=|�=YG��!�RDW�F;��cՏ�s?M��K}5?�g��W�f:ᄳ��ϟ9��_)�X��j��Y+������,pO��%d����`#��C�R T��:��m_����e�2~T��N\%8B�cv����ک�K�|Mg�L?�˿�/d9~P�Vc\ˠ_נ:��`��h �V���	��p�*�Z�"����b<p���v��$RE�h%����q��v�Ö����q��ܛ0��S6�F��fh��r�&�G�����__>,��BHyT�].�c�
�_�"ہ.�T�T	����AX��〥W3�@�n�D���?�̠K|�|5L�U䆢p�S�:�,�lu�S#i���H��>�f��YI�(|���I�}��Kj_��S|�H�x0�����l�Ҏ 닂��
���l���=8l����
o�$��z zl��H�bl���Z�3V��v�r:Q��ʓ&�Ek�v@?��lɯg�0h�nț�Y�ͪ����X�@���E���乀���i I�,^�: vg1K*�)��_���iB����N俄��(S�$�w挱��AG�O���2���  r֞���ߎ��ͩ�);��SO@M�r)}�*�ʅ)iC��MN�0��($�)��;�@���eAs�N�����Uxn�ڶ����ׇC��%beM_���ĮM}������]냯�Ϝ)�¹MӰ#������7�x6}q����2�� �`�CVb�S�� ���l��C��5]6L�ű���u!���lw�,+E�f~,�� �a.��6&G�pČ��w��,Ut��c�i��SxH	�3^���L���{O|�T��6����g�gzI.r�+��a4.��l.~#�hllCT(`�)�u4e[�/��?��Fފ����ef�Ag{�)��,�E����d��l�d��f_F�YTJ~�����e *�:�z<&D�BW�u�[�}�zD0��$1�t42Aϖ�r�1��/H�:�/����(+��� i��1��t�j�N3? {�����`��e;`H��N��M��H=�ߏ6�Թ�`1�ŝR���+����-"�Q*��Tv�`g��.25��$l�a6D�I�������h˶��Vx�E�gB�+���Q�_3�ڎ�L����p�����{f���s�d�Bc�϶'#"��65$�I�He:�gȢ��J�|�weʿV�#D<q��y�Z|��_�ⷻ�t����bj�t�i."������xCc�4�^�%Q��CE����Ex��5��(fccpM1��O�0/u��,�qJ@,��
�L�.���R>_�Ԣ��� t�I�Ƥ�j��S���E�� �Q��1#f�,���������jȢ����yz�ݛ�ro�	臰e��{?)ݨ����Y������I�]R�w��M�^�k��B޺��{���U��7΃�W<L����ŷ���~�xF���B�=�nWq�J)o�^p����	�[*j��0�MJ���7��Cb���9{�HD��d 8�?Q�jm�`���
	{�d9���FV��Ag����(xf�S�⌉��=�R������r�;�.�O�H�O7@כd�@6��ܷ��-�1�p�=q�P� ��m3O*fR���G'�V�aG*�Q�o�bbX�,����F.��I<�&�� \�ݥ.:����M�&R���.o�DH�q5 ֺ!�#;a�:ü�"nطz��T�
�;V=�>��!��<r4��Qg.�])����2�=Ά94�n�v_�V{�6Z�Ǯ����1'p�����U���C�)ϕd	����0f[+A���(�=�c��g��yb5��<��[��٬\�'����ki�t��"�ݤ�ʍ��K\|�u�S�F��9���Fj�	�\-�e\�j�b.<�����k_YIY^�@�ijMPS����O��5���Ďl���mz%��Y������5�����82�0��(_�7�U���\W$A?�ֈ���Oe�Vտ�L�!z��
��$U��.��h�x�Y'$5S��2��r��H���_�=���Xi�E1���䫓!M���"XV]���6���.Z׌���06����z?��!5��쟶�d`#L�ޅ �s���c3�&/���
W߭�X�<�(��i��X���Ы8�����D�l���pmB���oBJl�b�<W�#P�X�7�zF�l�W�6,�FJ}D& pm$nf�f���$�ti�#J���5�kP%�e��hhL0����Z+z��`���pd�n��%̰�l��#�==��:>J��]I\!�"l	���	'��ɤ�'�Èu���x�rF����zR��,�\i�+coX��7�u6WB�43�,�|��W���t�aW��F�^<ao���v*��s�x${�����qΠ�]Ǭ�p(���O�n3��lw��������vn\\Sb�~>fm~}�G�F�r��T7e�Fn9�^<B [a�a�F^�8� x}X��姪��17�A�ir����i�L�"oj�t5�K�P�,��p�^�<��(͋6]�T�l%qp}b�k��ԁ�&����"�F|�(^�?mwe���{MX�Ñ4�;�a,�[�U�.��e�&L77�'Wm��A���a!��_��B��I2�1S�b[�\��4�t��a���Mp۸���U��ΙP���=J��[nPf�'nmL؋��jnL�꿺�~O�Xd;kҝt�"������|��cU?OY�3wP_~�p�g�WM���pg��3��]��(�������l�誋5dUҔ��Nh����ueJ�Q�Ղ����+OYnp� ��#>Yz��]»̞ 6�Ι���_{~��_yZ8����Ay� �ؘ�3��D"��6ի��7��Y��������^L�(�����wH���m��	>־��uTM�EFp����+Z
m�`�a@i�H~ƒ�j^,@Ʒ�� ���a��&Z�,ڭ�a��_�.����E�Q4O��#_Q�f>b�X~ct^i�u��r�p�
�k*�M�Yp��X�l§za�R���k��o�m�)Q�d{��p��I��o���;5�o0U��6���q,��i@������.�`�ßq��JѼP,�Хy���_���%wȠV�Źo�}�0�������]YU󻟌��O�1�o�s�Ax���!o���~w5�9GȆig��8u�T�ʗ��/�fr��3�tR�hxH�S�Q���чE&��Y� ��-��yhj�y�EJdRG�?�E�Ĺά8�?otC��0���7��``���Xq���"�`6
���.��K��*s \���r��g���В���q"�=�A��)��s�!Gg�1�7k6����Yժ,�:{��,  �˧rW���g1�/ğ�nX�։�2��n��ÿ��SЭ]=C[�!f}�'ʹW�v��`Z
-/�nW�?�\A��%�~_��� ��^m
�ucAon)x1���b�JeP���Pe�z���0@G��m&7A���U��Q=/�ӆ����=���X\�vZ�F�D/�vXV���'F��[�u;�t4�$Ǔ��L�a� N̂*���*O;5�/3��ZDrJ_D���z�U�x��JD�z@���wL�%Z��!˰�ց�뮺���B��sGev"@�'qJc��⽇P��G����U��<��H�+o��h��cA�7��m�@~E{�w�Ψa�����GVԏ%@�l�+�6L	b�������n4��"��+�ԛϘ�E��yV?6�JM
uHNζu� �4eꖗC�)://J�Fd߳�[�V=���Q�~��)��H&�'���+#����zV�,��r\���Uhi����V��j�~݂y��H�����	�x�/)�E���筶'�R�Ĉ�A�o�v]�^��r���x0s�]�k=� ��V٦����8���ӿ��GO��]�,�����G�l:&��N�w���`7���	4{7�(ⷎ�J�܀A�S�����ʂ.�������VH!N�O�07י�g�j�8w+I��Ψ���S,�y%���J�"^��w(Q��݃/��l&�}��;��$�����]qf����LO'��M"�e���EY����9wLÞ?�?�@���I�Y�ݳP���^((r������t�ݴc؊�Wuq��x����9��q�_��MB8�p|�=�3�2���	����<��J�c$8��B����{�c����S �,E��r7�n�w�����R|@�����CA�{��ɬS��׌u�j�GW�O�nV"�IA2�{�(\u��qڃ�����!����K�v3�o���a�~�6��a�dd����0��\��ƞ�q")�*��b<�_��b�a�e��DP��Y�QH(fwy܄C�3���/�V����}��^����qf�('G3��`�(e	0#nE��NC�Z�8_��ɪJJ�m�Vt����8ց�^3{�p������O���B>�
�+��P�ʌ�RIE�������f�f�J�*�%'36����O��?��2����:�zNR�;Z�����E'k%�%!���'+��?�b��L��[���Ey���B�����+�~�����L
�ڕ��x	! V����I��2 ��NQ�[�N@�K��n_)�
.y�oV"�/�a����L �����κ_CJ:��ϗW�%�%`��|�����`��f骕���B����%ҙo�Գ2	�JO:B9--�l�8�Qkz:r���+�E|]�}���*O�kU��b�l�>wsA��x�h���-���?�!��gJ�y��\~��%\�Ĵ,�0���c�;�1X��40�u>�ԥ�JaPg�h�LL���(<�C���x��ygR� -N3�}�o�,���h8��
hq^CMj`@��ͷ�f<�91���])���j����Έ1eK���e�d����^��J�u 	ra K7�v\A��*��'O䒞���e]�d^�c��x3�������?SC��2q�3蛀�=D$<��p���6Ò�$J�� <�\P>�p�r���V�����A�*:�����-ܰ�ɞY�9��|c��$�z"ы�~\t��7�A�7�k���G� ��}�o��_�X�lԥ3�okX��>��JP�#g(
A��c?(Ov�LN%�֗ӛ}�g�п��C�3�'���=L�ˈ:�bD"�p�O�'}�_�P��wS@��%�D�@�֡�C\�GjD}����P̪��l�����E�`��A��zI��h|&��*�� �0��~]� �����Wf����ż��:��;��o�ۙa�6=sz|�6���ʧ]\���ZK��%��U�����	�F$��F������7�w�EM�VNJ�{֘E�V�߱�W��J8��Ũֺp��{:���6�)�M��e��~�PgoNQY��GNM��f+}�{��3bj9��������N���п����x��»�sWT7��k��V��/���ѯ�x�o�6�,s�DwT��c7=���b�KdI�x�	~b�J��?��69��j=� ��"�v��!�l�������s���Nt�Q=Įl�L�H�` ��*��ڱ��i| �]�>_��JL�XxS΅}�J������<�Ԩ^�@��S�u��a7�k�~�� �������@0z[�J
ٽJ�\U.&/��v�o�V�,�޻�+z�ikx@'��O�(ˋ.Vbtf��:H�*2GOR�=����b���8N��|�R4y ����x�7j���&�T�}�O���lTR�l~>� Q�:tc�G�J�V���C��t�b�i���T�R���9Wzp�L�^�H�6�rrي��cž��2I�/Bp�o[BCh�Z�C���4h���
��N����`g?O�!�����ZLgE�b:<�,B��R`k}hB�ł����(������чs8����NI��O=7�) ќ[o��F�������M���Fi@���
oUL���ʑ����RI~ą�8I��� j	#e V�v��R�zj���OX�W�{�좔��׀5h�BD\�4C�1)��S�#Ͽ*�{�C#늒:�T��̅	��V�*1�4���~V��/T��5[���\�c@%����Y�-	5���#�S� ��_OCw������z�J�:��Q�v*4J�?q�&K#"�Q��䬉��Ӌ�K�Z��?zN��랒9\�V����O��p���x�3:{�(#F4�SrGk/�'i������*� )@�ʠ���>gn�+�c��i �n�*,�8z(�{]k!_a+�n����R����u�����p�G�y�&�@�1����n��{�N#���Ш�=��A� �7<�u1�h�>�h��$��@VT�T�l�F�d���$�����)6���;n���-U�A#�}a�`��5��n�oݳ�#�E[���/,�V�r�&l6�Y-�'w���TF��O��i�wɡ��ԗ�\���a��1$��-��\I�Gx��e��7���s��I�A?Ӳ��8���C?��'p��������be̴���R��,�ZS�.���r�S����܌0e9�<�����ٶU�(�M�}���7������I�Z_��K��py�*���v�H)��o�Oa�;�ɷ�7Y"�ճF�-L���+�+Z���!����'��}#�9�	�iMow��w�<
k�Q^vJ��k�"A	�rɞ1bR�v��j_v��/�#�ׂT��ɝH���15N�c�{7	-/、a����)!}��C����FI�p���xQO�OG����̬^A��I��]��ᇰ���`�[�E���2�P�{�VĤ{5}DX�]iI?�ϙ�%ymԊ�5�,WI�՟������|�c옛O7���4����ibUԓ��m'$[�&7�F%��7�8�d�۬
R� �	j>WuD��,o#h�&���`���v_��ϗ!������ ��`���'�$H�[�W�;PIbd��+Sd���,2Z�;c8��3͗v[���Z���&La�pGr#�f��q��A���Y��Ѕw�X�r"R 	�f��B��<����H���.�H<�pC�2�`�_��w�B�Z�.w�Yu�#4
-�o��
�Ig���z�WE��U�̮��V��\��@.lM`-����j}B��HF���=rDF��oi�Z�@?��<�q j��cN�p��(+3���?�?f-ݵ�sr�7$r���~Z��E�-kx3}vR�W]eN�%)��kE�9&����2��;c�sLq���o��3�<ʠp�}{���}�S'$����sw���S"O�"{nL�:F����WIBY �!��8Ɵd�͚P��!�H���]� 2����Ru@y9�%�y��[E���N�l�rQѣ��m��
�ǉ�]������&d�ڄ����-�R�4r0b�Â��s��V�ԕ�e�:�1�)�o��>�����|��`�+��4V
�}��|�"VL�C?b�������!79��&r$U�<��f�l��lj�7P1�3#@v:P(���\yS�% �iv�;�{Dz�T:��w�X>ϭ���|3s�J� j	�.������̄��M�Q�Xudxsվ�o��*�W�/�6	�n�2����}J�L�����c�����|>u�g���S�ܞ#&�}<r�*�{jd��*x3ǿ����_��9�
kO�������i	�V5�+Q�P!�-�f��eL���@��b�v{y.���r��f��HG��AFf�QA�˭G:��Hz'eYB\C�����z}JT�(����ö,R�F�ֻ�h�Ѫal<G�����������/m��Xܵ��M��<rX��ж�&i��z����b��ܴ�����R��P��a��������*z�r�ԃ�������ӫa����f��Q�Wg6����, V�NI�@��/#�'3�����#��;�`����`P��O��>�k��5��gCP� �s� P�Q�5t�����jЄ5w�Һ<���Մ&���ۼ!� ʏ]�TV��%2if��W!\������7��رE��$�Dx�2/�eZ6��S�w4%�ծ�a�f�`��;�B ���|�Pz��6xvU#���̫���c�E�g��:[`��	4��($�lqS�U�!0b(��L!p��q�۬b�����1ꔰ�M�6�_�����pt{?%.t�?ZU�^�1��@�W�^��鷁#�y���H�K���26h3&r[|@x���mg���0���8�fw�,�u{g�y��� G�&t�l��D�r��t}Ƿ�v�pg+#M�1,���)YVI�����A7~9K+oJڎţ���KC-�I_~����A���:�=�<�A�ח��f:ذ"쌳�>��˪9����������Y&��ȭǜ(u��>�v�5�:�EDjU:�d`�."���!mA֖EU	�2'}L��y�Fp�"��c\r���h w�zcߨ*�Y�q��b�h/N�� k;��O���>���Ȗ��N;7@��D�������Q�%,�����r�"���$K�Tuڏ�����,�Aɕ���%A����=��*�X��y�Lȷ��l%�-��z����VP��i��ɒ��EUj����������'��ذ�.w=f��ܴ�����;k��5�}��K7������BzU�h6E��K�8�������c��z�pv�N����G�`�ߨA�1��j�
}�W�f-�?���5��foP�3ޖ%׷�D�I�',�Ĩ1_H�7'[�El/�ɀ��%ӎ�F "�������z�+\TF7��4q�l2�!�FֺLQ��%Щ��yv�����P�/,P�U�!�\�[����L�G~q���l��ˣ�G�����b�kjS�N`#޳*�(k�j��]��{�d�~�����90��7uaz�HlY��5�?"<}�ꔲ�fK�>	}R�5/=�3��u<{��7A6IQ�(��j<�r���{�@fBw��c�~����X��`T�x��7��H�򍵲(*�����dğ,�k��:1%Lw$U&���+�	s��ɝ�ȇ�Đ�}�	`��~?����
��j��H��U������=-��g^8�e��.��s�6�o�ݎ	W>��}�!����z��;�ee�PdwP2��^+iZ����M�X�lj�ܿ.���4��!��Z�麔.����~�9`M���������P7�h([ ص�D�7wɐ�
ɘ����зXi_,x�=�m"��m�R�	ٲ�f5]|��T��[�QN<O�����1Ca�(LIś�C/�ϑS�Ջ��v~��J(P�6�h��v���5A�����U����Ȉ�>�H�d� |����"l��g+��YV�2�Q� �k vU�.���
��BD�׳^���^ �Q#�y􅪀W��o�Fjy�X݂�9����)��H,֕$��o��i(w�����r�@^�q>ܹ�
�l��g5P�_�E��jިɝ5��wR�����1��T���c�Y�Cb\˿�.�7��<��� �C��Ŀ��D�8,��E\���i���t����XH�W{˒\��}k;�������1�ʴs3u�"��\q!�ϬN|MF�CM����l]�I"o��K��X�w�����v��G	� ��|%Pꃻ�D��r�z�h���n>AFE�zW���ĉ�;.h�}��:ͱC���A4��'��6ek&�k��Z���chþ«�z�@<��J0N��,�I|�{?�\(dɜUA��U��@DhR����anjhk��	;\\�Ճ�g�9�f�.R���s�0|�|�� J}�*��_,�8��
�Ejڃa!��;(��t�m�a��& W���v���t߱���M/��o��?`��'�G����㍨�D^��v�\VI���%�U3ҕ�
������'����Y.dЖ��o�+�o ��a0%�ri�����S��� �/�b�'�#ߵEF)�,��TR�mJQ��$�kY��rA1
�˲hA=�zQ�ƀ>�q�xLH��Cj�� �P8�X]+�a�>�L�ҏo�`�X�hi��8�����A��\dlb�/LKR�2Su��M�3���Ь���$����O .�-��d<�B!Sw��f�]�a�9��}�X�-�<�FUs�/c�����T�5��-`eFu��7���\�C+d�����j�UW6�9Nfvj/_9���-�6�\\���*r:�Rp�w��?���)�a��Ru'%�o��WjDF_��BҔ}%j��M���$髵��6ɇ�����;!����D\���;�TX�Dw��ٓ�R[��n�1����Q"'譝�2�1�"��+c�m���5��9�n���I��q~�l��Q��Q6���V���r�uКg%�i���)`�n�_�°�N��B%� � �����L�I��Y�_�� ��������+O��Q(�{�):ǈ>s;d��#�8�V���$K̺NM.|͉���\���;�¯�5㋹t�S�SbFZ-!ݓ��(�������B-��	'J=Bǈ����/�Y2���[^�I���=Y�)������i)U�憦g��Z�)C�u����7��g��!-y�����Q�p����Apcđ茢��h	"?-ē$�!j�5�5�.!��g�>
����0r���-�58E�~'��cO�8%���CL���)[e%�'j���:^�^�7m����z�24g�Z���T�����'�5i�A5#�hh�%�ɶ�%�߾�՜D0��*<dh�$�GA�M��������+z_w�F�\=+F�"�LW{�&�e�c&����Mh�ۧ�R�í�8�%t�W�\Oz��:��B�j?n�)6F�%��|��T��_�6����pi�f���e���֊Q/���a��!�YED5m1@2�5Q�� `�|��E��fR>[a9?��YX#ٜ�(�f�k��i�=�lC���M�6L��楉�Yͽ���y\�L�~�,v%j)��?�K�iӾj5\�T	TY<#B�;�v��V=�37�zt��2��	���a��Zૡ{��5��}u�`�9�`۞�h=����<��c���m��5����w�s��|�Ҹ���נ�t�p����XvC�n���8�N��� ����^�-"����]¾��~��R#`����W9��w�5k8UwjSb�=��T����48��ɺ8��}��=��}9V�;�e�oy$N��Z�)��W����tAI)$�R�7C�ƿO��M��`;,��{ �s����)2|#�j�Gy����19��x�m���;�cB�����7J
v|���Mz6-��?1��`�Ɓ�r.�E"�vYzo�>�B;��j�����������s2��T�����������'�F��ٓ�������Eu�c&!bؙ�#��+�e"3�f闅��Wqn��Vq���o��B!5�a*�-B'F�����d�]_Vʔ#�xΖ��&b�I�^�=���ȥ{2e��
���:�fI�h3\��E���?�`ͺ=���+>�E��VӲK��&	5-r��8&D�.�	=�����79��C��4�!�Y���&+�^�)r�M���-<���x�+J.�d�4�-���^��3��L��j�9���hf�[)���k�s1�~���g<|լ�O�vy.��ҿ:8r��=��m;����9���\gO�&�:0��M��[�2p��V��}�x.6*c A
�^�,nQ��WM=�~�� �R8��q�����i���)܂�Џ�� �D��X��z4�̶�>����)=t���E���m�-�Z~%��f�P����:�1�P/��Q)�˴n��XxPd2wbE�ľs^#�؊YH�"��}r R�:n��M�y�*L�0��>�CaE�����w��:`jl�x��I�Y�	I���f���D�"�����=Hb�42��`P�)#hE�6��w-C�=�V�Xa���\���.�a����[XUJ�\��H|��;{��O{7%[�l���)ps�1�r'V�Aa��hD�1B�l��r�ʗ�����߸���ۣ�E�@��#S����I���:�X���%
_9y�'��j��!�Fʗ�y�M�a�o˙<�M+��?~�a+��i-B|`�-�Ѝ�G�<��#��*��4=�ʻ�H�\�)�#���*�iI� ��$2N#�z����E��;�6����/~����'/� ��;��|�B ���;�3�:�L����c-e��� ���,y��3̞��ϟA�18�\�Cp��ڄ��<��D�(�I������5r����4@ٛ����ٝ&�G��������f S���L{�H�A�N?�b��h�[�#���8�ͩ3s�Gh�r�S�R�0+�	}�/�d
���9/q��0>���[ڋ�^C���`hz��-��L����&4���fI�8'4Xb��b��=8�s���$%�\<ӏF��V����plR� 4�g�.��F����p-M<��LS~�>�|6���[L�0ʞq���4��i�6�`cY���Qq34��FY�#(�e�M����<�/��&�.a���w���qQq%Zp�-qq���鯂<<��~I����/�s`z4�>nTd�j�tA��c��s����pQ�w1�;16�v�0��,XF�7[���u�V=��sr��J'�#g��Z�Ż��p~�.�Wѳ��l@}CC0M�fQ���Sr�{�LE
�r����zLn�vQ�X�χm�.z׿M�}>�ArS[6j�j� �Y��v��η Kp�*��uUsR+K���WD����Y�~Ȁ�ܡ�h���t^�=ث���uH�dB��P6%�x��|؆k�j��=��k!~*�ֵ+, c��G������U�u�I��5�*����Im%�a\��ړ�r�51���0'LZ�ZǬa����;��MOK��o�(�+$&^�p,����s���~�(A�NavU�B

	x��+�(�TU�'�������#b��Ýh/��m�j�>�+��:	K�0]'�R�;d*JB9�FtJ�RL���7�̒#PGC�*�9��w�@��P�o�5�ď3�P%V�աo��?Q����هmZMUn]��Z�}Gf`_�̓�N�F�mՙT.#x��\T���`�Y��?A��ΛRP	�a˖�ݞ^轫��Y}$"��0�j1�O����;#��ᄺ���Y��C�0��S��@�E
Ѡ)�.�W,1u?��8�7Fe`zIɃ�ʋ���6�}"k�3G�%�{ £�UE�j(xu<�8�$�y��s}�B3��|���0�r�[�8Ȟ�5
�������8~A~����5�Bt�.|OU�*מ'\´ǽb��@��cb�j��8��Rx���H@䉄*x�(���A����2�)j�u&<.L�,��H1��p\��T5ś�6a�8:�rՙ`n,���i����������28/�H��d��A!�D� .�9G:���*�_�zwiQ~{�٘����C���F(�����܉���?���3sͥ�e�	�o��e�M2T[lB�����Ǡ����d]	�pZF��P}�Aǌ���qI(�4D��gͻ�U;ô�7m�raE�SX�B����P���v��F��������C������j��E����'-�%�M5r'�IMu��v�T�Z��q�"����m�)3���M?/(�k��N��Rd�s����<�Xx�b���wӂ?�������W_<��!����������#IN�������a)���P���jG8 �L�q�� �Y����-8��Y&b��T6�&��/UEi��A�׷H��r�p����O˓�[ȟ+sab�Π��ry1�O��T�j�Y �w��ߐ9u�Y��V�C�a^kq��������?�o��:��?��m�<��Cf���,*ɬԭ�&��`lf��3��-k�'�W$�s9u�ޣ�Li33Lu^9����'%j�+Q�����_d��������	��6y� ����'4����EyD^+���cd��w��+�E�9�ٝ�<h���\׏��@RǍ;�oٮ����,*L����WB�։-d� ��1;	�4���O~�4Ȳ��%
}e�����K���r�.c�؈���CzK��x�z��e��z�&����*�2޾o������w�\�^y��E�ѺK�ў�"����c�faH�O��s�Cn�3��%���5˦�K\Ȑ%T��\�gP���r	K���r�0)ӗߎm�gb �~Z#�=w� ,i Pra�Į�g�KCl���i�6�T�p���(�*���1ҀV>Ug��lz&������J�8Y��m�<B�9�����@�|g��B���d̙���x�(�h[���F]M���53���J��!~��@B��ո��C�l����\�B����vUІz�����5�E�2Iy����=���+wg!w%u�T�hcN���*t-�ȫ�����H���O��Yw�z�*\Zu��=X�T�ޫ!��P�7�|*���\���K|,㙒!Ί��]6��������d^�	zˬZi�u�{������ie)ӄO��{iT�~|�P��嬶P�R �}A/���uu��
�@�<�?{P)��L�X�=�fE&�2_�1N.zI����C��L������g.��,"d�~
����W:3&G,k �zd�]{$r,I����K$�²o0W��dwa����lJ�A�2�X�ˑ��(K���]b�����?T�#�**��鸐��V5��'�-13���g���H@�Vgs�33�mp��nx���/Ì?���FSu�%$��_��WY��ip!�K��=B-�X�.)l=�`z%���eq�I�|Y�ey\@�XK���MlOi�Ҋ6%���d�/�zb��1P��q�$O���Mq jf�o�2�j�$Ol�dY�žUOv���]�ͮ���#k�#�3���q�\�R
%�>�w{�ۈ�[��j�����H�����T�4�!�a�C�$��[d,���/�_We��w�ų_5
�~��6�~��ă����V�����tw���s��9p��VFh9���#Hehx���H��<!@���ѱG��;���oD����s=2�p�^3�|��,`X�U�Pu��'x�Qr4��}ܼt.v���a@�g�V�p�M��foJ��b�U|~��K�OCS�� >����<і��R�3�=
T��x��W��&y�	Tk!*�àw����f��X��s�|� �k���QӍÝ���(�P�{ث��KB�U�,I
�[�و��'L�?1�+�V�� gM�>қ�?��1��g�k�kT	����IZ�ƴ7��g%����}k��K �D8�Q2�ƪK������|?���+8����d�b>�)iEp��3������\~{����uV��HѦ�y�����\R��,�����j N��|����!����Bl�94��:N��K�P@,S�D�Kv�\;|l�вa}��'�N��ĩ�?o���z�W���FG��Mpk��	��͆�]�$���'��o�����Z�(b:��ULQ
�>�#U���e��A!��n�ä��2���})2?���۽��e�9]�e�
<:Yŀ�:��}�u�6.�{W�c�;π�p�+�E��N�����8�<�{k��pI��KF�{71���u(t\��0-Y ��P���%�`�V�����d~�����U���QE��B�VϺ%�°$�⬄��u��6���w��`�?��7�r..����J�ϧ� @K&�N�TI��;�ۥ����,NQ�OC����{),��tE~h6�?�g�{A�vKZ«e����B�ɜ�]�1��Ps	4�O� ��qݑҁ:�z}�[�����D�1��h+V"��_���b�#C�2٠��Ƃ�b�X�#U"��g�5��*��g��w���#Ds�K=B�ԝ8��ee�9���o)�_���IU���3���0�<����UA3F�]�(r���)1���-1��%�經�~�Y�-ּ;�͟�:��*-&��-.O��HD��G~�H���d��a�g���=�.�t��W��~�M����e�,������Q��ԹP5E�v^��D�u�>]Z])d$pU\,�ݑ����TSv<S0<(����㇩
j�Qfݲ���L���ZQy9�4����s��8�D���U�����"��R5����Z�D��n�O�;�PX3��E~V慳ے�E�����F�Xk�['o��T�����G�C�j!e�L#A^��ޛ_|C���W:s���@�Q�L��gMh���b�`S�X�8��@��'z�:��B�%�hq�.2a1'4�����Y < 2�p$�R+�~ƀD{7$+�[�W��&��yj`Aml ͡�����&7f���5��j[��ٚ���=1L���5iU2�G��wW_ �N�A�|���sx����X�q=��:4:esU����6�߀5��n&4��b�=P�����s���i0G?��?���x�f�-lO�r�k�%"���a�y�}G���k���M�٠�n�:��LtU��pz�U�3vm:maĚ�O�S80�s���`�ͅ��+]$tw���qʕF�;�œ�s��/r��48&��X�TDsQ�Ĕᜬ�84�,��"��+kq�7K����a+�z���������d��jy�	ۂ\��c7�S�`�E☠�s]�0u�_$������hP\k^i֑D�7���Ӆj�	�}�L3�)C�ȨVĢ�	{�W,��VD~�{ꗙx�9��xb���Aݧ�	~�h�1�����~��jOV�d��	����g��g��\����a����bn����P�	{�5��-���jͬ�$|RZ!�@�]�v�k�F��뀠�\�W�.��:�~D>� n������H�8J�;�㶼�R�9�6y��K�_Z
����p�1"���H�/,6Fj���
ӧ�y��甭��
�K�ig:����c��\(L��M����ǰm����b��r/K���:MO��).��C�^���/��F�������Z���!^g[��#f���s�Q��CWhIߟb��q`����ks�n8><ۖov������9&ӹ�DӇ�H���o�
$���<�0xt��ЅWq]��~��ped  `�6��O�"p�*����f����6�v�1P'�3��7��m���:{v�-��=�؉N�B��Ga���E��ʚ��F!އ�--��G�Xy��+�+��n$�M��$���ً��kٳ�?Np��,�~�Ė~��K�q���}�*Y��αZ�6��0������ ��qjM���_�#m ĝ����^��	�_���.E�e����()I�Q�����s�~��6��k	$?�ͲQxQ7��b\�o��(�m��8��N� *P��Wz���M]�v� �z��p����jZfa.����-eb�m*�$�IŻQtƯX�. <��t�w N���,لn�d���-�Z��T�@��x�W���!���׭�N���ހH]G�����<B����$h��q#���k�5U��b!����0d/F�}�LP�ۄ�/"�S��������qm��8K�7v���x�q�e�Ѷgu�(�0�D$\|�ySZm�,k}�j�w*h?�K�>��� �a�'�����Wv!o[2r3 W*?x�����Д�}�AR���H�=q�� Q̈.F�qns�(�2x�\�u��([i9��z���=u�X{�>\c�垷^���F��.|�ޟY3�I�
*}Hw�8㷴(Q��&�#b
��?/nս|��8B
~{�w����dn+UL���l�y�V���pOKd�T��=���d}��G!�8�
uA�zcJptqD�>���O %ҁ�ݛ��?O��0c{o����~p]�D���ru�������Y��ׁ����FC]?���+�=��5ѩ���=�A�$��:�̗�=Z��(f�͂�#x�I^WKۓO���D�mD pQ[6^�|���};#�c�*�9��������ő��Ɗ�zmf�b�y ��S;�|xL	c����D��U��.l�f��Ki%����N �N�<�b�\���d���·�ȼl�`igҤ��3C��J�Ԧ��D�ރ$�y"T����,t~��tOϱ��h�Q�AÀh=R����Ɲ�hs���:qf|�7.Ў��Ī��+ќ66�L<Y���.�ۂ�"��֒�{��p����$�@�����������u�<s��_�3�U��JH���Q���^Baf{#�>V�l�ե/D'Ei�v��t@5�����DM�� �GHG%�2��́Q���h��p��j�O92aݰ����$ �����ŋ�/h\}���!l�&�)\�j��0ـ25r�OziM�
}}��n��&B�����4K�)F��.���cЧlX.12qηlN%$_�fr\
����V�df70r�~���q1Ա�u�QZV��p,o:	��j�\,�.�*7�&�Ơ>z���0$��$|�bl�ot��<0��}^�+����Pu �UL�׋�eۛEq�w��ŨL����6�a�{���$z���/�Xĕ�)ȹ-[0��U�6a� vUd-��;RD�to������:���)��ʠ|�fJ�גu���8���j�#Y��`^[�w�ƗU1�0h6���H����;n),{�SR�)7Lv0)�����A����v`��'�r��$DQ���r��*U I`����J�iw�����C8�΀O���F�k�vB�b�9�ʙ��QZ"*������)��T[;+a!|훮{�i���Z����uzZM �I���J�����l�49��>��/ڭ��}
a�W��[�w�]3�V��F�������G�����rM�~�3�WkOy�Un�3�}E�W��O��7�
�δ�T���;a��U��/ܔ)U��P��*�n|�3^��B�؈�O��̣pLx,�!��܇�<'zൽ�\�XWiX`�[Rw9���Ƚ��UU"�>_O��|���;,xs2u�������^���`g
L.)�{�9�ɜ�e1��rR/w���� G-�����Xj�/� ���I:���B�:L����.���Z2aa��R*��E̞��{��[�}!:�����?����ơ%`�P��,*�i���������� ;(�_�	�"��}1��:��Q�/��N������E�Y<l���M��t�rI"��c�-~��v4�
L���:�׫f�e�#E�r9����>���E�	@V��1����0�osoq����&� x�u"@��ST?��	�a�
���-0�+��鮅�>ϝ:�.{ۧ�X�d�,D�Ox��`�?�(
^�P�2��
LL���j�=-�W����i5��䥽��]��8�W�;�khC�ֺ�~�y�'�*Mܱ��@�����������=@�/��.q�LxTd�\8����V?;m1H�G�yH["��P�50����9g�R�%�ր|�Pw��{؛ �0 ҞM �&/�X��W��g.��O�^3+3����Q��=(����4p �2�ڛ����������&E�|X�E���e�c��8�b���m4�mFA�,�h|�Af�u�tRT�d9D�ۮX]��f���)MSBq������H��J�3 ��>'"q���(洽ķr"lb�3-��褠�b:��p�c�7;�oP˘�9
�K�ZGc�0�>��m���+� �o-T�t��+��.Z������ 3����t�o�����L����PJ�?���"�1 �`��C	�W�B.��+C���>��W�Dc�x�+��y��R��P�v���/\tH�$��[�(9L��/H�x����A�Q�:x�Ki�e�Me Sfò�䂣)Q�:����w�Z����5��������㸫@���3�'īj���|ϒ�G�X�`\kզ�J3��_"f�yH%j)|r6��\p�
�>'����@;_���iA�P��-G���R��A��H�\eV���C�\��(f�#����ER�*4%��ͳ\�I�4�W�蟪�YfQW$���Q���Wc�T��ӎ�M�I���>�h��}�����i��O����eL��&��
5{���W=���d?�T�ͧ?:��"W�(�פ���X��HW�v��3+�M��csP~Co��ͧ���&�	z _XOb/U.�n�����8��}0�o���ILdA���'Cs�<�fpu�Q��sF���	;�J*�oX[T�H�5@�
���,��Ė�0�*�@���H�n��-�γ4U��F��o�o�0nF���^'��]/W����A!��Q7���i7CG�o���� ���!�z��V�'$6�a��}�?{wl�8j(E
"������<�2'��h�pr�"�`�ߦ��y=3�mqNe��v�`Y�*��8���x��<js�`m�P���5�����q�v���V\]���������������w�:�/3���7�ƠϏ�S�P�&œ��d��h�Dg7��<�܊>������#�<�������z�<��yywblU�W��>� �pD�����\�度�ՠ[ ѷW\[M���b�\.bC�������Om{���ۓ��c{ ��,b͈��m`�������q~�[�wo
���嫥<a��0N:�yP��,�n�����n��p5X�T�U�q�T�j����U��(�uZ�M;b.Z�x��4J�9�VE3�M1	@�`/��`�����e����W���l�	��-M�_�TTTim[���a�?ի��|��2�����P�4z���[~��o!wA@���/0m45@j����|I�\D��m.�}�<��y�7�%U��z3LnbL�H@ �:�������#c$��=c��rN�B��_޴Æ�m
�K�$�������֫����QQ�f!���C&1�uc���u�g��r���t'��yP�La{d���~��a���b��*�+���rJW��,5����\NoS��+p�_�L�P��2/�&3�1��!+h�;F��S~��Q4�%c�V���{Td���OP�p�~g�K��M��mo���Ƒ9x�tW�|Q`�54���S�ˤ\<W�����7(����"~�e���S6G0ƕ;n��^�ps���b>6f���^ֹg����$���xy40������7��?=�r�Tʶ낚���g���8��E!�b�E�5rUIx�` ?��l��L�!��xQ�N�#2��>#R��k����K�����7iA&Ӽ������D����Z��bt��(�O��n��}�z�c[W����Oe	��(a,�B�p���p�j��6�����=�"�H�Yܲ��WE�$��SY����?Y;|��6��
[oI���t�-d,�3��Al��X[n��D㋱ۺ�\^�Z����tY魼�â �Xu�Ã�`�jO,o�hup�˪Y�Xhb!\S����4ύ|}A$�3�{<�Ok����ri�3���^�w�6��[��X1��r��k/9Z��S-�0}�p�r&6����H�����z�g�`�r�[#	tc��'� �1gp�<��zRA�h��cSU !&SH�?���Dt�ZǍ��|����%�����:��{�X���pR�(�.ȧ�N&���*6�I�J�0Iq<��K��qLJK��܄�y�S�|�(�C\{u��_����m;]�V�U�ħTF�,@��ʇ1�l��AĻ/�p�Xa�R�n���h��J���%��+P�2~0���zZ�1u����1��j��^�nt�y>u�"i�?�cS��)u1�֘-@�^�|��n�Io�ۑBڃ,���b�		��JF?�����A�(�����-����k��<��1h���tS�����=Ĥ}AA��^Ĉ��.X����U2!�8�����d�1b�iOe`k�I���q`{�E�5x�[�BN��ѥ����cͰ7�V֜��8�7���^�l_�?��D��<&���0I`��0',���F�]�8r+�r��`�[X:�-6@�T鳱,@�x��ZrH�mJ�J9�5�:����d:�e��><[=j�(���FԞ#�fLjI|��Eb�<M�RЛ�ٱ4.\�_e ���M[4I9{
N�ՏɉAh6���3#�x�Yۛ��sa�_	�Tvv�@/\�B�G񑈆����2#"��������m�9ē4��4:y��l�§J�%��5��S��.���R��u�^��.��8�����i �9����I>�.8.�D�4�>�,"�.4���\&*m; ���'a�)��݆�\!ɻ8ss�0n��=���7(N� �z�Ų` Yrue�%c��O$By�Ƒ�����1����	H��	��HO.o��h��0��>T�?y��n_�W�����
5?2?�K�z�^��z7�P\����r$eX��\���zנ���-}����d�2�BI*9O��w�?��c[�"�;K��M��3��x����d�����4T��kݷ2<J��c,�Y	�׵�#�5JOßS��� {<Qqt=45a���*��ȭD}�pEڮ�l��f�K\s蠛�e��2�)*Y׺N��Do,(��RǕ�DF�p��|(�T��'1{Lp��$��<��؟�_��1�8!�y	�����\&��Mdm7w�dsNȊn�C�4����u	��/�iB�����1��e.�����(@�'Ag�uۣ1\t���7���ˀ.����듚�1�MrY���x�|9X�0w�����M.��쾾f�M�F��L�ǵV�*�i ��PV�����F��xQ�7��0&/�/�`	Q"��]/�l�y׏C}�1�\�T��K�˗��M�Qb)�=\������,aw�Y�㤐�c�9Hk&"�'�,V�C$��]�A�c�^�e�du�$p�CyX���u��L/�0��^�m�
��`ƌ;�*;��Awb��CQZצ��?D�މ��e�M�s�a�9r�,�[0w���
��
�|�������n�p���x2UVcI���t枨�Ғ����������905[lU\!z�m�0���F�~�_c�;`��\.z�����(g#?����I�?���_)K6�#�@A2���R� �H��1 s.W�N��$>}�N�F/}q&B��)�F<��	�J�����ZV�Í�i�D��X��8�>�W[+�jR@;���ٚ���t��O>&`��ˀΥ�����bt��rW��q�2bn�c�$���H��6M8�ƉF����c���}z� �����`��W(�&į�I-
����ť�qxwA-#��G�30ӛ{GDLW��z��i���(kΧ��
���M�B��:R z+����u�A�HG�e&rq�~1k�>Ӡ�&zp������[r\��>�KU�݂�qU�/H�Ġ�ze>�23'|{���	��.�W�U�)J�y�8}�����se��/-6������]�+a�gU��fgck
��
D1 ����»KI8H�d������56h�Por����� ���.0�F�Y
�GpVV�ܜ����H��.���ٰ/(�Ji�w
f�8*e2&M*��9�2C1�m��H����0�P���gwb�s�9���Z�_��!̺tKjl�̔l����`sb=�*{�_��OfۙG�^\��8_İh�_�&���L��  G�h��lLk7䌼�X$�%���3]�Yj/ m5`B��Q���_�D�y%N�{gQ����V���W�Tx���;��(�0FJ���4�Ep� �9u�ט8�x�L.�������lWT^C���<ĈJ��?�Mx���n�8���_6vå"���ZnB*&���00q�)�^+f�����M���#yR$<U�̻����A4�cg��W���j��@7�u�9����5OS��lC�2M��H�BV��5��}�r a�:pum�ĳ�D�#+:�$���]���p�~*�QP��_ն�PH�-�4( ���I������w��]���n����$�xqM�%v
�޺�_�ʙ"s�t!]�YJvƣ������Fo��'�U�sT_��a���R�p��6u�0���΍�I��hkc�d~�D� �&.�Aފ��`w�i3���E�7}.����8-I��Cl/�O�8~	���'~(�35�X���L�Q��QK��׵��V�v�{���2����$laU��icv�����x�=0�����c7�F���y�"�s�:-����G���ǣ����cF�Ӗ���¬��o�<��S�BY���j���PO�W�;�ԓ0V� U�,�B>�M�Z?�AV��r���C��#�<�:�8�'�S���E�}ʑ�ߏ�َ���O�I�=_�/����{��`B}C��p#����	�W�zs��%u�5�Cq�����#!�O���ms�'�� �K������f?/�G/��l�P�����䧛�F���Š#�*!��[�P���^��?&vɃ�EnU����p�S�b蠩I���;��<a�H�=�Z�����^���b�*�b�,��ޘ������F6�\Zk톺�~���1T]BK�6Y*iٺ*L+��;��ax��"�z9Nq��ԗ�Ɉ;6����u�%�t�T�3����.b����M�'0��*~��2| L���
��N[h�(V4B�����2מL��D���Z��Fؕ�.�_-�/#R>c�c�� VQʱ�d�5�,�%���!��n�N~�o�]]��Hׁn�Ym����Ro���^$>��Nnry_~��7FG���+��u�"�p�2�u�)��o�ނ�:c�Q��$nh��$Q��B=�k/��מ�ɇ�F�p-آu�3�0]���r���Q�`$J�՞ᏹ.�eZ��}��B�Ӹۖڢ��|EȐ��JNd�{��m�͎lYv����&�^�h?���$a0����Sϯ����)�E���O����)@����{���hb�Q��0�=o�����PA�竜n*'���H��o&#|~O���V
�Ꜥ⎯��F�՚�мa��>G������"�ZxA��v{N~�<P۷��u &m��6�
�/���n���x=|�w��#��koQNy��hG}��B� �vu.,G�998���+�"���Y��	!����f�� `��Y���ju��I��@��Th�[�_Z�mҽ�LU�mGH��9�}��
��u5xV�|/�!�����Z ;���ׅ�.�z(�U<��>�whQ�r�(f��|3���Rt�N���~���e95s������"y.�O�FM؝<�Q5����^�x�:��e��i�=v�;C�s%�Vj�5��hŢwo����A�r���e��V!V�/�Ӧc�XN��y	��k��LC��Rk`!M��.�&�M>$E���٨��m��WW��iF��75����W���no��Ř9S\���֪�:�UɞR��ӳ̺g}D�cH��^�a��
���qe>���j�w	�HѶ4��|���u��Af���=���C�-4bN�I;/��"�QYRyJ�(��U�ms��`<�EW�U�e��[�:��Ȝ���Y�縅X��a�����i?ܓ��?8�����x��������e]�J~�l�Wq���N�O������OZ�I4i=�����d:z7D�f�:�kQ!��!sUs�G#Cw��e�e��G(�3=���:�_����PV����ޜ���nk���";��y\��0Kk�Tӂ������W@�"�� i�(9��
0dD[I���|]��%��J���ty�|5����h�)Mu�}�Jь�}��g�����n�,�ו�5�\�H^������$��ss�W	k;Ջ����>\��M$��{�G3� �;G/H�k��v�����j%�48w��ڰϘ_���^w��ex�T
~M�)v�L�6R�e�ﯣ�;��y���:���Saߠ`Y��w��<w����;���s�4��{%h����-����Q�=��;�w)�a�jN #�Zf�{�[N���R��� �N�(e_,hA_�H!�+c��4�С(p��s��-FM���|��!�=����- �9�w�.u+��c���=��ݽ����rc�v�Sp���*�dR�x Eb$��,ز�??���.m[�Eu� b��yX�m��e��Fa��9��ΕB��}��[$կַ���-�54N�	~qM�2�Mv���~oi�|ڭ"�Q��EC�2�H����eQ�0e	HPd���R/=�·�V�<@���*ѯ�M��K�T�OF�G�'d��{.[�vك�T�֓y�qo���c�4��T�^�]��!��+�WA��׷�>oLu&�L����z,�+O�@Nw�iR���@��mkN�X��v -�s^����~�%J"
�X�t:>˭�zWG	�b,�N�L���PZjA�Ɋ����c`t5�R�U��<+�B�	%$5����݈��7t[������P���٘��_~�5��:k=!�f��f�8&a�B,ԜuA)7_�u5����M� �@�'�jrd���>���"��,��չ�f���c�u����z���ä��Y�.-�/��p�e��"Jg��=I~����R��{�s-�Wi^�N���Ţ��SE�~�ō����n<;�[��Ψ"2?�H�C�����ˡ+抛�+	�a�����O/��ɍ��c�}V���xXͦ_H�$�pD<�Ɵ�@ֻ��s����8���w�i�ޔj�jv6@��Eq�ȪP��DEf@�|�$A�e��X�b/T��0+�����6��G���g3j���h��(�%km�Vť������|5ڕ���-�WO��9F�U#i�g>[؟�9��>*]��~�m�!S]g�9���]��P;0>0��07)��B�Z��!��ӭI:!,Ua��2��2���I+��3�����'|��*�t�p"��^; ^74jU�����JC�LJt��+Y,�� ���N��m�'*T닩��.�~,�q��:�"ȑ��v�`1"W�ۙ�+
J�QK)�|GD��%u� RAy%᫵K�.��z���p;��������V{��H�Р70�Q�u��UO�`�֡�!��y���bJ�q>���yE%ڱ#7��wN�I&C������YlA��hC�ᯨ��<8�CM|�O2�k�є�Z����U�'
�jk��j���C����蒧�ͩ�S��L�)���@�BJ�&���'��=n����{��� ����H�Q���=�<)��������ʶZ�2Y6���:��|���ȿ���4�5mjͦvr;��?o&��b::j7�4�AT�F�8���#Qk	c���&^��.�p��$��=���>��7�����6��-^JKǰ��4�UFv�F�0����,��g+YKUo�|`q>8ؾ��C2��Q�
�[ga�\�M��l_|�v�U��X5�4A�?D/	�gL>�����6�9@^T�s��k¨��9�8���]��ĥ�5��kl}�К	{|}���(HOmf+�n�S��w%�����W�J���u/�$MȾ�>΀�O���5�h�#���DF{t�ouBes��\�(-�=�U5=8SPe�u#Hs���KQ�3�:ܶ�OZ���$��ѾXj�BBSP����s���پ�AXMkQj �H	������)��e�4F�-�tBG4ڒK??l�/�L��������/����0���;%��������IO��=r+���
�3����?'A`��&&1���T:�3�4��g��td�>LN�i=i�}A���?�Yj�7�iI�Dfe���h���q%.���1b
`W�_�b�Y~:�c�yA\~�Xp��^��C{a��N��y���IS X%G$��{��������ć�6�s�iUu���%���K��_�oCBO@WD'����ư;�W�ADԨ�"���E�+������3c�cnL����X����f�]u6ڂ���0%�+T+�1�ކ �
u��bا���B��7�T"��J��	�C,�v�Q{����D��j����1U&�ʀ|��M����U�}O�H� �y�����2]<v=vf:�;6$y�	 y����
`��4���+��\�k��8WvD�c�P�D%O�B�?߱}}�j:�``@:��Kǉz?�j-r>^j��t�iY��q+�,�Ä��KzG(��;_�#\���p!����Z Y��-V��;J�9�(�qsP��pԬ,�%��1-�P8�}}2�a9%��;%��x��;R@�gE�1��f�n��dE�Frp
��P��>r�`�CN�Ew1g��j0*�'#ZLt�*�U�*�v�x��أ@,}�S�u��e��@$z>�w\�V=[֤t�a�Е&�$�C��I���O8��C�xs{�g#͚3�x|����ISI�,�f:ҟ��]z!K���`Y8�ӥu������P�h�r�2侓� ���i���!�*���͗�+�й�����Jr<_*�쐋��8��s���&7�����pl��Pˆ<�T7�Qg�^~��$���T���b�������@`2ٝ`�b�S^Cʱ%k{@�f��Z^��ϖ�(��m���Q<���1��N�war��P� 5WXA ���x�M�|fhv��;~����˓E$>Ҵ��Og��W[W��$�O{.�����8�n+n����X˿K���԰v�lE+2���No-���c��N;R���I�T�t�bD ��_�0��&��+ŘB5�q?	��)%��M�d[g\e	8or�3�^=�*���ˡ�z	T��i��C멣�v�Kv�����%;ɩͯL�{�D����t�S���q[��F��8����*�(6I\Fe�u|[؁8�㠺���܈�:�t��t|�n/W}�e*����Ja=��~~�=�?f��8ꑷ,�P3\p4^C\�b"��j�Bɏ; �/���)�ng�]oA(�%�ܺ�|���~Cwf[�^�+���4_�$-�����)읳?(V IN��ПvG��i��[����7�X-FA�4y)�w b�;��/<��/��B����
@�Μb�Vq�<����L�>�S�`��� ;׃����'�+�O�2���R󑉙�w'�j"��%���3��G7��&I�l����U�7��;�nɤ�������8̓���!�0�]�U#΄���&z�`MI��\��cɶ#�qe\Q�@�o�a�*�z���p&�|ǵf��.[|�Z��+��K%��Xy|)���J�5�ƉJ� ���RNy_��v��vĹ�|�
�n��QFݱ�~  7I�y��v	 ݢB���`�kTB�T�>�-:��4v�RuCg~�C���o��^߾�uz����6��W�^o�XAP�71|bh)�m8���X��"S�L�#��G)xWC�]������#��������d �>����nE;dܤ�L�}���a�[��Pu��9�Q�U�Q��V9�v�;/Yz�!�)�(� �!0Ə�ޤ! ��a��g>�锸�<��Dd�84�M�f�'���˿���XE`-�(Q��b%ޫ�yGdګ�v�F3dt��I����"2v�
Nfo�*���C�8����{'��"��'���x��5���/x��S���(^Z�Dp:��Dc�M_���2.T���|P�X�� ͙��u�a�S7a���?p����D�2�jR7��s�'�{��U�1<��C��C �[���C�Y	X��&`|��s<k��{MD�ح��,�P���N���;-� �u>3u�D��b��M\6�%h:Cg�v��O��o�ڭ���S�%��0�j�Q �(��Wڀ�PoY<;pX��;����qpl�L�j�g����%ü~�*��F���ٹ:��_Gt�
G�
=Uj�j ��ٷ���6��]"/������^a\�F�i.�>��d�9yk<�	�^Iau�EJ翚t+a��	0�+,�7ͤ��{L�xmJ���f�	Zݙ���R2���!EŮ�U��$'XM��#��7O�K ��T�=#��C���B��.��7"��w�0"dD .�Ԫ��{bPfZt�gH�T�>0���H���/g�i�J�K
�{^�[1U�5B�Y.�:��#�5��J���J�� ٖ	PI���qbmI4d����5�*������ާJ��ݪ��܅�ap��	�6�V�T��:a*pk$�[�ED�/K��,�Ab��u��j+��]7 �����B;q&spJ�Њf����ho��5ς�>���RÊ���RT�_��}���� �^+���?�T3����<��b�,0&EzA�6�P�I �[��2@�ƣ\O�T�76���ta�gy�X�/Ȉ`o��\���(�*���:?ڟ�k�p �H��r,$?T���"ךߎ�+W�jzI�t]�X�=ӨbV\*R(��ᭉ�ӻ��s��a��:�i|;ܮ�z*y�|Ip��-�9o�ⷞQJ������e�%�=���"��Po�T��w5�T��iM'Z�Oǒy^�3]Ԩ.��p6�����9ׅS���Ҹ�����"[U�-]ä����%I,.}
|�ܨ����y��0��NB����4��jF�?��e>�>pٰ$�JQbu"�v���c���Nʹ]���H��ПyL���
���S�/�7jڦc���,�6�Km�:�~*F1'���k��U�I�\����|M%מ����rS��we�Q�f5!�iބ���/�n��+�ܑHtI� �/�Ϲ���S"˒yc�"�q֪i�q��2�s�h� �t�*d��ɘvk#׿p]�kٞ�4��߆�'�&�:d{q��"��vE��?�GwZ�<VZr����.ы��X��Ӄ��e""r����P�!�]�"�&��i�F)\Hr�n�J�ط�{cv��}� ��d���ȲU��=����rߠROs��ˣ?�}:0V�%��2г�|J�S�?f+�!lu�}�2&��O$e��"_���"��^�{da�q������R���*K�_q���.��s�Sj�\���ic�e��
\��oh�t�x~8Y����f���2a��`�0S�9��)��?4�^�P�b�= *�X��J|\<>	�;��E+5�$�|
Y�`�}n)��&���H�-�o�7��z��%�c�zO�e�j���b�i����q*��96]��L�ɘ]���ȋcͫzˀQ
��9������_�s��F�^8D�:��yl#�ט΃�B�;2�X��E!�T�q�|���ҫ���C����`)�d�[��&�V�_T)�������!S�<d�|a����q�n'�g�('�׎!#���Y�?�[��]�0���2�2c*��vw6F6'���;O�^�mrŹ�x�s/�{���i����R�`��v��8+��9Bj�G�Jl)��V����#V!>��2�C���E��V���;ź4w,��g��2�GĪ�����V�/���$$ׇ���\|d��垞���ǈ���a�{��*�E��0-W.F��sBTu���0_�w�2UZ�1�(Z=5�o��v�x�� �wѓ��������!ǚ���'�
N�@�ﭏ�B;w��@�~���/f7�i��B���B8�Pw)����cN�;�
5�ὸK9��!8�/�q�?��b��;c&d�?��Fk�=��@�� �I�4�2���������GcAN>�ʮH϶'Wg��jf��㖝n��gv��<���_K ��:�tV�y�0�z�����Ǌ(�=̉y_4m]���)m�Ǟ�;�#�u�>�{�e��* �/�s��kg�|*�7�X����V%6�z�%2p�ʎ�\��� ���i�/�XM���j��]�̦[^dv�� ����7Ge��[FIL@LA���5�p	�~���*"��	��Z1�N|�ur<S�VShE7�� j��I�d����m����;����d�_�L��}$ە�!z��_�����r���=�v�0aL�w���>('�,��%�p���^;�TZF_�x(M�2�n�3՘��.�2��� ��
�R6�@K1urذ>����򶔏O7H����h�L�HPk�������iB��jj�3��&q���SRG(ᶏD�Z�l�'�Ը?R�6f�8X�Ӯ#�W�DX�����������+e����xҳ�N��v�[��F� �\i+���x�Ў�3mZ[)Һ��n�"��4=
�8���=~.�IKRK��b,R�2 S��!�ē��9�3<�U���/�s��\G&�B�� �Ko�s֖#|�^�\��MN �0�~���4��-����51i2����i�q�Iu�t�ެR�T��w_k���Y+&�(�'! 2�UYY�tllN~��w�� �J�sd����>�w_�~do>/@WUq�D)<�p�AO�X<g �,W���y�������!����=���2��#B��m|�z��hi���"�������V}t�e��7=ʂ�5[	3�d�i�oDŠ*�cZű�2&�6���{*B��l��o��	�n��U�G��'_���ؖ�˚
��y�F�G.H�H#��?%��Eb�B��O�%[Q�J��vl<�BU^��V�K�@��Λ�~�l��5o8\p���d�Ɉ��տo�!*��&$l���g$s
�V���J���P�I��yd��b����k������X�ѫ�]��67��C��H����-�� #�"��I��NRs�'Ʌ��ʹ�.$��Z-��jN�y4$'��uΨ����%���/����Z�.��P�p�f��d�{#"�y�
��A4�C��F �x�+�6����17�fi��c�q��jO"P��J5�4t/�a>R� �ꈄQJ�v�Ѡg��i��%���be��>o!xp�x����^�D��C���hpx �d�,+�LR-W��J��v'� 0Y]_�Q�i�����<�W�xܼKc�$�A��ՠnw�m��T]aI�[�_&�1el[[`��{Y����+�[~�)��,�����~lpJ;�~�ꜗ�l��[a�<q.��o̵�y[P����qm�~��"��8�����^��6۟����O1������x/�8�ɓ">�����D��}�j���J�`Ϋ�L4[�:u���*]zm�qO��@�\��ۋ*C=n�g�l�Nl����96�g���~+��ϻ�ǉg ��(���� ����,	�5�5C���k�������n$D�:������$*}�n���g�$ZLSq��d��粨��)�T�_�HЇ=�"'���C'�S�V(�e��G�לVo��8��ҽ��.���0e����@��|~��sa�Gw��j�݇�,N��`���X����Bk�,���9��dm|��E�w�Sp~�2?&��������2<��_|4蜸�Wј-��Q�)r�y�Y�	��n&
�T�e0]Qa�a*�P�Q���N�-�O�z}�r:��3	��f��y�E���[�(��Z�_���(-*5��b�kh�Rٌ���)��N?>*��(��|b��5e��iEYH`�IwA�Pw8�C���'F�K~��^�>'1#�ݱx��m���'`6�<*��
���D�盓>�H�X��T{�P)wt\d�a�ͤ�q�BVH��ȱF�\��ÉNd�5�RA<("��6X@HGNYT,R-��줒BS�,o���֚k.���Lu1W.iv�j��h�V!@�Gtk�#��[�N���i��v�Y*�nAp�Է��ڈV�m��5�J/u�����
�b��%k_T!�L�1C��zH���Ya��J>��[@��$ns�]~>KU��:�3���%�9*�K.Bsa?%�p��*����r�1H�xZ��{<.4� �M��74�\�MJ�U��`5���U��=4� C��K����̒�v�]^H���?�VR��e�� �#=/c�t8Gu�B���`�Z�S����������v:T��&'ȗ�y�	���1�Qm��ib¢�o�2��q"�|�7��}̯��T�Ǎx�+�_Xh���R�'��Q4,�?�9a����qO� ��Dp
�-"��g�ю�p���R ���JL����숣��bP7��޸Y���O��f8B���Ph�5,��+��l�9C�{�N�������	񰄲�2������D���7X�a c]T�ί�����>)�1��fqO��!2����������?�j�B	��V���-S�E�|�	� ��D*��5�N�+���&�'�I���l��=��RP�1�A-w˻pY�p0���Y3���)N�ޤm�z(<R�&����?i@p��2��#2�O�o�֯��@!>����_�o���UD�h2�ן�r�q6�ܕ��2�?`j�}zF��ςVtx���N^>D��{cC2�hT�a�jl A��2�?�&��n���aJCR��o�r�s���ى��v�)1�U�����;<�;�[�PT���n0��Kj�2��i]zaW��;R7���6I�и=�Ķ�;���\��q��B��G�k@l'@�T�o��ͧP�"��#�,�e.��2/�.�s�w yk���Ϝø�����{'�Vh�"	��s���F�Jv�y'���Sf<��x*l`$���sh}���H��p�`�6и��R+I�ʈ숓�����ܚ��:�v�m�ҝ�ɔ��@����}ɪ'f�A�P�gH�����7�I���q��*<e�1�j�!G�L�$��7�ߠ�ww�^B��f�ݫg�p�y�ފ�U����߹a~�n�ԓMVu��$3kh@�}#��b�2cDp�x\R�Ou|��[�1뭋uh����йf&/ğ2{�g+`�����b��4���%1O�y2�f�F�ib���V�F(����������<_�CN^{ ��D���{*k���#�
�+�C�"��?�x���h���p�V�輡�Nm[�Ԕ�U�:� �G�[�#<�qQnݏ�������fL\���� \p}3IG�q[rG5Sf�YcJ,������%߄��C�c*�)�L[yx}g��ӻ�v�*���|��8>G��?���b�Vp����/@n����q��.�l����MD=�a!��UQ��t��ȕ�k�8�P�?��a�W�,z��i $2y��c��Ȯ�����Y(�Q���C@��q�^�֕%�]=���ҏ6�_�����S�J��'�-�R��Kid �ܑ<tt����Kc�ޝ6+L��js���^�߹�8-I�I
}ɿ�rvm��h1:Qq&����`=g9p��F�*��B�U�FU��h��l�7 ����|e�0��+�f�`^�j�j�;������o-�G��@f:�ۋ�Y� j$��r��<r��w�@��Be�X�I���٣k��D�ڪ
J����~�߿����#�l5]�9���i.���GW��dl*��T;��!�%�Q��;ߙ��Wj�|bB:�TI�`���i��q7Z�;�Ԣ��p:WP����_Y:c c �g����P���G�@Kր&��V�;J�/d� dJ)5B�֑���|F{<�Q�@��e#��)�s��Et����\y�K��[1���Њ�����Y����T�A��/� w�/ٷ�޷
X�u"˲�`ף�BU#����{:�j{�F��:����:5�w}>D�*�!��1/�b�H�Ӽ�L嚟I8�L��o��Z�V���8�h��Ƣ�XQ��t- ��3 3�?�h�����Y6��w�����L8��Ȏ(v�^�v��R`������G'V&E6E<{C)\N;���(���9N�/�$��σn2����q�i"��M��א�1����nR&RS��fDy�pZ�e�%zs>1��+6�m���}�E,i��XC���y9>Z]�Tc�0�{h��K����Zx��ɂ�No0iX��~�)�ߩߥ�-�iw�w�;�{�D�	���j�tR���E���E��A�bϳP����a�!��R���������,;�y��P�Xݞ
�ԍ�7��j�~u�ꑪ�ƏXw�OQ���bp[�V/��������B��
����̎��S���(6�nt:vi}�hW Yf���=� �:_ɤ	��2�`�s0;ˢ_�	v8+^�������L�0����c
QM�!�ss�n�ib��r}��Ֆ3���- ��mq��jcЕ�$Ɩ�I�Y]�	c�B�!�+X9M�HPH@�Wͦ����7��V�%m����䮙R~w�B�{�Y������G`��`�\�-�)?���ˆ�U�)
Sq���&��nÊ���~�~�54�p2�Mg� ������l�u��?T2�.W�j�U������ڻ09�ǣ�f͗1����
o�e�%��@��wp��L'E30x����fp�=B�"�+8" Ka���ȿ��uu��?�'��8���G�(��֭�R�+���P�9�u�]Q����3��j�q�L��ȸ��Gu�S;g�b�����#{�~�o�f��^׉r�]�HT��r�ڿq��}��ݞ�Xkٚ9����mC�"2�=%k8R�"��7�Be�,x~;-X� �۲�����_� g�= ��pt�TFɏ(�X��@�6:�H���~��KpC+A)F�E�e	��gws�I�%�+ãN!iN������ŭ��r9��Os��T)c���,���f�?��aQ�O�W�4��w_l�׫�Zٳ�;�3w�7e2hc&���	R�d˵��_�� ��f;���ݟ��=��-�@�	����Y��e�Z$�d4����y� -`�юǙΔbsi���K����P�c�QU�=��	�Yv���R�qX͞]�8!�J�FSz~1�>gÅ@�����h�����[�_���W�Lҿ�&� ���%�]�c5ɇ�lEh���:[�l��rt�O`�L9��v��Ts���܃Q	�����b�I��7N����� +�(��z$~���]��Zһ���6���)<4����aB�Bա���&�J>��w!74�wy.wndM]�ڂ�Źȱ�趼��)�e`�crp�� f�����w7�쯫�Y���=��_� 6��p��~�3�'7��D���hḋ������C�gg:۬Yx�\r����J/�\��p�;į���6𴥦z��qtǸxP��cC�ƅ��xC߆l���~�3GP�Wv�r�w���2\`�䁨�����e�N75,x������:���h�)=h��J*m��c�{]�ʪK$�A;�EӿRe1�>^,�+��c������SH`�F.S|�`��eV4�7�2��f�Q!�m�+��I�T�ζ����[���[]'�Up��]�k#�q1�n�{&�
�P	ˢl_�0��[-�7x��zE��
uA{^*������ϐ/�Úd����9������F������>L�b�m�V������1�m�鶪sZɭ'넞 -�}��{R��3&B��}��eh�ZS�Kx��`a��Oh���a"�$�Pq�>�V�B=���Ŷ�É
Xw0��x�	����H��0��o�ڡ������[ j��E�m�|�c(�{�.�.\�FV���J���WKj|�ඒ#ҧ�V�O��悐ZO>��N��(T��A�e��jUGv({+6ÁqF]Գ��xͽeCo}��a+_�B�$�%���U�TG�0�����K<��(��vuS0P��n���s�f���W��Z��{Yp�N{{��
W׀q�ْz�tIĤH�^��I���Mj^��%��4q:?o[�"y� �uq9�z�|�;���%޾���	��l�e�g�������v{O����$ʅ���]s����{@��ϣ�&����i�	8g�e�%�B1�s�u:����%�L@�'"_�9;E�1�b���YI�ЍeM30TW!�i��կ���fcD��i�6K���[Ei>�5�P�8�'�&���ѕ�ض@�!�9t�$E{�p�-�i:�h�t15n1]7�t<N�	�v�u���d��Nm�@ѧ�=޻��.�W<��-���zN�F�&R�SY�˰�9�is��1�W�K�H��T:KU�"xK`�ESA���5�T�m��B����dlo���F(i�����������e��.��=��w�a�F�LN�Yܽ���Г �����k9%{T&��9Xe�]�>J�X3j�(�����uQx�z<%��� �5Z��IG�y���t��'Ė��9	�`i�\Z+���d2�z��:����9�w(�>ZJ�9�ި������o���M r'|���(C��A��|X~�.�<�6�mȿ|o���֏�� � ~���<V���\#�'K�1��R�+��9M�l��;~��f��NR��:un���]=~ɕ�@�»�p,��QӓT4���^�C(<C��F�_S�D}@���U-�t/^��~gPF�v�ʡ�.���ME�f�.a/�-di�ތ_{�m1�����Դx��'���<���nZ��W���i�~���Tr=
�K��ʍ�4֝N���lz���T���?q>+k�w��y�Hd�U�~ݟ^ ��2q��1163�~H,8�>�5�����|��*MM�qOx����GX)ҋ�,���i�|����5��1�xJ��r����� -�
�|iU�T& ���tK���¬f�$��6�X
�2E@$5�.���jW�J|�C���P�=�VQ���N���Yd�3bsջ0�}Q��Kr�x�(J�~
.��[A�(���L�oJ[�#>#D��`H�8�\�%��n��Ð�Y���Tƹ�U����7ܦ��
�Y�菗�yi3qq\7����+v �`f���7���o_����J�	:�G�k٧E�%<�m��:ma��kZ�Q{�d��A�����|�D��y�W�[�%f�'X�`���c�j+0ړ�R�X�k���FM�_1ስ�R�s}:�����1#M�n�@a6g���q�T�O+��~mK^x0a�f������� �s�/w�q�	WL����Q2�ށe��>J��lܸCf���ĥ�R���*��;-T�T�Y'�A�q�9�IΑ�)��ƚ��T���_��������l��\����'Ǜ���G���(�Co�.q�~�KCN�}]Z�;�[�O��y�O��U^�*�c��1��)}��*�z���
���8����js%
�B|V|آ7N������f �;@����*ڜ��,odX���D
8�53[\�2l#h��s$�a
����G�f��)�=��gF���`����8���� 期��w��X7�$�ƅ�]^��)P��h������ �}���⚃v:V�1����(Ψ?�>v��S��)"�|���l��_tx�=���zDE�O�<�yd���+y���
�$�t�§s���k'#0�,��*��e�J��%���Ԁ�-vK�",rQu�V��m &=&9����j�8��X��v}���=��K�H��5�t��)� ��hʖʶ����.u��Om?-x��3[uº���^�` �2U$���GI �-g�����j}ڠ�zSaط�9C� ��r%�c2H݋�<����9K@s!re��#��*�;�
t�s.�T��n��R�
X������=�ݖJ�}��5� ���]�����Vh�nو�1�O7�:$��u��3�� �A�X�u����"����؇�A�Y��;���� ����~�p��,�^T��.>��.��.�����AV�o�56���,�4v�7uA�=�����?��q�|Լ�{�dL��C���n�0���İ"��J3ŗ��<��p�k@2�픐�>����OlM=��P��T��}��`�h�W����;�m�22r��N�Ƭ�8���?�u��~~��1C��ǳ�d�B�T�mO���?%�K�hi�:���Y	��U��Vs.�)*t�4������y��e��.Yj��A	|-r�I�D�0[�MqJZv8c� � ;2U2�]����O%-�o�"-�0Ӷ��5�z�����Zfפ�{�%/09)1����,� �I)�Qu*�T�zW/P����b�/7{:�0;��E�P*l/rfgÏ����z�_s@��1���BE����z�H�~���q��P8*��0{��V%Z�\D�e�1A��[�r�te�w51\��p�R�C��*S��J�i��ŔLw�L0���і[/5�?2�ĨB'�h����)Rrc�+`6畴�:6��1����'�ȩ=�з#@9Wg��N�	}#K`�"k�C�M#�c�8�f0B���/��aZJ��Hzg5aKu�9m�-Es�U����4��h*�^m��]M�t>T@���?=��p{�Qe�"Q`s����� �'s�5��=1��O�N�p�Wl�K��׺�Pl`�A��]�U��*�@�+���d�e�WT��d.�����p|]9��.����@6�ɺs���Ts��MBd��n))*�Gu�������j��7S�zhW��^u�Q�];�L����Hgb�`�Ŵ�΀J���ȝ{2_A�0 ֦y곁���S�l�9;�"ɞrj��j^�!jW]��U�@����~e�;5�Cn��M��������1S�ɋ*�l�4T������{`YGC�|���e
��P��F9Dl6Q��)�#b�:5���#�" ����N�]��&�N���=�ӡu�?�fI^������}�Pø�����ȢX�u(���)ۛ�"�5,w\+�6}]� �%(�8ܣ�1��ݞ����ZH��s��
raf{O�f���X����0�YN��w ID<e�6����t��ђ�0�H3Qem�oj�Y$-R�\li�ݱ6����P�4'0�>���vsxz8Օj6�\�$��(F1�B��P�N���k�m�uT����C��Q����\?��i��A�;)i&�;��I�{}J(��!b8�����S�Įw��b�t`����׻�)?:a��ܖ�.�����k��#QKA�v� z��0�`�9��+��#V. xz�!+�CD9��%S8���:���$6t��A<���X`�=�>n�L���pz�A��T��ѹ_(V�x	��D1�N]�
]�>���cTv�	D?=���ʒ��!�7_#p�b+˧����墟Ar�h����&���f�gN��WC�{��'�ˇ�=xI��e��������T@'>�>P���������l�Ѻ����X�d�:��M��"�	��J��k>C���\H�[+S�dV�7�r�o�DS���=�r1�h�862P\
��/Y�}��=�G?9i�����5mb��ou�Q�V��	y:v����3!�� �>��S����<��~��ϸ�/wA��+
_H�2����z��C7�߼��8��:2�6aR���om+rf��E:Y�,�Z�~4���C�-�y���{C�(��������^:�/"�Y6�J���>�F��T�+ܘ��\��~� h ������;�J�*9^8�\�朧���X�M����f;D�z|��<c0"1�ðǖ�x�M�|�%�g���9D~&$ʵn�mQ�5�[.���j{i��K��Ww��|�u>�t�����5:�����['&I'0�dVZh��(�f�J�e��BFga��tkj|��z�F1�_K�Z=�Uv�����6�05���od����g���t�#��=��ʐY5���/�� ?�
;��^�����e$ԇ�X�V쉁P���A-~���#�"V)�����'�e�hX�tеQ��R��6A���4�VӺ­�Zz,�(�#���.�?��*��E�s�z�sy�@o�����Ã��	w�Օ����=����T�b�Y5�ny�jS`#��ݤ]-]�qˬ���  ���$D�*�k���pq�T}�6/��q�P ��Ԝ��m�9c)��)�F�-�{����R����3[Fn�
Ae�xB2��n0re]Q�McŞ�A�b:�n���Na~�ED&�ے���)0����&>�"|��J�hWU���,�m���%���C/�7����Ns˹����8{Q0����h" /��%9�L�}��#˝� rH�" �_����8
��#����oT�P�r[�5��)9���C����A��/$s�p�{V�]D�X%3ͷ��|����<e���J;�LVO��$N욏�
���O/c�8e�+���+�J~5A���Cy����&�>�#L�cj���p��b߳�mILrUo��{���G�Җ�g�1�*=��gX��O�jk9*
�%*I��y XQƔ��9�5�-:ԒYsG�
���^� 3�ŗ��C	EV ��M�tͩ��h��nr �6��B#|ݞ(�a\�ȯ�6j���>�K8�9�%1{����2?���O�E���'�\�q�z��L,�B5��H0���)/�o޽P�`�[c��GF�Vz�n���>D,��PB����\�E&���)�?�F�JI���@���ƙ ��#�}�֥!G��� �����+�ك��CfTL5�6%|(�u��F�����e(�'8�ۺ(����ٴ��@M���¥&C�_`�i�|/�4��LA���������h�g��^(�oǓ���vw�����dM��n��ئ�������i0�\QbM=Ngo��\��#ހ�� �=ϖ�6�?gF7���l�0���^۹=���>�,�"�����4���Q<�'�_#6���X��{r>�@4�K���	�i�ʠ��d⮷ӹO���%�]E����$�,�ۢ�9^!OP�\:�W��
�;��/�^Լh�\��Q�.���Ĉ��{���,��퍀�;�ݢ�f�Y�J���
,��fk�V�IwxQ'��|��Z$�G^�Z��O�`��o���갃0,r8�3�:1"����뻊V�3&�>�r9k�\��B�[4)�p��)� ��`��X0����R�2CM�G"�C!g��8'mB&ߜю��=~��o:�{�cu�[ژ��:��1��c��7��뢊lfS؟6�\a;j��K(���}4��kH�q�t���`ɬǸI :��v:�P��zBt�I�;c����wQRn�?�<�d�Z�	 �+�ڬ܎��3������w���܇[={:K%h���ߣaf��Iu�z��/�f}�([9V7��
�vC�{w���̷ޔ�k����W{`}�ϝ0J9u���ĕ�g��RI(o&�����C��H�e\c�N��"���oD���u%dSn�..�]	WW�2�P=�:�Ϛy5Ȁ�Tb����v�{z�f�ȇ��G���8S(^�˘@����/T�{�>�U��i(S������a#L넋}8H�K� ���9.��yo��;gQ�:��]tKγ��>9�D� �Yk��q&1O��Ƿ()��9j��y!�7��V����1x<9_�S�1����F��l��j1lf�Ɠ[�F���\�SZ���=O*D*�	�������cn�dP]��(�3���~�f�#�ܫ6 bӥ"��Z��؁� �b�ib���ʥ>Nv��<Tx
�q�ڟߐC��ǝ�y�6b�x�?�}4~�����'+���	�@��:=R�<Ѵm�^��i6�N������ED���EX����NE����6�~c�S��ٺ�,���B��� �<�#�V}8�{���u�K3(K��͙���|��P���)������;�j^���}՟��0�u��h�9�)���6G�� (�����`�͉���+]�����x��H`y����Z1�*�N �3����vty�%���oM��OmVVJ���N�#X�sL~�L㧴��1/�'����f;�c�*�	s!7�y{���}p^��od�K�?G�m�
)n�'t}�A����a��.?�1{�'�	7�����m���kߣX7IP[p}�6o�7��#�����2ˈ�[�*�u�.�������@���؁��`���G�h|�r��	�Xw3v�P	k�_���hx@ȫ�-���Dۓ����&��qE�dW�n!��S����L9��U��Rc�
���\y�{bo\�*9,�U6K�݅ �c3x�@�#wlwԜ��(�[v`����Oٙ9�k�o�É7�mM�FYM�c[�����e���C���-���ۥԚe�21��a�{0-��[���Fl�J���D>N�$Ӡ�Ĥ�(+uKq�����w-yNg�*�O�+g���;��"��J㷵d4wѮAA��G6�����p�P��1� �i̄��S^���i|��v�[ ���� ����w$�y�>v{`M�+dWl�$��
�eXľ?�t��`����h:�MV�;V�~�cۜ	|v�#"�/��!��a}�xvD�i�;�^Sa�S����rp���i�)E���3�����)�|�PX��h����&��r@��ǁ�o�R���3M��17����|S�p6�[��@01�Һ�wf�ZH���c��)m�TCyO����fj sb���>�F,&��嫴�F��u�T���n�	Л59�8"{�0� c�D(��L��D�hT.�k����4��k''L|�?4p�T'ۤt��������@�H�gc��,]1���C�iar�s䭇��2yM&�
��4ܥ�ҀO�<�=z5�.�T��pDsAKV�����|F���K���A��X!�X�ۻ	θ(ۿ���ؚ�q�Z��+������R�L}���m<hܣ������r�ݙ?H;sf7�z�w�ԙI�� 3��r��,�M�ĭz��G��cɵ j���/���^��;���S�}���$m�2�W]�I.YPw@��
@�5��=�h�I��*gA����W�ޔZiR����"��a�C�1�Z�'5V|J�V��J��l�W�G��[�t}�ʰ�8�da�p_�0�f�e�Q��7��ύ����C1n	�x�MC,\��0�[�A�}e�p��mL5�\*�`Ж�.,���KhAM��	��AѪ��
:��P����R��RZ��T��Cw!�𤽥!���adZ8�ߴ/=���I~� ��"Wާ�6��j�!�A���ϕ��{��7�5#H��j��ql;�C��XN�9�w��qJG��y�s��_��Z=ܧ�e�Q��"�<�Y���*�����l�<�)��4�-�-�� 鲯ap�mڪ�������������ǻh�ȃ4�6�����ྖ_� �����,58x�0)!ԝAP���SM���Dʣ.?)v�~ax�l��;��e]�컰\G �r���p�CU�ƪ��:�(̺��>�dŖ5��#�����%r� x7������Pz�~��ۖI[�ii}���z�O:�& X���ܳg�3v��ha�8�2:hS"T�u��O����!ƛ��AGN�+�RR�q-�ޗ�f�F�������vC���2�[�1-�T"�{�,�1WA�2_w&a��<:�{���V��g6��s�.Y\S�owl�a�����=�E�����v�U�x�VEm��ƮC���ҋ�ld�qt$��}�������*)#�6+e���_��;�Z�O�%�|buɎ'@�n��*=�D����B��'TN�cel�m"*m��z�����w9���2ԕ^��[�d{.*�di����Լ)���T�?Wg�բ�9g�v��z�vR�7݌9��/���"([S:QD�I~����t�HT�:�B���=���w�Yݛ��!%H9f��<e)�p��T��b�)g_��UR��Bf9A�0�Hg�+^y�O��Fh��m}5H%|Ӕh�o}����M`�G
��z��#��-g�����-��j�r�x���Om�`�.��t̺K��zjyA����;���%�hCNS�4\�4����*<�Ȍ���(���/�lM�0�=X�ms��P=_F�m�R;]��9��^D<��Zw���@�w�Q�N4m�4����8x'\��\T=O_�7��Y�;��_S� Ֆ�Oӹd/ׅ�����ki���}���g�E�>�%g.���L��<-�3b��"���5����?���(ں��^� �\��U�I���4�9��:�
�r|��fs��1�;S��	8�@m�z0���*�#�V�;�П�,��)�1#]�̜+:��֠I���t����0Z�3$]�a��o4ڿF3�&'+�ZŖY��n;�o�J�)ȆLo�i��9��� ��R�adFր$��?&�v�S)�6��)nt���kL 0vF�`l�Ezo,?Rt���. ��癒]@]e��l�@�@������˒<������N�/�VL�P�rz�v���&f�u��5[��:)F���l�T�X����*�mB�L��Uً� �d�A��Fo��O���H��D=�s�}-���俜\<� E����!e�%;�͘�6ka��Pi�o�����^w+��9ԟ"෕"�*��3�	��@ol���rWՏZ/��,�E������m%�1������r'ޕ�&�>���V=-�G����w� ��$���{c,�.O�)��	.����C��w�zۢ��l	lB|N�5��LR�Zt`��q�Т�މqNSښ��>諆����Jh�V$|uro�9N�Z]C1�w)X5�� �'зNb:�-9lo'��B���fx9�UL_ȳo��/�i� �����>���������]n����C��[Q�W������N���n)��t1j�4Q�`o>��yr�����������|��c�vmok��׾�un�
-����c�_e��M������B>X�s:�T���J��7�JQ�@��w�T��lK����d����=���bm��D���WZc6�Cy���w�5dz��C*��#��r-G�z6�6A��t8����T�I'��P��n�6�'S�aG9����{���Oأ%$����zl���K_�3�="��Cˬ�=)Xo����㼧�+�V��mU�2�Tt��G�&1�Yu��T�x+��kC�e�r<-"ˆ[��i���|��x*ש���k����������_��|�_�����h)	�!����z`�pG_ iR�]��G���`�m������j�BB��LG�}og�G7������p1s��}ka�|�:-J�0�xT�Ih����7l���������ŏ��,��;˹`\�?�V=���]��iz+M�i�*]��V~b��bٵ~���m?��'�V�?1�K�͈A� ��܎G��Z �_�;ק2���V�/��3Ғ���ts�#��t%�]��a:�z&�dR{=?����H�{>{�TC9��i[SQ>�%���;Ѱ`������H�j�;�[�9���t���\垠�O���	={�XE~���hF\�|�9�3�S�S��j���L��9� �S|#A=yɢz�[`���d��0�E3J�UC%�zB���TY!A��^��Q(����(��1D!Lvb��+��{�yqO��u�ͽ�Y��6��I?)�Ӳ*�f����ЦlS]�A�GU5I�07�/�U83s���(�b4K��w%�d��V��-�,#A+��7pb�¯��n����
 �cI��}��J���=)t�\9�U�>\�8���8��z.�����~���0���,�u����%�;$Q�jQta{ԛd�$$�x-V���9Mv�����Lq��������DH�����&oɿ�%TX���l�iE�ԯ� _�+%�{�o4�b�iR�²`��?�`�W�F>���P��}�n����9,;P`�̹/�R�ӌ��csO�l\��@K
/cRB,��DS�v!��v�9��C[��?��ԇ	�
��/�T�Nq]�H��!k��^h��gQY��e3�kI ��#J���G�S13b��k�i�3w�B��2`��>�I�(����k�XA%��r,���5��=��J��:�qp����tU!�WĘ�R�ҍ��ƅ��r�4�t�����" l=K!��:WP�B8�Vd�8T��W7��Էϵ�£�al�Z�<K�"���x��m��ak}nU�K�]��t/AbpKTd�J�+xq��zj.+��[�l�4�Bll@�P�Ug�8m�܍���[7���r/��XLۧb�<`��M�6�5�m�(�U�G��iF�|��$蔮R�R'B�"=澶�`_?��$:�M�������#4Q)���>�r$rt��i��z��ښL��۬�4Iw����F:u���/��^�0u�{��Ρ�V�����K�r,�,� ��g�J�� 2�Ե7�X���@����|���.fߔ�ӥ��������[KF��ݩ���"s��XN�n��cX�;��*M���2����z���Ȋ�]'/l0Z��g�TͿmU���6e5��R\���ð��P[Ӻ��:J�={�&RV.�L��#�5-����2���8ע\��=l(�+�aVN_¶T��}ʰ�"u ���+k��J�\�0�U�욶(�Z8�s|��R�dB�����gB�q�P̃�����[%���^\��Rʏ @�v�w�Sv2H6qY�8�MhL�~h�|�����iq��k^tU��|ҁ1I'�d\��O3͵6�fCwڦb_]�ՖQ���\�� E���=��ʙ6�l���Gr��h�H[Ec���z
���B�qv%wZ_w���hݘ0g݅�X�`�� 5݊>x�h�#D�ե�!��X�cu}B�4j�����$�yF=�a���;Oo�����i[�7��=u|a}�LI��jZoZ\����B���@єFXb�,��Jd�jϩp���m���Fk�Y��G �ρ4\Fo�f�1N@�d����iM���h���O��<X/�	������"�h�널y ���B�!d�g�qb7#;o*l�^0,�D�α;)�V^��򼞩��|��j]���yUp�O�+�T��T��.bT�vʬ2�m���
�}�D�L���zkFp#��~��������X�#��P�%FA�b����-��FxgE� ��L;�hKW�5��,�/6E]TP�Qm�)F���d/�3�Ӫ%���w8:����$x
71�KҀ�aP�~Bf��OA '�ػ�ΨDhLF���쿙e�IJց��נ�E^삉k�y�MjǪ]�iq��f��-M�HEyPIs���;0��g��|�2?`y0��D��̳�bZ%Ȩ�-t�l�c�R�����R�?޺s �(�_P���5e��x�1�a�t��B��YN�b�$:[�ޥ�}q4�4Sմzǣ�'�n�]������;���&f�ss�K�pR0~zj�MI\{ �yP� �Qߌs�j�ޓ��v��P0E��IEec�I[��h�>�iu��q�DG�'4o�arc-�#y4?�z�"kޯ}��-ؕ�|��m�r�m�4�.km�H�H��t@=����j��u�L��1	$q\�I�<l$e~�lE�*z'��~�� 0B�p����X޵��lm.u</P�9;M��"O߾���LB��1� >��e��� 0�c�kb����03�m��`Qq�KJ�T;���\��6(q�s�O9��h���Q;D'2��yD�R���X�a��P)TxiU��4�2y�az�Q�]��&~ `xX����e\��+�z��ς�ڐ���3�qA/Ꚑ�� ���7nG�&�y2�����Y�u �#�y���e���{-x��J�ч�4&J��$yd1lm�����r"#��#\S��ʎ}�FhƳ��L�9��7r4�
�0����Ҷ}1.8�!i��e��� F
��[�|�ڮ��2����ތ�M
���)���w����Ս����{g؇�UIU�$�J�x�����F���s��{%�~UJ������]���Dg$��O'A?��@���iv����˶Gv��[0^�ۏ?�G�ȓ�
��5�C��3�2|,��">��@���[��9u#�2��D�ēc��
���oǛ��͵C�JX�>Z�H�a4B��8��۫c�ë"��;' ���6Yt��Z�#5m���=��{ӑ���l'Z5q�)L��dD��b��D�o��YP��B[C�ey�_�4H0�~�F�:��.{�j���1�͞�˴\���۾����vZM�G6���P�[Bm�,���d��<��u_$�@Yͺ d�� �6��L'������m����ytm ���n�jc>ڽ�Al� �B���	*z�^#�/)b�
s]ɧU����Z�����^�<A�F���%LZu�6n��ey|��ĸ�y����|jU��{�q� <����z.��o�GI��`���w��^�
K_��0`w����+�F��bj�1�KV�A��s�/�m�Q\�=���V�,$Gͽ����i��XØF_��
���h���^��� �77�c�l�LN_P���vms��k$�F�\�tnD1%X?�^94��0�,�>���Q� ,#w�&�,J�6]5� ϋ4,l�	g}��j��6��I�B��d-��� �E����q�/^1��'f�l2;�m��ץ_���:��:T��L2�2�B1�����h"���a�#�qP$6Vtt#�M��#c?Oa����N����t3��?]g%2`e咒ۣܓ�4�d2�j%�3P �m�vx7ب��`��j�Ә��\^0����ױ`�X�Ϋ���ѻ���u!�e����po�����_���� �<װH��9�GDtJ�Q�l���=�q/�W�_��3��~ tz������ �3=�2cĵ���J2)�E0^b4gR���^�L����rB�e���-���P�-)M�)?��#��͉&��U�3R[� m���Uc���\}_>Co/�HN��-�?��^�T���@әw��^�i���t��D���_�Y��/��؛�	o�����o���B�E�.%\_�,Wc����������tF��Ni�y7'z�]w�S^��Ie���aFƤ�d�n�6@$r=��~�ᨭ�j�q[���A�x9"�//��\l7�C���v�#AX��,�e(&m�θ!��G���`S��c�#a �	�����Жy���f�ry���LɑJьY7�A���d%u���J���M�x[���p��-[����HJ"Z�����=�t��&���v��t����/�iɸ�#�[��z�7��\V���	rڥ(�!;h;�0(�og�is�/[;]�;���a���#=*�#$sp����_k�x�K�l*;W�_w%�ˈ^ȋ�%І�N��v��c���6gc(�j<յ�eMB�l!�Cc�*��QD.�Ɓ��TT��I�r^C������퉪5O�_��;��W�Lj����5�~�J�D?˃[%�A=�,�;������nFJ&^ͻdn��*�=&�į� dS��l�y�vAE�;I�W��ᅩd��V�\\W%���A�eEЂS�5ۊt��@x=]�ӸФ���SJ]��p�Ws��;sЬ���ݵ!I���f��U)�<!�ϊs�T�Cֻr�;64X��p'4$�i���+�����>�a!���#�O�ZJaS���?�Ó4���~�ތ�'A� k0�M����Y	�����(@�
�\P�<J�7�o�{̏�c�yp�P����SS]I=9���b�X'��G˙/ՐQ���2=���jn{C���d\�P��J%��o�m��Z��h��-��:��E����4�>Q�lǭg��Ͱ�L�u"� �qa�_�ٙ���F���`�i�(�!Z�s��GF�S��y|.ev������Dg��`}��C�r���i��	u���i(kN�25�-JM�����٥��K�힋�sq�M��'���o��_�e��kX�2+���s
b����Vn���EC-��R�:b:[����mq��X��%��7�O>���tm�Xy1��S�W�WO!��FP��]b#�hѸ��pS��^0���9���F�H�Y�&I����#)��*q�U
���Z&{�Um'���Ix~��&G˄��(�ԓ�]�!j	�-r\
���?��z������U깢�O��Ə�2\��P�|��wa�^�ܫ�&Ge����x��<�P�c���N�C�J��(8��0��J#,�ʄs��>>�e��P+�8�r�Ο����K��F ���쫆��ּ}�T��B,c�XFy�)�X=���5Q,��jQH�z]�bK�BB���V���pu������@}��\l�\c�ݣ�{)�����P�Y�W�T֨h-�5=�[N�/L�T[�K0"^�H����\~��o.b,>����I���Y��]@�{��K��[ΐ���h\ Y�f4!���؝�dT)�D˒���̉U��� ���>_�aۇ�����mR�#���%0�cl쐵_��d���〉IU��B�>88���t2Z�Қ%,V�J�W��m���HF�HV݄gHt�:F[s�f��.�}��TfY�� e�
�Ow��1��G�Lp�E<�ܺ���)]q�id|���a���c��-�/�4�$���g�U����?�%�5T��Tb�4ڈ�7��cFp���$�J���k������2�0��ڒ�(���４)�@�K��ׂZ��
&����0�rt�~��l�Rmx����aI�oB���8>��6���:��T�3����7Ɔ;��k��������,���������h`�4��e8�I9�D�a}��xj�!toQ�	��2e��!1>��>�"�2���#�в��!w򵀭�`�O��pN��!ٝ#�#|��q\S�����:^)�9ߐzwi��
N�q~�>؈7�wVJ7^L���/I����s,�r��:�aAV�Ew���i~
�{d5S3��%s�|�d�0�3&��N#U+e�c��8�P��ϲе#,Fб'�dn�b�JT��fg�sə}z@ggָ}��e^�+��B��V��ƛ���,D��;��z;� 'l���1��,=�L���y�%䯦Oz�8�B��Ka\�s~���/�+&S�u�+q�h�
�~"R��%�j/�E!Kx�M����$l,,"��q��f�#'U�S�C!��������ź�:�4�9���P|���V&�ɋ��(��c0W��l�>&]�;Üݸ�fG&]}��=����J�:�l���o�Op�����u�6����$�v��v���ϒ�p���t0L��H\X���1�����|��	i�/�}|i!Vt��"�`]��i18^Z��h�MR<�9��>^p���p�{q�8�q�L���d�7~�;(�u4����dJ��}ٕ1��)�	=����.�;��,$<G(���,��\ֵ�^�bgl��1	��1}'�������!@��s�??%U_}�향!ȴN��Í0D�Pi�q�%c��^	��h"�(z�O��}�[��fۊ�����HC��_�)1���]d��(��ȱ�}2ҳ��w�3%�枲 �/������ Ξ�J��	.��K><���?Kթl�h�i�
c�σغ �h�c��M��b�{�¬��4,s��`�	�Qz��C�ꑄ�
�+��D�����E�'�/��)`*�qC矄�CΑ�[{3T�"f� T~_\I.Yb������m�c���E�����O�-QڨJ�&�g������a�����幯�N�^t���>U�(�DS�����s�7��ߜ����{pa�$A��Z�b�q)��݉N� y]���bX4 �B�޵M4��.��6��#I"ٞ�4� �{֖�n#�m,�}��&�|�
�G#��'�W�$�)�C��2'�,��)(�`����Y9̰3�����f0�a�$���e/���5���}��j�HQ����F)�Z��r�x��"N[�˗�3"����I^��9".�i�>��&9XsG�Gr ���bqU�b"� �b��G8���j�Wo���v\���K9����TFI������/�Dn)-��'WH0�g�g^���Ӊ<ֻg��U���,Q�M��xit�&#R�i=��ϫ|�.*�2A�O�	�V�R���m�!�.E�,����jeE�u}r�ɗ�x��c�3>эN��V����靝�wY���r:�=�`Pb��� ��Kn�'Opv.��e�U�ɂT�)8Z=%^��lb����ƹ��	������4���N��{�o�z��-���0FK�N�qE�}JG �'�ê��W�'W�b.�D���F-ޝ8!�i#��f�~򩈘 u��Q���{O'����v��AJ�4��hC�"��Q��3VI����G.�4��zB�a�7FN�O��{��PՋe���?*�W������4<K�*줹*}�~~5�^�޷����zc$���3G��ݛ�?~T���V��.����#Q���^ǼA'����|�fI�PIq�.Z1-�2�'o�۴H�~j���8���m{�� �Wù��X�tܶ�}_��A��2=:1�8Y�xy$�,�R٨���]cU�@v�bT!�������o��7IW�.���o�ҝ� Õ�#t��������|�v�o}*�>5+�z�&/�`��-�5�5�����|�'m`�����(a�Ͻ��@�)��xF:	�lM�ʊ��ϛ���]�'�xFN9��>�;s���W��>+�=/*|���w�U1�؍j���h���p0SPj��Iަ���C&j8�sQ�5|äT��� Su�DOVC
R#~'U�o�S���@�!�Y�5���Q���n,mp� �v�������Va�r] �=F��t��ު8j.r�����fpS�k�M��B
���)�pYyJm��qm��2��8�v����҄d/�O�$;�
���3?��7�ࢹɓϮ��1=�^G���oMtl�٣ܲ� 4�H�3�/���|	�/C�[�g�O���-_�aͅw~�F�u�k^  �"&u����]+	Ψ��wo��B���CSi��i�#�����Ϊ-`c>��iěv��$���s��0.���2�*���J_�a�o�wMk��e��.�Yf��C����YA������&���Z1*<�֨��
�p��7KWyr�L7K���"arPdǫ R{a�wdb�?�|��h� ~���>]���b>�����/��R9����E�h;�)��;���-�@��� Y1��8��Ҁ�>��#�J�K.Ab;�¯Q�����d���~�=��@���bm���[��q���p,��� Wk<hc�86��;����[�ӗ&�l!T��n�pe��T�6��Fl��X 3���Tc�"��"��w����u-��^6��<(����ww ���ƛ�j'��re7����y�gp��T��'�&F�P�G3|���NA9*H`6�ǩ,�0]g��Z	;c�b��]5Hb���Ch"vb܁G�P\����$����!��o�e�+�W����E �Drt��S�>i�/��w���Ui$���[N-�Fk���x���	�����;A��E׈D;�C+Hi�������+�5j����yx�3�r��;*OV�O�,�r�o	��ɠ'���vP��������N;��z�^��]K��H��d]���hEP����b�0ˋ��N�m�+�L�u���>��KPNՆ��[a�w��I?���Ԃٍ�<��f��%/!���`°S"<0��i���F�-9H�A^=[{��a~A�=`2�}����?𦖍�Q,�(@��s�����:�3tҐ�
>&�횊�9s�;��U����FD�-_�	�5At�0�|�K�0���H�����Gj�����Q<�,S���	%f�1}X��� ������:���p���$i���ᜯ������=1P���`��/�W9T��s��](�����VP$��6�mGic��i�w�?7c��_	͘X���y&�����cH�J"4�4�Md�iEl�;Щ��lӚ��%s����/~6�(��~D�ɩb�66���Cz�YILUG�iz`KgMP�R���xۘXB9�fZ�,$7�� 1]�Cq��$/�gz��z���w��9;.�3�4�t�S��}r1�%D�1/~�
�)VX���țs��^l	$)���%,���F��Mx1�z��l�u��8���z���m���t#�٨>����ڧw���a�F�:kF�qk�G᧮ ]T�#�|�a'�U��ny���JZ�)����ok����ŪޙW<�ě����Y�<�0��-\z&�������XP�2���SP��%�L(:PV��`�(l hGe,�P~gJR�^^�DP~��}[ܻ�6��7}����Rm�$�AX]��M&i
�����lNuYPC*��cm��15w��Cy�l�AA����h�ҕ!t�U*�+�-��*�А� o�qF���
7���G0�i��gs+(��"t^���۾�-���S������H+$	)������;LMB�Fa�&���W�����XI�� Ww6��>�5��-����W�%��x���uw�aK]4�������(�R:��3<NL}���L�[�UON��O�:j�Ez�f��qTS	50Ȍw�d5��aQ]��#���N��?\�"�#K�%e�������>��!�O�g��T��n���פ�(��� +��{}�:�z�q#�k!ς�����/��G��'�e�@����;u�g��q�j�j&�