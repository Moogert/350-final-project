-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
15+MG+qYcE4kefm9CNxPaRL3Pp1wkVNIQjF+xz8bgQ6q+SvVbb59AxUP8Wb+g4q3iif50i5rgDfr
npjMzNXH/Qs+dgwKZ2gOJ6yhqnW4Lku49jskd0GXlGGXA7wY7GlWnXl2rYCqNpPWhkK58dbQYYDC
rT+WgJ+/B2OFE0lEGCDGUOoGDCGLIunrC3xLEnFib+axRN2I2bdFpJx4efWxwckz4xrqbkvPbvMO
MBLqv+oBOleKRr3qRKvjGIfUdUewoZdEgbglYxz/kjqSRtu4yy/wFBeBaDYWLVersx0csoz1WXzu
lhKzY91v/+aQ5EvQgbCZguhUIU/aExTf1Nt0ig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
Hqbxa3cg99N7hSNRnYSoijAkN/IogwvUMjMhqbfbSQgMpTCJJOZEJinddxXCGkop7VqepoZJ+Y2A
lv6WETfvMiqgtFeRRi+Yl5Z4RGWYInaZ802DiUf09bxA3SNnN+CQnK4QHP42rvufBZMzS2003+4e
09OeAKk/luZLXS5STJVhiuVFdou2zPX+m0dPZCuUaCcSOkK54EO6EOei/Z4Pjn1aA5axw62V9u/e
INSLvHqkra7EzxmLyWzUtd7/+dqxD29S7QiIO7Yhlie5EKMiv8flkRnzVC3sEdc4nQ1MqTGrVYp7
5lbSFWGUJYlGbAOysEcfamaQAW5cMg+lUF9ps5PtKuY0PYcqxQ6DSb/N7tJUwEfHMgBVfjgyEnCf
1nk6NC1AQlGOu7UZoMQKzFhhrR1Tl0FCKgmHGN/k08EOQJSR0FbXyZEsYp5II1xHEtrp8hvv48ov
PFOZGbZT0XsZMTUvHutzBWwjmQaWLkvGyXDMKLHtV4oJSt63sO95ANFlCaZEqDGnIFJKsnUiiyAk
SlooVXbltDTtBqoVCA1rmLqsUD3AN1ga/Y2UrwS5q5KF1N+qkWAFBTAmEAPOX6OigDiUa7OTAo5d
Ee2NvCmW/QzIESCwa9anSVN6P9hEL8Lih+P715fpZzl1sMc4KdsQJO6/nXQEbPcQY5s1lLp1Afto
zWL02CtFIHv4B4/Y7zsNuDUfkhHdo+7VfY6Y5UXLw6A6PQaSyzW9x2olH7fZoGJLodimyimss20M
nc+Uqyiq6OxdnkZUmelDjzBJEkj8wwR/SLn7pdcwE6JyEftYVuh9Qbykn+16eJoWmsln+cEr5Q8k
8lsyCOGeIcMoad1M6lnFqADUz9Oc3b2wVI4osN8QPDTo3capxMvCxcZms8Iuyzfl0w8qyEP6d980
Ft1vITT1dwNsiP4XkPlnARTTt9gOnrycUhFM1pDig9TDwXNiSsSblrXveTiTlkABpZxUxg5NlmWZ
IxuA3CJdxFGrMLI5GOAaSX2wmBYmaPI+PLGpeitJ7sQcuvLLAB6pNXOdu5zMEHbQoZ5lqRGaKbje
Mf1HtwbUIkC3JPEwSYuJExrjW6yRSBbMoNFttp5Y01kxGhBJvnnpp34B8VCwUWxM+rgSJHSKv9+4
w8A0kOlOiPeDae0vsx31t0cygmMuYxMKsikchu47MSEm47v+30JGEEfAVypFuJPh+Hiz60v/zu6s
iEiyvBYVaazgVf8CkfXxyxdRp9qRpGpGU7Yw1Y3QmzudeRkxX3Z3n2ZyBSx8s/mzGS6s+aZy86Z/
pxJA8Q39U8OLXh5ODrJvFzkfkNylc8pTt1EdyYOQ4oFwYpETl6AY0Ck0g6rTbXEfHmuzFJXGMeE3
rICsCAWfGGeYEWucjQG7wL0yTbk5zB46sCsydkoX1YFB1LedB1lf0Amh+D9ca7A+3gYAR3Mrh97t
GBRWEcrexlAeQ3bKhJBUwSddxe2I9ApCU2p5LUpeyA3yzJHCLyDRukYCjiHqXzjQnkq8EPYmXe34
tC+ry0mxkbKQHSBwHIP8/FUShLZiygnOXX+HoO34JGOq9fJBxEV9KZbloUcr4yfHGE6wDAPpgoXM
tiaMQyB+Rf5Jk2tly6IaV9JmKLX70SFn1h7Mq595Tl+JXO2LOdg0LOlpH7SrJjKRSYEonJOIV7yO
Sls4NZdleawh8vrNhMxub4aGdcwIrEBus8P5eSlGsUkW6nJ6YELrtti/cfBhPdozAgIGJNXi3jI8
UyfD2/5SaNodOaPPQmT9eoGoB1NGnAcOYxDgYdYanBa83tC4z1RgVWKB90FJlAIRj1k9Wqua1C6B
XgoFQGNa+mCpDcE/jmdpu+bkmKtmArfTCss6kGtKI8ktOmKQ82llPBhHtXnKFXz2EA+6mP5plLOJ
8nHsIp0kGgGYz8v669fBj3MEJQTQcFD+0hl8hWKVpbHX9vN6W3UOC4/3WdECBW27+0NvBIfLBiId
PfhBqHYgCO5qXXnmGSzYGpM7t5UhHVQF0VZ75RtB/n6cPviK1/ucNXoUgwndVr7taZyp3gagbkCD
RVyh0ImhtsBuFQiTd7D1qjXJuKTFGvlGEV3qRTSffrc4mzoZZ7fRldTuhAD1p7aG41X8RdGRa68O
3jI2B32HzaPCHSL4cO2KkxxxEQXctbfJwDpZRO8KjdeFCqg9R1/PV6pdzHfxBtVyYe5TbDRoT+Uc
DQXUoIESbEzRoMPdDH935AoYpdnF4UQp7wHio0ik4o4wXybNg6F3DsrbfPu3/Jxe6Sd2T3KCrYuN
+ZEbmhVmHu2ciCQQqFMB4pKwlM8p1C3lIqo73IP/TP8TWAVmA628+AlS0hZbKcE2ijGzKBzvn+JG
VAmQwWgj2ixPQ6MpR9M/3TFgCwkcgal0Om7wKixU+uPkpwITo+rlIMZie6GVouhjgiAK2RMvIp6P
xuUAfueDM3DryxvhVQPIDEVu/NyFCk1Pygo/IZU5fjEr7ZwMZfBUH97Kee7q8GClz62j0hkRKa2v
7ERlMw8Dp/qteAOMWxTCEiuNqTCw3qx0Bi14Jj+TJ7VftpBA63JVM0vCsK0sbftz4YRiMxydPTJC
O05PpISdCOYjVUInJmyln/xyyGjVoNMuJeuNF/YYPt+mj5uLlH8L4M2uwbiKzvdFSYmG0kiQXCWD
yhaWqB84chFQ3IXQQpWDRJ3v30YKx7Vc8k9zJASR5jMXRj6q/sRq3bzy5Y9SX+t5o64Zyxa1Zdwf
AP9D9VNznEcRhd+ISRmUSWSsBfv4PiYXmE6okeyWSIwfk6ZUg33u1Li1zi3JRttsAc86t6V0z5ue
/YPjjlifqXWvGGedw4+iBHk2HFKQTMdnnKQVen5CYhzO1CoGR28RKtH/X8aMYx/6+2/hYrQItWyN
irvHYaZGC7xS0pvk/Rn72oUL5ouO6HjSHOQn5g17BH4GJ3xm/h/oiUyAwWCaeWMrXMXElHJOyJvY
aTyOiPmUdBW/iAaobMbUhKZ0GjVeQKYDYIG+qO0JRs0Ikv1LMbtc9Ox9LBEd3mys29kAhieHc+jU
AoGEDFui6ZlphdARf0I8sEZX7HguZ6PziOw2chVMMrqIf1LSdizOm7Vt71y11vWVF8K/SS3HmmBf
ElDuoFqV9NpbXlWluoNvMIJFXJrPGMfQuYBAHb33TrEAujb/yYRriQ3r+bKTLtSoExcOTmLlvT/w
ReHl/JdeFyR+RmgvF4F4oEvGGRgWQaIf2LjoPI61gaFVLnAliyofidz4WXghBtgmLDz96AajecqR
3wN9/Omq+c8+XQgSUN5qVkYeOBlNqx3q/sq7NefKuzaEnQLHrBGnPJ0dz7JiXsxEInLiXWQGkyhb
1XBaGJtp1uv8IdJxfQ00kRQi+mEi2XR3AEe4x4slEy4Wk6qx6+MGPOvOtM+Z4Ibl+2/1XRuCHHDu
GNBt78fCgZZvZpL5PwLMuILBsL8JoVcmgpu54TepqYhhy8L2o92YNTMkH7Vn6Z4HIwZ9nbzRZ2xb
Icdhv7tBUscuBN/d+GYyiY04MwvahwSvAN8z9uZmNWGDdfENvtHZEYyC5iDEYjoL4DqGOAHWUzTf
3RwhpjX6KJSodyr6rwZTAg5om3fWla43lqliqS/YGi1E1L4n+X5HyQPzXcGOkqCkclKWFeiXi93b
2Ro1i5j7JHvBOLL7jOrI78mxhpfEwCt6UNzaNVK/gdwpujoxsLBE09IMY77dJcmDjDFGbSPRRn3Q
K+ViTCQpp2bbAO6cxJTTekGb/onyqaPi12tSre0aaEp+rJP1FHWCXqUbc6JD1QyMSK6sptzIKnlQ
++wGNAg+5yqbTJC9OObtBJyhCofjGAjPImfpOvcp0f8B+Vd6iBdO9Hf/47fSvsVmL0NetZLseVXf
EcReDzcDwG7K7TafoEiAObkm2Wwgq3qJD2fpbcNX8ucfAXjCBSw7AY1UNZqTnmG+ODSiKD7RY8HC
xVhdGNkBFSs5Mj/ahlkAQ3t4hZSj8xOAyryBy1FUVfc+tUg0S5WUeWM8384+wbE5OcnxsynV7XjN
h8mxpKd7Sm/oW3ZtVZk8BEZom8HF5np/W4GeUJnu99ir2dRlEfp7NxcFl+B5h8hXn2VWPYs/iWQy
ymK2uA7+eiThG9aVAOXHWMtg4KeqObsT7tpM3vXnrBpyJtoExqcJAD5inAy9DY8HvyWvBiX15YRN
g2JxVN+K6UMX7QJTx3PX/KPtjIPPJmTXsvH4mR349gJCIxbwv7U598lzoszjmT5LDPdmKfz5mZ4p
5a1b1asdJZB0cDfU+Z9BXGDC8ACQ/KwRC2RMdE8mVX2WghEJ35VZDf64NYLco9TbqSPqzjdxOv/w
wlFejUPTtXflTo9P0CadnUfIp7eX60YjzUd37eLKpMIDxP3kA/a1MnT/Bom+vJrnrip+0cNwf3kF
Os29vJrNFaHyo33G21eAit7vNeiHSbseRSxhLCnDkvMEHk22np+m3znriKN9969qHW3XskWpAr6Q
0K1Pgz6EoKqGdQx9HS6cTOfgDo73Fm5pw8g/a1Svw7+L1YUFG9MklWsMnWt/uG08ucMYSEYs+ZXb
pB5VdbtOx3GiNtt3rnGjQ+oONgZBCMQsmsJfuZiAWuTAHJOQfQDThAwBWWhIePG2FTkwtaNUSr0S
LuuG8nF+GOrGxnkOQnP9SycJ7UWGX0JQBZOTQyHq6JomoCMSdZsdU8xdL81H0F7XPzo2uUeQF7gO
ohr+9PHyMKC7M3U0/WwfsEdi0/BM3+sTI3VG+5WqRkI+4cftayACCNw50r8hGxFCVFnl7WDKUg2O
vxuIeMHJmcNVs7hcMC8iHrb/Vf1HjJk1RrFx/970xGspd7pn1IQiDv/XXEhHtfmbeJrbfrxlgOF0
vGH/GSdSSkHm+85zngCS0D5PBLPgOTl2ci3NU/MS0zVeTC3+/FrvBFtsYsgq0PnA3UV7hQc5S7rs
thINFXsTR10Z+L6DT5x5SR7TW8fqQWvbr6P0oLsD7Fwy52IoikvD5jhwWLaB0s6keq/s+ABNM/1Y
LcQ4NyX2kyXM486ldwJ0mmqoP9CVD8y5jipdVFs6eSWxZ9EfYczDz9TRplAeyvsYutbi3VZgfvln
CZlf67nDPLEt2eo9rGAQbNLMNBibzgIBkM8kVe7sBkb2OyC37u1Gd5Nu9hbGUCqbqiWzEdMuBbuJ
g71/aHaDhOl8oBjbsSuVopPIn3/GDPDMavRPJNT72LfLXkp0wuICiOnf67ZOGKKWaY+1KghdxkK4
3gIuNo3M73vCdeajBZjrt3GRz79K/YJUIgo4feBLsehx1HoLpwhws5Hh08uzGBv1xNDiJccis4FQ
jB/fJWk7GQaKg8AbDj1McoE4nioBfIePxtVrVe5g+dmdZM0tJZszh6fkuVcXiOvUozD85qKSyY6Q
L8Vta1o4jy1J/6cXypaT7tthj8ktH+KhttOzM2Yekh1ImhYaCJH60cIlfSf3NdvyEAxcdHXJIJH3
C0TSvy8FY+ju+f/iAwaM9WbDmvKxJ6dhmnWxclKe7nrhpxBWaOG0zVBKlKUzDGBHXX1qJHb+M88X
JTSi4QHvs/rmJIQXKji6RLiA9ISKNYY8kr0vkfBm2JNMPVP3khXBD5DRAikt/3+8ESgO7GKneU94
cqdHKpoRkrjTnzRYzilwTIVNYR6Monm33avbAkH3IfERALE0tBhFwjo/iXjXA2AwyitdUGwjRhrq
91Zr86ko6SUkCDNkwLPlebtUO5o01pFNea0699IsuihSK063EikoJUEQDH3WPEzNb2zhSCrUDcly
Rhgpwsa1kx7CLdXtmdft0c4LzkIYgPlmPYn+hFWlzBTFbES7KaXeKWr188Tyn59qXA1TA8aj34Rn
H/56WSMxxBiqX6Gpnl2VUlepoBioFJ7v3o9pYpH6xmFTlrEw9Zs/6NltOHNafS730POZzt1/f29s
FVUCd7eN7u3Mb2azvIi53+tw/wucnGTBPQt3cxWJp5k6fwVtB+t+0WH5IrW+9yDpio2Xfkcv7hq1
F4koE/p3QlJZ/coJm1PzRq6+NYtAvL8BNqddVY8nO+10VPDDrNeZGd7aWf+WrWiLmzibwuadV+QK
HX8eCN91mdWzGxONSNQqiP9PAg5dN4yi0D8V4IfB+ezPlTfs7+xYcaJPPFEBwvRpg+rXK47Grttk
mYH1h923iXY/Li2SV0R8Y3ze6qmDq8jHMmw4XuYZv/ZCbTNxOKD3n6sd0iXLeliVEEseO/VDYw==
`protect end_protected
