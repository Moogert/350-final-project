-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
G2K+9jff2liAeUf1xhrliVltt/6iLnzrPhe2SnRF8BbhcsUzUIxVHMUq4zpZPLDe1/AWLlnIqG3e
6vmm6WhBdUj/3n0Onlp4AGUFNQJxEi/i1sLPYn+T7EcJV3Ra8dmWyNc/HF3oI0ytgeQNFCUK7trM
iELwlrIdqlZ1PjOWoiR+/rgnN1mguBm4bk8uJgVSVhfWnsxM5m0ggPWg1HoP+Cumq4hKqTGqqi1O
cu+dt/TQMNDw6tBOpKc0YhaQAcLLCRAyPnuDCEkAiIxfXfoSRvdDLdJ+clGvD3ndvcMui/We+WO6
DaOaJtpWWFsXlVEwSc1dpwmfCy33bGv5U0xj/Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
aJb/YHyzpWfPh09W5udRdIUc6AMDEL4SLqggNy+eaFT+BkHxkqUz1ihfLiW9Ldr8jV4GcExVhOit
psrpuoKt5sOyEfZWAzKxcXuijrXS3vm2vK3VsDf2/NsRLo55Dzn18YAI2OWm6kqAxJrwIAByueZa
JMFoDRlRnHOQw+39+np4miwTXiMunQLe2Npi2Fun8P0Y38qJnTytdKH2dHLhEfH0t4wkox47TFKr
87s8uDlqVm6ldp+Z5ig5EWV7bOwhjewos/wQQ0MPsQOu/rA0qC4iB4UhDsaKPfsWJORaulFfWHmp
5YrjUzs3GBF8gpMA8Vh/dm3Hfn+KSnlsqIiJrRzJDLaR0nnerRkbRfRINZMhYIOS81xVbyV+FX58
EaY+g/zWJylDcKQJrxd2rhHBAjg8HDdzxNygLAuBrZz127zm90R7E9YfhFDDncvNzKk+G8R6TSpD
L3DTOyLbx3CW5xaagcUHzIjth7PSlNXBVevgMITAD8GEFp2QpmXUfY8j5rSslEljY+XMdX3Py2VX
4ak2ooK7blVohTxxP3Oxg67pbWQTbP3qfAydDuOOSX5wPU6jEru+Eo7xKILd52vuTmsU9wWaLlRi
ExZbyQCRo6G9UPgGJaGz6IusWXOagby4iZSlG2xgTWIT1upcngjt2yN0BBc0SALARkJHNuouI45K
xasMhAnSI871yDib6RRFJJtMPGtHm6jtpqVqfjP8SYnZZNHJ/P5EjvKsBtd5CSiSPCMzDYsWLtmN
lKwtc4uCl0mBtDoEkKaCRmf0Domqsktd86PXrvBelKUpzvMYsu+Da1+a9PTDWDBmUzwvUhq0PIVh
0is/uwHzMBolWglpF2rvJ6kinQFz8eRuqvd0+KtpKoLJdHwfAhteXxUneQWgSajvKxOB4yixOx9E
XJg4r2sA+UX3LFHrIDlRz5uhHTg7kriN8WjsmxHVIVkQXoEON89l6L5Ik0i7gh6T7ybt3pfYY/Lx
FmgsXJIeymGNjqq2gl+hZC+TQwFDFrXV4qfnrroVbK+TeMSyA1SU/VCejj0cc7bU06vx6XuaGacE
Z9haSy2gUrS8iGbTc+7PwAX9ia5yEBEk/PTG06gj12WU4Abqf9cesnD4GszkM7wQ69DxDJ9i4312
VOT+jPxMnBG0S7LKj0yuDgnD2ghtSI4txYEDjlz+mAk+TeENDBfqxBmEWOMsSLD9BrFC+x8WC6ZJ
O6qk88sAO/+QbsBp9VGinTG3INRN9U+OTI3NAyz2tEkwCPCWEJDd4yGEapqo+7uB6GPKJpwq3WGn
XH4RG2MxR/em5//qBGrWwhPEzbx/5TU7TS7WF0ljIJmadwzB/PyF+bGHCgHkzOglR11/tjnykFx+
AMFtDbdQsf/PPI5XhH0k1AWAJ7bkXSjBAvU1fSpRsKySDR2wDdNMscqz7F067r2pzl/dR2oVbqvC
AwDDVjrXLZLdAtTmG7Okad8jEgUqyiovkl3UIAoY5m2FV0xG34kKzY0oSG5nNgrKwovsFf/UNCjc
lXG/aKuG8rhUAsZFaBszQ18bqiIt20YPq2i8SzyUs5TUmZIm8o9asECNvrHJNwfK2KdOWyG5weZd
X30T0OnLx33NcihlhghtpCwG/qyAi3w7KUH/MptLDR8NegLkyEIkmZSoIcml+xnvvcWqhMG0RDDW
IF9NcvIP9XbcnPN8mlGeEQ0HfTUrTfpQ6Wx4oSOp22Dpru7SagogtM5lVsJ5bT8bNxOsQZfXyOEE
f16Tf7PbR3Woyrf2m+t0cAHxlzHjTOD+NLCi6DumAsctoU/W+M1GXucdTZPLibgPZArEGYIIUg/n
6l3z5YuTg+sSkUEEQJh4oqLVkcXHN5AwRGG5l8ciXxUYOf5RnmWw1hkozBk4uk6jQ1QnCjjvZQLa
0cgTTGXBhN1PFDToI5eZlEjqnfUOYMCrx+4AAP8uNtxqVYiGbSj7amM501wMHMQ0ZTINOoSni6e8
upmX4tsC/Y3cepvhNgpqaOz3E0vcRFrsYv2yIKTGxYjiWLQjoV2UyKF0VsFSSzUlU1tAYvMWIkaw
5yjJp3TF9t8qafZw4opIhMAOYdFEF2lwmhaA5OW+S/OtTLLa/G3DP2i+Kr+Z/XirOprq96TFkaMK
cqhs+e4xm0UBdYn3CnD9zCK0Zg8c7Y6NmPoTUbZO/MwH4M2tmT9upFSouQUq7ZFQmtWzGRZq5VUN
XMC29l99ovFgba6vg2o3NffS40Pgu9gZILCFtU+Ax6rzXZ8ADhJ5HL1uCtYYKWwpXOzA2ft79eOx
Deiw9TTqwVw1XAqtQ1BrJUBjYi3QDT64k4pIdtmvn4XITUbBgWcHKxc0uUr7+pZ41tCkqve+bCKl
GNwT/NiFa6fIUottgkPZP5NmI17SyvFu5XcUrKfXdKCulm+no6f4l/nvFcOmKfxFMvg5dqLbGbB1
xV7HluhcnixsEbHuNTZtg3p9GNvTT7wLjTUPMuYvWo28O5AtTZVy0Hl7uA3sOb75DmUpciQIX9Ir
vhepGLNZN2KcFth7VJDY4jDPfg7fqsGajlRiFZxTkAfeNGRRJDdUxJmuXB5dVaW+sazMdVyMHzbL
9bkCgh0bU6pCa9BltImZA100SVPpiYNx1wOt6LyAKtIKJW6MX4vmXYjGO6LxQxFCOJd+ajqHsVHm
n1XvkauT2m5U0Ia4CaSfYFRHTOCNLj5OykLjs7q0akYqoA2kQcK0mqLHeYP0+C8ve5hlkzQiX0Ai
vsZlYvQTkxmC1aNtMpAbg7O0Qp7y/AcqfGLTQsaa97jaDNL20+Or/EmNlt2mqD4uLrG0jW0GHpcX
TxmOf+5MLhfTcvwzLz8D+e3IJiqdokNX6EfYaGN+8yCivCbaILIqLBx7aIvdsip9ywM00cuFel2R
sjduLGKsNVQc59DJoXYn3GdjssepFXsYMwo2aWu6FS1XttdaWUz5WsQSRmrJR69dl7fa7TFKJgqP
lZbT2UJLRXJZJ+4ydAnJ0cxM3MdvTjuYWZrcZt33x/CVSYbtUvsVInxPOxtbsICowPpT4JqcuNlU
vQv+nuMYIEX1J99UGHzBV4Sq4sVxbPyK3l3hRBdzC78NY3wiDW+GVQmFaQj4NsiR6L8rWqfDZUVD
Hq91ySU38o8SZXg3nM4+ISxdt/Iyo+/6r0iIegWa4aNBqd+2CcIrWxJqTtdpLAT+LEG9yMxIz9gD
RrWpGRmixt+QATfaXjBYCMPj8VOuYf9+9fxIXS/oydXXxes+Grl3XYbz7RaMrNOLLccKg1BxksP/
IbYy/AvbzZn7ihHpN7YOyRhCyUs60nS0Cg91paOh6PVGr8TOHzfFteEoSNnLNJUJzRXEd7FHRwXd
6BM6rvIIK6DiDLkxOCF/W73lL6k+/+ELP/SDXIPUsk6PnRj3rNb4bwN5cwg8WSVptYNX50PQ5oOV
lh/tWiYE4AMaP6MJ2ASGEUsInZtKlcnT12FwYlvpfZd1uYeKkk7FcjvHVqXx05SmGSmmt7OGxJ90
HsD97Pu2gjQdjOQqp/y7MgXyshgAMKhZpV7JHzE4Byz7RH6Kk+qjMnUrb+pU2tjLdSTTNgcBFenJ
kmp11jWQz/Iz3jDbJka1UvUoYpQERvYUj24dQ5oQmbsb5L6GoyE2xgQbyWnzTg2NlNVH3o9oDbtA
kBTLb6vFP5r5yDLwX1BEofNaYzbqvgI/Uf2AFaeHTBm4fWz09CBWq1td6EoefByXV6vKJ1KvcHDn
U9XeFNAiHylFclrRBqhqGWyGdo/wCJ8JV6kBCuMBhYnE/eI0mQyrMAHpF6kHnwr+s+7ZuKnrHsm6
3C2HUd6RlheGHTBwzywknEe5Y5HHDgrE0Coztv5AOUNycLIbWiJLpW9qmLF6SigQHOfWeCShnENY
K7bJHUz1892XSXFDKJtBAEVR2nXYu6ovuZLnKJkaOK8lyoRd4tBSChH6IO2+WdUiQOt8LdSS13U/
IG+PAYa5+wtbv64CEZlwlQ2xSlW7EO8ve9fqkfgLPmU4I/9/V+Zm7YprgnI6fedPPd3jB7orJcVd
GZBfZa79ZTjQb4pBj/gGGtLOUHGlh39A0En9Zj3sS3B+qNq4ff5kGfxpThl6CELkxWrlmyYjgsAs
RbICSpXffKkNaeKRgzj9xf3BXiZMQalTofi6Jpl0WfQqySP1Q8+O4q75fx279eiAZo4O5xEkcqv+
i7yK/sNX54g7rkzeZtZ4ftHpYmrn7TrXS06b7TSIqmkGbpK6y27Lr32RBNIeycoRed8qSxEjnD5j
bfZIuZsntJD+WX3T4bxCSbDKhiJHxgSYA9mCpqvhENdzWmKshXUJXB+r66yTwsJeU0ngabGzf9Gl
I5nSCZHhL9+eAqbY1ElCZO4dm82WIW8yzTDpBuLeI6PqE2o8nYMwWzARtWbliUwHaS5T+xmYBnp6
TkFHWtWpmiyEeRIHWG07+7ARBWHdE5IP15S+MZYhEAcoJe7ppdoZNNiiILu71u1xdFJ0ET/NbqeL
wkI8PLMGCF6SNReNvWpiFLU33c7Kv11RtwwV1zKjKqQausFiXiA1J9gGm5iNrhW0slYeHo+yA7F/
Znvjux4l9sD/dy7EfZxJKCxy3nz/2IoMPvNaeGm07ySCO7XztjdN0Qpx34z+AR33KRhacNTjI5Bk
AEy8CS0dHLqW0I2YvXbmkPOCng4GoXIygfXm1xljYU6kpZfHgr+Qz125jEEqPqFL8WgTJaxLyBdE
E8teIBlsyFfLrE+neuiiYmaoNJZV5EkG4uEtXdy2u0wcoUtw8ahVPe93DWlR7V4uGaVBfvcMAdFI
fQ40iKlbn/LOGZHNmdIWwNikV76MqBT4Ip3a6zoZKKwh38LmdXGqsT0IGwNzzbsAefeRSlEKJ1td
cZwafVzq9XmjRk/6sYoFhzIR+9DjuEu0t6SJJxF9He0ie/WCNHo5B/Yh8TqPPGzbpapxMonrf8I2
ACh+wgNJx7ghrwbJlCSzkBE10qnCoEHEAd5npBQ6k2UsFHAJ9MibhipjL05eM2igCgJZiYXZHekf
nxI6Ky/F0htVGV/OmIieMuG7Uf3xsbzuivzQvDu+CRSPIU7qRH4pEK2jW05Y6VruUCplwS5Ltv8C
o/EVyPcnC1vcyydSwVne3I1qcn0BqbSVHAz2iUsd1pWb6kH7OIrPQI0iO0cSDEqkZTfr29PPdel2
6TZW4B70XrEb3eAOofSLrM++iHU1dGZLhK5MNNMavITPDtZN/URKnPRTYrGp0ctQ/uwB5MfksSnP
8ez0qK2HvTty4NGErRtfwYclv+QiExolz7ZahAnE7k/B/O1/EwBnaKVLVUEe4NkwUOITIeCrwRhr
R97AtQ0Pi4trkoJivH5++LLNd67z7JMJl/FbcCFBB7lJzQOHCEQOY9LwmMMwZm5D9rtQHYZ44EkJ
L2CAcLpUARTxToeW/3leIJbyzestg040R2iN9VafW0+n3bopsnseVsS5ZmRE51nhI5Cr+fQwMbhJ
cGQFIXXXuNNqSZwpA14vY6HdhBixJmsc+ZykPMEPOIYzOAjy5CAtOEmqOuLg7kh+x+YVYJ2rBtq+
B5oaKVjd5gaxnGLcsHLwzlKtW/Mx5i+YT9uGD+56qAkQoLYuJasLF0EQ2k9IcWplF2MmbWK0LzyF
cfdRgpxY3AYwWrABnUs14/OjKJo19Ph6iN0YCnH9VR3B8s6amgbZaTXCjAWFfvWsb0to1dkiwA1O
L6scw4wrc/1c5c+p+TVLRMq9RvqAg4noLUU1MbkCC0jF0RHA38KIDJqQI2+5eTDifecak9BugnFS
87Npgo9ZZjJdkFfNMHE4aDf3u/noMbIWtCzV0vPvkedN70PHV1j6vZVR+OGvRlInVeyOhoWYjDon
ywoSQ5gU20lldzjLbtGA3bF4PpW9drHECPY/hrB9z6l5NnID6nOhbTytjD+9Ql4jWkZF5x8Gb1ud
QO9unmDXr/LqWKGdNAxEIuJ7+h7/DwhfvVXkTyxUpJAk1NSJSX0e1sfbuGPUk9IeJQuUdJA7iFUZ
PJM8Psitu2VyZtw00h+qbpWY6RayjtzvLm4Gr2BE/8tiRnCpOIzi8fuwO7pHOnU4IUkP1Tqip1al
5ZcB1CyPLWdgM9PVYsD9OOs8Bp5zuWY888HCmvS7kxgQ1FkIX3tpLNhOC9j4ELUSe2gdXd6X6yZ7
CVX8NmA4buPeR3xiGPTfSo94aGpps+f4nERZ1pCATZPbGyWw7Il+SsUo+rH/1MRM2Hk+Tmtpof9H
JiMBiw92ljrhkBHAbP3ZNkxMhTjBwUUsrSerQ9t7vPqlT23T8Adhq9EAhgRQNXKCjO9ylK7PXmo3
2lj0iajnUXkIaK3oczvSfLaipsCcjIbKR1/kgK17+0SdVVlocWrQmmPuXkV5xQRuzpUnpDrtq87y
RSKTk2stjAZBGHj4o0qOu3VMeG7w4sGyNh+Xfq1+O81f1tF66vTxYSidmSHw0We6OnBQOf7cl/u7
FIPPLe/8tUlrXxZu31Iy9ILe9sbTQjpxh847puvBa8B4hdPP2q40xUVjSv4ti1kVW9vtdS+FKTNi
F6OyBGe0Dt1iuQqEfuRicZrH2JkN76xizpo3mhER2eFjIwW+M8DDiC5zGMRXjuv0gfkPqU4m+7aU
K+1VEeXATJSzKEQvEmoScZXlf3A5mj1/k8rU60NEQb1WrvQinxdMceJRe/sZaKx+rZt0Fg3oKKXW
bikEwOUlIY52gTsGnDh04fBGBlGgJmI3MwhVkVysUbWkj9PLhos/2/39Rft2IR7xWH5tqNV1AqE6
B9zsUmmyRXNYkPpVkEMGhRfMaveVR2cXA2mSZKpgBGsqieMK3UH+iW8oxtdz/OI7xUDRrU+kHAYx
HHUAtOWcmSsASfaH/zdyyirafkeakcF+93H035gbOc4w7b8+Zy+al8hAZ3LRCAnNkR7ujDaujxYQ
sFARSP3gSm9tlcQg36W63+PoEal8R+swB1Pv/UbdcWVsze3ipUZ6O+xqxig3qwkFNVoABLWROnMz
9LGdZzKp58/5m4helCicxM6r8GC68crhN7W8nZIKG5mvrHcaxLmdj99guCxZ6xY6QR6Q9Xj0XpBV
696UmExTOT1128LwTVPxltn5rIiI78/eFnVVkdHn7CjaUMInaFumZ+KtcCnoDAtC1mvsYFIKGlql
nDYAp+q40mWjJDOupZPXpUpYnQUQWR4ZuQg2PQr3Rrur6HHmKr7BgMoZyjkdC56xzPJVmjaY0ceC
lka50Y3NUVdf/Uwa7ihV0b8fWaMYzlt5CaPR2XvmB/iEfRGxVb5QzCqpE+BJIujV8AhGFkKjDM3Z
tkLsYI4iOn2t2NjzuDYpaS9fCsD8RhMGjnBm5ls5W8yL+PP0FUBtpatNHtfo4WFc5D5Dqi6NdYbe
GRhkDdm2zBQjDUh34dJLhLaKGKDwQFJgzQKKbv/Fv5OyJoLfCL7nKLd+S0mAQkha5IaQUbzaRubx
kIaH/RuZ/OMiDoA73oSCriHW7MtGHrrr4USPtZa1yvx7G6bo7QTx4gk6Fw4RKxQnZVYnHFujQoO8
iGXl0opYyLY0F5ocho91qwetqWQ+OaTCKtHcuDHmytSb6BNvDLN8qBP2QmEDR1x2+F54bYfDlNA1
+0TLs0zl0rIzAdZIBfkUu+RJawmJhafE6y+85YGIBYqKH4cvN8yNHOtjOpLGxlzTsB7NEiU8uz42
Wt7J0UXWy8erIYorEaRRHthxgpWvrDmgpxYvQacV6DoFlsYbh2j9xsvyG818MWGqsR676IeiMaOb
+Js+9285hcX45H0oqERuNXNGE+T6vNdGZ/lAnHmtWo1ceiYpbeevARFeb9ildP5HAU29pGG5V8dZ
8EPMMXAdMjTZNv3STXdqeNqTLU9FeuRidwHI+mP41FrYV30+sQwCwppu9rfdOEZq0/zp0FutbyQe
EvM6AuaEdYcYtOdH38EeQBjduv8vMVIZBTINWvMMlkhnJks9lmmdwra5z1/j6AS29C4W3GFZlELk
mTK8LwsJ5RySP+xDDbCL8NCbgYGouUvCAB/+cycMGTDQBrEkc5pwnnjVTCj5zsx5VBeqaaI6tZkL
L6Dq94I+stUYcQQ14I1tAOJ2yYrrJKi6GykWBodDvMj0Lk7c7r1qEdO3jjMtNpgLsT/dkOWKX8Wk
AUS05HngYaZ7qs9NzxelWH3y7gQTADL6p1Ygquov/mBbfK8o+89m7UjGzQGnyswOV8pVR/F6jtic
vV8kBgw4vOiltQCwpF3U+RBOtmD/FP7E1R5NIkhy52LZMj9VCUFvcIAp55cZ6RhxCOyBjmDFGQ79
osduVNu7p93hDBJPzECjWC7Z5glc+9xbK+7r47Sz9NTW4dEFtSUBCfsdnK/jrp1NfNwAdIY0WHAC
JgT5WUoir0FqVW0WRzLS7hv63sdQKSdiXitX2tx2llFf1QlsbEkVQVoW0b1ofwKeWW5afUetSWNO
jUb4JaJQ7zVfoL07IbYlA3j5riY18bWotjxf8r+9bKpHRBgJhWPQ9QAQzWsYxt0bZEQDfiV+W5Sk
2ZAvclocwhXHkth/rK5coorj1FuyuSCGTXlyxxHVL39SXcraFa2Lh9q/gpWdglGSDTgGsHhLUj9m
DF0LRWz6Pa/d0S+3uqenVoQSJrzFxZnVQBJegwt4oHe1mZvgVG8Deeo5JZCuDpUny/ThkhzrLkww
fTSTs4ktreBfHV1gU6csjtOOtrWunYTM7+4c4mXalrcGPTYoeB2R5pixtIVyThnfJhz24nDPluaW
eFf2BLXA9IdtiRCgXCi8lhmOO/Nx1lIjdtwQrGhVH0AdimrjQDoali4JBDFb6hi1LCwsn6N+qrl5
fvDenW6wQcxBovsLbbXPgEWfxsaI9vEx7yvc7kTW+XoIwPqH+WJzCVdHklKCa0ceSvGgnahWrUDs
wFmk6jSVkveLTswFkPQG8AwXGyIWYNBKsFrT4HRVFfCcpYCVLmLHLXnq93XutvqxnvNgwwD1j9jU
bJq3f0pO/zzrVzWklwxN/QlvuGcmFL0EPBzcpxDQziLTehls47AQfQwX4BskcnaGARL8jt6dwg0E
ZSsb0OeiavBD+ZP52kNP826TtT+uCTp7xL/7pnGpC1hlOWHrx9xqROIeH0Oh69+atIFrRYZ3r0P2
atF4YwYJxzBEee+rA+wTCwdA2TCldnElDTJUSrdos6dYEvrOShx9QZeXluwDDHJmNebpEuSL2vOC
YyhLUDQUa4Q0lHSHyRy+MVBCujxa5DL0Na0iQhce81QPos462gFMOcyNrhRZl9aYRtmFtRM9+yDO
JGcwhAIFkOhkGP5iy1ArtdZcBjaMQ6psEEJmErVFkldesEZNp2bQRNrNgE7XUheRVG2tEHNrGfzZ
1kJQSrNLJlp38vLP5aTeQ2Lnxbv6ZhdIszTD1B9MqT0/SDxhONcUwTmeBEioDaetvYb5/RipIlOy
1zVxTxBewQiafsMWn/Y1nF33X+5DEu3CwZuGw0cI0oeLiJfBhSobHJInvgWe6+WHLGrShsJlb9EU
WQiR8kxhMMkNBNjfuYgiY9HG89xzudSkN2rZ6LdRVTyeAEnKnpxLot/Yx3/hZekRPqySBtHyF2D4
HEX71gKNWxS/6sWu98EyJbbeAKChYDgoNGNj1XrN2duvi8sBDEOkQsCIOKQ9CiDzrBO+d9r+NoH4
ht7tHi2W70t9pyZC80W1wlR9CESNyPWcxt7IdbbL0Kjq7TTdVJmZLX+6osgneZ0APEyHB/frnlJI
m923I8AiY4KYmAeEfrXeCPWBEt/2XDrWZkXLc7+4Lt3ipaq9jpW5BC+0eQqWCRJ+CATm28Ny5ucn
PTsu9ZyDUmv4zin8MnVKDPGj5a47Jl2tcjqPEtAV/ETUT1cDUHJ8uwXXkvTXSXhUFMaB7gRLCZ4Z
7wSEiihaUmtuCwt5mWsEwit/Qd6NeJBtEomoRbeaYM7Lv+WfuJUkE/SD5FyLpy06ZGAghLRydU5U
22AjmxVcf8oxWYrvAFemcKokkNfal+wENHXMcVMcZUW7RPmPhMxJQqyyuoA394q3Oh6skOOjofWt
g3NQX6Iw40AfnJYJSSMtz+OhvkEP4IpEmsPYNvAeSzKrZjf+FlL5KjFVXzEVPU2/tVfAFw2/axXk
Cbc5UIW0JplPlWyqH1ENeUqRFZ3vnLJcz3auMkMsvG3DjxfmcOQgNaHsm21jrLnYNi9y2/G6kqUR
jd9z58L9kkXiCmTtWAy6E3X23yHdj+eEZ+wnrIQDx7Bmz1NODG4Z2Qdu4QdxBBTwwTmjWHyhT1NB
eUqxoYRYEkpDzIgdw0e7xHUlSMThlp/9gN7meKk12TJoc5EeaK7nuLtd24Rn+SI3DrY0ClW5e1r/
kLbbbo5bvXbM1Jo8sHH3CkU83NxIA0K6ayKyDU/Z46GiWN8x+bFms7GAzTGUH1OXEw73zE2NP/Jh
IfWLdBFT9ftyOJT88jd3TtORQAEnkL7t9gqqz08kbA1lQe3KSAOzW5DKOFukA/cHOqB0r62wePTj
dq5ha5eMJWNTg7udYQLbC3Kc6f33b9QldPXfv+qzSdbEuFlYfbUAIcWpU2b+t1k27ul6WSWvvBvG
RsUNovmNDzbrFPAssvaZC40lDkNLMyMfKvdBiujoZ2DxMgST3cVkmb88soF/k+SkEyS7Fvk1tY8e
39dUn/SgVDmXb2hX2h143kLgdek8drROGtndO777QnCN9GQ8ju+gPQDoJ5qifr055t9BipS857sa
+KnsWrVYDltzy2kVN6BUnCwV3Vj68otAOuUi4t+JW/mQ94qqn463Y860qUV+O/MV9TXaa2seM8cR
jfc3btSP/v446lQwuLTexiN5wE7uHVXM2jkz5s1psx/BOa1LHSAYfDfTaUhVeUDH6zJuH64EGKZ0
Wo3xL0ylsKvOACjPC9Jj32nR4nESPqHR45ceob4I/UZvQ8O6/bLAbkYZK1EEnQS5+aEnrbb/LFPJ
8jwBdnpMRKsYtaWDeOFxHA7IFJNmWASo0gjgvqQ4nBOqbtyNdN6mijvUFtqw7D+Vx7oR3tfqwlhs
b2DONUS7P/QmbSfbgf2NXW+f1symsdIZ5eCbcYpBHl7btdxeCaSMze0fXzB7SjVS8Byd4ZSdjw69
DONVuN2GX/AWpkc12GFU0AqSt+v/snhQjLi/b/cbKBPBjXbcM5rOa0hSp2vUXtijLZe5LdIEEFIW
IQw7bAosrThrWr1J3c+ZzGs0jRQiIezssD4AgsmaXRvS+Im3M4R82KkgLyzfAZSK4MF3adJ+5pZ8
ZDG2uFc/MjXyUW4ADgBrpw8u1zWNlriR/WC9fF8GA14kc4CuGga+H4I9Tod1lEKiVruEP9C3ve+o
GPOaAetHbyJjqMK6KQF3MxV50Ij7QBH6BpiS69NHYfGsOTnk1zuwtkusK3GTDWgMiGhBU9Zr4ZD3
np08w0G0/+KcfKZc56knZkSztu2sSzbmLjjmboCwwrmfSJIdnT4NCmNPQWH2gOLx0TguW+UQCLGT
fKrHs7GZESiec4Ub3i7X59Sx91bpSOaHqebbGLPqWrp7GNNboEPpbIfWAuPIOXdKIXjr0Li2/7fh
NkBNXsS2FDobgoq5VzKf942irgeUXvJws2drVLgHo7WnPiVfayPGjbFHPNtNbnLSAs/9O/NpKZ50
1aDcMfWcQsml/RzVXdZDWn0SalAovP//sK/PcplqIDp+N3ejDmenaT9VWSiGGz/cqYYfXROmUGvY
GhwV0kqvwKnb04bwrvO4mhxXXZpqdezCllAGHWg6JEkorfu9X/Exk9bkUAzhP5m1AGwb4aNJoJVx
EtUi2pvhWQl+RrN9kT6nAscyceycBToz3WE3l0W024VtCK9NYJxcyfRdT+kIgxi8idyiHMpxITCp
GSFSlCJVRzBw0WpGyVh359g6b9PSoQlG9P3vpclHBNIIPtF672L8sIzwm0+W8cLeRyFOiCjdzHoa
z9ozM8GUOfwSsq3J7gGpn61KVA1tkFgiXwy2Ujf/MFCymrD/DjLqBatP3W3shntjWSzqzt39CTCo
/W5hhoTagyMUvIPwBEpLLRaJvqUrYYgh4/yxTq2Auisz1fnOSKT+mr9iCGMDqfucvohH/clZlO2d
mKEM3gnF/AlpI6WUm2NpG7CkN2MiWXb3CaMKqAnjg1VkWbafj3HfT2Pt2miHx1Q3QzaS9Opt1FmT
k1Rbb1uz1E4os7hPipHIhAbkw3yVtfKZbJ+zqJIPF3Z3Fk63mlVrpPqsY9TWKDtNUXiH2bD/Am/X
WCzaEyk89zS2eMFOdjSVg1rZtQvzF4B1llGi2JjBWyfT3mGbX5Cr7CBWlLlhba8G0DGT/EA+XEKo
MEx48YFtD3bSPvOPxgBVxRXWgMaXMSs8+EbGedt3292HEpJyojtp+mYzs9p4oYdQVwWyCtntpN14
raN69MHAerutwU5HmCE3uSgiQlaW6vyWMtfHGp9+K/Et9GONxyUPkTLDURAz4hK/z8gp0j6bISKg
72/Ex020zdDJ+kNSYbP0Uwbt7Ybf9I9xXIDKmA8LEnxlqDxl8/YTSFrkKyBtK3jW/UmOuTZsQ+m5
26Kho4fx3ygeY+1RgfUJdpQ9NCk7eaD/2S/DlhlM1EbNyNrT3s+22kpy4CUSynH4cUCTGoSwWjI5
MEmA5TnZhLOb0wm9n3suvDzPQRLFhVUEOxnscsQeCaZ6//yTtTG00f/99kUZEw7PbqTPJv8LWnay
gPWhpQqwjrGGBKwjzseOjCUctmkFOXN8f7sDahotIdRjG0sPYWnd0UHRGlnSkzy8aBZqTj/5bMYT
x0M+s9RqyDsNEKmbMylX/EBB5ycBV7U+U0BvafhIE85fN1FaxTI31mvF8zzR/Sf8q0QcGQpNlXH/
lXyPcULm7bsQ5HpIOWuLQvjFpKbk5jwJmb1CceeKbpRdPVuE8pJ/3o2IQ4n8gLgN90yVaZR0UPcU
QYq7vSEfS64YxVx8PNDYVTI+VqkNBkQc3Z6mwQcozHDV9YaMsWZ4DybghAoIUKQM2Gtz8RK5YT8h
gxe1ryH6w6uHHrU4yWdgwkyPJwEv8Qhx+bI5vk3unQlcdRIh5+a5oSgmdF3GjZzyqoqDhHKRLbae
JXuBDHqtQYsPXiAm2cHp7l2GZv/JPJfvwqy2UkmORmz/tJ30v6/3yXvxaD5Qu7oAJr6WKnjqmQFy
AAr0TX+ixoxpS6omleBFuLjKyyX9w9eKVJccvcdUVOFQZuGyIsZX3Z+zUJPte5Wa4u36mOdfiFkK
WjWGVTYwLNzBQIuUat4J0T5nnxlVEYdpmrDbcQ2EZz8w1+SiW4P97m5kipzDpndajVDZymItne31
4Vv0WjHUDho2aAibj0CF7JZGk+mTWrDBzczaCEAkyygVw923A205HvsXFfqT/IgiRb+cQhB+jfOm
NFtBIKPNxkaTk9YmwxDvSabiLXe6ChTXLBFzfdSFjUYh4C57KQyPLFxRt5+jHJ6cRGXcMdnflfMj
lq4J6J8vW/tbLQKKfsksA2sCuf2RjE4Dzokgjl6LZzSsExGU5qQk69ITi6H/aqhXLpW35cAq4bf1
2jpj/cq6kvnJL0UWw0uRiy0pRaIEiHEm6OoU2t0PWIoeFEZ4Z7xyICVzeVxxJDLMfBz+4bmsoHPb
xCLCG9Gi4TtkAYWgWJnsQYfcEtFJ8tCwzU5kgrHj02lbwvvSeJjrdjsHgMJho+Db8YIlYnHVkA37
g+9R0PPqP6me7bwlqFp7IRC36zNa2d4kxNa8WK3gTKkJ7Oi4rnM4L2TyYwF0z2xhInk4AcjjcHX3
49vn/5DFoRxaGeVWoNA6o72gDPn9X3xuEoIdx18dCMFZH2ZtLXWGLUz0K+V/DNMuD2I4QiOJwxuH
tW+BO5sDMtzVOK6u5VLSxDjZCXsqsIdYJDlmNhytUFMUjHWjCJCWF8wRM5tonreXhOTTJ84VLGJD
hM2h0K8H/GX3sKApyDSKZhu9px/1k9MbEy9j6HQN4ekPjpNDbmroO/mGx37On8EkCOwCX2VZdHG+
+XX81CbrX/7VvyT+PmmbteVYYamNCbdsPaQqO8IPHNkvc8vS61znX0U9f0ais0zT17/3tnFIkOBt
22IPdUCc7AN6/gOFHlndFZcIiuL35emqM71DkruJvNIcMDPLHs4KfIoAVBkva29DrXaYXbKE+ZQY
djfRtdP8GQLGCU82ncYnj86h7KBQu22QV9FAoC10Taswzziho0aTcgRdf0u7aI1NdS8k6Kr7I73k
rrYvKHO9neRoMSTjqERNc/Zflwe2dEdGiQBLPiP5+PIMQJYScjDu4/iJUqWGEoA3EP43Xf/MSkjF
eNBz8G5lPYr1U1P7W2fY0jR6CwYHG00nBaWc3d2rt51GjS6+tax6pvg++7phjTS9QNkY39J5SAcG
wP6jEwPUyJi6HvyRncbEntwmN7MH4CCS700wEWsxDIfQrlJ9bB4m3WA+Go0jadMWnyFq4L4yx0Zh
sb+eBSzFxPY/CE2F5ZARuqgpTNhuEVlgdCKCWqVzK3kBbAGZuLyxgMVtu73uozIoplewfnufyXUv
rRfk8uEADU5TRF/kj7/z+zqmDYe3mJuoiWHT5dRruD9zGsonaNG/Uesebn7gZvh9uBmf/gsYkSbn
FHiqNsO+xIuxbAaBJmqBPez4NIOOdH7JbLGYvnEFbliBLARqvlTfoHoaxZguqjU7olIjCwdj1FGy
vv4eLGnn/ZXcM1LPpnKIZk2/jccOl9t1IwtBgBwDPEKLcrumJoVpsKppw3iHDjE/0abZf0yRsain
oHA1KbHC6iBbQqWyA/Q78GeruxGIOJMnthh9C7FddO3e7Soz47oCDQajOOk+PMun5g/1+DYglZQR
0ZMK0Wd3VVKHs1nrzVRHefmDHjSkCLqRaRFPC7b7Zj3Ta+tEVCARslmk4dICkHv/45/03+HAxP6d
ZG+oEHhxBR3eFj1AKABkxOaXEGRtlWURk/QXR9H261emG1w+6CtlTVVKlJF2GDCDxRLUxjVFSVNF
TtkMNlwB4VFfugyvZp+3M2mlgRlfQMq1npTonXSkyLVlrULx+v+lyMGRFPKuWIBsWG2MTpXUS1Du
G32yNR9tVem+Nj4TSLNB/VKEWoZmelD7igYpoJfEegJA/a5WoQfYL/WOGDWoUb37lSW0IZEFeMKN
yQ3JngoWaUN89zLdA0X4Ic8CVf0sv1JOeOYoq8hO8DkQKLAJ7su0JdzdIls6ONS+6BBIh6xpHnT2
QCLEBYDTxqArzVO244NfuURkwyqROPrLBzwh06+IZY10/v6CkGdLyIKe9uFjw+J4lclt8voFamdu
mlojKom4vp9IioCOcToH65Ym+uEgYiXPEnp0mdSsi+JrZ+/RXkO3gx6f35OvZLmYpn5wM+QPtgME
Q+UtIjD3GtMDK2sISL5NOtORMLyo44GGM0NhzdydBy1JSSDdWyY1oLSXVkY8jtKiw8w/pPrJ2e7/
PD8y4aBQ5+X5YGOvSIwXXa37KqrexXQWPAVRGN/ExMFDfFuDaqHqLQp++MQmP9whMhcRD9Bgqvfd
8ceRSeHgu0noGtd0gGglKn0eDJHk07uiWFyvYj6961rMON11v8ODcPHt+mal2xDgqayeyG++ToWp
gGK7lDntikT/DbUkBZH8qiFG1biHS6/NzdMfSZJ5B3xljKLrbqI3Mtj0aia9Wa3aRjeWr+4I6hlw
ioTGeNqXvTgRd9D4Vmg31v4ujkYCYeBVj8AUm6ir/HmTKu4DQnCWbLItRRfaUdDt+sZJHCge5vso
HntHVGYORRSPq30lrRhySUVSr2koQ1qKcQe/TLqSQnLWEJPUNSV/3fT0Gz5bHZ533oSNq0hq6K2k
QrQmAFV2W0d4NhcPEUUdqpqYUVGzW6GjWRQCtZVFBg523+pEFyy9J+PVScNVBZwp+xtjEBlCblSL
QlEOfbPbmF/Yf289wOaLWbDN/38s8fFoid+6BvByqwEC3uv0eFrr7hjCtvA4tOyVPe6px1oDea6B
/naVOlzZpqPlhBxAPdsuJUUAxxywOyOo3ckZSYmcPOP2PkeuQwq2VzCn5kCsKX+GWafPKHyB4nhA
pEDckq74nnhTxIkoO6qP34deB+485hIap140x5vpCYyJ7a59Bi9tidq+ITSIkAvGtlpvEo92Ov+C
ZhA/UPRKP6+nM8SD9p1yU4kE6f86OGCjavHoKZvdjvHMi1pTz6MtWJbVvE9qYW3RPzniwRpWRw2I
aGqsxo567PSjfc1wimyvC1DmAqaCZC7CZ2PbnpbU7k22pTyqT7PinrkhpPV+sNVfE9eCYQKIpaGt
dr2L451TTa6x7UwGJtNU953fXFrJtwuvdwZTq6jonqtVr1pwZnIue4vQkiYwzbiP+P6KgKKVZ5Jx
JXsqyLJBnTBOsHEvPelGy5K3EYAAPoTJQNrKhGxYcnXxelaEADg6SrVPpmASIARr+vVebwtIMaUG
OOtq9lGmROLQiKceKCTfoXTYmgzch83nZTUSM7jI5XX5zN+vl1kfgqgz3DZoWH8VUZE7mXzNTOk4
Y6gxL3iP0Wrkvwc9LqlzwDoQMT+FrkFrYGJjw0Wy2W6aalkexk1Q7soNk6KJE4wJIWs+yBsqKknc
zreI0V1fuoUVad9c3U2UlmxPiVhyS/Gii5ivjhO6DbnsLwpP+hBqKypQmETx0krCPdDltR+CaGYp
tozLc1xsidzM8oERotK0tS4cJtzXTK4unsJK1qfTjxzyk9lG+7xw+syH7HbvFxI6cDsKr/T5c7yv
kalMM9CARiQU4SIw+547RtZl3LQgcH4O99XXmuiPZlQRiGDi0sOAETeByi2D6RI1hjMTyr0T3uDI
hQ91DaGob2mYe6LL5lcEhmmTcSFgbtaPg7yizi/475U7P73JpmySbggNr8iRQ6uWpPiBVC4MzzfR
/Wh23P0622v2jHw+q2TpmYJEqtZmiI/ZnjehD9dQKXLJLrc0nH9dMTQLWwCxm5SxnkLeblbDXXoX
F6vvpA9N/dHvu7oYAnY6BsVtMNW8nTgK7dcXo+HnYlL8c5eEjz9F6kFvMHJG1RgdfDOyaovoaEy2
N0OoBt0ZJnny130bHXOPs5Nne5a4ObOmEWOFtJ8JntGZq5dclb6m/EVXWhi/J8TqLJJb9bqF1wsL
C4tkLV5LJkDZ/HacqaZz4bKBpaD6f7Kq6TQPBza9L9bdn1dfUswqaza4SL0XamcibgD5onaxRhs1
fYQL96H0UvRa/iqc/11Kx4jPUebi2kqhYs3K3NZ+jd39F5+oDU2MbcRNJF7ClUCAa450LBdtx+8Z
SC83sHnonk3UM8G13+h9e+ItmGEIhAoA346P/5J8fXa1/qDGPRArr09U7tJoqkygUVOADIdw/ByC
O9L7GflB41xwDeOGhswSeqWSjMVb52k1NA23arrCJK7zFxvqKM7TL8GTk4RwJF91K/eSM64WWRUi
jb6gBYoY9n0tw8PyliqghDmDypwGVf98dQltwGqSMOTxMTth1ijbAHpmPsSfvq6OR5XiuTw6ZUz4
uDxQlLdJ2Bl9mDu28Rsmnb6NucHvxKfE9G2d22e4Xw5/xZF+gDA2CR3BbY7hwzdZ5eqyiOHKZmLv
g7mQ2P0fYMqs6aj4Tnvhk7JzJOHU40DIxLpEQQPl6YHWaFcXW5wMYBvDbJHtYia/7PeTBppgGY3G
15SxJzwBMj2fgtsNbBG/2em0mVV5KP57PkBH56gbapZkc/Cr7p4ELwQpdgN8cyzHh4oV9SDZGJ0w
9kVUU7S5qyFaH4AMXMRHMqAtP1IxAdiBeRkWufWqYm64rObTgjvqh6ySg1S3rnVzhI1kxTr98V/9
CsTTxeYTI9mnNZsWfmtcoxEeh0LOhhlBcIV5UWvomDj+8TzVqTcc/2sozlHaO4ObHM7nwuR8oJG2
r0kO+p5s4VJDV2J0I5NTcRMH7G8iAFz0vcQVfUChyCrmFEI3eEbo+lofWjLBAw/v/q/4DdrqVUGk
k2q6tB4Kh5dos6RlWRcqnUijqnF4HJgHf52Fe+pJJfxjEYpeejXc1/E27roXLAbnAYFBsHXHhO1B
xDG5YdivC45fNHPR7VRVGxhJZbdLQgj2t7XaRtNQCoaPdKjTCFB3qPOPKhuJGiJREkrgfwlC9S69
cgG7EvIr82lpzJudXTUnsNsDVn+cxz8I1zboVW7zBB1RAjgcWeFKjettkUgyA7CWYlvf6b8yizxQ
/tPqnv0CDUlj+hBTDqc2WVlKPaKBN7dyUGfuYmTWcn7KTy7SAVxuU8NiI68Wqy64yK8uH8m8478I
JDubuOoyvZA0xZcAIqcYLS3uhO7wwu3GOfdsYr44O8kbLyAwV1IgA2hBN+Wuzp45H+axtheOBoBH
5cMHA6JFPT7ohmgnRh5KYYNvplE+IoCAszedrhQwzHyqMGEp3f4IXlZFrHMEp51ElWbOBIJcIo5R
xgPE97dJ1FYWvrYV6ioIDpA6ZRnwmIPqiA0w43JvOtqk9xsnkqJILU+dH2s1NGcz2iUC9d7ll8b2
bPq4YLbYtLsl6tSTNlqQt9qVbwnzit/D4rLan+wBu7QvLisOjw+Ggv6mNsianPeATekQA0xxQQbK
rFdOcce+jZed7R06sQ82kbvPPbdc3S6rQvHQjyT5wQHPoQdovZxKQ114gV40gU6kqHWGYnIlqwyM
lADPq3VES94nXXuWnWGNmqJY+BXxWUnUW4njTdwgzMRkyagtDQ73u3pEHiB0NQBtbUK2s1cWrmi1
bnqpFs+OI+kAdo2zUQYYpFcv7EbuJND56GllwH6/g36pFhL/jen2DXXO69XWdoB7eQMt/DMKW/qY
d086fWdc3uykoqG59cxEeqjTAPKa7s6PNR0Kwbj+PJrm9KMT54nc7Aql6AcVgL0NEmKLE6EKgG1p
/YaB9P7rP+qS1wYngLk86RwXeMe/4bC3T5CAYHJGbq0tnzf2O0ICcozpgkqZjavB5BruJEF9ivkh
5h1IytncB7sTvZ9U9ri+kUYrgkioGn1Ul1VpoHE6MSa/aGRuM52OHHNJyblGtwpRnLnY7M+egTWh
wkxYPdaFVZLHXxD334JRAaUUfn9lDBtYrVaIhai555ZEJ17uX62+OT/CX1d/UwBA2ivrXg32IXR/
PvgC8BqHKkkEGiys7kdqXNTIl5aJbgYbK71rlWUpuKzYd+Vm2TdmzwIMDI9pr4Jy/1dXfhzNDAny
iTaPAtLNwmtfVDSa3xcZxvpv187rkcFaJR2ROenKUlrd6nAIOIMZg5FVOcz2PXtJ0gATKuRuSTeu
1Vvhfb4OeSLdl89AUWzyjQENYIsyCYZjTcY8uSyh+gsyVH9Vh0xOSemEU4+4Any8/6iP09i1livI
zVy9rIPnNLh5xgXei3f75a8G14tBekD9lrTjZ4l/Lr34PtH/j5Io9qBEMQ60p+FkuDTqlts9fpze
Z+ydW6lt3jmlqwj9e+wXEmixxMh9RIa6mt/XFCx3ZKgBxtWKuvwXB4qaX0iOMCCkWdN7scbfmc9K
QQK43H9oy3s62gK/ET9wsyoeKdchTstBsnUOO3tUTA5qVJSsRewcUv9YgCIsCZjl6utNm36yw5us
y7c1bZFPPIUNrLIqSI5getOZA+V9EIFKxAnAfMjqdfG61FtxlU2/DMzuYFQQ1BUhbT8/eE4V5Q3j
xWFqQno8XQMLAckFHNDDvqW0l7ZNmhlhdafWHSLHgaesJ801BlXgV+x9AQO+snfo0wGxaQV2cw5D
oot4NieivlAeDtDz87X/UW8fEQFNTpSC+IMha6DZLmePYBQhGcqyZu4Bzm4jWSpSOvnMZXKGP3TQ
mKNxsshiGfc9X960n0tMa11+VyA2wq2lH3UZ63FBFwuOIVfuDx2S4j6KnBbl0pLj3JHBv4Z6MjEq
xz0QeM4NxlZSIX8YHNjgU8nN5c6JCumEJ+d8XK7pM6GfIdKSMlk6nfSYbO13XDmj2chsU0OYct31
d0+euemiFJ4zfrsk3weatgmVuHCLn8AtmKdFJ3LuI+LETx9cp/oEGMS80fBGLYasH01x21aYJwLy
0T1tPO+otJDMH0SOX+R6OdNN5c3INwyKe6A/R30Rqcc/kmimyWHtesNq7ksx3RZHP7OyroYHKu99
obRtDL0ruZJ9JHx06pYVSKl9R0ncnEeJ6T1C6208YW7Lb7i255akiB61H4EO1LFl5uDBTq4u4LHE
uqUSoHQDVPvuWPuvt7kuzgplwZS4AmyEdsKpvKLzYXrbe+hVyNDaOaAsuvCsMqxvjVGkhhJ++SM0
AKf88nr+SvXRSqMcNO3IDvuvORygQPC2yxbne4HF/s6RQ1KEL4fv+qPQXduLf4U/DGl5e1Upbvub
3996b6bBPazUhZIqmFlViS3DYS2UhZrrVBP0BwRtd/VTxS4OlEacFXebMZ0LM4tCZIUl4tEIr8+3
YDZIN0Ff5GHLiviF1FmqX/EbFrqq2TywjwM1dSFH+0qSB8rmJD3+J2aniN/Jl7f4Xw19QYRQWU7P
/zXGl4fQU1Ib4HSj0q49Oc883Hq6RHlF+afjV7o1GqHiUu0qOpPDqFQLV9GVzt1pBNrFPi2Fn0ao
wQURmjDsodOGgTGAC+32FmUYN3zzHY9Up59YakSs0J10aRpqci4ubhTuQqyb/aOrrazjavnHNenN
FMZTJ6MGaPaYbFT6RaQK7YdqkabFT7IPiL90O48KYn7ALE66p5GUNtmOEXrQnH9Do474XHdD7d2l
rtXhe4HUX5L3be5cQ7vZjx7p4VC1ncEcga8FM60J3jxYGRlTzJjA7CHGzs2mSwIxFVzIj27LlDUG
4KNqzyrQ+WMgJ85+r1x2l005WMyj4lvpDrns0oH8mgkot8SevTgMfAZtHbz3Ky/NhcgzSvgWobB2
XM+lCKzoUtcQeur7stlRyxhQbbRLVrngWfIwCtxDhtNfVKGkyNeDQXx+c+Eg/hUncCuU5ZjluwJl
SiUba/wkcgg6NN6EbJ6YogCEGMglD0RvGZfUDuQRBOOT/H0u0GrOZQ7L65TfLlkHnnmrd3CfFNQL
vYWShD3AZcIH6bBE/E3mIR3N8IRjowCLKOPJnDwEPlHv+q4UJa+el2JUUs0PZdbgtKLLxDrh04G1
XV54/I/JaLYGy1vCqYNduyZDfQvKU/aP6ugp0+x1XCkDpuCOYLxbr5aDjnpXIWUuDyVNqGTZT2gx
yY5AcHjdHq9NCBcpkyot7LpCrNgjyB5fMH/TYor6beGnsxxUn7yQzZjmmXR57/QdmJ3D6RQCEIsp
IcfK0lk15an0PbC50Hw3e7xM2i6oDh051/EqY8dqcL5xzKZ+h0gnTSjjlxykmVq1kfbAc3mi8Ija
1pBUbvB74OUrgxrkHr8TWZjQfx4Z9bW5sVWafwiMQKZ4pXoosjcHwJWT1jDPi4c6f71HlrwHx8nR
PNnEf6kgsG8vQJCduJiGJ3PtYavgpBwc6jwjJod2+TjGslqgu2teLWHXICXD3PbGIcrfU3ZlNSvF
cUXWkIlX5N3q5+NaPjNandZmcj1dCmBftLJ7Us6UJJ7lHP5+X+UeSwQm88suA0DDoSAQVKjo7CGT
qfG96N/Pow8x3JkH0tv94JIkwa5f8VV0AWTLDICSId65X6WL89rCtzWGh8CKGxdRGvm3OTH3MS86
2yL9BSvBT4XNk9aV7QoLotB7ujYJ9ccU5yzwg8i6rFMVGoR85snoPZASlDtxKOTma3UoDIeIdjpu
2Cyh7zjS8eE9vv/ePRheSJFm5C8jbd3u4ei5cQ28vSItPTbv5NfZ/Jc2isnHs7M2VgDVtTei07db
n7J0G6HBqCeh3hPI8ZKJcEX0UybDNoL6y1hi429+JJFf6iISLC6Ly6pBXH4m4VJ0qnEusIMrn7OS
GaOuGVQDUqtdk9pHWAf5fbn1+SWWMRPpPXurCE0x+tTMwoBOWhq4eB1pikZ9R18ZZovVEX7Tu4df
M0I4ahJuklao89yTr6ROWbBnw3svGUSK/I+Qn/+Rkx6lMRrhWBpRgdGCQKx8q0pDM0wuWKT2AFFK
cGRBL9qvTPZ0gMSlgwQBqMhHh+O42NANo1QRK7jREK5tafW9NgsV3Wco+u5uenrjIg+A1Ss8LtxJ
UBCRJ3NzG1AbDVvD3MzvBfYIVPvlq1tgqWCZPJYY0lwKsxfvsjSw3BAY3JDmlbM2C16OI7clyY4J
iWKnDuhSaY2ey9MFROOtqllsbzko6VPCCnF1qjx83O3x4XoMNHHw/jvqaK6gu+09FzW7ZH7j1Dl5
VZitZCgPFZSsB6B+l1mmBqKF7yjS4vH9w4R9HEzBtkFKEdeySoc5txZE/zEN3MKHS+iwwNBiuYx7
b+XiETVoE88MJrwkmBD5h9Ur6EiCO93VK8D+t2YUYI4Oldt8wM2LOFhl6YToLyThaPCr+CFQXf3c
wvZcDqHXY51ClKhW/AeUZZdQeToOXXBArh0roL0s6aaTBq/F/BqeAnO8BjGs+a3K4hMJSVg/hQT6
U64rJami0DXD3JyqbbewiYz3IIjd3K7vnPTU2uCHv4s9/gFWktw24jCQW2aDIzMZo3+D8svkfj1p
Py5gSSVNPEdnT2P+orPA36yMPOtsb4TzkOHAoMqOEVav2RmsgE3b1sAZQM8LjTQ5/mNbYAh/AXJw
b14gdgFz3U+F9PQpWpGKObWBI2S3CBo2+pJzpIZvEBL+G+XX7OuJfviEpw9xf0PcjXuSl2BNrW0n
ryMZg7kT8aKUbgjsHH0GbS0B2/4CkWBmff9S/ASXiIaDlyLqJGOg2m9sKIWAGVYE9IM9n9C7vb9/
C6DRXOOfjyPtbpCOy8AWUM28oDueB5vsUWOwFGVtRmqG1vWWsbhE/vqgOIUkOPqKAW9gtib7hsBN
f6WSNLa/y2iRfsPhuaTEsXMw6xItC4pDT78xtZWPU0nXr2oAvUXSdF+xVUa+gCag6Oi8zU2VzDdO
4kLzpOTNzN1aYpUK024CA8bjaa3ZTvvKOUIS8YwJM5oZcv7aq5d53bnews5h3jvpGcR7TwGFILti
933QwfzR/QJkfbhXidytpAb6A+yWFLX0BMY9mZl7Kvh1vpsoOaT9fzqhSMy7RFoGowobiTQOcmgv
nlxgdnNF3skOe7oBlgg3w+B7x+OjTI3fyt3UvAgmg1lTZLZHA+r79/ASjxbwnPwQBqtZN+lq3sgb
n5R1J8+DHm+VYqA6bU/LUCR7v7kdiXLXwlHi3w8HXiAo6lOQTq49gIKRnPwZ/vJPQ8iO4qJ6mxp+
YpOExQzoNz6wxiSDGnbg51AfZEnkrxY82p9JaGYHaEuJyMuD7zp9dAEsyabH1icNP7ay+f7D+CvV
x5+EeH5tltxyPl/r6RleCeXXvoYq8QTVILjAwo0D8u/uGggqnzzF69PhH1ZnuLd7kMo0j4hKJB7e
33hvqFBWlPTxC3r1G+dAhk6QLpMOddcP81NvlQYsTItYpqAM/jWt446mRbCYquZpdTBhnhUW0k3t
WS+f1H8CfakTG7ZjkDfyjS7fQG/Erx4mfRGbozKuMe5UIrTMkCIdN93HsMi1SVEeRxS/zpzDuWW1
Fg4yLaijBvDmHn2wHdkl3u7dBdqpelZXDrRF1RZlcPfNnsjcCi0LAkNP50yTWqM5P6OyPZY3pRfL
NwHdjZ+9RmD2dS97QNhfNZ56oD8Xi09eFPu/iZj9YDzzFtLq0Tg7twU9uceURWSC+xCJPrsu7wyY
ogFMhoBQPQBnRk6v0Zxs4cjIn/U7i+2c503Ayss4OvxtBwa3PCbwsNFVnEI6su7pLcOsSUR2I4r+
I91k+mNZ2p/Jno5qfHbKFECXuJKYR1ZnyfsTMXrFkWepos1x8e6+Ghub4W+vghEktkiSGykPAr9p
gWRBVO2WYJ9RovUiW/g5+R3WEIAJsx2/XnovJmx96w70ymDviGXXUOhcw04wiYgrTrnUsp2Rfhbo
NpgujZvW5U7o1nwCucvk1iCRGvd3ira5RZvc/wsd3CigbRqVMld+OZJ8qUhrXG1InGlvKAynKFGi
3nUPWgJahybcmY9WMupPP/b4dyuF0VQ5xQN5pqdVeprZ5gC5BHkv1gL/1AIitoTm8Sa9Nfn4Jj2Y
hfqi/jXDc9pD74OO7DKg4k8JAb0nNCyuRJwzOOi6DleFndPbCvBGopW8NJYanhpDmBx39oeHv7rW
6lvcRGLu5qNLqO6jTJFqCpMl7DHfenSNg1hOtUrwvViRhkA4v2/GJrW/Pz1LFtm5Dk1sqYfOQBM7
jvIZWzkDKHr5Rl7glPP62HLIehai+vhGScfJA8NtAQkkzmmVZT1D5qcZlmziE+KWETs7V6PeFVcS
DjodOzirycGYJwsA3FXHlPJpkILo9F/tDGZH4kaXvvzt0qAgJgnY1/iCmczqOEDENms3pZ1aLVXI
OvDaT0b9IjgWH6vOwXf1/65g0qNvk2kN3TDFkl1JdbgT5a36nLhX5pErKAcTYwn/ACoEqkrnMmhf
2rzF+Y+XNi6NDFD/81LcIsoWSlQ35oihUFTxkvcSguOkVZwC/W7DZWGru6BcWqUqgiFcbhbiWQc0
/CmB5nvEPo/jX9UFVkdm+QL8gGC/603Cw6Rhf36QdtCtKRnFbM2jmSdvzkCUFTEG0HRFs8foGiV6
f4/FNYr0jw4a/4fSdITKAYUPEQ+WqECoREL//jcg2kHGLJtKTwc3WZqEytipZpY6MLqfPAtkmgP6
XNi1JpxnqXiDyNwWY0jw1m/XsP3vUU4vCzAzLSUDvLc1sy6+xHKtC0pxgLHeF3/KVcbXSiKs+fVe
rRZjPucDiMrUPFLD0k/Ng6jrH0DIvOufIOEZfA33a2UVHFN9oLjZDpy770B2/Fi/slAaT5y26Tb8
HpZB06Ec61xJljVy0iJPeY8pfhsUOVlVYFEkwt7PJz6Etf9Np1ag0ZDAdUb3+Ca5tKGpACVRuBAC
lxEist79ZuFO2vLQss9a0Pf63XZH9xZIDbSPYizeo11HI6M8qV5Dwsz2p4uQiyxsRbtj45JkZvxB
Wuy44C8qerKFd1+n8jUCS3qHYOtTJ3VwqVZaA9zEvCQpkJspYfNwpS9lcrX8F8tqcVRVQxLxsS0b
eq0wGiwwf8jE7TX9pfkZNojk+kLzIc7/0rTRusTJlvM28cZQKjUJJZeRyCbGk+1FcmdQo7DE25hF
jgCH2XZ0F+DN/fIbAhY6fYvDwyPGKcsx9WYbMQZj71rWuCzWTKMACsjCZSeIqWURf+ENlN0no2AD
t35muZQonw8n2/1qD6VQgAJfRUwgvyLCiyE2NHxEFO4CdN4ybpLo/pQpI4pZl1pEzC5kpCUIoiXL
mQ9nyUuEIBl2kV70AImNNp+UgT8dZKiSZLqcf1gCITMNtkg3vAg+W9q0Ah8pPvaShkjw898apCTw
GG7E/NskJyOkD1wJ7Wpqs7IGDFKvtRJ0qw7Fr2npGnSLxTgwvUT6g4kobbHVJlrivDMsfA29sg7o
RLSDD6DZ7LKQe8mpmVUr2DKV/OWpDcrIRQIoApOXGynNXqOAbwD2p6h5roPMgLo+lHCbdt8mr85y
YhadWbKJIur/iqESEE4qnC1ZtC0kHUafKXGX9J27qVdgGY3sV35cup4gvxvXOctzIXn1aq8F6nC3
ITsQNSm7HDpw9TkVLW2vbqqqxkB1JhaoA+uLSfF/rX4j3qk4vhLaSuGePqXuOAOdKcsw6Yzb9Wby
+BFu5xvVsL76FZu5bPzP/rwUkWjCt4/uW1q6+QQzcRP5RkGzNfoiH4QtJHSq7vtAZbYHrhUbH00i
VUdH2t43x98Rc6LQ0vcwKyr/e4RFcmZ/1HTNakr0hFtfDA+IrOXiqAzQff/RN2ZPRnoAZVn5potj
oxpKbzDoXx+ByecWwjRqrKwk/kFooSza1sNppCsNeZB/VfO8OWNu3rN6nn1DBchOb49/sME7xRMp
Sr8KaM7GNf9UPGW9moTZnLMtiNI6q+4REWmx44zwoMKkNivxasyAjl+43uFXCNtTKzDa7D5UhQvC
LpNTOKp9MxLnGGkhBEbjNfXLzaA1RWxZG4LlJdLu8DI3tHR8YON15rb2mufUH8Jri6TwX19IN3xs
5MnbHfMaSB/GPL+BA9/Wh+bFatGSDrkDbmeDOdLJfsLWM2WLCgL50b1XOeFkzoZy97Nz/x0KWfkW
Yp1f8lG0iTBNV1Urg4uajaE3rvpFXuVHZJkHNirSZBAL53cT5EIVzXIBRx7WVA1d08cb9cxoqBRq
67h5ZHTv/294SwNsuVp414T7z19ZO9xpiL1dyid6olG+1ee+t4PvGyUZBeEhPdHd+YKuzbunESc7
M09ASywo/VwzcQTrfejigWa+Gk5aKgqV2OOKctgcAzmnFcYEnHfeyUz94tTL0JDt9md22O/jodbP
ffqziSFweSN6B1ZkzUnFCKY4KZl3tSM7Dglk3looEwUM5EOIwM/XRdKHtHQ5a12dUYnVHNZwxKGG
t+xU7wsHZDdq7AWF6zM6PnpGaXWNON9SvEOQKTUabL/YESLbMxCL0vFDJ9VRopWd4HE42XFWkw6N
thvPGkHszBjzQp3JIbdEZNQhtG8Zm6VnASGNRF2n3rJQg0A1eqTr8SeYE/N4R27eLYKZYJjqbP9N
HffUTW2CqfhxOQ+NpnmhxiCokFv93jz1QzC/L/+8KEf/YN39BGEIThWbS4QLXAk8HQXH8YROk8ij
c6GkQ0W79O5t1sxhxrgGE4Mz0h/yOGHOKJpjcm7HPh6a3TgryxU6SJaG7CmWtC6uLDkR4xHTzOVQ
IDN1Lts2UOf30HhVqn3VPuxuQQ/6ee/kIMFreOHCGc0uiDE4hpwWxuu0U4CoreaRY6LJwPdzjQXd
2HaSTD2RYhBqG26J9GJKc8Qk9TDd5tm7l3IQGPD1UgfbEW6VvZFr6o2wdUGQ9WegmMo63zF4W3QV
/rshXd9fc5k/fNHirlZObxOpvILKwMlzyjf99klLnSZuPjd529zaBPkh4PKf9b/Ixn6W86kbwk51
loDDmthPJSmitzI5/YKq1uSqY4OiLledSgSNbbViNsjfYuQsGy6IgX06haZxoJbgAoC4BMMBROWD
3kgLvcyOLWutAKyZfOzeOgL4hxC8AbxwvySajvTVSNB9KlH1uuJ7RVO43rLGiO/w5b2kJYV8ErOt
w8q6m3i1k6DxD+hkjmZevJNm22GGXvAoX49IrELJq8IOAAG59tY6l77kYkzZ8gcORNwqoxy6zRSX
5vxpgo+j9CtHHkBtbfs4JRAbjFRBOKggOU5Hd+XAQv/n+ctxCBfDZOfAdvLubzkouXeLlmaI29Qz
a5wD+WcaOL8puPPBzgUxX7tLXOrbLVwt2IDNXmLHFNpPCrGqD8qGhRhC8rY7D03ZqBwYnjcvyg50
nTn+MLgtxhvUnY4B99T2CPjVvUbJbvv5cj5HVYQ/ciOnt5ozMiq/maLkBK9SFXoTZsYDwCK11Ant
KSKut/OLuWMIDQzFpjlSiyeIA8+O6FVB2VCLzq6bvS1nC2U6mGC2xyMXdiemF6bzYqs9tRr0FLJd
QMbD5Wkp8DTzWOprNA/CRckFvHYbck5YxY+5Q7SxyUutvLSx+cpm0d+wcTm3B+hSk6vcq2cQhVA/
VUnFuIN5QRDnvVCh3jxpGjeNyx1+ekSEMVIaGKFDQhSIdx3rqXkSHD03SVhbRTS0SM6WT3DKf2Ue
c4YCvC86jzreIeGloO6/zIZwL3wwj3Dt0eLPl3NRhUmAF7SdcU4eCrHZfLw2N4HvECBqYwZlIStB
gUMKUcNL61qHTdd7xQgIpCatinVcm8dV7mlWnu6V+pCKB5Vx3WIIQTGPRm8/UyWukvuUHRrr7QEk
c9yA6SVyBOhUPghmAVHCEo4+ap0CseIrs7ilu7Y6hKafeUMrgzzcTl8+qNoUZpjUeZLNyjXBI+nm
LIRAzQi3NnOKBDEhiuFG1kXIYgp1hP684QWRUSI0Oep57+ZeJo/tLRa+FekV45dgOKI4Fuwq2JQt
RMzHnC5n3Ydn9vQJifgFnuVCy1yPmPkpod7HAK+4Sui+1wvtFMkEIpIUe86n+RtCbaW/gMnPnONU
zQ+YjnLkKnqILawx+AxMX4qZynFB4qIMmaUGHNCsz+xOUe8yFhLMxatjb7frISrxusAhr4o5x+Jv
1Bz7PQbYEnrlvwkfwLigObYTKYz6cpHAV4vNGe1tbaw8FrAhjpcrWB3GiU5VaqP1oqTTjPcuD1r8
bMS2SxbmWoSp9/zgZNJm0DC7RdtQMzRuAxcF9x11+cl9pd3IKkGjRwcSvpw/L0KoNXwxQ8bsl7vx
ntGNPcTwnrFeh4cFFmkYo+mZFVZr3M1R5G2kmFrB/CMRq+i6AVF1FaDXTBCtpkggZ9E0vyFc3VaC
TNGklx0TFMuEUpQkyk0pkQKPnBBsPANbjsGxeWJCDcOhBkLG0L4PKiJOZzGOwe4Sgo4Anj8+ZX8b
77TUbCW+6DHyyRpFcGokGwoumBJySgNIutqNlXlffyF4dc7/zB9voLI65puymobw3Olr+Gha5O5I
x+gXbGq1hEcZqH3DTp/jRMiEIIhT+E0gKqf9KyeYLxiRNd3jqElo4saSbNTzuvpJR1mwjhYCQv0F
YdUnIWvzlLssIja3beFCiRUq5ZU7goi1bSBMh4OpGFqP1bx2tPHCCj1okfV3uTt1RNJitZj5oDsY
TN465mZt9mC8/rlkapf3QmGzECdzPhe0GTkg+Kdcs670kMQuATzNEAjWmHFjhZNpYkVEhXm8vmWO
TtT+F+wHzbl5GbahsCKqACcAlai3XiONBzLPYMx+TNDHHBnCh7oLLpZcOCb86TbiwPUbkCaCFreD
cKnTpNfraS0zMMCQfMb8uBDeSzCqHhKANbbyFxa2SIrpzckSj26NtxfR5qu300AT4H3/GossDW3j
ARs8LdGUDWmSzTtDXskS5F5QlnjlVsF1lrOhEtwL47vRvq/Gpij/VO8FhQETlP1Vvz++RNZ/weeG
shf25HedMBaqweXwKy+pBRfgNtgG7r0/pevHBVIueQyQqkrF2wwh7oxiYBTdVJeafeQPhjt2bPiM
pCMTVM/GOissKpjn41Sds52hy0MR9fx3fWCZf2uFo4gL2umakAN1BtBFXk5nzAZGxYky+gZBkFDi
8AV6NU8Mg/4vorhvQCEBvx5WoAxSmwoTIqRRttxK+rLJEwNeEQ8a0OXLpQ5XJR0MJvXiIT83cfLF
AjTeJsnCWTQGCfe8kb7GJ7Zogd4+b8F539sZiuR1AMKSF8RN5ojC3OkI+5/xYh4/kw27J+teobSN
0is2Hxa3Ht5kp4y2cfj1/EQCJaswKCtiZJy4+beAxE28gbZzBZWm/2jH1jkq2xtFvUyiYycHkwQ1
onw35vik5DDDFSP3wg+rdo1eNj7qt/HvGz8RoVEIDRKbHFUd9QNq8Xa4QxgoHyjBiPYHTANdELgJ
20q3hK4i0Y+bjoVe1IVl5AyUlzfRdKd15SnzEkerXA8oLthZ9QQlwtMExTZ+BNjIqSBad7WsIGAU
fibZiFjqkqDwfMbT6ZvAasrbZlIfOLEhn7cGjrTiAfmZlemqwRKUvTful3Ef/rf64qj5x3ep58kx
XW6cOONClz8MbpsnX3Wdkc3l0rXXvn61nE6hRWEqbMkNUvSUarA0SSvCfKk1lldi8CqN3bwDHQcn
2xdOh1iMUiWw0kAUg87GG9FwI7JoQAenjLBKrEFO7N7y4KJgfMjB5vGM5ImKvR4HaXkTFhIT8e9w
0C3y/y3ydf3lMmnd3Rlc1ANMQ3Jo9k3LjH6OKhLvbJ2fadgiITMpa1yzWZrZXVIL77EHLo64nz6R
i8VE6e7qCJu6mIjdgplF3JcTy4KZosqrwNWcyzuaLDe44Vs5yiR8NpYLGvkA3uAFunsJHqrVUde7
bTq/uVjmcoeZW91NICRXMrS5Y3nTEfMVmoXqViTa8aaPQde3AwsHxqOIusegeMePgX1Wgpq1PUqK
Kx5oaxMQgo4C6YU/J0hHal5wOTIYK8hAGLF0cUdHxApv9G5lBNN7LNh0BcKhhIWrYMm5i6tcA2bn
v+cz/VMpWiW89pA4H4gbz56U8N0kvQ6kc1DBBt/gcYwxgh9PXuGhmvjLt8nFEpI0Rh6A5RH+XPzY
4v0lREdxtINGsSOHYy9j8r4Jhrt1DZX3tTV1SmQdBFKCHUWTX1edaCmXZNtCxDGCqQZ4c5fjetzV
f8ddMezd9Bsr0AhTwdwxEnPbAUNs8xyjvLP5vLpz8tY6hfATjoXlm287ZzdAfcx+FYkwvWRXqPeW
WOnuN76/ekrh3jV4/AgjW+cAyKnDoFI+95vggBNjwRkmLS6wNHsw7pt0Xc1iXhKXcVTZmJe8Ivkk
wzBfDSGEwN4dgqMGq6gEnbw3qZ542sPxifAnkgEs3vsETeCzfc619mhVl06b8eWuj0svzM59rtig
qFAL8RrC/6le40vH9AZsEyXFApYRnKvXYqgccOZyMjxQsxu0Hd/O27RuSy3v0NSHNzLOdGwDx7dH
XQD8+vINRKf96H758wFbD05h7DPPsUE6OHgIrYgk2exNV/vQbEq4bA/igfBf6R0HmAP1HknIyI6x
5f/fqvXOPOI+g+aA6DZoplQN94XmRQiEox7QEWIwk16aztHodcJ+QPnkZws4HnXI87HVfPpGe7hp
xoNLHe1bnMzWyJQaWywOhBQIsBV0tKF4uOxvhIo3rYJxZchZNn5k8N88edu5RypCVW5rkUWRLwEU
hJytTEJBTdWDCtvhaqmmzdV3XJKCqrel8T0nfEfi4UnazwMafaYbrSplPrft1eWm9K9FSs71ObiG
F7MXaP4F0+1rjj5zGfdkNORDSYrBj5mQtnBAMtGi1pS6z1VbvLBZS11eBMXgffYbx4/dxiNvUsu3
vhUdnI6kkK4EAH0NbNtmIhjeUT0dwZJLEalbT4uAJqHernX/FYSC0sS+iZBvyH+ZVAgp6ylVepLe
MnT/ysgEArgHWSm7KLHLqIukSFQXsCMaRdGEFXZhwohVj5Ufu3cu+urhUWyLyrPrMDFX/1+Hy1S9
NHPchCwnz3pQ2KMXqeUV6MdvBz+4y1kurQ2VSfNlgJXGTc1UBbIOZ+RMqdAOp2nukVb+Fm0oyc8o
LhHGXdZjTujn8gUJhihunGCwugFeH/YAJdzWr0sJtIjSCY0vi+Fyy9h4WQ8MTdj8uZgVByXhzC2+
r1hIVfq8dlk2I9VyCZn3rRcfPr6omP6+W2oY+KLPlgEL3bhhWvMi+jo/K7t8Smsovlq9RCnYbI5P
8FAsElNI/PRBsEcS9Q5pL+SX4yLU9+L5pHVv9HER0uv0/NvK0X7hp1gVrX7jh2bCKdM1Y17UzdQV
JLtwdPj4e86xk9nRjgDBvr6fjPrpurJSkDlTdLjsCuH+1uWU1cSZzfwAQgv+eoUG5QfIMZSxi/j2
vqlX0ItZekQnzcOIAJDUWK9u79eZgXBY9gFCQH6tVpi3Iz7++JqR1hh92G+GOlXtQ72Q1xkybcqN
nZQW3GPr/irryCzjtGZ3rCzZFwwdTBcISLoOUOmq7QoeG3asQY2f3M1Sqg6r1uzUV6V3yvrIsCdh
zK8I5M6aN9oW+F9HPH83/xizCQCnqL8ycbTz1M/9SVikYtrGrU0/pNXemOU5YrvbFAmDjiYxiItS
HEkV+Vxt9A64fzrggtzJoGsdk/TrGOAfSkXlSh1dt/B+EcocUW74Z3iPi9Yf4OTGrbTaCxjIT7xw
+EuBKnaTbrGL6rpoR5LjuE1RyW8vUWa3ns1yGgmbXOq6UEC2DypIMHYPlJ95Nt0nSXLQdzd+qui+
KU4giAiBAuZbpoRgNusOntP26dvaIEA/+pxO+1jt05lqtB2s5lhlgRxS+kd5gXrWFvDJclb6Vo0B
HWbn7pa/jtnhVABvDw9Yrk1AZVKxiHs7D4Uv3N29j0LQsygwlNy2x+Y7Y2Vgnlg9RNCgDL9Q8ZEc
kXyXxUz/Ikm41HLS8wYVMW82y6qpgcvfv5K8T/Qnefrh2wq4vy5MmV93656vqLlozEkqTDBguVcp
s9t6FnUD75MCN9k8ApTNxHkmpBrc7Etl4sNrmoRfraJmOMgVqfuXCpieACfO3b+swdXleWEzp5hP
sB8Gc2v5tO59IRZwjiID4joNPvG5goPu0/E7OlSOJF4R69XgkEI6uPFO2ngP1g2CiiQcn6BzYr6U
5BGOsNUMochlDlSC5noqPAGxu2MZo6HnQVFIAHkBTJ0yky9Is7sfzAwqg4MmsWNNid4YS8gS5vfC
oWgs9cBkU+B+c+IiL+sXNGoypKjB+MzA3K/Q7ywmzO7O+y+rxRngQRsjtHsS2blUFSMuuYqoNI3L
UD32kqTD4ReXSMtt/VUraEXiXfDvDDntFK9wMfXRRKmcgeM+iYMPMY87SMeHLHB2rV8sbtW9H6De
BzfHzH31gZx3b47a6d/ArGu3JbqopcojdFffvDe3sy0FTFrCYZLWZ/cX8/W7Juf7Rmzfnks7S0wi
trEnkM1/e3mmg3uKaF4qPOCdItKEOp6ym7XhCllz2VCXHYOAf/mtz2bNc8TkqRsPmckq1AiqJawd
oQjlJjzXzpc6cLzj9VY/ABWdXSFrmoHJH+ik0eZP8MfRC6MWVmpA35edvQImkTxe9NVP/X6TwK6D
VZoCsaMshx8LB+DFFMxGT6xPAe0jeH+/+seODvHf4ApGVLckh83RMjO4UECgZLVLWWxRi5BXBAR+
btcbiAnVbFLSyi3glNI8fVz605XIC9UA4RDc+rgBUpZkIK2qfMA5/GYpkebnjRcu6ZNGk1HkkwlQ
GcMRO4Svaxl9Si8BOCkE4+caOazNTCSBAoEf6q5XBIB6aYl/nrf2fkzZdMF0dngNiIUXhPIDLdew
azaRUZ6rpygQ1tdfQ69GIWIf9WnWIf7YNBz4RfN9IcxiUHQU432JhgsQegz9n8DQQ7KK1zm6Vgt6
cjZZWoA/rFMtg1q7LHXBBuAEq7xUxKnkPyPb2lOQ2LfDCotz3wKc6RjmVw6D+am6hHNqc8pr59pY
GvWQdvwD7WTZzDT+t7UZEcocTisu2AJvuOfkY7kRwBvRaSmM/K4QqkI1ROdrakwSqNAJhDCiyKPv
T1rnPfMWGKpNTrpYnh8jwPItp2kFXO3dSwPFxzteQLlRBfWof0geWkh/GLW49NSzxEcvJt7YhWTG
TayL3IhSs2Udd926PYdgrCv6NfL9DDZ1bq5wiNI7SQ5tqjd6ZUxdzrgi2jB6++XbXspxLJedd89z
UjWCVHwAdzGxnAps2IWIyo6I2Fx8aEVrWD5LdMffr7/Im1KWLWRixwmzR3OLvf3ZHAN10HDGQI4D
4m17xDFbJKMuKkECuklIxqNtPMAjfDF98kGn1NxLybnI/q9BYcKUfELgSeCOP9ME/wdK9DUclQD9
ueAGxBVzlBv5u5rbWLCymOh5WqIRrMWJt+TNefcp/hIPS3b+SMwPsL9ecSABm/BP0yYZR88fXCA0
q1nytfFwSuMD56sw+JIyEaY3O3DcRTofXF7jr2r328zQ19dUoBu3/qyhGzvLKIg6meB4J5FBC+dw
sAaeZZAfTqF5qRd1yZ9HbPjShzlKO/rNgkyjoe8k8yLJFE9HreBjD0agKcgdEnk8INfPVA1TWUOl
EOL07XT212Ai6OBV/cWpEVkp1Psvl122VUwOtZo7HbF9MvTMByb8eGQ00PVd7Zx4RhNWFOxTZRJM
51NJzdTNOIjL3zXrOVh8mnalE0jxFJq9txO/HmKLKNDOTNEcjVyCy4k5vqjVv5a/yRFPj2LnTSWV
nUwsz7QdBhDxGAi50LbzXr4tx8IAAGRJl7ypMzUEwFrKEITIbXhJJnRXxhLQOaElq64zT/ET7x8G
X42ufb95l5bBLx1XcPlHXGDXK2QYCXL76tC8tNaXoNQCuW3J05GvpbPYmRFE2hcPn9iMU6D4E8LI
hcsHm7z92GE1Ng8zH4QkLizQ02uClJBT7AZ6Olvi3tWmw6B/lQxtevd8NCmUtvoIAkQu/CDttYFR
T9LM9oAjUw+x8NuECCIvRDGiZDndtu4QL4PF153wxV/0zO7+6/F6PCN9eB1XnH18iesLut1516Jj
BC6r99I9WSEFy2m0vZl86lka8IkrZJoXArIj+A6WiVs09N29CtGCAYzgPOqqCB5vThfBYLdshCWB
csD6Z/Laumc9/OyM7dH9Sr2DmbQ/aP9i5tuWgPIiUEO/r4kwE6D/K3KPFpZFXdnqczoi3wK501G5
x1kcwyhGEQNZJKHLTG8BqyUV8bYn+zXVjZizYkYo3uvKGMuyql5dAdQmuhjxu31urFXsnn4R8c4Y
pypn+H6fPtNCiv3suXDiOx6nFZCxMVlu2M9c2MRyZtpryejvqbg+elMHs0F6b5zdthOzzjxofKjO
FiWHNcPDmLKsh9q1n4CsNeV9mJ/+sx3rtq9L503Vt5OVBUBIb7N9CdJh8hXKfYkn9L5WbpG8yMrO
pdSfVUQLNgT3ujz6sMXci6A9ze4SCthwG+USupOT0rVACMSgZhXTtB8dSLOb5NjdT3rPpb3ClBkB
fneXQxv0kXBvJUsTHJOtJzJGjo9nSvymx3AirNUJ8tzpy8tONthAXWyImuYzEXeYqpUpAL2TIp5y
PrUsbA381AcSTldpDMZtqoL2xlpv2R9Y83lI6qg0rtfBBP54XNnuR1DEYNuq3YYl1yVQl6xJhJc0
/35vnIfk3PDO6VQqCUeGFBTWqCP1Ir4llT2vuAR1CM05Zu7o9rA5KcwkMe6aww8omFE7xllsKRgf
MS7yjIJy5orTNVXvMR3XC23T4fU76+5ewlGf5HMXXlGDRaxwtG0Q1bDrgeDR4Lbwq9+mXcruLspT
IFg1akieobTh155Ord2cejRvxepp5Vkv/EbIEbTrxgDXPZjRj1YDS9ywpCl0eKjVlTOdPTA24+lx
n6cEn9JhcQBZf2zGyMcMkIMNndSam+BPwR12OvH2nsa4xthxZDZt8KSQfcCh4zo8WbzkLhP9cSJE
DgONOPq0XZ/FaH3vf1gAMoRtFCQkgNsKPV3X1z5P3gUie4uxCKUp/+NWxYPD6vi4Id/424qaBqox
A4/Rm963xcEjSsmDgDn549yIda1JyRuzPKU8KwCzYnZEBYB+UyrD9mq7q54UeLfud9IOXCdE8dLf
aqb+DoCwu4LZ2no6rBAPyCkN4k5vSKktFjHeftsW8zNEeEihVZEfvn7sXuv+O4Nx86wG2et/Y5cY
fNTThejnhKXRGw/gbivRqpSZ/67fcZfF594p6z42/pPu5Fb1NrDV53Lxy8VN6l1Vt2a/yqZUtqie
MlUVjySZ32GYpFS2NaK1CbqdxX4PPula10O5udM+4dj1TIY7cK9U5EYkSrBoUQbiHsZ3LSDwqKqG
qjWg3T3Tt8xqV89tRPeFzKR0QNSQJ9/laU84k6F37gcHVsphlPPy+87JblCNGUxYX+gRulnske8u
0HMgtDTUANlK8P39rhw43QfELBv3lIUW61klCLt9PLSJzf/Y/0a3v7QJOlAjPjimJx795qTl3+xl
NCuj5Sa5TaHtemQEwN5jRLPtQFYZ4VGC9hbX7IEWRFnX62WSE95LPDYIhU9poxo43B78w9AYEvvo
iefIiSQugZ0xajio//uOkWmkrc3tFR3SifEWiLFTkzzgKWrrV1dpDXppa2WCXZiOj8NDvOGk/9If
3ZChtfsIZEYEo9dfYHSFs0jyVkUqHLw7HUoSFR1H+9lUPIHkj4WBTlb7eNpeeoxnayV1T3a5pRQX
nroDizwdvU2gi/AjoXOEQiRdqatrzirPYEwQM7LeXcHQrv16ur3mvekOwZjFkIBgnkjcLPr3W95+
1m5mCiXTKW53JKtMPNlsckNkVgZIdUT3OpItfVzJ/+zZKlA08EMhe9KumH/SxkiZ7i/0SPHSmtpR
FBbKWo7yCSm6Kmw5kHCvUhl7cG/pIiEhchIl/AFYuPViUCMZV3cU/Su87CpBbr+5UxM1R9ckQyT1
2DxvEjl6Vnx3gW7A7HXUyNZediq8Fr3RR3DGWpAYM0QbP4+6OohpwKTyiPYhYSXV9Qp+ccbMLxWF
j3H6oOtuzKqwuKjoDofkv+KVmaQ0PM/sQaNkpjNe4q8juIDYVMcHpy5WopadzANzJu5Nl80lLgOW
5MSGfkZ9vqNepJJ/6v4Y0rTXCSvzhMfr1VeUCyZb9Ml/Cwcx6P5Blc3zCV9xPcv3XtvvDnA+MGEs
sHDBl/dkGv/E40Let7r2iu9n2KpaJtynmHS6OkMfAEFRhL5VfItPlRDy+xIWJiQyo8jt6VKdAvbW
IIz0fuZvMFD9hFwY6hbgYxHvwIqk63yFc7XJPLX6ffKEvBGi5GXK7Vwhu8pc32u+YtlXcpBHyPSp
j6zREx/NnYewLS01CTSeWXztm8s+XbTtIm+aEsmCaZLxrhknJO/Ik4eCL/Uk0VC0iWpliB6FD1di
tkDOeNL4M03Uc0jlWFZj2khgvJ/fh0ueKDvokS1USOyxmkfw1K+RgjVRzvXfDyi3Cv9PzGgrLA0c
oiefoW9EgmHPZ1X03JLZ6xsCtHZ18QPtnau+DtIIsaCKj7ua8DCXfQOOqwm+jtGRuV6ZVd3JRrl6
PLUWA6tI/g7JMXD5oqtkcm9tY9FDRZefF2gzK8fOnEgW0yWhJdSWMyAXLvdBZ1wJwQrL6fwNXIBg
XHGhOQxtkyHOZ9x9Du422A9W/222AkhV7OlPk2arASjk1vLF8W1GTR3euXyxnA+6TfaTF2poDAzJ
lm+pRPpVcBH6abyY0gRmYp5cS4jWxLsCWbLU5rJq9H+h2vGvwzJrWQU/V5zr7GYkK7yI1u32UJAx
L5Of86L/JA9aU8clA6PxjOt4Zb4PJBLdhSV5FoQYpFbHtbSzmZOI2b6qFOcLfhJ4gjfFZcRxuX4j
B2nMY0tn3XFwe2Z9Zzvf69+EvHLysyIfRuosIfVitN8t/h8IfV6fxfKZvh+Tg6pNgy5BsGll0Yfj
Jr327XUS9d+F9MDhl4FzBHYRSWY3pxCavjZsPtkFVe4AMUoM6nLXWFeu61I1hWgMjsiqVmerK2Ol
01dKQQeWX3Vn4ufvDYmbfde083LWbpAlJ3t6xtAxw/nDxTaHuq+QghySSCAV/THpWy7gMbEd42Zt
1XMENArYOl72qOM2cjnQNuUsFa4tjRHTs8Vn4wu5OknE0c0mXdkC0vQ8qCtL1/ACzVT1ypkCGii9
6fMX8M4yP4glDh2ppikL9RF0npGzcbvnnrMiPvW0fad7ccCbZoxg2ocUhOg6kgJ6dSUrVkbRz/sG
mgItIYIM5mISuanR4V5F1COc6SIncVI3JANQ269p/ZqMIxCBu5jHjJn1fNB/pEGMnY+SrxrOAh1Z
o6GjDUcc+qDew0mIlPYmkW5Omu0TjqKonKxNw9xoJlchhyzIUBIrwK3eewY70eUgSavNs08danmt
qgDZ9SJbiaqFzl1YxSBGC9j0Akx+qEVX+TJf8cjVU8Kp8ZkUqapd//HzdlUErZnIFIbCt/VzLFJP
wZGX5H9DoDFgjPas/ZhZ1Pj6qBYmlJvTbPdvEvRpL+FB3IQ/x54WP5uZrWN8z6T7QsXHR/p3LIVn
zvZrNnxfP57KNQ3gLv/BkR7+exmUhT5cnBBdhvvpMsnstLFFirVKBaEfkNTYnQYEaBo3Hlgi/fnN
e4lVFHERHeQkrAImrqMNdNt/OdI0tAEmQBvsxFIe3curWOEfn7sRhG57T2BBjMW5Pik4PcjSsZlp
wHmOE3ziKr+Jlfo1YBEY0/D+BoVD7JDgAE5bM8BrCjp07HEcFVFpxHx6JdK1xzhuQrmaSXl/1vSh
KUit15Yck1UEZZH7j7ImqitO9TVxCWvSaWwi0B2RnfMdURBPCzB1aN0tOos/vUWlE2pvsz0z25oy
khBe1tig7A6ODXQQS21Lb3we2ZFQSffqcVZJM90T01Fl6hXr+fA6THLsigpu2Kbr10cH1dmpbLu1
GWN/4ab/V73jePBQtQwzMs49eYmYkRG7z0eilU3l2SyYLVLibzmrqA9bS5zrdyncaGV4mb0IxeTx
vofcdLZz2/0yB0ldBjgfdmIlsh42LOuJd7ndfmUdO/6PksODQymw62L3iabiet6bL+yiOWeHMWPs
rQVIQ8408pRXgvs+QD3jzdfWzYqmTd3jul44EdyAhRVStjhFOMRLOLmTe5G5eL/UxbcUjFyBx9Tt
eljIosGVok1awjGHETFwp9R2JroxhtHwGVj1PdfBq8CKdNyc9o1a6nI0+OS/XRzKcNn1NU4D8ouX
TLdktQCurHIdyPP7EB85+J5ub36JAdwpQWrsABwNMgRDapWihZYOKlG4CUk78d31qh7DTERLZ8W1
fmG3fzGBelvGbZ70WG329/h4dxi/2aPbuPP+H/OsOjevM6Myy0Pq2d/tk/P+pvViln5746Z6hNEw
ZEW9QTUDzR7/9P2AHv30DRM3btxWSpsbEAFCO4U68RQj44x1PNoOnCjKL2PHDP1JyZb+GUZpbgVw
rKL7aqHWIwlRfFxwS2lsJ0Xg1kwo3//MyLOBmrsLWi2wzKyBVqkVC4npsJjvsBdpMCCA1/5byQOr
86VGiov+1DYEUAiCHaV0574q2Y9uKBl12d1j9EHuoTctGvb/F0ovqDqW6d+7hXrCaibg32UAAj6o
ET0/dEfc8/EGR3ku819xhdJpCRDy+ROUySVA6y09UKaKhXrUlXKEHGrHAz/Uw5sjyP3urZTL1pZM
Sd8yW3CnDfjVBnQFmIbasNDj93qoo0b4OHKntluNFfMD9VcwQSPZQoxd0ya5rJ/zyWqrT2C6t+p0
I3nWXojic+MjsnhDOkKxRJFesh1GBMwPAiJKQGXO6Th36CapiT04sfo8BtjdD3gnc+BAQ5QU4uZf
pq254oqJhq31nUzxDpVUTuAPe77THSwMagBTNkgn55Xn+X84qGft7GuVBmecWyDQjRiomap3Jl9+
HfK8dBs992NtpixNBtAE713m+yf03uus2J27CKiNvywfrcbWENiOLLYio8OsLEJVlReNFFbU+Yg3
TIROyNXdx7qSeeRGAL1OySfxz6XJ2OderfUCViFL+hqLo817jRgZ/IyItxixHL/xBDPv+cfWOyn5
aSUJl27TJPmQ27orMhYcc1Mki1HGoY8shRPuqHCcIjpwkuc98/diFVO5e10PhBdDcYXd8CaFtojH
ekE4m8DttDzU7DNasxI4kg65l38TLEfaS6gZuK+UiMBF6kg4QTfZbI/k+1qhoy0F8SSvLI67S020
bcAIteUOoQ2UceFWN4R1yr9GfKOmBVcD3IeIChVt5YnkxLdQGtCKpVqXhLDsG/n6EZdnWrCyMcUu
ateKizog8BTx9lMpCa5SdXnIK5TKFOblzrG581U1BIJumJM3AbA8zz5KisPjPtVKeAyfFoeN8TV7
JKcNM+NY/YS4QkN/T7pb0WtwSZkdhOVnaWSkiT/8tTncl1GHh4hFIty6lV9Lh2xVI6p9LxA0gwhG
WRzS25WUSJ46ZaJmQhPDyGztdhYsX5ELSyzjwlA5ayi08vAUF/YzQhMMIySHKv7tyEvx9NyZb/Yk
AEyFH3VSQtEYmpDpGR8nur2ZPUPMpXx9fJpgQmVzfdm9U0gOQIi7ajOs6ox+N0VIy0eEvHHQHhwh
dxVi/UMk17sB0NtXX9VIMX5KYG2Vh0Egfmp1cEJ7TVcOL5PGmeqWLGCp3OoZMvsWFhgtXSBYHNq7
AjecVFVpkuE4hXR1UVUJE9iySaew1kGz0w6FUwETqg0ZFXs9F6ANb03RHuDhgyYGa/QpUBmJYIT6
7dMocB9IpRejijk2pVu1WSKZJ6G7BkjsuZTAWAVRWBWVbxUzzlSgXL/14urLOKgKJ+9bl8Cqfjg+
CL+JHoiu7GVOuf5ODa2wO11EFLD7mV/nu8UmsV0WGoSxFqawIbjAdvWCPxoJ9n1GDvFOqKfN+vVa
D2dEnbxx0dhCNQnrwf8AzVRIBABOXzWuv/WPrApSn53PnmteiWlH/EKd2Tj5gaoDQlnH5rZXcPJx
v8PlzGKFOLi/h6IV7COjaudLb3Np8O3MTn9MgR/0g5lm08LH5VoFIy1AeHabD03nMTvKJdYiqOC/
vEL82ZSet5AC2qzhkkf8kcmZC+QkEW6kQ6NX9UqUXRu6ot8fkPuGGesyo3/rmVwUqZHVmHyY9XmT
rJKkaVQ0wo/9pshe4ILwKYd4YtpC7z7mm1r3rVprf7t57UUTs3KRDf9Ag3bj3SXM3zY3fXJg/X1C
weIa6AsqOhRU0+4kc271RBeKVeT0dt5H4xJwQb256uyJHf/XnDsRPzWVhu83OE1uaVj/ipq7pSBi
zA74f5r3eqZXQ3CwyM5TwPGVKHxtb252ZoGiJpxXLc7kPgngJiYHgfMjyfgmv6f8yk+oLXmB/11P
uJfKcI1/r1RRZHsydisrzGreOQhPCjAbbI3et+gSKbOn7W7QykCNw+tepC316qc+IPNufvBJ+fo7
a6oACaqJtAYErGLhczVlgiCHyK4Thn+7/ew6kC/lUu6a/2z15FEhHkfYKEK4cKJWazR0O4Bh8Kse
3zUd4Vo8NZGkCLx7e2cuDU78KWcgVWe5r+tdy3q68nzuLKqja2jze9fnPzGa3EJWKj1vgdqXrpN0
Gvkd8Q9KY7Ke3JFrHa8KPkKTocxlf/+TSR0+ZfgYVWRiYKy35B7AXcNvEe+vlMKG0LvOIiAga/XR
nW2Zpr6X1WXllRrQN2+pU1h/+RcpxXQKpn3/tsZeFvVV0JDrFaYQm4I6yTvuxGk0TRB/x93vXaYb
SdFL2JuI7ULLqz9Dk/axxykpoEQNeNk+pvnIujvWQoeWdS+Ux5nU9bDTgAURTkEY31ej4TPlwtCO
Lu1ggUl4ZlXY16Jufgh0ttEKaUug6pnqDJ6AZn+WvD4Y8jfu1ieOvILZqAWiTO5uQTZ6K0rzQyHi
m/AV9j38uOtl2/xs4PhMWrRPGgUdXh6tM37ofKdCoMfVDKohcgCpZCzt6WmKlQS93Ei3cxCL1Fwh
402+XJcheOIOYzwZQG8iNUvfujHDLO19sXCt9KlX1xpjpr2yG5dxDXH3P0kqn7ur/BE1smM17BY6
DBhkYYbt/6tyY9hgA399zUlfGcICMLAn6W9sdgUs6TY1OxXtC1+kyg5GEhBV4o8RShDieWpMgz/x
5qhvsJ2pyDgb4fV0r0/82mhoPlgP8YKjKec2uTKAbLKCI6BM74s85onkP3JoZVJn3PgCB0X0u9IU
tYxhDNPbKi+BRaHG7LbRGBeGeudNYnsmKNrZ9avO0iDPMfWXYXiHzUrh6OjZi31/js3+mBALDJb9
9FDtbW9bq2CFCpBMjb9JkeyE0a0MdV+xSlPs8TAsJTYbqH30pUCvLjtyjtiKaXmHho+A+DKAAqce
D7ymymvZByN6Me00N+81yK1T4divkhMkUMLHJh3jnJ4vQvS91X+63RjX3gWT4CmvnmlVqlakVjYv
nTvEwhLucWt4L8ridnOfhMDZUrTTX7uSOz1+AEWd3M9/X9MXoEdt9un1ztIlDn8JonriBcz6gGah
opYfa66RdDOeOl5akgss9bOEoVxyfu4pWqgnmXXwkuWzzSjsC5qeS5eoq/zUE/Xm9VwVw46liCju
2aH5S2vvK9jPW/mVTD+fH/lz9UtLBxhUj4/BaOdnOPnjH/vfDQ+iaWiEopt+vy9z0V7OdoiEuz72
RlQvW6MVh579CBDR7Kxn7rRiPvRzOXhSdzX747Oaj4hAR4aEpqfa7pIal8uZFy57NQVCE4ts8otY
ljxObEsZPd78tP8tjb3lZYldYN1G/aEmtYZX6Ec5ARtiOm1MQYx72AsapERk3eywX8gLRgGbV7uW
ylXyYt/ZZR5eG3oY31JLteSEn6Jjtb9KBtXhgtM4pOILIUsm0T0/M/kL9+CCTyC/wjNEDlrgO37w
TnFDCNrd6y7XaDTFSHyAqJjLrYulcLEgeJgPBbUfuScKuHhFKUqFGQGqYlKvSE1hJPrkuh8cjfDf
eMBmZebRE43YQUJ2FomUW+a+fLJsNttwUfUqxdGNE4de/lXqwg74qXhPcgG3lAJE5uDizFGfb5k+
vQ7uh0HTEh+I1+EDpO7eH6346HPz3rnVsOCxUyIlSrKjULIT+JUhW2qtSWIxMd/GrliHAovR4zMK
Gc06NSzIt/X+kbHIxpCNGRyGqWgH+siXY0J73CKGhlcBwW2vEcFMtppWiESKnE7Gz52npwXNLgZR
CPt2TvrP8Y/BHKD1HDcwTUJygldx4lVGU1JdjLY4tC594cV/NuD9eZM+w8+0eB4tPmVwSLdDgwcE
C4tBhTM+nTQ2q/73uS4mVX8g4NUQJv88j/MQfjIxqMxxXQTZpeKmI8vjf9aP/KHpOJ3CVhgV0ozo
SHugUDcqth4Edmzhbb3he66U9fZA+ZY7WlCWWndbarpcMjpA9G4SnAnY3GhnySZcAObNnKNH8VIL
pBPkONx4b3vOsllyYIOOno0HyvYz3M4eHeO3dhS5XVumzS9kC6IIXrdPFw7MBGAFs9AKwZ2tM/vL
vkKtm3kVSMLUk4jkAvE8pDIt6rb/5816iM7VqVOYctPaZ0L4Qq/rlTTCOy9mfvSxZBbrVPX9NGa6
vc50MPycx41z1FYqUJsUVh3akjVCrvEMCBaG1eSOTdvP5cajdLiZjxitRHFwxBjza9+naI3oy6uU
IaQz4PZ1EkC+fkuKT9heNl4Ky6m9jEaDMIHDIPCBdfQAauh3d25rF0Xd28k6lGWCPeKF/UjxJnc3
ucRIYTse9xw1caEmIdu6EzgW7rVnvb4LKyc4ybZJhtIUK7KbEoQsBrhbkTFt0MMN50T0T4XV6Kxz
ay8G0g9MhdFrT+D5qrHqOYZhqWp/t97ZrrC7GBFxeFjbucDyZTbdC7ZqIyYlRNdxagu815wBD0WC
h0BUQK3HHNYFaq/IW4wEBviU6Ze2+rmyp966ctjxwUUqDKTw1Z5EvRAsuVcrw1C6NobvVbfWBGAP
5BXz0KYpeuKyp+ebXy4wF82lSodAT7ZG7T0MZkv78N/xQwMqli9JLO+1xrxB/fwGnIsmdNCrYI4R
NjA498KcksswesTP3EAx4gl36DX4zqmBVDSZ3w1cxStranma65vJ64pTvwRbuwzt4jDjnq6YCjfw
N4rUe3OlWISj2F8YjuarjTsg8eSD8o2fCtBqoiwiqchCu1boOJ8Jq1sNm1Gvwb6AKBgqIW1+4k3i
PRD7pc3fPISqbUP6ffHvVCPp4p/ntW0bTaj0TulvyEABCl7ptTp/q1Z3CNQUC91llnNfv+FI1BaX
RgyJYEiXuUTLXDJ0WxRTW0XFSGM5xJSgQ1QnAfYdIHzNi5NmuLhs8UI0pcc55/8TkE+hKuNBmFBM
oHYF64foUM7pTDlB4s7wq705NttCLPD/Qty4xXCGedC2zqXR+tZ0MKZW5eTTmaISidpRF3I9dZ0b
lQh7c8MjDdzYatP2R7jSa9egv6O1WMiHk46fRRXoMrALcBW/cTulDGrTwc6h4Fj+lpyTZzh5Cmwk
xBWfILUzsB7jhwlvtoaF46L0zrnvcKoYrmNu62mAg6wzLYFheecLOo3UuS/s9eVrm53lN1jEbMZW
apAiyJHWM317C8yxZ8qihbf/F+dAGwn9kErMU0wnC0di4dMWTyP0Dk5YceOBMiQTW0+j45JANzVs
PxScUMNDyVSj2rzYcShe1EMErKgXg+BY5a/lXnUzot3APCDJJ7wwQYTg9tHqBGpw2/5m3lckQU8q
JiTpw2VFxA5nggh9HwrGo8jxICymTqAvUpGKTCM/Gel/oJKM+qQPt4nL6jpvMXeogzVmDW6C+i1+
Omd/ftD2K/JwF7eEZskYwMiPVVm82s+pHBBXBzKwjx1rT105oziLp0wlbjoReoa22TyPLk1WXBej
8h5xeWdqSoEQow5ajtzMTxnpZz1vmgW1TUaTclZQbMbNLE63zYF58cGLo8UYStQfyC8fZ84jriS0
UNTgMZT60Sb1MAaor0rps060kPbLgsQ6hCaLpXr9e9sG79Y2FYmGFex4znxQNEel6KZVu8JNkjR+
fKpibWZxdO8z40RsGMRQRpf+j23Auw9lrbUskhbY20d2yHtwGvP1upf2zGElgnq1B3R6DULANgoF
mMd9LpDZSMkvGSpqmGGuOs6juRAVuqWogaxWOtOPYJaEbosrA1WQ1GGrevP4Gl8FOdaKhq+iTQ4S
t9us3wll3MTCToL39i2qzkMu6X3MyJ9F7+YZy5vFo6yfP+FtimdbI/HjB/n7O79IR36QzOvsj4fZ
moJCLE7dMcVFvP0zCELfcfK+OqjAvXlkPoyFJQaEDkYD4bsVYpU1zRdRW5qxE48lBSiHBBqarWMz
E6pVUXZgY3ZzL8OLChrOOo4aAqArnr1BQbuUurQMpDb9GXrUBgNj7Hv2vb8gCzH6fr+9ARsvOxHx
RHMmErXmc0FNTC+wpz1yV8mRalQxFOURxerBZhMVjuRbgdPuJ722DzI9OG+hV9ZQmLBbyht+E2QV
y1dbh1g8UBFvCXVFTYlfj0LcoTcuc1I3yCDgGQDsWbiOsfGLMeBmqGndY8DVHZTIJBXIHoa6b5fS
F5FBkt1hyljAtmJeBoIIaKXnmISCg4+lRGleetDX3RgDAhifg1ONjizGV2tY59kfXInLsTh559m5
SZ9utXAx6CLfN9LEFf3HtYdxy6F/PYIGeKLt4qZ71bCRgQKRtKP98FbCtH+TvLOiUCl6epyQgw+a
I2OKn8XoUh9QUwygFbKNoBh/E+et/btwutGCJQJ5UfbhR9RBBFokL7Li9xW/nMcbpD6G1IP5NUS/
E6AqeEqLWT2wxUxImN6mOYajmLrdjNRCsmTIfJ/+ymRYymga+Fv9C5Oixp4xUM255ejDtsNE/hM9
DhYZi2Lxyz479GJz6IOwcdiz0APhU3Q1aqhpuZObhuCddTUGPhKstRDL6YMKEXAztOM2vgWWP2lE
f4oXptY+Oqmw5+e+jvzT79kXHxDEK4DjhiD4ELEnBYUWSBIPhIqQrsu0I12gg2mnYA6UoHq63KmS
fp7u7qwASDNNbuOKwjF+wbh+/GPcXD6z/GqPIAV934lOrEBbxTcFwH2Oq5yAMBgbUta6CO1/iErp
FhToKH5D3/8Pgl+vS8wmy+UMTEGzdxwNP7MZrZDEiQkLqlrWpwlHEjSHTjvW3vAVUXQ2Agpuz7kI
trNaBihOJCBB6KxbDAvEbjfBHk1cFi6x0de22cIhfoWW6sYIk6dRzbW/GeV2k4towNKBUBBclV2I
I9opgaQTwFHmBjKrE1OdhTCQI+hfyN+/p2WP8BSzTMA7lkEBvW5T7wUxJjo2F5TX79GPUQOL6hlh
nsMjmvT9MDrSOX3pxge7jBzPWntENhCQuqPB6zzKAcIXxlBOK/fLWfFb0TgdTkinMAAZ3JnJzkKc
5fOFXMyxw8SLxbct0TeR94ld6l/PbLXTXuEXkllKtKX5NUq3NCt1PqOAUyw6s9V59WnW/ydqwOQp
iUvYl99AGOqlexCIogh0z++SDIEjHCezcYZsqVQm6CKL8cEULzAsDlRbYDsr62j8FfUaEjLssQhx
tmvE0XW1DhGXzbBOcBwFSK/AzF25jIJtEUzyvk/SZHFEMwnrXExD+x2rYfJt44BbLoL0aj648IvW
UIWCCpDUQ/NxXyXq901wdcqbPBTSK5R6myk8Z6D+z1BhNG5m6gWPel7f97rYzvp0C0EXbza/9/gC
cdoShLDojejl0WgRI06anOmnZm0Fn+E6Xv3WPB/PPGdmBrEUfsZOwhvKWOcLde4IbtDt+a3AVyUW
M76/gEJBilT+rIWFnXTkvN5Ip8dQXZcOG8qM2RYlNg0Qqo+DvDHgyNX4I9DXsMZ1mMCDeQ844TRJ
Z6cJwVnndvcyazs2AUV5i1lFvkwffXtmptNxO8e7gWyah0v2247wFT9tVl5UxEbntGuATmf7yr/0
FReRnJAMG7VS3zgZfwkx3PX6rACckKKpwrJojIyOkk+pG1wcH1XRR+RdctVEgAefYyH6bmv3N1js
d3z/1CiuD0F8QL0x0QKu59FWwu/WItAQ6CuyBTGBrojiUK64ljB4Ex4wcICBq9Cs1L0LmDesAt9D
5zHEt4ZOmpsfk4+kH7xP+qKEsXZ5BLWn/vjAYSJXFqnn+ib1Fw49mRHjtN+gQWNa7ghHN5XOeTlQ
UnTTVdfVS8fyz+9fhKXkxH3L4N6p1maXL40jBTroJ1QtOw33DJalHAVRKIEEB5TdYZB/FugcRyTm
wVzncDSBWs1eBHk6OLXfA4KC0Q5kgoloZdIA0SMgp8LJAibAxOSht7z9EVHu9kXFHroMDDvRp0PZ
SvtEwYJ2uGkQGUN4LJHrxxpJ4kz2t8Qg5m+3+MQ6ALqTXyNXuzZ8fWeQBJkkR9wFYGL77V7VpdDx
BfHyFG3b2rJnEfk8JDEfZ+YOjXGccY9YMmnQCy86bCWCjPvcpzUfVa4xffQtD0fMRHLDHcAOhvPB
lis8XsZcP90rRuYxVQ9+Cq7FpHtf5B71eFMojLmXaB/hRJRrtCZ0X+IIuMhQ+MrnazA7ltvIFBqI
koZFz4sOv2Yc1DOuf+N0HUEq1/w/mPpWsyw3tlvIiJI+U/exF/xIgAPw4x6eRkVT+RZpD79hyKpL
TE1vDm/Cw1ONHvzFavh2P1FZ4fNmeFgiPn9MOB+doTJUnoB8+bPlsjm9CKOPiQ2JG3poyo5t+azz
DZgtRqDNMwJA3bnJyImuSoSd3YEMCQF6dmtkw791/QY+pxj88lxoXVv25bdSXcHvtP9XrrF+NS0d
mCYp9rC4Tf/ygVGY6oAD6MttpSf3rfigkhO888QiWOf4tlVGgK+kvigMw6eLjXJY6ACYynmWH4SP
NmUq0ZWVlgtxlxiI30B52wxKJBGh8BKb81VQrkwgT23xai9zs29LD/vDNaLTQw3JwsN9TBB1xnFK
gLjjteSAwWMq2Mn215t/n2XCqYd0MyJlCNMBY3hDozA/sodhArBAJZ7PpMF6BbWd9JZw+zpaMjx1
q3pR86tJEojNkSontQADBEAxo8Kh0FeYFELrw5PPV8OWXb646k2nJfWo9NBJGQ8Nyv2mLWfiYb4l
73I1sJrFaau9sAH/ycRAp2BH6fhWNVQ2umtAizZSdZ8s4RiHxEimjJP64DwrVEn6jkf04oCYwTdw
alE2Uu3T85Ytm7hXYPXCkOS2WjEE+K9aIUg/KsZ4i09ufbkn+lIu0F8Ap27daoW8mVgay8m9N+kH
d5r1+r2EEYFXIGx5bYowq65TM5gGdaeiFIXVMrmj1k98yIiXiI3c1QRE511ZJ3wuex+z1SMTPN3S
kFsknI9b9P1e5KrBcQ5gJptgfRKBjpuawWgDkY49KAd6gHHSkv4Xq642MxDi34T1TRoHkPdk5sg1
2YxaF/ptcwr0V1eLyQlV5N8nBh80QYhQQ+1WC5Fqj76rVUgGZkspc5lPG8AX94BFzkoF2TDCmOCp
etylb/9uvqjxNaqQz9zKlJyuz0P4UdyUw9X70SsRAPpSqaFjGNluBXNMOtYKfOA0Uwt7ADkJDSrj
0HTNz9CMj+Pc+nAEgXt124siOi8k0PnYQ2ZUU6U0/kHfJUZ0/FWLcwBn3e/pzEv8eCXQcsGURjyC
Jj8cq7mTt9EvqEeYwJdLzUFGLUOqAn0OflZZMZPIoqEjsZ+1NRLQKye53WWVdSNTzl7UZmaLo6Je
eC2PvMSg0Q7XdmnxccPTxkp/aqPZfI4oWC3bJ8YCxKDZwZ0mAbhpT8UK6lDGI/ngNNKkDz7VEkg6
8oYwxth0/lDAYezxSJ74GVImpNMnRpFh4wLzwi7T9TeiK5sB34I5b0FWoDojqi1vzmIGeQmYEuhQ
w2qsgm3GvrYMGg+piQ1uV6pBZrLgYmiBrq9IN1SRomV6LL/9fDV26JWFyGwC1EKdZ1PnMMn7Ixyo
ZECv8ANAa9ZxyeW2TuwX9VAK73lAfu+IOg0Mm7tKCju/ceJqmY9jkkNsnahuv22yDBg9z/HmZTV/
0UdZ6QlLAv5ztKz+Pzulwfcj29elxdVRyaQdP3UMK4fblAE3jniM+q9Za4/QokVkoJHmUGHSjmne
yM7P090uMoRw+Wq+L3AqzxFgma0gHnZgo4POQGyW1xWwF30tXKLiuCVayg1lkfCVFdUmh6GbKI8v
aUAjw5aK3FC8R46mPN9lherVqnzFvRkxMasbT6gH5aqCkEC5HisWYOSVVDavwJHor7ukEQ6FABay
hjnTbDImRin2rtqBiul8oZqgVEjeUWFMdd9aLOWn4Dbhdac5LHqXG1fv2/xLUaFdK+RXn4DufJ2W
Qe8kod9K9PzAaTtCEC7eSp+wrMioWnwDDu+XFYGhIXM9b9rZdwlf4ws7P2krmNdclL5TjQYC4pBU
M5PXvfcLCF5fCJOFQGpZAX7ur8OUv9OERWbmdDwBtV1WRwizwYR9M82Aha7MjCHdm6G0fQ+KBUX3
LLnnKgfk33eGahs5E33JJBm/vSl0zGWJz4ANY7E0/Vlc3k54Afxlt5/IZ7ePIZ2NWL9XY4P3faTk
Xi/18a3CZR6BpeDMQP1YTwnS5bbtvHcL9OX2XISVQYjriyaAwhN3zH4/H66xqzhI3NVqOPAmEb2E
5j6n5Rev1TjOEKhL9SMKe4+2ySvTulZsRX9hdePWwtFB8+raFoVKngOaF+ayNxpXH7NWGpOUcYj9
c59cb9QhPmtk0xAvPNBLk0TSD1KNiwDDqPlW36zED6wDwx2mJPyUs8ajyV2QZFOxDNSQ464TNICh
tvv5RVnyMPEBASjyMRSCvQj8B4fgv54UdbePpzdgYZAbdAgjb1t12rlivJ8lxfSyb4uUUGsjJue3
RSwmaeRFgZx9Xz23x3Atn8/Yd9Vc22INkDKdleiUcYzEZKICd6BE214/MtrusaUzNMhYAYGfDTaJ
G0OdBTB8FJ/40Yx1IS8BVJyL/JUOO1MAckjG0qFZcnO/a0jHRSyrmYXeQyQ9Y0O1+h0HXISd89YG
rYZ94XEvEJ550rwcPKXRrplBaljFwpM6qdU/2YBfpJvrus6GXZshY3T8MDaZ66Ikq80rQ+2hk9Sg
AZpxVulj+LgbtfoQXc6rZ7wwWxjPr2ifjczSFsgPPSzaTlVsLFviXmdfbT0dFkcMX6QPMJnfOuCH
llDIfvK+jjalYK8Vpr4z+UKli/wgjA2jMPbpLfpEsdxi1SUdSJp7yREWCkf9vUO825CA4t6090/k
R/noTH05WsZdFlA61xsUiKYYgk5JusVihErQTD6UQxl5jsov9XG7OQ5I/5tUQGoCAPTwpGloLjGa
86qSNX9vSs2/bwyudiQ3qPHlhrCBSvELFZXMAqwgl8uOJtTVdHyHJM+en6GtIOYXPYK+6otX1xJ/
gbt/JrCM1+vMYZBb8SrGO4CAfJrhoTbsRcKpFYN9ILgVESkegZSUEWQNkHwe1nVVix/O2bw0Aj38
sXGmkSA7GEqoEUtBvK+SFScRSON5ypDkcTT8jFN8e9nShF1vpfN49kV0rx1QkrWBfYqaHHR9/eFV
gNZ0MUSGrwFTVJ2XEHVSDre4LZVbd/oEfnKE5JCklVDMfCz+JliqQtHz+6sS63Q+4c7xFI/ihWwt
KE6McQHY6dPvl4ZIOBZXkWbNkQjIQ3vvhxJXH1xucWW8pQiqBDiH0PiGqosmEunQoVotUnLVM74F
2OXBX+c9H4lPbWueef39kT0JJdx+00sIb2lD/VbTNMI31Mc4DFkZrhipJLpWsmCi3HATIOwmTnJT
tn+mpPL7V3+Y154D9HfsLT34lZS6VAlaUTJMmwimIQFQWcq8ZR3o9cU324QzuCIICqsnc98rahsc
xmYSPkpXhP1vm9wsvE1E64DWXxh1j5j1Ws1K27MLVYaz/zU6mo9x2m17VkuZY4Jd/Sb9pOJVgK2x
usfPh9hoSTwNwhGMxfHbkk5UbPoQfCwvmR4Tw+CBLH3npYUnNthD5ppCxaf1xzrlezLiwKchXYh4
Vo4bc85ELLoYmXUJhN/hqyIu2Ps6bomJKTqXE0mIua2puGj98SCKvBIiOr3D82aCdobjGHd7uDcN
9o2rHGGwKBDco6FnBfXKkqoh7avt++U38x/fv+f7E8W0Phd039pDCPqvFxtu7ZhpK0YgxKBYKXgb
hEq7hmebHOaT+tkcTdhwZ+L7hYNk3LO0qlxGZjFi+vzENTxzvNcYnxrKjiwyCxlvX64zsAu51J3a
bNKWxxwGwJOtVT7+C83G7eLjZeUVR3rW/4gNy41/wpDeKzHIwhxdz+Op7Kf1gdx9dFz5614a3kJF
Wn7DPDxGhXyFvi1RpDRR/yHL2axyvhBFRwzdHlvaaSgJGH1FeDk1udF0ykduF0tbHNcQzZd2QVkH
uzoLzanTxSkuFd+ahmA6uPMxOCQWBlIHlubrCfoV+PIiWkg6ddD9hQm7itVyogIxLfvC3stsroPY
VWwDUSqlMxqg2iX1Um+KEEErJY9AmkzK19fXoAchytvNwKEyiS75KnAZjKQb4Ymclg+CoTglhOkC
D3pImSB1T9EYPCP6taEPtRVPdgZQKChUvdHu7GIdVf2MHPKlMqCgIj7Eqd29BDhT/3h6P9MOG0/y
nTZe/pZJddeym4DKVBHAFjbSUV143z2BgQRfd56XnAijmYXISGIBug7ufh0GUwXroiXe/0Ml2qQl
DKyb4oP/sBzV5IlWGYyA4D9RuIP0FcYUKtsQ9yr4cJPdYT7hoZ1zX00cftUEiSiXzTAFwT20egWA
/vytKo+avGMVKBtVMlkLNuCuFXbGa/S44xQcZMDIoOb4k42GqAzlYxpQ27T9Y5tOIexhklXddO/9
N42WLETlRIDBEHQQYVQ9PPn1n7DYbs18APzhPg1/hsEw9iXBgipdClebU6uwIhb6+Eg/y7EGjBy0
gn+Ioi4sTFk54hoc8izsvXwzhqLSD4YSLbq4HYAMlqBFtftiHOfIGuT/31JmFsP5hqB00g08KP+/
gFH1oWWIEcrz34jcffaqK+lzpjVtyIdLdXCk3PzxoKy7sPM88+veLmUB3ZKCeXoB56onR2D6PmUy
Z7vg99/XwCFKcfoYcmDL20sSqfp5g6p4UtXxUonrILERsmFjHbHEVvq8voKd2BGHd+enWylqyKbb
9oO3Qc2gaTLzC4rIO28VagAlliYBQkTDB9+kZ9xp5qsQ+GsBlqR6sp2jd91ot10I/cK6//SCZr3B
iPR9WwsQZVA1x43A3hQ54Cl4cMiALdeFUYp+7L9MoYyqZPHzDZqBOncwKgFU20ZCPNQPsiPt20Pg
t9RX4X2YXVGmQL0qJulf3bUCWUdPW956+y7fIms/aFacoO4eKXy9xRfwwdXpEscGC4AurBPHkID9
xTQJtmSpZh5OBvZE32evq/+X9QLiyvZI2cJ5CXFFOZoSjapB8ryQGz0MRlbgAltSOcslYKSYMUHh
wXETDwn/hTd11H9o/zE6Mt0IR/FJgEyID2ykSnI85wppuJLHnYcgYNlZic28xouD8M9zgMwSo+ep
MJpTze+rqpal3iYi3zpR8OY8qgNmnGMvINQr45T5Iq82dLHXMHQHMcIhNBjGIP3xKrq/Jnw03Gwv
LlRlN5WdnA5bjjg1AnN3SBs9A4sIw8EzcgQVRapTPgPzBeRdOckIdxLsRzNqX6tkvzZZKvndqFH2
zUftDSZVlL4S6mvVuWZAe4g9Y9BWe3S5GwONRZXY5XYCJOq1PcTBfBuqofcG0aGap2cZbVZarwgV
eGjFTvdRS6nN4ihw/w0n1e8fg0gS0uuBcY2UxQIkpamncUvwA3p8w3xMkzRjjpWQKvJGc/qURGgK
K2Mzu5zBoW09+Sk+Kfk5rpWUXkkw39QiAzpT+mTdgWHldbQLr1FrcqJz+C+dULd1PSmsZwHZiMwL
ZjBBpFEk1iijFOYfTNkQ8hWiOiIv0HOWcr5E1KqpY/rqDf+G06vFjvNvAZaal1O0xg1wwIDRgqXE
l4t+9pAK1W8gPPABAl+BPl7l+IPk/A/warfdhSa2n0KOTK4sI/vPGvXuZJasIADwRyFxfjc6bxe8
qu9v/eE646rpdfUOAMX3Ge9tq1l0eCgdP1vo28TDRcP/AWrLp3aU9vT2N1luhnTKlPXlRC3cPhES
VPwqrsah9kuuErGpkYCR0/nCUN2DoMTifk4aTuGDWYLmchBJpmFLTIHZE0Aaf7DQLKKB5BnNF3be
u1XVFwQ8xp5CEZ90t9/ZA25bT9kdhw+yI08SLRZjViEAy31ZWj4BaK633RYd1T4KIvnWlY6citCa
ro2Nh4ballgT3PAnEoqbP91Dg79s5lz6Z6voHJ+GtT0y649BfIJGg4ZxdyleqajjIsDbkXYcM9Wf
bAx7x0bv9yGdAVnIXar1iMOUuz3Qd1DNcwR2/MSQSzrpaN/AgnUcqjpADoLjIUJ4sovRWmyrxwGq
E0YWRik/T00NCHv/oHwdD+Xw7xQr/xSLKAclkVgJgwbz5XPmB5lJYLxdMedsDpxgLeOWZeOBW3NB
lj2x5bL7pLaEVU4/E6YFGhSHnXkiO0ORG2wgXzgvH3+/GL2npO+Y6tMpq0SCA3JjMMALXznQAXy6
HLRSFl3XcSIGGosy0FSCzdsaKmzF2foN65geZJEa4/kkM7r+tPaLdHzVpr8H5gZ51Gtei2K3r8eo
nbyz7XhuQg62T0B+d6pDnyH+hKiHIN1izx6w9XrxTS62b2F1RQhzI1s9iDm0sXZqhMvkY+DmUyMs
aoNAtrUuQF1eJCk/JJ7ool6AwPcBCRXYWnMgmv3uTPoAm+gLE5+WILgGBbhSQZcac4hu6OLOGrSR
3PTrd7zAauLH0nWhqswNEGfXwpk3Ol71Z1FTcTJRafSin0zPQPP98rDLeQxZ6mzLjcc012VqGKER
jSpu24B4/9H07Xq27xTj0wfo8dsjjgImKlUXStN9zcKcAh3aDJf1AuTzu+ZyKhweLMOfiowCUokL
U3Kn6DtsQ7OB7pkKLnpfV8J7r5yju/8dBdNNUs5VFUpseJUn/kZzeEVvJZnV0wgfyQZwMifGP4pP
g083gIQcYxDtMiRp0/DnPhAW4zlVw6O2mPQiGMoLt9z4ZNbqgpHwRTAfJNttvOf3E6FzmuxawdBX
1jKah70QAWy+degdc+WQAC++N2q/Qs9AmAeDDNR9pKozeVbEy2k3nlbGd90XqG8IbSdzFY8H8WCJ
t6d9w3NUjrRnVOH7zAi3UebOhJnWpY8jq1wDCWxJFJ34ACckdk+9LjVbbtuWTYVZDs9uhDcBNzNo
aMhWswu8+yk+2csQIsFf6n3EyKSXRvhMQYalGfq0MhWLp/bcqZhU3K5tvsPo1zFAMpwNVyqheYpF
Pd+wZbRLHhuHAa8fRAoe5+KuJm9Nkl01JdYdyQ1bknZxscNO4Scdw/SvorsYG87i3Pa98pgYqUA8
xvvU1q0ulGaLuaNfbskKvSjDlKxXVLa6waVYuifzLtYcdk3FnEEbA08sToW5L5XrOzDBJr4ghzjK
SkthWY/B76398uL/T12suMAz3/6w9wATbH/gsnBhMcPEuLNuNgmMY8AKuxXR3VUoE+A2HNYkiYVi
oEgAEe3cKRcnoBwP+9iUruPe2svBKERQ3jgLKLnNaVjizzOuttJX8T7ciNitGE8U2KvTg/hWbvMo
rlcOil/wMoovtKyrgrsjcBYdLoIjsmC7lzRukme3EPnER+pQ9roioxLLjcdRFMQa9p/MADGv7Nzv
SzqQ7PU4rR/8TCBxMXMim3sA9le3+jTDvlAwp/xadkJTcqEId6y7CzZ2MNbYKsw5RB1zFxsj5ndQ
qW2l2ZKtroyQVlneGqHK9XHtyQe188APETBexri/8a8G/6Q+5A1Z5/Z1vOQfjTvhygFVwEWVuet/
tgfZfuIk7Xxo3kWT4ph4vJlAHvB6kQFXeXJyrw1remjj4A9YY5o0IcFXnPG9IR/p4ZcMB95Lkw38
tsF7FYkc3aVIb7E5iF4fyn0DqFQo4h1ajEqXc8ramKU1wz1iJ0fqos7D5LHHooKRkoM/olUbTu4/
6U5wpN6QtL4NqmXg4BzB2MqL+uXn1YrKTJp/9wUPw2gEmOhyIesV7j8zJ9UZBgMeyxp9gMi+Sj5Y
n3XWDOHYOL42Un8YvvQDopTc7WETJzUDw854oUCX6nymSp/ntFQAZgdDKqS+leuW3Ixrec4lcZrg
wpUU7G3f0vTYpYJ8aqWx2h4z2vYrYtYdoLCVvAoaHLmmiryG3sC5pzEgZB39+CiI5GkTXYUnss2D
KN6JK8pmCmS1xkcOqYnnjnQxR9wF28blavIfhM/xvI0bnepHH7yExktCspxfMOLlRg1LvEHBWMeW
y6Z/y3TsmcPweOKbLHL4FP1wX/fjxshhcPw7GizcNmy0We8R1JppoceB5bQ0T+HOkVQbtvq9nBdQ
fb0va5NlJ7q90Opbl1xmeCS3iSdyCEeyezEmrWKDFlfEiDTZ3YrDOwAcW0tvqRDF6BeHZiJc/Mmi
Xe/CH7fcUUru+sXruFAOrSLWpNd6FgwtgKGzsjy6BYPNqIcyW5wFnYxyEl7EvGnkByHk0YWwNI/8
7m9wV2cPOCwlTGWVlZopb8YnrKaVToKp6Zr8eM1tUKdp0kXPKpsHbymV/QgzC9dNiq7OVBMl8UV2
W2ipNfkIAKfc5NcmhYIjv5Na7S4/JZdcd5wSQmUbLQR5aF3YfbwBTeh46rexbR/Hwg1Z9uYlFfob
KDWKfjw46EXjKOWbqRQupNs1MPmJNfmP6j5k2lCfHxRFmGJekOAZ/rx3z9BL27jWXO9iMz4gpJO5
VzGnn/CsAOy1cG2UHevM3mkyhp1eu/41INk+qSr2kLxL/D2oeAxa6aw6vFDnA5cXvREJtGAk9IDC
VMTYCq3+zWSNiE8Pi0mJhd0R/BzGl7jitgTPcs/FGCN+NNasCNetAML31FqaKXIa+8UHF2cPYMCe
xP7lNZmYaXVRMU6RcJrHSvhN1dL+opC5effsTfq+Szg+q+5CnQHJlkVuHFEYAu1L2f+0JUY/rnyL
D+CbyLBJ8nLHLc/nyE4AkGpaL8P+7a+r8SoIDLw1i3M1tn4xJQ/0r10yGV6DrblUectHcEIq0Nb2
wDr3zINO5ax3UuDDbrSXJ6DgU0cygJRUdOitQ+GhJ7IWDiI56nlmfRvmtknP89lgETPQGPN+35Ow
zuii1EBY7wdj+hfpcXdDLiRRHn3lbYNh9zlBcXTlhly/r90y7zzd1tV+QCQBGrg4+XoUv/yHnhmM
rxa2265bjdXnZ2WFuH4u4EejfOjdbAvVIyaRn30739Wzv4rJyxNmK0EKcm3GkchCB2VjFANAZAaA
ErhU/3X5/OvEBCPMGPCiBfGz6DPc1QqGVTgOEoWDoWyOBQR92OkTSOWlJb8JaBy1X96diavefDR/
ad+2fZwteGBM8xo+pO59U7JWvvqzOMcMU27tFNnXhILwH0k9EbZlibzNjl9oARcjKWyv90tfvtk8
GKkFotTDbLAdumO77ADntDLp1lskFYJC+YyJReeII/xvxVzKxqtBsNi6cKOvTBbvH1uUDlfb5fo0
O0VhjzEvoqkteX7dKtiiP5yuwj0KZm+sdthjK4uzeevqRq7+2obUgnpfvVQzEKLKtoQKkAODQj5O
AXUkTD7QIG9HKPbVxvBqIQVDppiZ9TghFD2glzyRmJ2Nm+1GxJNGKrsLFe6FwQ+b+eFoPSm9fG15
e1aOoHe6tb/A3tCgwa65s3imJ9K385fWs6Zvv7ufOMr4LyTUyBH0CsMzOAyn+Q7WvocTqw73satt
pEr3pYqsRgH7fWU0bcEIewvARNYGVGMfdAeUBdIJ/wcUGv7ynmVK1ECU9SpAnYMRyYFxcwGxHQ9R
MA3BdnnJGQc+oSA5mh4/mizFlyQQ/mO7HC3k3nAhPdNsMjCkvLbjRl0nbxbC3XJQHKbDx0SAn66A
YKZbb8Xcf2DpITAKbaQaSRlOadOPIlb0tjZJu08p2j2ZG0a813+pcvUTc80ju4xQDHNX6pef/sea
7oS6AhUzx5fh7EyOcg8/uumPEZUJvZ60eltxU5Euv9jtngjjoR9s+rH0SL09OT87OGBmIY8BbQNn
6OrRRGtIUjLbScPPl3QvuJ3mU3cUKeBySSYM5qJI2z5eHUQHpncxX50r0HBgpe8oR09fvwvLtEt5
ND2bycclC8ADcjprYIfi48hCCcRs8YBZFuoa5kWMAmiHlqTxXR+/Pq9bdAZKWBBYBj6hs+XYoE6K
Tp054SiKEwXxzDyzki4EhjVbG8X+eJ8V56tv9IVElw7ij5tmCwVS28YDvvrnqAhLFcEO2o2b7ibt
J9dRr/IHch43a4DCKQu7wQK/BSUpTegx1enY8Hn50dfsWYKAyqS72pw/POHjufFsvGX1yu6Z3d71
XEMqTJQyTiSYghSAHTFhArJGqBfp2jS6zWE3JqxCRKE/+7BPQi3rdUtZlaDtqpxIFq+1Pf5hoxTk
5c/Dsc1zpEhqeg91i1QF52Ml58Se+LJXN9hrS5K/78pw10HYx9qzNsYHHHKBccQUKPylYJbMtivE
5iv5kvFxVJlw7GwAwCj8yRDfgcdRWd+3V0QHq3dAcTequsd4BiAC3bGOLY0otthzSl0yJWoHBIaY
3O7jrEZSeMMCYhVi1bjkTCy0yD2hKqrDzVhQE9FEqDitOCcRk/5VFcaLEzJdgbEYo3tqj9YF1SYB
jkZ56nzQQ6CEo+npQWlggebb7sas+IuLkzm2FZNgkIjTqshIUuZaUKO8S3x/jSEt9FMA8yAXFDFi
91bcoGN9joXPxttHRETNqEw69ZRXJX4T6lfPNHfVrZXntyQcqvThaCQnAMcny8oDockM0OA77Lcw
WM1+Nq7x3lf85hvaTuyksgOo1WbPRs63Wv1OIvR2d+rzIPBe6dhgrkwZLiymEaOQtp4fd3mMb5d1
Ra0pklBIR2lENYrLMPF4mfULoB90sfUSQCb4/SGxr2+vMdSl8DPcrQZHpWU+kjogZwKzpXrSRAr0
L6Q4OdgqAgR+OykGK2OTqHsevxgNguKNDQJd7o5N8NS/jTa2JHTpNdyCOX+UGiHPK0fxA9mkOax/
aovv8q3bDmZB8HmvRg+u4w/bjQ2gtaL6VatUoOQeEJEI1vxLeBIpj0Cwrg1Ln/raNn9TCZFdtPyt
123IjWz9Nhi2Xh90jhCewjsbn+JAHdEGZEsVSnEFsMp1ci3XPin66UgIGwBIYTLTv8kza5lfJJfm
32/Mw4YmGHIqTaQcnkd4ZxmrhwWai3xnB/lRUi3ux6lKI3P3fje9crMyIgoxbsiZ8RHkofCDWNEo
3z+pbvzrARMz2GkQFhbF+DHkOz4a23/d4Ych+OL+UNyx14IecCpKLdPXa445bzY0fYV60gi0Zzde
00CGISASB682uF5hA56n1CPfFnUaZssI41be6bhc7OnzYIN9E/McD9IF7G2yUxHIuOksw/4KeD2q
TTVWwQiwLlv6aJ63TfL1sCJ1z9Fp62e6NUwPtF8lYadJ1ROUP2HebGf6v4ePb5crB/E/aAIB5bHE
2gmLuCJBLpEkDF0OKhYSsVRzLiy8NkHYyi0xA2ihkDwB/oJ0S7F03jTTGMthF4v34frn8qaKbLqJ
hqVlqaEUQi4SjRF5jM7mbhs03WjhJu/tDiwRCFImKfjgnFamHE/PW6h/na3zHH6s3kEjfbB2oNJZ
GIbjbTsLeDiKpgqnLj2xiJw4R08Qkn5AaO1W9710ix7KQW1wfj1kthqBqZ0AL2Rawhn68fUwId3D
n03jBxBqMwVDkWd9asAxVbpO3N+8y/Ai3TMBOxJhAS9v1JN6T46fbigRcrYMgVfYl6Oroa8qrMtF
kCSHApaSrjyBN6HoZx90v9MCjf+kWb+8l4GwkbMKpuTw6ErYpcdZ1QZGR5ULwN3IGJd7GsBpx+61
BQP8ab1FfSmUJlD4p3XoycpAom8xrdlBeIpy4Qqscxrhj5dbhE807x+sjZ37qn6zhmpL4+IKbMWB
4O9FJ+UfqatdsJwzbOdmZ50E0xiWMHizDLAzAglVablm8ToUBUNztOF+GN+4+JDS/Z8T89eQpsiP
6n/qHD3qa7kXZp6r15IYGe3eeVtGQ1OPT85XxLy1GWajsUpcLNh3C17sFA7Fexl4UqsorVqqaBFP
QBGS/R38V2G7Gdv4u2k2sjRkuXCearQefDkkOBLEd5d/T9PpDNd23nrO4+fCLYig/Q5LPqnW1FM5
XEJ8HhaZdkPzEgxyJkVS5MO0rv55h0Ehl5HwSOvIb33QPzjdoeBpylva4era6DKLd9R0y0ilO/D0
H3Apgzeggt1d9tg5REYzi46xQWov0o83rlSkjOJrdPSb9JtfAhLCePd38CGT7Lfym4La0M31iANX
hj7IHXDnDjLXNrla7EfvoZ+Y/fbMXGj/RksXDZaTnW7HBqzoe/NRUkCAjKmVGkkTJUSpMlckzyxT
Coc470Ix3e2BfVrxD6XbK9YTxirySNBGZ7hsroOoOCY7pIr0FIBHFEiwdriulzpBya4/zvhGcIVc
Db4LeaJ72VEINXBOTs0X+xxQ/0DeRjt8gtpE1MidM7lJ0kFUEbn04Wj6y8xdJ9im6UNtm7j50z4T
oqqrjYNN6b3nNt8lnRhCjhmIwzFbb4icLjBkMYQLVLiTY0uKlWCl8R02s2K2AyKHZXsw+ZExt+30
jmBJ0Ruy+95fkwcc9G6zVvtvSEvPG55MtzpcBav0OmyF6BSEHc4hXIsvTE443TIHDN4YTXVY/0XQ
zhTGkAa92XDxP96id5hGJRT3fIRzGHNZRotjoAIRVMfS2S8EOUPxoMY6UQB+tq+5isuYa6a8Uha7
+0ZGBT0BTP9lRms+ZXO0Zui/jUnTGZESAyHnWY5Ut734W2gkmlSRmggH94PPTy5EiLMy9xdN6Av8
BL+iBMvXt76IwLtI51j1KXJ7HjKSImwExCSmXXqMIzGoqEQOvG1m9arF6ylwDqZ7PzQuDxHoMDM3
EXLn/ICv03o2B+N4gY1ZUL9VpInickfZ1dwge9xgtD9A3s3ktXQsVFJkGAXL2qQ9c54S8jm3TP1/
GVrGbKoVNDAHPK3P0S/+tHGYRtvkvl/82Q6qrzGqmVKgcfWAm//auMyuq52/YwrMwEYCMO3CdZgj
t1HS1r2pAfzJ9VhDZVIq+f7InFljQ4K7hAeP8d/yaHGd8I/4cnL/PIVvRMiqGBhP5g1h6WgfJdiW
cjH83cy165JsYKl3NIZW2iCkWfmGenWEtZgurLvCaEX60fT4Erco1ZwT8/3P29JCHsamVGqAXsxy
9T0tfWvVRsw1yyRfpsKzJazlXTuuyjLcTLCd2+Jmje16uihCP2WFW7m8+BRls4mmCzJPQwZ3Rj4d
IojpepGGbrbHETXih+WmUyIcqMgJYINmlGkIL1TONM/SgGfYb91CO1WdYqHxE354iuJeErKnQdUg
EHD3jt7cuTPQ3JxrlZAO6ftjf+ksVEzsvdhr8F0P776dKcdxFFRuPe0mEtka+pPfm6VcqVW3XHgT
ccDbD/9yiBHWoF6AXqGMV89yjLcw90miJ19qq92DTHb5hErxMNQwPnfsIPfNWR9fJzz49FWh5Cgy
pMsSl0mTUfrVx9fTAqkpuB8ESkeq9Xv7fiZ97pUTYXeH0QXivJF9zQGdv1jlKUAs3Btg/JGmQgrS
Gu2v/BxeglliqwIDJiUtOFrBz4WAdqPdKJV/q83Z9KHLHH9zCIUR4HtIAVnjOhYbYmNbGGWHiE61
clPeIqUzcSQF3fnZJFJikNig/s0uXCConIy7Sw29GN70UDTVXzEPDsv/fQJCBwYfLp3kB3nvZGz/
WUPYDvsDSVRu9aylJVvAkJa+ZdtvXfbHuJWS0r0cclbcM3JUY9jI533fPa5U4oj7YwbElCC1zy2A
mORnBwjhzkemB/haHnmrHFJ6pLMC905iCK+3Hcb31CiOvDfFnemB4x3/8Cv/d8ZFBqJkIfB7YEg5
04A0gkJQkfp80dAiogk8ZMrQNR6JouIdDv1avQphJ/WkrfngYWCnf6aOZ7UirdRPY1BtZxJpfj68
HZRTfahfqg5jjfZXUnK7/lmubDpY9itKw23658qfyuqGxTBtcDjyuCBx5mlTEqz46lMywybwy11A
vJcAKtkGbrrrpSo4W+HSHPrvs+Q+TqjjwIYiir6OFU5r4qVw6pLDM9AqoWgLsAbubWqYZ22w8+4Y
FvA3xdS0p9U8+EGWvjVZ9Q8BajGIKcTHDZiUSJ/BCurAlk8D0OVbt5kE307mUxM39Siv+80Fc3ED
hz4Lv2dgUmB1p629KQbCzFxpFbkw+8sjP/B4orVWP268VzRvVtIz7LuE5IeHB7Qk/0kqCK2zQY2G
Y7B1GVntg83LzivYm68Ejsl/0ToJs5/e+1ievOM2dL7xGSRRAqFrThLA0oiGKUMjL6/tCSz8do5y
Fz+4ptUcQyW6J0Y+yqADFSBB1xDBIekncuwTUT8vyHEMqSJZQ7abyyVWxPzc+vDQi4oBx4bOXHrJ
7b9d7dEgEZmdf/OpitNc7FeNsP6v+kGYL51CWbJhMN/5JvQvMgnjJ7VegSpiv7Y945rQP4fuEiey
9cW8Vh7GZBbe6jSw5KYP8vDTLBvqDiYa4BP35wnEU6uMkW8v7eVY5HJtijLCNAhIuRUzxSU09BFy
C7NHI3JcLBK5BpOd3cBS0ZVmvO2veZcfyndfopiXrpvR0A96pIamOlkdQJxE3+eJW+Pw01N9AxGF
41w40ISJVOC80Lhg7uOQ008I88N1HpEavvekRIAbe3RZPXx3xgwslPXQV5Ef2vVrHqeIBz5T/CMt
zCAlWkuR9AJgoqe39VtKp1nfMvVBCLQWAK6TWJf1Eclsma5+mS76uofEjKUzwd15YQJjXjPvKThs
tyYEghLxsAiHfnBsum62qlFU+LfxcRtheFv+3plSdmJRUCxDXTX5WveuC/TsAyxbGhG3O6CNDs0k
ipqjT5Vbn7Bp7AFW02ni3gnnnyXPUYYZ7T4Ke0wFEfnet3cgnhinFuEfNTVnoS05bxMKFSlwAjCI
970oUfshdYTGhj2cJnHHfn6G5VZlvBW7ABkfA3r4aJ1Q+wrg3p3dlMtBZXW56Z+3HddeqfoUJDOA
5ldu8ezXeGQiTcpiBd3xbDKrgFQ63KKuWhmyq262Hg03p61DtMyBLYTD4n6bcdJbMZUlOh/GsORS
9UXLEghN0RdsBDh+ZHnI5VW1OuJXRPgE2hjai8XIKqs+BqpCtagcEjceguFqmdAH8RjUz9YNE43P
uF/KCpD+k55lAYDOKcepAApbpZy4L1IsWJV0M3v0KJZVyjSCdxSNeLEiPJJMaq9JuWI9+1ymAkAU
o2WEKGMpSs+K4ZbFV58EBt6gaqGZAmRRLVrByGApHlU5idSPwphYyzGRSE4gS381/eomM/XFZbz8
mIBj2semWFzK+84ph8fTcB2nZ5UbbKm38tms4t0l3a22JTn06K4QnqvrptL8tY/SY37wjx87T16k
+KyYe+NSSe3fQAyYuNszmZeE4hw8qUTJz2U6+2wq7TFEMjGNWpkDDj/Wv484NKJjDuWHsv0Rm8cu
2a5ft6v4m5YZPtTUXk17wVRDx+sUBZvsoGCjR2ak4fDnfxfycTlKMcl83eRXzvg66ihD7izCcbsP
PFo+OF2B4sNV5T7IF1EjoPK57va3b0ujf90HcubuZhnRrTlswYqEe3MfsYIUilgJBGK8m7d48VlC
0q2iWTmeKyXHWWc4uw+nP6VlbzlATTmbiut4xtNqGMEcYtoA04K8m8BjZjMkSKc3UjKCeFJwkgbL
fMrGQ2SPSu0jrBmYhn1ZqtjiLUSrQPvI+AYzUN/MON6c95AG+EUTLPtMfTrC7aPnYJK61ierHdX9
Li3SVyGnuPSynfGpJaqew5afSYdeW0zcFZNiY713ZlHJw41SrSSVJ7Jq45gqHahTd2t0dh8ST3pq
PML8ASz7hPVSsgIoxg4gUuLHyA443GhMW8JncXg7n7rDFeK+4lPDLFWtIcMRzMF8vX/PIVbOmXdh
GmTeUX+3V9J9stnnYB3sBaK/EreuEL2o/kqPX3CLiYmjqlAmdEeprCeSst61aG7jHeSDDwqGpKCo
kFFHfpVMxi1KC7Ii6sKA3WZCpOzwkqa3Vvtj/ef1On+n2XoyrMUu0W8uhtp3fG16xMGpUIMDMrRJ
h1i/i+fZeFAF/nlOzcQxbXKKrqpObkqxwAgphLeLucF3yBM0JUE1H7KTwrGzntkcK9lZm1UiSIpv
SFr+F2cGJkMaSrw0DwppFapETAltdfKi8cmc6gFIxwSv2b53fhe92MG5LOs+uuGqLtWUf+jDeGum
1VMymmwue2lbrGtsm2ItzEEJPmFzeZsFX+S7Ho/zbxFY9kGtzm7w6AbvH8RJtoqngIO5h82gQjrO
aaozVTzY8cUKIb0XmABO3a350G8QB3PbJ4bASahszpMwhfE8Mmzr9boZCyufBm4puw/G8u/qDpRO
yXp4lMYVQ18r7kbD9LZpElKDWf078s8y5QxTSBlOTCnfvX1sLYliJXoJJIdvXgD/9lMf4C58vlOb
HcxTpt5Uz5XN1L6VIkQkzJpATe2BzFWSU2nXQQZzPzrEH3Jhckd6nPc272tTanHnG76qUCapsC3L
zJ+n+5PcxT1ExrlGxjenjflMSvWZCMHjq6EKYFvFWYYWSfamUn4iMhliyEK7BArEOceVMZliaPS0
WDRD+EeXti0JWh9255xZSiMGgkWq0BTmDD63A3E4T1mnG/ay+qIyqh7hR3KLm7sOekRtKOjsWSah
bl7eVUeMpzS0ixFlr2B1RPTKl5KjQd1qkEGeOCL+NrlmypbxVLVXSfsA61emGP6Ljc4lV6Cfefr9
aGw5N5P72BnFmEt1gBcNJTlzdECbHWY25IuAdH6H/2CtuiuLaI9D/VOL3x9Hb2yZX8qgtuAnpJ81
mA9HDkZSDWzS7BWKcMc7UYgyU9t/fmxvXLdfVtIBSqKV3NM25DzLzI2UaRd3nz/6ssOKgVIF8FXk
qVIFZK0IguREHVTz5MsRLx4VeOLhPB+5gZvSeWLYI4pp/R/u8dPvhbylKUv6vxvROvmEmrIm7tey
2FBe7ZwzvI7rCFylA83RbALca/9x4LxYXBFE0XgIpN+hAya4OXIO4LprsbW0oVvoHzi+hy2LEySG
rGoVi/NsZCm+dxxir4XQZxcs4LrJoempjhEuhg5H+G4HwybBiWQZVsTqvfXYtuTbXdMBRNZbzQ/T
RYCuEpHyZ69VLKdOw1hxgt0PtS7x94swHH7sjf7yfDCtF5NR9CJi4+rvbAalwqShs+9z1EBQOCSc
ZIfBH3jb4UrC8+hRBLusZ2nw9CarJ0l5reWTKkgYdazwDlweaDNTcYv3Pb3sUubu5ht6ZMHw/O4d
dNXKL3ShkOJX26t1yGHqUiirJH16ZMMnbn4MM9R4YH2XozgHbErB9mIPyCwGzV8Pl9+NttNLRNlA
MDFHMpzVAE3EZh77ZwFQckuUakZqsIRfzL/uOIVyseKadvlM6o2cYLPvF8zcWjrVoRVGqnM6v3eT
DufeIfy5gv1Q8q78P4Ev6W9L5RgMd1idRkZi9fTbpvsPpyuU7+Kr6wr6tAuhN+t9rNXCwpH6qJIt
CAcsDQn5fPSqmcivQieyOsWP0+k1aGWbzsrWXlxrVC7TGO4Y5h0kA5DLuT48kjp3+MRyaLPuDUty
yfEmTS4AOePAG5J8zCn29GvqzbKJzmlv0Xa0IkNeRl+3tuO9Uuu17Z/qTUutVtH2wCkXremPbmaJ
olJSvbuAg3o2Uu3FEMD+Hf1trOnKVbVjWmpO7WSLFeQE9nYvUxPZgRjbR0Hkb+3TlPXoLBeRLbSs
824FB4UMZpX4DTl/o3aZceeLp2FUj6gt7YG2TkzsK9VcRqJWJNuw9g8sc8zcXWxqZUlhUIhUfM6k
M0yR7h8e9BORBtXgFOHV0L3bpO1OFs74Rm9hO2noh55MyQ/AS6bk9HnTUM2Bc2fN5ws/yLzGb50x
WyVg7IlbJZADVc3vQiv4/jpKGF3Sftc3r5Y9qXK8t4XLGPXmiaJURDsvfIyR8iMrNNJCp9YO2A7t
XbUhkjDLaCK4YrPOciHah3OWGdN4nxZqEYLyVPZcfvVwgbjq3rE8nmjtUx2/IQ93jVQ0EiOi7U/Y
SBs1A+hUNiTSVc1AFQs7aSTCUF0e3BUQvWfgFljeCriZkcemBsrvP503KMO1S9EQ+Pg8f8/vJxXM
A4HBw5etvquo92jVWz9rz3F3P7jNh6I+10QRCFV5PJRaYpmsPp9YS3GBPi5GkHO142q7LoAm2nrj
cFJPrlLc8PCwsHghvf77TYrvPtdvbhLE2qfH5PmvZzt4AJ3mx5CXPkNkTEnBb7xZazrt8Is0zb2t
TAAfDfn3N8UvbXgR/clHjv4CH0eJUPBkePAsZzPpVCIRPDbJtGPimsHcdOBRKhymq8oRgzxgccZK
1mdyyOxJR6qrhbz9mfPABT5PvJoLn6HFCpihKf/ZMd+8ZzdyV97F3uJ2D81lF5eC5cz/h/PLdEo2
QjO/12SIDKj8TBtHQqmTsVRXSXPwlyBp+j2vz1n/3k2JyjQWZtCvCCxd78p7wsOyoR9e1ayQ5cOt
+REjGduqq21WfwwBWLMuXg8MA4XB/d8eKCGCE9Bat5lbqZWt9B47z8X0jKxRNJr95cVmf1Mx0PAY
Dp1oUXuaJNC0YEMeHBuZAYoDWsfNgw40oxMHTorWYYja+2euVgCEdMJpJGBwbVy6USf+QMEgIIve
eb/t0WBLI/i4bmntuN7n2QYaB8husfAGd72XLsNg4NIgJ7FtjdMQL4K0lxx1YWtGKFkFpCjgwt2d
/32kv79DkHiW5f2Wv4/b0x35b0WtWu/FDOAkAMe78/XeTI7uRrVMqWrQO9t2yKe5nUW+vtspHROr
CBpACwIEZXMsMXrNY9c7S1kpMVbD8tDE39wCAQPhDnz+/7ktnaFeJ9bbP4+ex8ruVsAf+AYeu5O/
hQqDf50dpVlJhh5YPKfuZ7dwwZFoxQ0VNQu3FAyGiTJH5Wux1jTE1ELhSR2y6vVAKsObw8Ho12is
EhcY3bh+fuoOAjeYOg4ntzLWgqxCEMVrtFEG1oQMx10gxQjRsPC64EO9xLALE1FN5mdJ8NSb0Tes
pydDP7uw71QUgmnap9OZ9FEpLcYN1aU726EcDbAduuss25JeSnenQdPanpWH2xlFcx5GRTh9OYyE
vnpAupB6HYWzLWEJGb7GB8wkqWm4HgyVR/LRmHcFOj15B/bgT9yj87qnwpRnn5zU1kDGJp+irG6t
BkiEb+D0BPW6j1BK6mslNnSExLv3qI8LrYD7MHQTc+0dkj1fc7Py/rixE1vk5BMeB7Ii5lwoVt34
phHZt+1PbHvfXX9ATKvEdAukqdbvLK6CXZ35roKiVWpUD9paUzS9dgGL8tMRBzt4Saft0/TIMCfb
nt2/maUZMXk3oAlXTRz+dYtkblkJyNZiuf0JV2WYjThkSeXxCQ3RQmuTCmGvsoRCy4vMyddYkwa2
IvYiLOn19Own73qiAQRtmERe53kQZ/u7ZyVwqeb+5lz36jeQs6iyl1Va95daBPqD4/VbRZGKrJi6
tizQPzJQsR1wIKDlgk64/WyciW4a+9HGWFy3rWXrC7NwFiuqkXPAxHyezcFPJ03DYDDNvp7ZgOpY
zDcohWdupFZ0bd54Lehb30tivUcfmPFC79NGr9ZvZHHaisYc7afeIZjeKQd8Kg+a5w40hSHuhiJc
5sdo+pbdxEznvfGvWn+P3qRq3K21HjF6DuRgQP2MDNlMPMzGZto83M0YeBuiCDBgoEEUKZqQ5jTW
rRB308W7NZYxGPFBYRgp+7kPxk2/ITLO1DB1N1v9AiIu2FNslisuRYJLSdoI9aGecXNsSO2+lwqh
XI5mS0m+OonzSzyQXc+iCKQ58l20Rc02c/BzRkcWKoche4JxeLsBMisigpWmhYWBD86kd6otUvJN
poYIs6WdGrw4noggDORBAmTt8pS9ycgr9A0HYuelwKgjj+jE9Wa2r90Ir3SNxIl85iMWzkQGkMrs
ek3rL03USKemSGh+mmBmpoLex7j6vvf/tX1y7ANdaQ30LOdpV3+qnsO5sJb2Q0Sg51AJo4fyCulV
7abUxymBLMoqTTIiOUVSoS1aE4qDfJR3biHQ6G//6ynaZ965b7+kJ44EvSvLiW1kSlhip5SfmFSm
+fgAsK9krvNprgo9z4nqriyEpsJeHA57T/mDt1xMmxTSAe/earVuFtce3xX4TFrtoy9bUDL+87Om
zka2kCt9JQJY6OPGEzn3MT71v1FxqxfHOiqdiF28aBDDaeTwB7mXGPnZ167V8Z8X8wMSIXektO27
xqJJ/TyYtd5CC9EYbHr1iytpSa49yWxAl9Wkobq6jP3Gztc4moGJfK4L+auvE4EeDvFCDD6oIb7q
b6VS3gMwmNLcbL/jLuQ80hE0fkAv0joBBi0Lfuzit8vijAz3HwiM9t/LDi2AaAUOGKF/ZLF/ndjo
+fl2LNmAnbGzFnlSphufwrOSC0h8YrY1tYU9QIabmTtSbLdfa/bk476N8Rj8e8yzRZciVu9LXVUv
kudvsO1qZ0KsBN7tEJNZkwXbKWM7NNLdudFIatO4dhXwBYK/8pbfC0fVt70il92lD+zInnkNkUNl
PJCKgZGRTAMRgiBWGkcT0ByEUX4ttMbB8CQmo8Lux7CHiXju8SMOzpZ6avRGTV3elb+gnbIbaGpn
5NMFPS6uC30jDDKvEM9IWk1hoIyYsf0novkc21SHfmVhLVdK+dpSUSlx8dndWI3LcLQsagJ5dDtT
JEu488snajK+u4FeJHgPgeXvF94u03sGEmu4sPJa34LPlsecW4d0lObhEDYw+qpqTv5WZIYFJFvu
TLQG3c52ernSTUWA90mFfQeXLOfHRurQYym///G69MUcF581S++MMn5zuhVv6qQCF5/DjBO64dJ9
T0+HbaF3sU6F3hM4e+xl9xDSO2zw0FGcX7GHVyMVli6LhMVcpmDASaz221rW8SBYxwJGagm9y9Wr
uZEp9etS2AJp5yQkv7hXNkeb2Wdngb5WhHz/mFDukwUF8q5UnJ5U5LujVeREviWjytfNwyVrmGgj
VhNuEPgAuktKblmSCsNUcK6tOX+XBT+M0soY1XhjzZWf6Y24Ohzf/O3bkM5w7W3bxgj2I2c68sbB
PjVW03QHXqT5QVFF/j7Gp+DN+TxW2XlqbiHAoIhNldKz0c0tV6pw57od32f6RzPikKyMO8JMYHKB
RQkwFynqohYcEZd+kgZqwYbL1tNvWk4dwfgveCn8KUQvEr6CSVGKbYAHFEL7XdbHOICfAsx1nAB6
UdBM5IPbgVWV/S5haWcmbkU46EBYLXvMfArZ4lynL7IJjNPrv49qhF39MRYRJSfHAk3IL27x1vv1
KhBrBJg/R92hx84kuqkVBMn6b5tLWRxzKE/6WFW/rDAnecf3Ti6PKTLQB8XBo/ywTq1riUgQruQK
SfXQwF7vPPU7YHcOYsJ+6wBZkqxz5Onrf1GF4SJefMcJYO565QKLO6QADFD975TytUiuwRDV/g2z
2fVUp9ebX9JrzU75Mt4ub3rfhr3cz3erFp27R7zwn9EbipUE4Qi1kJveqJTw2jtYGH+aLQZS6sdQ
H6cgB6Y5cQjIXg1QHD77co0zxzS4//P4sp5wel+4uwOhqo7/E0uzaZoD9fuQ6nSSew2bhFDMuvSI
TLP+ybnovNKCAcM9YIYyZCWPgqURVlY361mTuoNyV3H0LDrtrOsnFbCSePWacdcQGIkyaDfDojI1
fTkQVrfR02m5y3F8IjCjlB5S+pUHQ/eQuGegl07Drq9DLlK1C4mMIMHCKOcEmZkh2DFTuJg8TOTm
iCY/JIGfGEH/xcBupzPyHQWyPPJ7u3BkUMO+40sTz/JkXhYTFNcdpcq1krcNu3SAo3AXigMv0I31
zB8ObiEND+VNQhnSP+xFcCSdu5fiifvWx2vPGKbdOpncg3jq3kQ0XiaKj/YB7bKFXbKjIcNLJkWA
68sREOZejS3SbDy6qBqZGcC484BlsIyNIMRqiPH/LAGaizRD8pM63SbUoiOkBFf46rWW/LreAd36
SwIqaEtiqo9GMdbHhV6Xhl32+PqQubRSHcOAPisbqw2TNqHJWRnsz8yCrElNPZsqRhLs4M9NUcOz
IqtpqEjlJx6VP+5bdrWjWw0xR7UkiAy35EDgzyNKo3dfSgb7mXLeyZfadtQyOXepYmHa1qOpS6W5
xYOy+Linz6wGStT1Lcj+DofiNCYZb220B/lmodGG6wHCyraRtgCtbTRvwzlbMjHSS5eujtH/ibno
C8J5V7g1ZpjWx9H+NQzd7PKBRZRpj60x1bV2Lz0d4539ILGcAb/NmTjr5ACpsK3MD8rhSle3yAJt
ipvQteQEvhz5q3BhsXc20G9KYUsN/O6ly9uyub8j4QaTkgdRAmbYPYZpQlTnQ/Cz21G/c8T2Jxu5
1eA4PX643GmgD8mRl8BgQVo6vOtoXmLblRzDleVZOefMRV1Put3tE6bB9z6gWNxH1d2uM0vXV1DX
Y94iKvqJshFrCpaPGWyiQr/7NAmdJ0vgeu8vzlxKZ0+A3HDbQzwMzsT3erIXAmQtwInl+r5ZDLMm
Du3W6GI4sNlSvC+LO3D0ymdRxZPk3ZRaMO1FJpQ6otbkHyJuMjq3Uv2/s4vvgK54F+TBzcRpvY2l
vsC2KVLZ/rzNbhT9AuK98MKNuig0uM2/XBuHbC267uO01fqQYSln03SZ5Odazsetcatm9uU91GSH
kQdrTwLsIvQ0wPVWJE91QEL8lQqHRIVjIDoZbHiJeXW3MEbdRffttMj586HNC5cuIXizqVvvSplx
oy86Rr095U7GF2IjCVMEXmlKJkmj5sSkFa371FDMLDpC0uN1nH4J3DMrrZruo7fVNVwn4hdYC8MD
/iI/kJ4uulvWQBvjLH9cDIozrU0xaPsfJkpNUU5RnUx7jvLlitkYYD4e00xolEBMAMi1FqwZRTrM
AWGSmrVu1bvQSpSHiOVkNxHnIm1g0ecVeJsb83rhIhzrFpHennXX+QJ3rUoLQ1SGpIJYo2M5GvIn
wUjLeJmfln+FhcZqzeHF52w0UhMan5WJyDAyO3f+/jIfZM9YTcH/pXxekw7apC0f9PZFAn18e9d0
LRxWkbAnzx50MP2EKAE6y3WHPw850WcIpcxtaVBZIBfMQTJeDpFa0ssY2CNXpwRoQA+LCFUw+T4G
3A8I+NgqyMQXTxHRip5dt8x2cSknl2uR/fAB6+ZIA3onHqwbPOYZo2TblWvmfZT+Ukd0XETHrd/5
kbv67Q31C/E9F6SpsaZ8Fe0iyl+l1YjBQQjeGFHwmIy9Fm+3Ew7IIOcaPpPwbPNybhh6a7/kE7T/
7ab6U1Oc0+LcSwfB2onL0TsVWE+mvHzBCDzKfaoWaSpuwWB3Abr6Ss5mYxxwkd/pW3fsJR0Ym8v/
K5pWt2vReU6fnESqW7e0vDiBDIJmyeEjK/rMZmkFt8SusyZCHwQsY3srkcxWFJrsrkrmyM7UCt/6
Frdcxq4Q/smUO5G895RVUVqT/R6DGyRgflTXHb8IvEkxgbbo9EsDw7FPeq6NRBHMpl0Zz5WJsK5y
LStZNiWP+m1IZo/Xufnh2F8khEPX6EXDKrQB1mcIU6AjR+EZ3ayWtvOYf7RJVtjrSo34EPPoIVx4
KMx+Y6qiOG/HbLkMHFlCSsYXeMKJbzmh5PQo5cT0FT39oGt1gFlb2Bwzjf1T+1lr5+U0Xb+sZctS
JfyUL3VdyOciJXse9CdErDVVreU3iZMi/irk/Za1X0sz/L56ELKfCeBGGyOL3eZK1jqa7IQ+Pau2
tWrtc9Fl1NFV74uzmop1zI+Qx5krFEW/Wf2BahMEPqBzMo3qVDtbQ580LnJY+rTBpXb/A4gkK0Vj
wpUjtvhPhEno9bOrzMqOUXrOnoDMrIuyWN1EOY73X/n+GmrgCq0p0x7bjxYbez6lDPHT4cgoRKuu
9M1KXoul4q4osLQtcbTJOYMgn+Uygf6y/+6AO1v83k4gkaFLt67x88prP5ZQU8yvuJhv48lAKh9h
rkqc9f04dMgSO8c3LLWiwHPfdLhdQbDYFmckhPi8kEznRmPLc/GNh6Va/Zz99OrGmOXZ+09kVBkp
zwu3YGnOoEym6xSluyTBOt2e550g3tCRAqgqcbJchQq4+f62S9OabRwmDmjHz66M3B2uGtlYalWA
HZ4yKubsYrtDByda+LL9dnbxmeLpfHkCEZNbF5U+XL5LSQCqmQ/S8kxTMrvWILamuQFrhSKxj4cA
7hCLgoBpze1le+Wz4lY5hBI1sUFQNCHrfqRzEZwxb+48KtjdyuTjDnoQgFtZjq7PboQeQHUSHCqn
4yFTUoBa2kDXPddIKrVRUZaj7s48NdW86Wci9+MZUjhMO66zLpfBQAD3USQ8DdF6CCHlK6/Sntoj
q1nVeT7rHNaHX60qrHwFnXIjT5FOxP4V4TsPWHgd2Y5USL7sCBxfc6pgohN1L1OX75NbZsl7ZEns
VY9PU3jCNGoFfzzCn8iMjiTMk76MWanPxDcO7Q4i6GU7AA0HmvC6DSGPF8Sx8AM+D68opeBBOR0w
FXYX4VtEYLLd5tK3HINO7UqQX7rZm0jmwTyRzjJlMKxCxLL/KjD7AQAiAMYB3vDNtXEL04EtGySO
52P1clRgRkuSZ2jqL/or8VPNhEuQ00ctHU/DgDEU4GjMBg9SYe2fJwLQorTjccgyd0NrvwGSo4e7
nD57wzplMw5Uq0k78yNdYtJHvGnGhzQVP7GkcF0gQtuQvU6TaCjJJQiw1BY7zzs8hV/lqruvLHWU
onAL/e3x569VrLgJdPfV6H008PR6cjPuWdvDGJm5gn/FjdGh/qfzZ2WwfokEOXLfJnOjhWEEm2xL
j86fAfEEdJEm9Be5MOM/MUwV7b0UKXgF5CDVch0wXTAZqSR5Rg0shx9HhlFS1YHSlwkwoUwnB26W
Kso6LUdvzpIpP8hfRC/+pZy2zZHhacJvEuWPcgMeMZaPDjICm1sFUWOBmKvhIzn48AQ0Hv0g1BUr
DKE3jHyJiSxHEdsZ27rZt9pCKiCbl8sg2rUbm/bmwkzOl8CVuz77vdayvWphf4ADDChsfd/K+NZR
vfDiMQjjS/NSy0bYbZQwVaiq4J29PyaclKfVk3R1lVqhuP2y33suqH9QbptiTCXURlApaxr6nSmI
mjKdrNgdwuEgeTd+LC0T63vUtheh4u5BdP5iYC8aqjeuDx/XOpLHPQ/KpvM7Z1ueCRAAxzWkOqzH
wfcX8VqgRo/dVDWEz9vdPoM/BwuUdu0BV27vRvyTNcwVf0i+l8+Dlua4irkXHgIKIU4YWMxSKM+O
DwGlZqvxBPTWMgyUuazwP3M+83HGSf2E1bEUtg5/V6Xf7tTA9mF+6qLGwGaPJFgPBLFJk/YYTOYO
2ClzrX+ukDprlW8/OkECl++PXD0THZ21T1kU7NQhFWlj0MXNbPr6TnvtYvrD3C5XoGW9rtEKpvFP
JFZuywmaN0ZCWzXx0bouV0zmnXUmMVHaOZJFWT9NfMGDwpGXP/IXipna/T3btuhQfOmDFvwnZ/OP
zMpFmCVmVIhNyyWthXfEa90542NxaKoH1jEwOa7tDsfa+cqgq7jzF0zgVDpOQyfu7NJDfIa93Q7X
R0AZ7IJbkDpvhSYihiHBnpGNv9dmErTE4zgCyS7ItLnd0RJ6k5QrbZ63RPcAigMpFx/WBV7fQLZq
nI0bbzx5VmBbxhRSvhQci0LHKC8juN60I3g7R+ZCTJ3vnd7DnC9veXD1WlgyddIlicndoUxe2fBK
I5a6RrEouQHSLvsPduzbF4MM0/9i9Hb0ed39K+b7tAkvwsAwd0oazCmJEiH0kGHUmKxZ8wHGxpKu
n26xcZiOKeQwNn2T/KJKmV6Xgsz3gR4PJzP6CoLs2Cci0gKEM3rHCzPW+234yf2zFWrLXL3v5OF0
3bUScyTbF6WsMj0McHAibB6xRC+/qaRfxRjEcuekWhM4gL03NnIEdQjpyuDaiyvm2WbUxaGJQq1g
VPsdu1jsvkVL0cMT0qXhC2nUpft2R2yf7O/i0fvNVr+hnSTWNooX4HOUJu9O2Jr4FLIGqC0WD+t2
w+1v5e8r4jznIWZ65JraA9ClEbMJs52EWrXv5XVL9WEF6E+D8IlwZJDGqJcQMaKgfKlheDvOPejA
otZeJEIDdywrM5EjhcV4/9TlwshqSrjCfCosu1HZ6mJIKRvCk+FQBGQQxThUc7Ey+S0vPmCz0iUa
lc8ALKwdbZy5ebn4hZS2kD1Ew0tej67Gveldw4qQiFLkhwdIz9l/IwCux/WwWzrjYgLw9/CmvqQE
zzHEYPlJ2Z33WCESc58UvSS6pS9+1YFErRzfUYsk4K5hVyeXafjVUk8C0HGq9ukFoaCUFuE1OjZ2
jX1ep6FVjy54ohniMQXIDHutYrNZ8igBngTw4Ep+/MTPCSgz+6itGby3QPQJSWv3JvU25zFj+OjX
YHPaFYTGn3MOMi5g7OCxVH89buLRON88ulSsAzkd0QxoLVbbs9yun0Xi1s2qHsHneHNRKODqltkt
hqcQ7V6C+reY9GExvCeUD503bpPS4BXPsl9qmOsUoOceYnGxzI05fO774nV1nD71PrXgAPdZk4M1
zmAEwhaJpGLf6BY7OnnmhvjfVrhWbgwa+ydTTZt/txpkV2GTCo2ff2Fq2XvgeVtHuNJdOdeBNcs9
hHxODS35n187qzYDQTUBd0gLv1VZowCXrh7rTG9TrxDZdxDDkAVfGHSdfv4Cnhyxr3I6Qb36WyKv
dAY0ntiO2vl0DPVUoANnUBurDFrtft1F5lXWPmTOCjqwbQVr/38HPA5u6PrQMt70t7ty20p78skN
Z1U59U8fLhGeD+O4O5GzYdT37ONN+6IKG4+bo7av2Kz/W1IgMjPctRLiiXnkPAy3RwRUGkz7U6hm
YUoisniF/y3kiU3wK/3XbNUHU7zLcOiN9peI1nIuub7Xil4PzwK+2ocdbEEFkszL2rq9s9TDVztJ
HabCYkjF361cW4cv7kJyDZ2yk7ifXsILnA6pkx5t3DSP3wx8NY7sVoNFzfRK3Pf4+CJ06hEPjzmm
cxwjJR3wbSA2/x8aJgEW+KAm2mp81Rt8d7LQTzmN6XdJdTZFUR3gwS/kCy9Y4kILyH85BMZtXfWJ
HVQmPvU1qJGqoIuMLQ6wOejsKd3JXgkVW2Pd0HrBqRLHOQySbtPguNHi91zNyA1Jx/gZt8Caiexk
nNNwPG0wfh4Da791v+s8UQRzuo0znrFR/EK2WhuLoacUvJn60UYxb8uoMvgiKA9cLPy3IYkS/3rk
NRx+TbEr9QLllJqP+GS9Vr1ZwPQa//rLj6LyUmnQq/SENC7TF+thSmX4MF5R+lpX4SExIBiENzAF
7yxhs5G3Nvkn31CfprUDVkRSxFa7FPnQPmG+PcN9xKgO4vNDn0Lchut3wh57b7pmrD+ZCPrzcj6G
1sjqO2X8VSztN3BlDkfDnPGLcJczOf1wm+qZUUb+zJy1O/0at984mYxAsdAe1PqDo7YrEpCWEbOS
qU0uYjk9ZNrkzOFcxp5Ke2uzsNLsQErnArWP3V4nJtgI1DRyqYi/rcSgplWvcPOFXrW3DJwwsX8I
4Mda5EMEQExftMVpVIuZLSWj27GwETCPTdTAjVLRtQNw4Dsihw7e81Dwk4VLYnByP4nRAB2HToYZ
CAwZLHnaXE2UiXkXK8vlQUKxgPmg5KZv0od+gEZTxDEfyYvW1ttGoStZf/kCLUbeaPeCS9kA1bcF
aGB16DHIrDHzLgLrakuRZNf/1fbEJAxoUSGy4xet8yJVkzlI8eap7ZsWVMGQ6Z1YjrQdz2O+E/LG
1BmAp+elC0DwppuoPdtwOQry1JzW84l1nP/7NM6xUZBv02QjPswYSxWK7AaRrB66L8v71pMiPpoW
Ekb562YNG+rhanZA3rS+IIRr7aJKe650G2NIqZjyJAdL/VMZB6JG1IYViM+fLe7+d0r6HR20mG27
DO0Fm9SfqKFpcAPSjXNP+Axlti27gKQGBKhJQDzlGHY3q1EkPIg6R/x8utEz2+XVq9mEpezFym7Y
fiJW6WubQUFHDf/ok1lukX1NXk1vqWFyHoM4HBuKKwW2NF0QfVD8IvE9vKd8Kyub159vUXluQ/A2
6vXdtmql/rtU/Q3v7xmUSN2EikpxawzQCMD0kZTnF0s9FkKucqLf0kg9rA12HOeQ0BbpN3xz1qfv
bLI5FqEYPWnthxFK7PMpS90mNQklzdcjs+fPh9fAjR44yiAP8LLAhCpUCGEc7mezd2DStRYvf3kO
jHkmQM41X3v/8cvpN1y57wTDuGSOgs4HfnlJmFNkRsry/EaxiNS/P4FqCJcL5kw3QDUmzW51egVZ
JVC8NMBrGyJ21+lUsuVF1I8KVjEQgvTd7x7uFZFYuC4l1NHAu90Tx+3d3RaDjLzAYS1eprSCa5Gf
4SgEpf+HJBYJsK6ebSaEt/l5upFVPjlB0gp3eEyuFwgZBwlBonqBACC9aT43xN9ElpD6RcHxNcBE
Dm7qTCeKiWNDFk8ozqnfsWPxNtb+ChYgXEavkaZV2FBbFDPSRinOH+t7fF/VKQSKKVp70ZHyafug
/QmDaY696yQPWIYF7/HTCwzoGV2y0+ncoits9mVEqUFLx4yRQJwi9UJr74uMSUljEVbp5obPbPIY
cXRWs0B0O64BNUPl816O/wBYCWrMcw1FWxmyjmBLLiHGQIQ7n9adGwqf9Ds2FKfSeIu95pogQjRN
3pO6l1opBIXfxCfCO61t8nO5NRXlh/Glmb2guFG4tLzeX1ObPYdoBE/WOPsELH99mzc4IIeM6Zzx
CqqKk+ghUukfcss5wesiylUUXcuoX5bZ1ZCBlusjm7sArhtUljYJS6QlcSqNm5OOgkib64LvcgE3
5ukKZ2q57O4814mcQTMhCOFaFDG5muoj4giSdM7dVr2eLAEtPXloFaPmOGE1LW3zGXhGt2D+0taV
VwW677+fhZRkivEk86GiItg/EdNUzIh8ctBUfjVxeBwOWprT+qtmSrouyfa56TBmsBUMzKvbS8yy
Bxk8QrFrVET98bxGVzq1yKaMO9u/RD1N1H4Ipja4lkMwRnTp4m2shfnl/DtpUpSC2EzfINX25cLc
8D6016KiY4ogK/C5YU+/0I+PHJ3Tsd4/jDdNP1L1pw90QjLGAjF41xVTAPOAvvTe1KHmZ+bfDCFx
Z86lT4W4qPJrquRko33Sk2KIU4Ye4Z1OsRA8F29sNegGOqrfI2FGhDzpeR7ixOjbIi1QBgt5r6HP
oBlh7xSTZB059zxo07Bo45myXd3pBbtY3Z4wz2lP016C/2hCIA9eA1sYyKcLy0ZAZMnv4+PBRtmT
64Am0nhQhH92rCjvmYbZQxr6+sN2XErg5L975anSa71sLsvRIbtje+flj5R4mgqX4rAegVj/OG+W
nvzFCbtdm1yjyWhYRu9EPb6eWnJWo28qhNUdrGzuziJhAIw2EqWGlm+IAN5DL0Qg3NdXcDHpQ82t
m8AqhMTUeQ51g31xo1buZumhdCcMDd2Jc5WwNuiZ0SPZbpP+vZY1u/ouWTFvYmmTrkxo5crMw/8T
uCmhKz8iccA9XlwIqq8SW9hZXGyRwDokE3DAL4QkN7oZO4IxIcY1gV2dNS/RT31accV3VJOJ3WnL
3WMgJmSksB3Fp75b9VY06340dc58lX0Q+RTqWDHG0H2S2T2QyHyk0KykJxk0vLyn0DJK9aPZ40OZ
mRPDWIpCskLInWkm1gagC0HApjdUE20by3Qxs48wgtow/uwQcLcwFhJZt4b2LoUU3IuH3HZbi56s
FTBTAFfQ+PV2mV7Xwghq+kG84V56oCi11mdzHA1bLFgGkZvNrVJG3MYPN1l15PkFqNWUAtqGXhb5
UV4VlT/g8iS2TiQRW8IbFP/WuvuOvO9AB3k/Nn4ru8fUccIC+8SWDsDHICm1jmuM/1M2iCJVhCTu
PRE+vfEweXpeivpgL/1VLPi/JTgumFMrVlZyWiPhtoQ/gvLz8NVPsqDXqNxBgOQh3r+bVfv+sRhd
JevVichmemNuQdVTe+sup21qwQxgpXCyKQ4gwxPyMM1A5McxLmg8DgVnjmKweW5EDnTeasl65ajj
lcX/GAt2FtsQ7Vw7nmn+lylBVy0Fl9kqJEguUe+B0q11zCuMJOWu36hRKMBpYsDHsGOCRe9IxbGy
faszE1/M+hhZqY18dSov3mlywPKnHOxIooReMk695xu7u0q2ygM0GQ0tvkKlx79WiLi6z5edEhOd
/1IfECqyeOdIuzbwWdWE3l9NiKcJepLxXh5jyReQRoAUIvBt80wAuStN6JhAGt0eCCTqVeuY6I1C
9fXtTiRyJZ3ONx0kJ4X0q5PViaI5W292YZSNs43OiA/xf910hLkYG6CBPh8ef84cm3k50OWDFmTz
Hlnbk+OsWD2Kfjls9xIakwtb1NCUWbfRtJLwHa6b2h6vKX/lt4sRkoRjIjrRLJvIEASDafnRhN5t
01jai1HeaxZdoubLR2WIYD0gg965I1hvi4A/VvYHbPsRiUxMMcqaVeJnmf0PUfLx6B3y+BX41E8e
7PPqVLock8rqdKANKLuy7nBedzXC/oZeApMYq3G8BseNjNbtUxC0rj1c3AsNHPP8yytujt/aDYgG
I6LygTMKlvvNCRJEhxybnX9kx26FKCWh9As0wDNnLF92EarhIRAudCi4FNUCz7cysEv4M6BMyLiw
hkJnojpvhRmleH2K4ec6Z0I145lciSgUIFerqojeD1nV8j9KlbE0kMkT8ZS1B8KUcJIF67quTa4m
QIm1jMbqrppn9pby1n4rF5FXsJTzo4vYbOfzw54Cut6kzNAtc1x20Y0zC/fv9TaFA2l4saTW2YVd
up6xwypBODQ0nDDN0mPCa8/8d2nVZMrlyUHNgnkfrTtobolDNZNf/E0dXhpUIkW4D9itEFfCzZT7
dNAK4pO/TZ1VMMaNYR/pUEWj2DX9cO3DHAqWlxLT/OzzIURt5/P4RCg7lkX9bIQMOGvPC68keuNI
F9ny8U3DTPj++gDnJHYZAi+0aPmkqytnSvZN7u0yKidexrvDZ00Ap+9+kBu9+84nuASwFzyphuK2
wae4rNLq/4caYrjTR76PNeKE2fb6Ub0+H9dLR0YiDFSsiotYqZgYec0B75+sxYS71m9KG6T85c81
/oHJXf+CjJ9RNJN1l/B8hjipRbjuDqB6a5qL6TCFoszeca6vHgxk3aztKTUbyJFktgJETpOUbeKs
ZnyVmzGYd/YtSFtXoGP/FbVDodvQnla3RQ9cuwxXwYOn/ceByXS/TyjP9Z9rJpxUXf0DRdnWleyk
1CnnWNJR1x4o2/KYurmKTXSefiJTHkNpSqTTMBWMN4qPkwV/xUPplMbxZg5d1VCzTdXh1tp3BiUN
6+Ec8TvLzfO4HLqARCydyd57f0r791Tkns9uW3r59NLK8o4L02/WRVnTeQhNlHP+ujh9G15ctYf8
tCobzSqj/4NWhyIfXweVImLeYHEi86DkW5HhV6egBZWvFrRzoAaxI64w/KE2I3/lV8VzdCfM1ydW
Fhl57f+efXq86gADxZgE6k3YKPCrmme9jcz6Udh/aEwaSP/r2jcaNejAqXA+4C/BFMaT07XV+L6q
oc8+ZidlfwX+q+RHPTitbv+evbI+0T79hkZ2Eu43aSZJ1ndbcskX8v+7M1ZN+Ma1XCKSOmGZLrM7
LLzMXtBH5lhFEQTJCiYnC5ZQ8b/1YzlcFGqUA7vMu38gTFVfWb1/eyWbdDlNJNv/8ur4ZF9aU9a+
vv6B1NJpJEW/dtGRQE8O6UlYtzMuZL7QRodBU79ULyXSdvQd3h+BBfMGmJwoMHgnqWUw2M7HciYa
q4VsHQmE20VrYJRzjJ6CNNTMhsrscTA4Lpneq7j08McwKm/otofczjcd7ehZTi3Tv9tP2WXwdyIF
voGPS6jBpiE6tdUFd9CyNS0CQJA8SWjl48Y16NuabwaMoqv6H+8LnovAYjNPZmkF6nagIn9jESP4
yLzi1H6nJuNxN9rxmtC26TxK+oYKnat+BAeJ99WHwXKhkK9p7Lhi8XCU/AiQVoLY4Ni11FeicGTn
DJ6rR4Wxjvu3FVHVq6iMLFT12xug7a4Jr1Cg5tonFAmDpRVVTlwhO5kPrsNm93Lg8KZJBB/bIaPN
gsNfPkjHPCxW8edWA6iu+c4ZpQtur3AABHxMwXFRnGO2elNFztpmKVMjfzmdWybpvw5b5wxeDGiT
/6mwaDhNH1+4BLK6vS3lESEwt/9F/HoAmQmjW1g9k+pkf5mXFdlXbkZEkmpE+zJjuby71G/esm5p
Hr2ETbI7e/E9f/PWgp2kS+Lt3Ej33j18uQa3IXcD2vtwIuT0A+AdKjvotP2Su4S9j8p2np8YDIQ+
8sADUaSwRkKQJHV8EbDTAF95OhqXatkI6dgT8cdJeyEk8G8RAkwbpjQ8NU7OuMqyBiSE8yHAaafL
IWikyZVno9OzuOjyyMejieAtFnJohVxN0nhGdbqqTOYvoDlHO6N2KbMbsTdnVogO03zhhtR5CCjp
hWxqgtIO0E3djny9MwJhcHhVxJYZSFG1M/zlFt1mPhEvW/XomokTmAN8L/SjlTe2sS06H5eOyhDV
t2ncywTsRnmDqWpemACkPmp1BaOY0K4NIdMr2fZ6ey0p5TYiVStxN7gCWxZ/PQ2NxKpZPuKq1MFP
sOsT/ADYaD8AcfYbTtPgWcR8lO8CJ5CiFUhkQKzzA1A7FP/RURqkFejc3djo+Up6LfESKwvmo5Fl
EIccm8atbJXrMxc+LlaIZn8ZseRBVE1gIgk9kcAOv1cQQ/Uce6zwXeHNDGlGFDUpZSF/7YwksIA0
tMw2O8+GC1lwDqprNA3vxlM4kZAD6n9KGsaVV8CeGKEiyOWMPQnZyS4CgnjG3BnFkvVgmhhrodqu
p+aDLehqvV5eFzqIPmrNeEOFcbwn7wIdv3g9c+lWX01cjr/BngGB+GH+7nQUCzdZHH+ukWefdRLb
ZbQSZrvv8utOgzq/uDsw34CJVnWR2BBjCyM0+obrwx0ZMZmT1Sf94S0m9J7+R1fKQFFkLU/r4NT0
BpssBAHAvoyM4+IIhjd/A3zt9XhWgp10nVLK9Ziv2rnVS2doIl7WLXu6bjTzHKAT6sTrGJpYjygv
kZ2G1c1I+li1/iRfJpttWX8VLVGOh45hBb1bKDVPlWsudZ+ERks0FGL+6XPqXaQcsrGlHM7Yla4R
mxmDVNZ1rZ53HdAZSSSrjkN6YDYjttYv+ezDBX6+Mwr35eP49Q5sY5EO5APd4FlaRH6SQuzwlXGp
BnldFRI0cQA53LzBYWO4zHp023W3bi9PR2yDdVQq4H469g4gB0Q0qh0iFwiC2fsUIDd6QL65WoW4
qf1wR3NBGLvmEpUGapTvCrDsl7/qmowb+Vz481dr+LKtSkk01hL0efV/WAg+sTg0kFXkPfE/hV1r
o9rqEVuXYcND15W3jKYbsc76eHlPjz6MlddtsK3/OjnekcmKKJXbwI0cSr45nIvnep8kGLUyg5T2
KbLf78ebOI26U7ResrCXF2hdtA+IHWr5sqjIT5g8CLeUMzBTog8VdbSRknm+R8FwC0HkLArAo+ey
SA7mWJqzoqDzPMkm80y6pO4YeAvhWyaZ9BcYd+370j6D8r/M1uSiJjTMGEF3Vq8YTBH4B2orN8+/
AlBoy+8t2Dkwvrl1GSpnvZEhDHEn/Saajbno4e+MhNxGlBl+E/EJLpToCTkkl3HX2b6E85kDR+Cv
/JBo4qKfJl14dXhpsAsNihF8xr1Lyo1LM3jZLezjt2wEvmiue+9765VgnW2CK20AS90+3aE/X+ZA
i0gwgZaAlJSHJDmgGuF3oTepXj80EfesrVijfHFZPUvbACIOigki0aavaLRe6OeLx1vg4X1r/KEC
EET5FYZyqpyfQGioD2LNvtxXT3hY+i+RGUg7b2k8r/u4H+G0C1twQHXM6PbGdaAsm99wrTRAQ1/u
if9RU8ygEnCmLdievr6tPPnMuJuq9HhYKSkWb1xBprQQawVpRzl/6F63EkQifyQO+dqDmxfcrjM+
Rw99+lgFRKGChz0hxNyzuEQM5HTHmD3nFEypOvFaJc2qqA+DTNNaFL65xMu+1mvKnLicDLw+5Duh
YGTsDD7TAIrhT9CNwtmUHFb4kmsLGamHZweQsXqv3A2j1JRFlrzMnBAbqODnNZLULhp/6GK685s/
5ydqN0GU3vRhSRTaKnn0oEHyVxbsenn1JfyKylU9JtFJT31AhKiB5ezCPtzMC9XTERr0zyaSMwsU
T5FNt0I4fGXnSZvIaQms31M4TNZJ2W+5Q5qPkK8fhTd5DI0gFLhVLB4vlGrSTPsNMo5OYfuGkvRt
W//1h16zTq1o8Ms95iLDBZZzWojDhYcaGQsXQ8KyBIKBOgrrc6ieakQ9JUTI/FAcwtNHt/KzxIxE
L1zCWXEKf53hyWrhc10VpsXZWG1rQJI75oB5Bmcc8xdPT3l9Wbz793tn1NAm8HQtaw4WeRSIm7BK
022Dp07avY92rHuzvnbPfmxAft7AQEfLlIikCPyGeFUPr+dreqvYkFUdG23AjSsTGhfM36Ms8V/7
QgtTHeli7wMJbkHCYagiR9l8NSj3nd5lfLrGwUQBBnZCO6HhZkHdTLqLjpgdrRfGr6fyYHqtRgwF
6JWJ+Yj1CH2ayM/LvbA9IpOohqFnRJR2PP3MLOLG6LG0D+O05XjdVz4cyAaVTK7LQsAGz7/edI8f
Fq2PY9UO03cj3dW2CPwozyUyMWLTtKFPcniMJPK712icvp0ZcarAkSgYO6tmMIhZMF/ayFU+li4l
bsbYRPgUHHLTzfTRIwiwCO7nFIhyKJXpTNMjBbuVn+WBeCC7h9ailHN22WpqT1FJqGBUazGmKWS6
WwAVXkOKjq5IM07UKf3pru18PsVEopK1qKKDsQK2sJYgeF26T2ce51oRI3RZBWM+ytPi8jvHNVMk
55zOtL60iCUp3S7STJVtTfv5t/ogzONPUzXBXN2CwtXzqzU0UNf7iB7CLqvJkCZEgiWMfftYwps+
byE7t4KUcp/a/u1Qe3qJy4ouWCZm42Tj6THzBC0uQha0bBd29XlRRhEFbd0AzkCxAugXWDDH9KOK
IPtMQwjgP8urIjIPwwSq78GePKMRUjXSoiPARMO4Blg+B5iUa3OTDOje1/NwRXOJ74beDutOrYps
CuOczNjlc+wX5AGW/BjctvCVFZJ8ZTWS+d3TKAX3hgjJ005J5YBZkXE4DpnRrl/VOLSryvFk9zlz
GD89+UJm1yIpv3Rpy5Pvv1vJxnwxtwVZMpClJVlvYD8o9/MDYtNBPnGs3A5pmn2ecIndtW971mkx
/INJAqXsB/C0MNpVoNvy76uACHN6P/mubMofQk/tkv4ObEtcZzCq3AEQ0TuosL+R3gIu0U/pgV7B
VHVWxV+vUzhSvksy/qcqwQgZpM38G00RRIcSx98q3MX5feiFtbp/CWC4hMLnb/2UoUwVbWXF/orz
kdN6xp4axH/+sQxq+qR7jbOnrX9SQIu9m8hOHhGqNcWgYJigmIfnqsx/HNZtpVLjolYfmMQhsqyj
EyPqkMdtAUlE2Z5+rtO7XT9at4ZB5zjAc5IUpbcgCMD0yrot29vyCdBu4weDZslIWrIBPbLrztbI
cSye7d6EgOwRfK8qNpDk+bmV9jJ1PnMqBtkycx98JqFgbdOupfWt5FrR0XWguu6G4Zve0SJBllo0
RGUn3zIfccxfHlGcO8ewUZSGLqyqJKwxeZd503384VsGOploM+nEinVCNeNFo6sR+gNICslw8HGh
sgXfNUa+SOpW7sSMLdU2fTeXaFYVBBV1sjBAVTDzofnSNqVSX4JeUfefrq1ZKkRELO7Eeh1k/lFj
lXPowC+9Cm8r/Ny7mNYnZqAlIoGiQDfdwW4o23Q2m52O2f/FqeW4YK2fyKXfDTCPzS7cNvdhFF3R
angZ/7dzQT6SZCbGGZfl9Rp+nczND377PGbVgq9heSeUkkZf2JqDV3OG1K+moJ29Sw21+L4Gd7le
wY94WkUZ8iMPVIzFqJmtyvlKZtyWyAsdke9ozEwTOINTKAAnis76l5ZQIMNvadj9GpBA+TA8yNF/
4JIahWtAzh/pr+nEwF1hoVG4mtWoaK8+A0qK4oDG/hgbu7HL8U6ciPN15sqUgFRAE2QtGRAZBFDL
3dT3XqDfvhHG+ybfwqGALjK2uXe0sanCsHyxcjK0yJc8f7taGNY0RG+vQgkXr2mxY8Q3sgRaed4E
qKKs9wLmIecQr165SiAQDki93iEKSP1wKpQgeayORiJsVwuoIZG1A+d1CE+An9v0iQUdgLaGidNI
ypIKlY0O07zz4KB7hgUuy1IY4gxZLxwxvkGvARFjXtl+tiTB4kil29HBZQpx20Rjjvfx3Y+pjCSA
Txt5dIvCjoQVfHbKSbQjewLWAbZJT/ZfxH/X4z/YrEvyVLfivPrS8euveYuZpEd3urorFa72NgsT
GiOrwBG7G1jH2gpVsjwnb+im3bPLmU2rqyJ7YV5uQKUMGjEcZDo2hK+ynbT6oWH0sidEnLvJmeqJ
WssI7C2v5L83A5xtdq/N3Gd7jwh1dzli1v9HJHc2t6A5asnv/cnV0mKdOO/cf+Y1otYsvwofay5A
F6t7tF7bWxbntzMM+i5gpSddG59gpr++ojH8fHwoPhCGtpjSlres+uuTkc+gX/CJS9cikNbGw8h2
pVevHmIq9Nj8NyTONWOIXz2p4BHWHKKRpiKmoYqW2RD+zxdcfKayyHv40UYuIpoYsFI2fx1F+laM
da3/ZrI73biLD/WS2ihPCfBl8dgGDc17pDlvWd4XxML4YRK7Qr+HheCGYFxoYanwPCW0a0piw7ms
fETYEBdoGaB6IKkkIuAhJmApFpO+YQxRUCymLHUvdx3amwL7OKnRWDujcdu3Ye4AXoxb0YTx9YMZ
q0pcrRgEPwXaJSnj+rRrSYWaa7nUTd9jrQftS3oQf64znPrAv+vUG2l2gCD4QCC6aDu3wpyBAlHy
/Em1Nawsbpnvp6KCrpAB5E5GOqSoKqecJ4K9eN73Zh1hLq3UT7SIEdMXCHs7OL6hOUQWJkCV1FxU
IAsosqeFacp7uCLvlvTvEwEpaW++RMSCepVHRaMiAqloPl1R78iu1IMJw7O97JHLPaGwmz5PHLDF
ZvvthkiIHbqSiaA6GRKO7ZUTwKXiGYq2WP/f911J1Ph2PbHTRXkOf/75etXTpDjzNR2eAVmBrhGN
LaCCO+NWlP2U6wdLLZbygnhvEzynYCLnMga2Jtq30IxuLV86k30DaAymdvxCqHaC3lWcVNetuStw
GC3HIRGKpkjEtvy+o0Qm+JqBlopuzIsxugu3AA9GPuVWpZiTKYkkm+8ACFP/LXOFxb7VRQZKJj/l
g4jANK6/ayfk0NPqvuOtB1CemhDxp8i06aJ2jgwH5X2LOU5PTxZXELvfrpx1L9YeIjgTODXOmsk7
5BHG7nGtG+JH6lA70sZrwlZ5cUNBkdDwc3jdcCDcsiTON7wS+e7lcITMnxfrUAjExq80guiRbN6C
PRs2JYZU+pZNT/JfwWSOVAZjJmL4Lq5ToFhbfsXc6kmntoFA7YMqZHxQfsUzBMZFLiyvq+MOyNi6
lJGYbvqYMgnt0TKSuGt4L16GP7SB0EU3WzVRoobchnFDS22XEQtvU6s7lz2grwJBqM/O+lenGKun
pVtsWoXazJyTIp43a128RxHoquUq1oFpkwRqwlzag93AKvwvkldSLrGNKKm6Uo+cgawjFmn1YLYY
K4YJMQh5mpDR8+UL/pM3Niv03eW6qYEAABnnfouQraKAVqEMtHqoHi1Ha+lWIVmNWbE290z1JhwW
t6SRtDFbCPKzb6R9o2VBJsy5zsAzW0R5ahO1WmWqSQwoHw+bjCSQNTKfr6KbmTtNCtMLKh1AEGcA
iL2Fpi7CqJQywhL+CIvYg6q54csosZ9swvWPY/8kDr7huSNA4o1VSHjpTG0XGHWkcsDfTKPrArhm
tLjmoANosr8R6JcvQf7cMH+8Kuk1YokV5jS3LYYtlIpyD7ZDUx8g/eHR4of9/J4v5ykni4lPZF1f
WR2qkpWxaSA9d1L1lFW0YDMJvjAxP4gN89dmijyFA5TsREJGI/4QLLLG6uEX/clnGKc93e2bEH6E
sz9jNlivvR7er71PDkffsfXQEM0C8aho5uJhZZgo+952cF3NXgvo8VwEq9oh4ptH8r5zgk7LJZsB
s1MQ1jWiX3ygw/PbQ2E/7doNfmp7h9+n+eI+k8asmmBvDGlWi7gdUu6ZhjjbZdWDHM9lJDNFPilu
k3rsz+yXI8mHJvwnHuaEUUqbXvoQy5VHOv9G4yGV539mgMgl+FCmxz+2mGxRXD/kvXA4IWXB4RHv
4Y5W/AQXwcbm81urmLGgztvpQN/2sQwCSFwpuEoLckU5dNmVLDeevu6ON4ROpn6ms2/DDbQyh0If
v3g0h4MGlx/oe2zL5SGsMBOtBeM8U8gcVUWV/bWqFzIaE/YjG9UF0y5Q5HQOQ1vSYtHoDtePOp4c
/uEqngt3wr8n2x/AuDHGjjy619qcvRl9f+OAl47bwbL5lKrKOGYwxneV82cBwPorGNGWTusDtrRt
I9cf/fuAMHoUJymOqr6u/5SYv6duW6sPsUrVheVEbSphaFszjuV1EG33POYLK+smPCIrlxoVgItp
NLb8HWpZ71ysFXzoHscKsGCU9C0Zq/xfs5lv9cvbZtgQS0EiiXGu/ROkK5TFXZfxwh6dao1MNo2/
LtPpGs2E9CIEmh0oViUXNaFVXECQqVyxu3s0EkKyfE6TI8MbYlEsTVh1hz3rSzq740dIhUREHtpZ
w7j7cxj/W7HDvLuJ+GRxQNpKLDZ34VYtRs6+pB8kEQHHWk6QjHIuPGfHCVRMv8KD8/3SvugJlEq7
Jg06OANEKe3IatE5bGaNKzJzbuR9tjkBOTj37HMx0H0uUPqbuLSfq+L6JCtytIM6f13ibV19w1Cv
pMKX/NAFTPLbVCAWcgXpCuhHUvPNYi+vpOPf5rpSZALdfWU33JItySf2Q8pI9M/B4otERwR48KfK
ov/ij9h75rx+0TDVXM0xGECuZh8FzwMBCBOlZtP2Mr7x/G6A3xRMEf/MkibWly3Ph4Zm7/s7RbFa
koSll50Q8nY9UhWj62zAwWmjZSgEBdIBVKP5adkXs8weL9LPy0+TVKyH0GS3o5MY8ztqo3FesfsH
YdK03FmKFOb32y+T6YD6FBz3Q0B41laPa7EcREoJELpkGUDqm3XvtKHbERXk6LHUDfghweslm21j
o+0nfRvo3rzTVGW2nqacQX+vK6J2wFyAZVq5ordqrUh/15toTe42bLeb+BngJoJ2SV+e5dSUcgrL
OfWuBfwPYadRIHllnY3FLtZnT2jo5LZ/4ZvWA0NlJ9pw8WFMsroPJeehjDesSvIW1/0rOqG/hSBj
l/j7UutcBN0akJUSzP3EuijQWfviLARNonPN7SPvRpvzGoXIs+8bUp2tg2uZku/vbYjAsgSSjtb0
iUFXz9wTQNPFa6GmSxWxEN+qoT3HgRLvGnYU3Mse5n/gG9VtSAWmBLoRRr+vl0KKg12GA6SRL/Ho
QjR4wzGUXkhlGREeBZadF6ugjpNAep6cPylmavGlPf/XqFYjiqrQeIaBZG/IN77V8Bqd4ZvvTk9X
BPl+gtnR6lHNnlrOwIZg35GFujUN+5avcB5IKK21oqU8/4WZfjBxFPoey5kmN7rnPnW+BXaXD3Fy
fCrbjy/A1RN+HWE0ctBbzAlZezxrOJ+CAs66w2HwAsvv3XigBWczKrBXePGqaDuk8KzE0N2c04cG
Y37X/WGVef8N+FlwMuxg6zuLbNn2Wp8S8maBAuZEyJoQhmwDYg/XY5V621LxSPr4AjEANqZc9WB1
o6yswjcd9Lp1DyBb5dIfEfDXGDuvI0SFTe0gExVL1xHgYQ4vRk71lUcCLmLNTaiIaiqt8be+JrqU
fteKizk7pnJeS0xAS2dhS7lfKGGtVBKCwK99mNBGHATqlcqZusCxybi/8zA1Wgp0JouQvN/1vu+y
pxSNjEJEKcLtyG2fawPp5j/TliXGUKx70/C0Uu9i0N2Lzlam6I8IUHMAIMiaYgXWDYdpVw/qeaXt
03Q3BzOMOYHPxKk/3FyqmRotECSzKvcnIqxhnYRLdcoTMAqEb0Zn6phkTgOcXrCQiYRB92DS6NKb
X8gHLifZFwQrkicqxSEOGWvUE4b2y08LTwdoN75IVQjonHpX6k7woxDbk6kAjnB1LVz53GI94ous
Jz8MWZhGcCxCr9VHm6p6tYxkhQOf27CDpSrzYONe1zqbvD80u9HrsN6ZCgssko7R7sjEuZobLdGq
Ow+AWzd7CqVY/js4Ew2QMUJ1fJRK6riALAWO+UREaNYq7QESwqlWQAc9G/eApMVCqIERq0Y3NOQt
5ljHkg+K7ui3wdxVXJvtkl9WO3vYFi50eHjhtiqdAzpKna1AyA4ow0/TsBofhZk5Tb7eK1krhIey
XSF5UE8W1JkBQjXvA6ooWIOmW5yLTL46wzbUIROAXwnh4MAbASnL/1RHs6nlvNF15GAo+BpeV8DI
Lg8tBETFrcwcrjWMhJxtrTsXLJ2yyOlIJ7FHkOpGPXnQiHjqdQ7uQRltkMtb6e78vOv+Xgenr2v8
dd4gh7/RK3kLbVtudIfhZ/pX4UT0o6yanq6Kux6IcvJjIlLFcBpJFRnqh0X9Hkk9YrBQlgS7bamC
RsWjwPfNJfLiYysCkpKNFsXUIrGyD8w6gijXqXfAvOq5IlvyJlS7o2LgU7bUG6ljkC5QqWrblM8c
11uxPiR4UmC4HpcwFCwHIcDLP0zoM5TrX6SgTpb93jGdT11oAmKMNP0pgvXC6bNIBD8nwlayACgb
EhJ9lR6qc1WgQBUSD/HkH0T5zwOYOSNcrqPPD2ZrJBv3NGbVpKy2yzvmJqb8+xhHzVFh/AbKHNwn
42DSudnK0fLJ0n48WlPMng+s8J5jaiH/KjgpW/0gmdHfJLCN+xdXUmloIsYtziIcaM7pRULUMHWp
YrQRHp+7VvZBih21s1UyCC2UFjPk8DYJvXZJ0ETs+FICj+FM3CGRU41OqtYkie9hr25GgCpgNrjK
pQsfMd0Hq+rMxGjuEdim5SM0BsQC/BDGeVl6rjHt0cHh9LVL8JwAqDDi82HxnzLMiLWbTgs7465k
IGxna0e8v35OGSENQ7i2MdSTbK/sZFGh34rkWMNjaJQhLbX199juw9NkfkEnmqHIN8hSSdXEDJ/k
O62lpOM6Vml1OAEjcDLomniIY1SQ7IjuktpFjYw5Yj5dsFgG+Czp69zs+smsfGGsrGIZIFx1GdL9
1LKVIZGH/upk2+U4vP4o7fniUmg2MneF+nr2FtGYBB3fx8hHyBnNAsjb8XR2ChIqWcyBl4RVJDll
qb0MGWWRyFUTGLbs0ThgJj5+fXiMl+CtxVLW0ufqWFQ9SUCDRn+XNtmiYM9OaMYB508XZMwqRBXp
fva1c94fezkpsogEQrz/Y1Lt1Z6MEngIWdETefXnxW5en8PpgFUMWN9y2pi80QlRCOlYSZHYgiB6
Uzcf0wxRCC2F910J1vwlapAmTeV9Z0omZGFaKajm9qyLrwY/iLpRhyCq2Ph26EaNPghOyjCTZvHp
4vyMKo0j+me/37fhBaURos50m5QLcLfCdXQStv4w9054zJAP85Xj0bxm+uTGzaOL+7J8gi+U6Fpf
6NwwQcbPZYDpSlix+x0nkd7QBIe7Jp+ZkpijLiKhu2+eA23xe884AB+N4TcuFSX+nrTPzlbjXWRp
LDjKhMM/LBPy2X3Ky1uj/pLFG0D5GuzxGKAsn46xsfPptrrVztUcUd+IMolMF9B+DsCdOwZ1FVU/
hZW/PWL5yoUAJ1UakJuR1H4thIwgU+RTssVIJmUGv4JpV/KBBw61arDH9PCesOTW/LSgcWbgMecT
sHhXBrfNMpJqavGBT0qIdV1+Kcx7U7YG6KAHhhOS4paTMn2Cdeie4hc106KKGN10EUqcXTbc7Dr3
L2GiSoxiRNPmoTI/UAjBXppmn7dMT4IBhRYEP9ie0chqBvdaI98MHna9YvyXkpvUwfX85jjgOFfm
guMEXeCJmpf96zkfMCJbmnS1VhYrKyu8SfjtDcELkyERJ5zo4dG5b3uW6pHBEPDH/o3+m1LBjetT
9xS6wCfwDc9vyEvSD0G2RFh0VbSLA96hGMjtyhv5mbXqb7NttAhF1wKfZStRVwH/PgYZZaj0A/7F
2/vIAaD9h5TbGGjREzAD97Y6wbXGUztfR/cxvppg/gbmoaX/XS/XzHJCxMJRvBLQaDIk/4Wpx4iJ
DET7YlbmKBo6pxTTcCZ9P5yZsyp1fDN4yGZxqsAym8MdFTcYR9WvkSQyxc8jh+lBWbVn6wrMguJa
4UHvkS5fdDcOEaiwfEJ1Rw2DSYyaFLqBN3GjAqrvLfA1I7xwq+y7qviXZKB3bpdWOeep/FZher4E
eetoHMfYi1Fp6qwFBePrA7nr+eTa7L9RKqUsyFqId3R7cKHk98i+F10olI2u6ygtlHtTm9XheQoc
9sRmpqdBmRHLoyMJeR7/wISVxSU5srMzQ8rogKwqH+4Uf3iGHPJqJ1CexiWG31Pb20XtCKf65tlk
1c2etzVOD8fQQwztYBFuYO3xQoxH48AIHZmpwsnyKDM5Yf/IoWr4UjkCq94y2Q0qH4zO2qliAeQk
d4IYkDfaNjQV4ejOffDppAb8+MAMokrTam/6sdDt0KIF2k298lq9xmK5znxdcT1LSv+TyHz83zSU
Ix/qZB560gFuchQ4xgXGB3cK+3GyqeqRC8bC4z0CrwFnTPudiGUVQlWRhH1LXBMDNjtFEcvhmqhe
+rQJzcehEn4/4fdYRSDhaysSquDFm84L0XgKFFYV7PGJ8Ma47dR1XlcOjdg6ZtPGm0l8ozezZiE1
P2UGfXiKwAdYk9hzTPeDKHrN75Mf2tlUZgjVrchyPdQVsuVMkoDrAKv6K2P1NweQjN0hLsEr6zHc
CH0o395HSBfcQIVY/7C1Rb+iISAM5JrNdZtE3RUAPFEhbUMm90TaMeM3vADPjpijv+ER20+eLTUu
6+0KIjKnuSeUx4LntHS7QKtWeQbyx+vQM2Fq1emLlGL5gThy0ApgdsOA8vU5wCahfFvo2oyBWFUd
bp3cvJOzqSnHlnbGtSY1UGNE9Lexab7FGdaLJUImYl3Oua9cO+gXzdvr7Z6qtvTn29DKhPvCyCoh
bifCfafzVH+ZUjz4+uGCXWWbnASH0aWdWLK/SEWhqyh7Gx3QFjpOW2cPsgNqRaIMAb5BDDYZJIdK
Sr4fcfThPG8+C4qgdVJtmHaZlgVYmDerhmHxwnaRT8O94MWtg5mJGUDOv2Pgs85gMqH0bopsOd2v
shZkrIsHJkPV0Dbrkn+idLUbg3FusYNwV02bsDYt8+uruwK47V1BndGcZuxnGFhjEYe7eaUhzZez
WbcGFfqatpq1G2cRaqXS+a+yIj2Nn0XkpMwvI4Xf3DcAAJLlARzo52RBNcGL9GQOUFhrTxmJPvDd
IYbE72912HxjG7QuxtLqyRd+SzM74m1lVO7pgi0raQ59f0lgIrQa9XdZZqBhhkDUBfFaK5Gx7twt
km/N9EFhuoLO7f5iq63soJFBK3uaoO6TFoCIIfPK5t00T8ia4U2M4CNevE/VT8q3yAR1rfBhIjVH
4PdaKmVs+/Y6KTWDSn+DBvlrFvsPEjWdMw40xq2zo+P1L2bB4T22mlrdr7OAJRAC+ZVb1I0vd9mL
ra2X8Ev0LK7ILmS7I1PiuqFJ1gKDL5uHk2Z8yBGU+SGZbGIJsTmnzt/ptT+M4QX4wIswLLjCQZFO
oRUgLgE+rVX/jlVPwtAgHh0FoZnpsZK5wI3pCYlcNelwxPk9X8EDJClQpGZ4G0DTCNUEP2TJZIMm
sRtuRXXe1rOFmd7MytSBr0yZpm1GlsPzOAZYgodAOoE49WP7OLWDYPDLqsWtBEj8zW4Jp7zskm/B
AubvIA37llZnnJU2cesnshUlha4Z+vsWNBS1ZCDrn3lq6ipIXxTcHDggSmqy1eMPPLTyb/ltiVwf
yp3mkKPO7AXkUmYeIZn7gG+lUM2V6E0xjgnAMaod9rFCqxeJ6dU0w9LfqKcN8d59YHaK6InoghOb
RnytsSKZsTACcxYCSQduJISEWubg19c3jPGIggq74mg7lbl8x7shPc28TOKFiBIkXalt0OFt7d9V
p4zXVJn6Du3+4NVMduljM8ATE7cP2n9cwBPLYHmRTAFM/RdXoxAgvxrPgr2etKr3fXsnooSrwO/n
1oTw8BbEC4EUoAK67+OJ31uxgbeClFdo2BsYVPqtb5g9/VYE+WowNfGXjB0RMgtquIasCYArvknD
d6OZl6U/roBJvQpUfy4/OuHXyN6vEZchLdLOniy//qALIOuy0NB26DS9xwxJR8sBG6Xi2g4/59z8
Aas0HoMdbZcdOB/YMDYUYhW+WDS0ANISzC4OSyabeaLMVvFoE++wAvcwtNW4Y+NCfECtAg6UXiWW
FdQgNeKzA5/o0Hb2IcWdZGhaQjRsK1gPWEBEANNC96JEc2zHbxRU4vhIRZ9AEzZqPklbcslSQvnO
+Ntk93/xwrezB5sRM02jrq8KnzC2Uw3RgSQfRKrGt+b8IRY61UGcwGZV3zkupF/LxRg4P+SRQccC
m+NgtVGKPnFkp7id1AMrQagd5DAHZpPylRXdAuljz2gW8RI7hMr0Be/5ELTSe4wH6oHSAi98a8hz
NGYx0K8mokXZhiIjzUv2VYHi9cs2EgEKxn27KHjAPwmX30y7TUDDOkNcs/l6bvjxpNdOW3cbHKNJ
EB2Y2jSTAPGqsBYdgLHrfqKvJOr9kUz4Q+9azXKqRBHk1QOmqMT3IzOK+B2/9CyXK1w6E6JOM9Gj
4+otg+n/fqaYNRNbLhAWYk/6pGCbm8TsTd0927/2q0JJjOm41SyrCUFQVgNrj7zZDk5hJw5sMypV
eZYqZ5MI8aoRM73LWy5J+m0gbTcFUM+6S9TCWf1l/GwvIFDXA1UZ5YkIg4kyzsiI5oyAK2t/XBDy
/bqVeY4+FaDYAj61s44BbvazqnM2YEkD9eIo3H0pjN6fQ4anBRrsDThsGIC02ce5YVPcl6jRYOe2
xVl2i2XtFUgpTMVjnITUhuVdS5IKuPdPmSMjuwkyHnbkPeNQZN9nf32IQ20jN8z9BYJDoAe5GuIu
JFZl1zNmzZprWN/G4/C818jBIQX+DJA+FScEDBL+mt50KmQ6Kg8vybPTdcXTR31V9r8fvQDbZWfg
o3sF/w42RbLC+WNIg4Figxokhj8XpxRffw2F77McLvwZXZLzgcbdi7XbuE1me1vLbCNyhmxaDJH5
cW/OdnZjt+tAbo22hkzaPhvCV/WTfbx9Nr5gCjoU1r1CWnZArj+HEn8f3CrAJ51e+KW6HFAhOB2Y
52eQ6WajBapjtE9nqFrOTttYspNPUs6eSmBntpDwGgRtgC3CQht40exXVjRoU6huUJMhCjQrk7kx
/8jeIXY66utpcdqIpGnuEepmNicUXd0wkIrZkrIc89R/ZsyfVpezpijzKO5eOrI5HvoZDlubrSUu
Im0QckaWK8aErJ/WntKWcNCBRZzx5NzWgFgFGFhD9YIrnTEEynOprafCHbu6VCbEuTLVNtsmW+yD
eyfu48RFbYSRq/XsD5qbCrPCCvHfrpVpj5SUiQP9o0FbudgQEGJY4eu2wlI2pgCEUz4ZlopmsILb
e0VeABm9UIDZ6w3AwoUOpUjAREYxHuPIYX+sHOPisIp7r2qzWmNBO5KW5ilYkKllZNBEGN2360SG
EQbfVQgENojELz8ZyINz4BQfMXhmPLE4qVjGHTI11FFDaSg2nrw2Meb32c8mTpvrfP6Ssu206tPW
/lEsXFsiwJdb2FF9QDIrAQD7pJk7Vz1mYCH/5dmIPodLv6CRbRh4SsDOIl6Yby4+1RljVAwq6WQG
y7NMhdne+RGGk0oWTYNubRqvp2RY9lyNTOCEzEyxukcRfX0z9RwJ4kDxLzs0aE5w8q3rdgsxWpy4
5TnF3+wR+RlizbqlPwIdO7UX40dESsSXUQgmsbm4/EkfVxsJKQ5kz3unfK6dH9EKONJWvAiuGF1p
jUJX/FFZV+OWS7KNIVMAMyWEMljS3yXXqN4ALu1oRFetQpm4BGoXBrq8drgOYRMrMpNv0BZvPyst
dCNA/7jhYkVG/mXg/d1r3OrI2NJErrT1e8ie5yzbzYA7FNrnV3SsSm1C+Ghms+v817R5VECTbudx
+VMaT5cYvddtGdITD8XdUMNsX7hCaYgO9uXzluBF1bng37Ligdvyk7kYw5ptQOzvkYkC1QY1zcRe
UO1N0I4Ll1+XvS80JH3KWRdWvczgwfJ7gZrS4KRg4HecgrIXMcy0MMNTS8sXHRrjF9QrOeC1AT2S
XWEjoFOIlO7nhLWy+sWiRN3N6xmieMdfx6wbRzYTL0qde+DvUrsebd+3kcDDJmkaLSzguuwi00ZI
6MynPJD2YIo4y+HjLlmfJkv29ZQuwr/sLKkuoH+B9Td1VyqjxyMzUv6jaVNAselW4OK9+w+yPY4b
pohehHTAHfDvu7iklC4h9AbAb328Hr+HvrxIyxu2RmAdtJBXOGg+G0LMIPRSIeqsVZcaZLQTlO15
7YjbpoS6WVWLR2OUtAplFW8vCQq4alUXnlT8emFbCm7fda9iQ5N1VDIiuAS+CILKgDU8zbIYYXuQ
BlapCjwLscspPwtnomfjrqX0XnlYjP5383uEISdqLsGfl88u19s8HyArhJzonimPFPbozHaH4PYh
2TSwLvGGxNKT+22lTfJvBbedDcKHFUNUaWkeKAHYagZ8bHvzw7t4/M6Zy5zAR32DPvxvRY6foSF/
xj9gsjkwrAOr7Cx/nJOHvM13ak3j031S0T4J4kFg4UWDGuHjQH4pbxyFqUjYiJDGbm94pOQJQQ9i
oRTzYMBK93srez1WKs5sn9iNJkHkFffMb9ptYHWPcV98XS91eMx6cl6OoPDg0W3H7EGuoGsc2T/B
kfx4FKdlAu6SYeyN0xtExHwqu4NDnhIvfFIPPfj6eQWYROFxtRx79vnOC9/OvOuOyxcMuuCzCnMz
xD6l77ogH0ykmyZeUk5YxCK4AvOKUbdAdcu0bynQ7g7UBmQdjVcCsabCkUxXZRnfkLuWJA1te9zP
clDotIphUI9IyeiaZy6WNVSm363W2fjNWq4CVAxm5S22DOvKjqcHjjH65F85hq40yfEjxuYTKy94
AZHUuPcJ2URemWcYwLbxUDJEB9hi4dpDR9+pwJOoICjkNMKJ2/Ln/5NpoRCA3OjV8KtH/vxGXmBL
GMES0BLNXbi2BqSWh9iEGzIcctse8xVaOoEQ2iZmfK+FUPBOn6gPPaVYLCWyECkf+MorIwmqE8YC
Q/r73jLLY2bQGmLAEFOhgRF19dZCwnXnhZ+gSa4vsPFfaayDCBO4287k7BWDAq/Gk3XP5BHDi8ce
qj4Ij9VdOdPsuYgGxPDlzoe6Jh2ibGiEtSLQtcJz0+0GZvWYDAQcAH8wNVD0uxflTcwOXIySHe9X
ez3ULKlgZX7OshhCG3eSDA4nKE77oKqLjXrsy4j97UBk7UaNDmQ8PeBmoeLtwTSUSCFirCAsiykS
CQNt3hVVeXS9VnDY5tiV5eUO4JtEsIrW7GIK+5zfdAdD2Qlz8kAen2GAHnY94JXLCxs70MuxmNuU
6nD5Wpllm4Rn5Pfnvx/YgP7/vBvDa+wRsqAUe2QX26wCHMqiu6Ia6fJ13g9hYGCb6fuR4kOLZKGc
Hmz1dsnCwf4Bu3aDoRTGq1/2KLwhmnLFBbirmNvhtNuBo2esh2T+iL5bZzQt96vJdd0d2WsPrwWy
XBqkN/sz+U25qYbTL7mypaG3Wibl1Iqpti3m2tRFmxR2rLUZvTWOGojw2PBaS0qrxG/2Tt9OEKqx
Z4IVe/USFCktOqAzvm4xd/wpxa1FvFOFPDVWRTztFmvpzjkYcEgvFLmlLixCYj58b6PT8qQUI3i3
BD9za0baZONtRBXC4sGX/FNoZjuhHHULJBBhxerdsTnY0d0U6wgELFJNWvjZ0TM6MMAE7q0KvYUR
HV9a7q83K2YjMXWiEC12rp6bPxZXAIgyBgxCx4zq12lLlqs/3R1Ag+TZiwLHEnY8Q8KnTEWSRqlS
PWWi5E1lXeUymwT6/1L5AP5xj39GdpjDskp4wRzOB62ov1ku050jC3A5/KuO1QzGV+c+60lgvKZw
isN6FK1AqUI32PI3zpdmUn2kqqItMHiUppAb3YfEYNBdnCMJrs+6dTziNhYQ2GLrrcx14TtijwXk
hv1UScV/XyRcKGnEUMOhGiHugkIvi/vy8lRRontklp1ielRg4Ggl334K9BDY+oPFq0ODqyqOI9ci
10bG/QhTY5+n3OYr8ARkA6RVJO1WCv4chSozdXMAMryM1BPuclQo5gKvvRVjHCYEHBe9PyllXuEC
pPwsFKS7a02FKNAMFqpNHAWEIxU3juMDSEx86IX3Qc47JQOKhBf0BF8ZJMlZ61cB63OlRs5M+RSO
0dLXCogrSBi41F3OXSA3xrF45qJJCqy19bZ+Lxw8hHbbw8vIgX5RcZfzN7IfIwRPWE1iGBgJ9Y/L
lYEPt1tOMhohHPo2xE2DvjXLdbEVKfZ0FxgxJ+gUVkCb5Tf3gXEoOM2O/o573+PiGb/D9y0Cf9zW
fOMX+f9QqoMlGiyMzT+MV87OLAAk++f3nghEsfMpQKaqJEnt5osXI7EuwITN4jphsy9v/ea+DrM1
XQNCO+WhRuXLb+6p3Xecb58AK2d3hHzWK/lMT9YgGn23mnEh6hoZTIc8KIrNMwWTK80Bqb5CFXTj
LeI1kokW82oOvASHmVniESQcyOP1IlgBBcb9PLMT8lFsdIH8GhPYEcaGx9HqA580DI2IfPzEONHa
qADwGb4VVOyKddnWBIR+RNlgC8F9DoyT+YA6UqyHGbFn05LGdQzaBNbzvQK5vDO9aqrqYrFPyC6c
Kt1NQcPfjSo86fl/JQlqiLmuzmDi+FBlXezivLEgYNGIJvlREwu3I+bFWFVhGTcsjVSPi3yapDoB
n/pZH1+ZiskbIjCoG6+LzjT8dlUFRKEWnC4PnGO5F72rjUDfRajyAeZGiHF80ib088R+jvCcHxiO
cP2TUmvkI0RdOSWHf4MmotRGXyl0GqWxLp4nvyH5+f2ghAwRvjQosbJau0XlcRKoZBp5IlJ3ztl7
OlaEX7UnSISoCM8PhzWgnA0Jlz0LZU8AQ5FvFMul0K4OHhVvNsYAcGVjl/1/aTVU12nbr1hDGWLX
8SavEqNNzHGoOrg5OdS+GHmSqIbLOQccMHNuvJ/7oKR55BAPnU9NlIKpDNM/xZDf+cRP56C9POcq
/MxO6K2XDGIuX/enzriZ1qz/ouL2aUeGoARpg7URG7LvcmBtrOUdrOVqyrN4gRAGxReC7E8vSLbT
sCQbb4FTkae4Q+E1ftSQEdtHiGMMSoZ1a4KGL8sRn+BG07or/yhKTg5cLWe4qxgocgVOB5DWzFHe
GljvadQs226Tmam2GuLqeCa2z0zuoGi+s8Czs6umQJlMwL3RbzEj2RN8sipA/CFYnEAwcdCjLMvV
+r4sLj9pfr8mWfyla8ailoOpn+zMNYgLicOpKyFQFINWnynRVwn3yNPRjNjOVQ3wWft1kHeZ4WcN
x20VBvD5KwSMP3/LsrpeRO/s3OwMgDzTe/ezMVXKxJ3cbBubWMKrqJKtIHxcNmBM5F3haTEjGtMr
JFIbFS6+rptu9zKUzLWrqDH6ExRr/Fd9NX8O37bFRZWD/rYHETSqTs/CGSvewytTHKC3htfeDgE+
3STUXSg0PbjkAiRKLizFf5vI4B4TbmgqWx7X/3V7K/Elk7fMd6hrJx+J2K61AQljjDXmqCntY1Yc
9hrkC49RyHr9EmMUnQsYW/f20F+oLNXu3Fv/R/7RMqLh+YUE9SmY4Q2eLqTu74yPrOSpFXTT+mY1
fgLdxL8s+WR78wZ/rwfO4kotb1JjNlE/dvhnugzPV5VDlX30/sods3FAzc+x7V+Dk1G8BsiL4a/3
2Owy5d6+MPpj38jtXEbXcpAHbt8veCplxy8WeBIIKn5I23/j4IuGjUndeOrAeFLQwHuRpVG7RHzp
9ClE9tNVKtk1bUdV6F6piPj1qyDqPJ+TV42t/qq2aPXnSC1VcFVzCqmsW0WqoIH3BFUXgNYdcEZj
piPnme58S9fwCJT+XCxX6yldQIoA5v3IbNGqJ2OvvwmNolxhUx/3Byqko/ms6qx/SFtLecLVsm2i
zYGsAQYepooYWLd9sv69LEbp5mxpPbp3Ur0BTMeVdIV28V3/DtiHCfHxC1EUJd5hSaPjjV420jCU
OXCo77Jdi7d2yg1vhJ6+9r4ep7mChxzibomdDdJ+wkkL1yFcr3yvoZ5p3udCJjVQGlq3egTy9ZiG
tRFeHqWc2EhQUqb1nnXqn65s2GzypiPk1ll+edDONTUkjGGdA2gVqjTsfYcpv1SfZyLfDUgP4NGT
xmg5/32pa5W81CcWMgjCZiFYluZGUcFg9pI/ALybc0mGWfDytYVUVbeVwuF1k0Aj8solwzEDT1cG
pd7Kh5f1W7ru1JFmQ0DBNjWKpukS+egYU8nGOmyw4J01/ma0YlY+WlOp+54JRqQ9uXGmAY0782OO
lhfIrvQ/8LFZdXXRWb6/Q4Qtb4191Ni6V/5qFne0c5E35tydRZ7vjFMRZHDCOu7Uxg0lhhM3cXs3
DkYAF0U1d3U96iIjnQ3AzZ0xYjmiPj+wc8ahEFuX8xZYCfig0q7dyaL57267h6LD4uwjYGIqTeZI
cdEDFjqOp3DzXv2eDM/5NafG6X5o0rxn0h/JHRVrE9tmIzT8hwIA5VuOlN8lIc8n+h2cXn75PKxq
DufiTsgKdSiF5LmQ1RJL8k+WUBAeVMuIj+RuqqgoyJAvk7qULV31qcf350njTtXq9BkRVaiexVY9
9HeGsD6GJ9OmvwWxvau5GfFVY45DrsVFZIZRia0oYTyWslRd5xKjh0FwGzSX8Hk7xWC2nFpT1oJe
7ZEXW6ND1LgHRGaq0ZObi47kXDhJOclxKnWiV98W4S83fikNkFvsZwYK6E08vWjXCnYwYelJMTdR
4NQcTa1b/VzvyT09DapY/uQZtIgVFcsDjg5xysRwIpKdyswvxCzxr0VpzGoNNjSLkO+i44PL/iL1
P2mG7aCCkvIQc8hL/AOrw/how6ERwj5RUeIpw16Y+sOIg3CUM6EAHYDfyBoKJQL3kgNXwbPCw4TL
0cIBlBu0AqFU3pkXnQjSzN2VIrf0ZhwbZ9aPcr71FVmNdCl13tlreU/R2fjkC5u6KdFRmV/utXtd
CyBrrcj/5hYJv4B7PxdsNT7S/XvJx6Yda/WqR5KSu/09oQAZVUNS4LCJPDq2CrFDrAmlcjeDXbSe
FExcCRd0ZPgOLWSCy0akavUBU8YeMwLo9zkZF5XxN+XQslj6LNOf1nhXAO3QQGQbdaoDft8nhEH2
fcLDD9B6fVhEoZctlYhlAFHI+raxcrh3/ok26hftNXLKH5Wgt5aGFSSVPv5wWghN/6JVfvGTlm87
zKi+UApANRC7b4riUHq3+gfqyfG1iChub2zsfyLHnKM+gSk2uHlma4luZJSb0wEgtHp67yO0oyvk
Fd+Ys1qi50mnNmarD5vX9dXDtkjBfSntos93a3tQVdcWTWvOfY2wZJVfbOe9oANT1SY5rhM+B/T3
T8cCK39Nz1wqh9ugB8TTtenIyskTzCyX0wiSUTMDMBGC0QBqns6H+1R+a5mke7hB2J7q8bzwLLk6
S8rMIm3hT0XqSu8Z7akGlrKUXSHX5URIEdTHj9CfSwKzrYrgnYLcIScTdT1loOitHMmGs9vjwZo/
kubYS0Pqc0fU797pliddqYzY8BXj8G+6ZJ286QhzJ2UIGSt/FRR0c3TlDJI7Cs/MyRlWizNkGOJ7
xZa5EBRvhw27Bm4agXnixIdpcLxGhGDCBgBchOoWd8XOHj2vmNKXLw/uEUvfPXtT+Mj+K1VBjNbG
poKrsqwtIVU6UIJMFSfc/8diMq6w/ENRa92otBohTTRitwSVTNDETxz8PmNLuIfeGBKX3rr80W94
Y07Ddkssnu/xYacTf/SBGvrLQkhrkgZmzoUfsJQhD2TIi5mNV1oByOOklFN1a87FIv/+t7q8z3Y7
A4mrqzg7PpK4QfE8AIsj48uNOZAhd2o9A7j5U0yYamcNyNAM2jVJW6XLx+5lm3NmOFM9qqEG8yGf
p/m1AdeKXXrQZ/EO4BE0+MSQ/MwkoNrw+8EUV6uasHoRTFG6iLCUF8uZi23yT0m1ihBc+TZLLoya
zeleED2Kb0zaBpweEXOxn9uHggaDspdoPy9BDf8JNlThDPpj4A+pF2Aagf6QWjRkbyFTMuzbNXCu
edZAI9oNprtE7eBoO8nIs6qPX3ilLPJlkrTRs6jYbpG1YuGK5GN7pVkBOPGmNunr6HR+AQxVcZC9
Lt3HuVsHpXfpYYYcuNZfYgF0665Sl2l3+nDVV2HJvMmBKj4fCoWbGtjh2I7fyO688IQ/E1NaBjM0
ZWF+iYjui6Mk0I6ty9FGgmljhjcCHBkGDOubBWRWeZwQJHU9MzR/Set0ub8hXn6zuhjeRB/6nP1G
igwRbp7j8FJUpImrvyN9NBMFNOfp7nzRvPN6K7Vrv4ggHzh366zGQdVE6lFhgVBAqAbV2RDY54tR
miIDsBkkyjJ/drCkm0NgTHX9g31179kuuJcDshlWjAQ72VHv1R4YtF6kfzOl6RPbdKYR8Fe/Mbdx
On3pp0/eTK/3zrsrdkXVgUm24xAbCbs40urYBK6V3OEhnRRLfdwqc2bJwHCPLHj5314O6CpVJCdw
BpA8QmDSjnkxhRFqSOe+KldtpbSeaeixtVypOHpFQuwKx/l5VIyo8q/Rn22j9f2ninwYNM7auxEr
tDS/ZS6O1ZnJ5yydGbACLqOxCIK4fQGOEC7rXgD1CD13b108rFYhNORlx1DaQadXRWMGzIm3eEW4
f89SXHrqno8UtL3kD2JJ487ImQYYN5+aUpcqeCNDcT6vtBHFgeFbMKSfF5l56pOad7mKe1ZqVo11
H48wlFtdpm5UWuGQUk1V6OTfDf5xR3WaDor7n1nxsSpkf9JXGHLNqRvVCOFPOPc0OLItZEIBv2A3
scVwrPNJyJ/IpeNesKObrmnOBuuwgCRc6/B+PlUTm9Pte7xJMt8X/HH/sySuLuOhJP3bPdtSlf7n
Ba58Rs2WrIfrYvXvheQCAVloI5aHnLGPTerq1ZHU7EZ+uYMR5GwsvfdAhUpH1ixrOsFfR67kMjFe
S9QdrIu6Yh0MS15ADxGOs8U/SrabmqUEFcvC1rpS9tVmIsekCH5Dq4qOhddp50SK6D6o7V+f1s8P
AgPZEH+8shrTKWg2GP4XLrbaLdU9ml2x5KqdoZHkngP1EQy2Uc8paDUs+iHspAa/XuUiwALTFpT+
0Ufv3tsR7ME9Jyo0GHYALXv/rZUJeRb0x3dzddoOHJVoP92hvpYMV8Hs6Os0CjveCMqa88vRTq9d
A2Ypz9sGAfNFX8LsU/lz/rI4I0tuIUxvo3wfeMJvErmQdcTXajMUhiN/zAay18mAxF32HIjINR9M
qY394Yo2q01roNJ2Y5QGDi+PHdNZRpVLJLoSNcTy4uBRqzeOw05jK8I7SwsFdzUAZd6FPsvO0zP5
bFdiRybZHbffEVmt8n9tcVpZmfGB3gWIRgSmtaEElD2RtJiqzjLlSxymQ0afN25SQ0o2zTmD0pWW
UgQoKUG09ChR2rcpSNJke3UedMBrUE1wKn4TJvciAkBR+2i8WU8ARsqGIhy6ATnIwcNVU4iY9aDb
TfzmMtDAYYCXdX6ni6abA6m4Bg+wLytHVnGgpQ78rjSBUGpyr6HxWZeAtkc8K4QQ8cCLizLmr7V+
Jb5JV+lKFdFKXeFbJj6sm/fDaSkj+pUZHOsZ/O2a7lYlOgYIVGQckiJjen+xkibtBJqLmeTXnFIo
MpES09cUuhw6UlTbNAHPlw/kG8+OOOxdIvt6UxYxjiJyiGzonWOQPdo/1swM6LtNBl0OGVRkxJFy
2eVF/QJFga57KU2TkYOAe4ZUlYUYUuQqTHscGkrZk+pWnl925PuRlornxUuGDUudeBiqzfWUu20y
wB2Pjv/XwcRna9dVgf/DPprb1J5IV+g7dsrO/ovr8cbof5Ypzm22Bsma9C31VLaXo050fVZNFn7p
VKe+1WqEscvWcsYrwrFcSKdThr+C/oLiCNCTDmxxhqPEdt/3VEinpT2H5KmOKefUbPWWy2pVtgRu
T33fukEAlF8Zsapnv17NyyFuulsm8I0WnQCrKLahOsPIisz4KfS8NuuWr2uekdOaD1ut3XHZ6pAj
xEnuLcbNflh+zEBOJdVRAaAL/S2G6reAS0Ss7vLN1kE0f9O7ZaIyHP/tmxbUiO3YxOm/EBXYMT7z
wCW18Kr6YQDgYxyZE4SYiM1cMjSUDR0JLLUETtYqsS5H6o26LXFr4nhbN4wYnt+FUIwVEb19Bm4g
qIhRHvOHKWlkzkt8GEyrgSsV534ZN3TdoZedEzPCsF5BDmOg83kHi8w18bRTitfY7Yrg48JOQ2P2
ROI5VMqSyuxwGuNs7yqECP0EsSyuRCyDELtXV2it3IFeQ0xxlvK+e64fN+lGfXj+H6/DmUSexWBd
t2AqMqgj7byf9A7kFV287nlptWzSd4ZE+QN0Qxjgxq1JwEnaCoFYVEJkMB+dbq3W2J86xgcMyWQD
D5u9tB79COi+/qcMDXOqfHApeMGYXPZ7CNnxyhwFRfg8ZP7ntTcRICYjGU/a7HIJbHxJbAJN8+lr
S0KRqwM3brFrsxAbg8tmgaG2cdgiFxcnJ5HeMI5VSo20Mb7O3vU8tmx+cHGLIlimXsTk8QBi7VcV
mMIDtS1jZrW+nGQ55W/nZBxH4q+gNtPgp2IVvWyqbWYOGZmbjsa9vuFisEk6hae2jnhypoX2GhLd
nbXGR7ZycdGhFjmnu2YiqYEZNBZn/dCmDVj5OJOb30wNGAu35SYblVi1BWdxUf8nLZmfhMdnFO12
kySpYsSr14pJzkUveu87CeZFv3EMHHIV7Au3lUqO3LTYfEx9gCurrVIOGrJMKDkHYUwTwAC+R3Tm
N8+HatulOd/aiZvONt2Jgk5qenKQE1Pyd7AyC/kGDZAWK1FCPQclF2wSSMS1evz1JZ9QI8VWOHbi
hrXqqT78qffvOhZygnTBtBnNc4VlyW73HNd+nNgQ8pDZxi0GYoRp36NcT6nWIjP2JVgqBRg5qurW
VwtBQqdEPkMbuEU/ub/00qkSTgisrI9gpiFKUbz3/GIBU622lu31xTIuWMxVq9uKDEMVDwcCVyPj
bMolZe3jfLzyTS1C0VhqOx+VSrKbwMTz2R+qduqZs5xcVD76yLhlA/uQ8ViLMUXLoFpJFfoz5aqB
KE3/FwWFp0oPyx5cUkbQPZCqDaTAHLmoh6fg/pyMw3c3lKT3PEnyLouJb1PnQ0qZ2QroW5obLdTC
ytzL6birXmciyS4/zdPdxczA3TPFjMr9WhrkH8yTFMbod3dnZ3XcWI5f1zVVIgPFDwQ+W8J9tZua
xDzi5H3DpEST7rLSn5nWnlevylmlJQ6mvRuUm92qfTSbopUDpG/vtoVb90BWyxz7Loc6TdLmjARc
NK0yBzKzy/bYRbji5qXBpoYP5yh5Ls9Znw8c9Mhi4d0qUhindVYjg8HVbzs2ektubkHZhTYkD3bj
1nxH1cI2c40rP13BYUv0NyrU8xMKqjBVJTwMwV01ZG3pAzru3Ijh2zFDKDYvGs7WMY51CCdRJ65C
HicV1SJjRuRkDTPvB0uOrMRKg32Fb5fFFfXsm7aTc9rbMtMxCZ7sepe4Nga5CVFMw+Rndoi+aCMM
flOZHjY8bDmyriq9OKAkxifUW0FnfGeNqNGvUa4DjnRxcdPL0piOytDCOJ1lSgm01ocGwwUB5t6k
CCsj5EbShMxkcqll+OsbFi0M1J/cHJKQqfCm+vz6tFBsE9c6yk4Vgy34XWl/DPAM/IRkGJ+VwO3e
zUHpdVp02hXaAN40IzHyBuCBUgffDplZuHLqlR18/Zi0ZBzF0m0QCsom+iyGWzvK3YtXDAvGdgyr
aF+1ZOsZycRfKsbRjIisdqmiT3S6pLjJzXtuYgGPrmVAhYcftgUqEyYOXDKrt4AecCsqMjYcU+Qm
CpKkiXg3OUy/Ehr+Pr8v0xlwHeYB+yJXe0nYkZfbZdj3XYlEafCJM7gMcWuGzBRQE2F3qpSdW0et
/+Gtsdj007wyvyVyTvJfcdEvWZVM3Kqxe+77FbbGQkqD/BoDpO2adHeBObvbSzCLRjw89tU0NIFQ
90jyiE4J4IXv5/EtZcUROm2z3M4YilY/fp3HMVreaqOfIpZHZbdR+SNGXlTP7zWP3yHJz/Oe4fZD
H5d8Q7uuz7z28EyuwJOpd6DddEa50qw4KUys5m79Da4rFO+sPHyi8SUShXDc6Nap/IjF09p88MrN
jZN54v0gopUwhPcUfOZTS81UUx44P87edrWKiVQpvQBUk/S05SqX2vV8NXVOrb7UFkKT8ypwPXOj
es43ztAegSklJelkBwGo/I1yQ4zO4MNYOyj0iwR6AFToFe31cvvNgqv0T+JYr4EgJ0Z6zuAoMnB8
HSpn0AAmABAUGZL3lvXXDK40VYGJFeL5MSY4vfScas4Ud1AZY32Q+5Oo1kopijENwnTOEJwYbzK0
HXIU3EC7ofF98ncCLVAsTxyICmqydU509VfVnOg4e4tCE8Ivd1k9029/GqxkpSwjtBAzZuFXAyBP
Mo1pdL9WcJRJ5RNolsEtHGDZqVRu11e9Kg2/LJDB7CWhUftegwGmrgdM1TUhZ+U8OULX8HFz/cqF
RRjhTPJIBgjSF9/zRldu/sdhzwDGQ+DyWdlftVEz+6dv4M7Pd88uXBDuBaRK6nljujfmg6INnTmh
G22BmZl7jV/gH9YMkkDaDBmChHuUf+kz8Cw/JoFrGr5aB26pJy9wrutA/RmT7te9NziS+Ec7UH9e
5BcrTSEDoLClhl0UsDSJYNLJhV56MYEfRax3G6IeUEmB+O9HptPWWCEwdin0fFyYYoGk+7nfl5Si
2MFA50t4prcn6uxEOGxKPOK3IgMlOGkAIzxtNP2plDqkqOICjFN7m9f8qvYCokU/oVv5KrCoPDMo
eFt7fe286xmtspjED+JeNTzag5/Sb2auzlXCyNcrQBwWfpUI7dRyVa2W8RP8RVca2Uttf8Cyjyki
6S4zYfEkvdKbFm8EIrY/VVcr23sn2zlx8Ac68o99M/FTdTcs1Lj4Ustfyh1QtfRFwHpkN/CAZR59
WDvvI5WpdUcHkbiN7UB2CBZfGH7sQQWLhPWLAgeeEd+MDqJZyVh7axXkTFyoAPQkwqRe8+JXmiXP
1kIp+o9ZiKGCcHe/Y5COpaGA7WefyP5MrOTKJFUjViFXXuECE/nGQhH6cG9w0wfQx5zO+luGozhT
yKy7RFMV/aoPaqoKYNcLJKkHY4xiYCotIZ9M9tdaFqWHVbIDgmLnIOIqxqN33mLLqAHTzLtEz83L
HoePFlEKThuMxMJgbevMbXuSQ1twuAo9UHGBb7C9vyAZpiken2ZbazC2VpbL3vnbFa2OUzyMgxmp
lGCoUfwou7utRap8tvGrla56OjTqZrkpjC61VvhmOp7Tr2WCB1XKUM4f1XPuZ/reNpFMrlLVlV4o
HJjsGqhrP/PyaUOfkOyBfjGsOpFz5i5Cknh2ORY5tecldpJpf9b5JVPZC5+wn68g5/6TkXPnoazJ
3VAk6NvdODgx4LMFq+rgZFodwShQkVH7bnT8VZHrJxZeSjLnrS8cWb6qRCNgys9sIuoliebVxegB
tQVi626kA1uyyS/f3MV2dU+k3yK/JCd3WzW33f9RDYmspdDOOQP7CwVt0CxM7wQSAj41FTUDwJol
8Zd3FRz7Fjx3mUXAM5eoJ8tsi/Cbn1m+rywNuOxVQ7cpo++Z0JByIM8zh/cLuPWilKYgvaGCMBlr
6uB/aYHuyjMb3g4KzLZxZ37b6n8usZZ299HkOzG3DtwmeGRV24LRmBeD8AH7LQBtYm22mrjvd0MT
zhohSJaaBSd0wAzgJrQENI9/NkXQQl5fUeEoSZ5af1MvxS2ZodtGbKa/TwlUycCUYQYfMW6fLx0l
bLcNVGMdubAKepncBCxhiln441D8I3T2lmBWOTWyAKMU4U1l32nBqyFQzMWUSEppVyuC3T/B24G4
7GtcUfLHCtBpB+RO9P6T+B9Bk+22uqLoId1jWzUDMu/levfbHo5Uy4UgLJ38zxCDTt4uUGaLwUrN
p+lqge/DBLDEOACv+AK0G+LKLysT3Q20q5QjeLwQAxNSi6SGwTNYsLpkg2NGiMlyGoQUBnwpuPeE
JglCkkIOjDozrhy82LvMfppALNgakbttMPnsGYtDg/B3pQQYlNqNOrM52svu2vcOxJ4V0WJ/7YYR
ayE3ToNv2vVX9Mrk1JJDQptqeTGItV8ObXr9x+6XLeBZqA53v0p0xln/3VGY/Cu0kQDPCS45Ku7C
4yD0OLIEwZETk0y2YOqeDtDbhI2GtBS2DzZlwmHnT3gOnwk19Q8QThG2cZe32n3qU1Nl8PZgQ/7d
DxElHkR111SVEORzHDyQR7468XQvcQfnzHkvG7fr3CGJSxPcTQCYl6cB2GADNJ6lBH6iFEuZZXcr
jgCl/oFKG9SIOjMdudDSuul4ki6zKGOXsCqoTvKUkd1U8ZTe0XBej5APaIQSr6IxxXJw59BcdQ74
JwUH5oTtLnmnesTT0CRQ3v5+OcS+CWNXuUAkuaFIeJNL81SoUQR0ad42vT4RnoKOWkskbZmGZVVJ
XJ1ncMhC8e5xUL2+8hCmD1dcEJBCmV6Aawrnq8I1q05/NNco8bEBpgik1z/55REb6aPbgqtDlm9f
lUKcbO1NPmF0Bm3wxYIaH9VDimBQF1RW64duQOHvS5SM1gBmPOZLsejimyYJ26oC18Xz5TevtDNg
XZH1C19/9aDh+I1N/jkcy0xGBSN3/aehZX1Q/Lo9hYMKtTuJYWuPlBFHggOzw/Ikz2vLQQbum7Gi
gUuhFO68PjZxvFeDeIQlIfrwJIgxK7r7cW6DPaNb7r7TiA6g3+F8WZuV7TJDeCKaSJyQNPsME+8H
iT5DVNbVnj459PXe8hoDfKuBjkvNLbdeZhGONFPa/Jx3vgHJavJU+qHZdCoUwwRc1i/EWcu+eyeT
oT1I753UNfSrgZ3CYV2mxfpCAyTMwWfEIcpJVV21s3u7/OrU4+5Rrz4c7CPPc+HgfvFn1TVxXSDc
Ac8faKw/UPTvoc+RdSDZ9H+JftNynKchHqgzqIUn9Mxrg97W/pK718Hrj1RnH7ui703nC8BsSyn4
cRQygNeMZyIfWW7xkddrwjrbWTvkkWSMjN/ZxdR4I+eQgLmiXeAQw/30NjDcJ7th49ZTEHfoGArl
6amzvqM+/FqEBXmgWdxSYbzRwOHBwuPdNeGVGAcfZINzrKbJsw5edziaE7PLI+JbApR9FX3sUrbt
OcBlTd1Uu8uz14q0N3yCmLOzIkKqNJNAb97DdBbUmtg7mk8AsGG9qHDkPZeaSslX0D7cO7bn38FE
3dZQf6LJKyQAB5I+RQp3q9E+hgwno/1vUCIm2L8gxnn1hxkJL/ZdlL4uQESjoqGeYAyhJaZDY/7W
9fM8AeypHIzISH5szwRo5vUDsathHydL+S0yQANEwRIcFV/6e9ApHP7u0MkiqYW+C1GnvR+KYE/M
qkmWf2d0wSaJzNSC+feoSvMjwTzwaJEk4jvKk/H63fX2O1Q8igFGqCvE4fFaoPYkw+CtntNYWQJK
Ob47mhqyEJuXmJSHxNgj/TaxgPIIpspDryeDNckAOh7U4f9PnI0zaeTKxpjSZ8lllghCMSZO5XBT
Pq76lJb9joP6iFAgDlpTQjtIaBQeY71omDwWwb0gHHzJx5QY0PNOaglSuABjqkfxCPCGRB8WHXWe
G7QeGVSPUCw9osea3nzchs1s1J4AGYSpLbzAYHXMXEv6GLjGnoBG/qwo08e/LKlY4bIrMqbpEjb8
X6RtCcLkSjYhCv6EaasNkCypOH3DbdpCFxc+h0iOpRAJ4pbXq7j7SACWZqnqy2cd3e21BW5dsRfe
nWLfKeUsptjYZ7wOYZqHg653DtDohenTuEtaFaR0r/HGdSWCtldZbGQCcVKqv2TwnKZgzHivG2de
cMNxsXi7bi/Wf6gn0vDyokdzSMUEt3Cn3ANEMHWj+g1UgA/Nx1lr6UxVMBMEbhdfes3S70CF2EHa
r1l+P99CGXaQH6AyDMKl1zhsmyX+/Ha/2gAIrKTMAxC+X/rEQnlyHuOj+mz9a8yd1fc6ywyQuwyA
GLAishlDYS5ywNjcCzyOwT2eDC02vzGfFJ+7bkXIZjcDr7a3+kOm7GNS7vGcTlZjz5Dp2W8dAZqA
akVCFmVgH+Kc4dV5u5yo6i9Nlf6MEU8cxBjn8LHyVBQsOzm5Cgzm/5F9l65tBniO7Hql1YU0OUeg
Pu85wRBZu3Wa431V1XuyYPUFnXjcI7o5hOcwGxJqRHKNuT7EosPF64/2GYBWy3alFtnW3xtvmYyS
O+E1+8XNn6mO+yly2IqzqJ8b0qvyIzB+QFRtY1i/ymeZ+eLnMI6PeOUuHdpTvA8zWsTqFdpLB/IN
omMh1MlD3o/wFCkWHZ/87hnPxCpnbwrm9jyxmDrGGmsLPqxfkdT/D/oZGi7gP18aGAxYJp6MHa0M
L/N3KNPmzCQweDdQDFdxmB2T1UXG+2qriOaSCOVyp0rsEU1pqJWcm4nIdM0AOGHwTwsz+bErgI6F
9wF2jtRAwEtmSK+j8CThReZUdj1TfEV0dmx/bqVBptaqB8ujmEUB8sTyhVRVGw2xKWCg4TFbmsA/
m/s6hg10Y9XAmVmAW6jSBLkjby/f4d8Es5kv3Al425NAtwmVv20mgDj2rBaCoQQPW0cxKhrmfbap
KonX0LSo+4alBVVbig2+5zHab8mPNAm2I/aLJ24ynJF9nOCh4ypk4UkTkka0cbIdomt47clVNCi6
C5Le+GwxN0L+xJJIOdsglZ4q3AWt38BGJrJPs4lk7anWNuksTMAD1DwoRprp3VejgoGrdXWTvAwz
s+JTi4dFh38rBhfc+glYEQE/G4z3B83VUkybjGZYuk4lr8Buxk/YRMrJHXuxJw3/AC+of8Nc0PyW
WH4cBWWU6dLLGoPI4tdYI+yXNqIvr/5AI0HQ+C4c3w/is2xDqzeCvt9fNgHrtnftti4ZGsSUO8tt
BEdvUOGT8tHFReekenpxExSgCUIFJtnBw0khRtFy0wLAzX98OHUYkbFZ1hbTwEykyYby+Q4OCsl4
Gusa3dd02s+VDn7WZJWKYk1B1Mn/yidknT9MD9YFVhxA+RsGIWoSUOFUSN6Bz2cH1ReMfpFPLi1X
gqr9HJ/52zMwbLhCNBkfmFQVZsVaKurDdjzgUVPcjsdHwHkLG8KOBfW4/vmp5bRGbOuQItL+N7Nn
5d2mTm2ItQ3Kw1EPVyrPsYPsNrzTd8odKO2YbgyuGYwdgAxljtLHS9wUlhK/p6htL+fd8UzYWTkP
wuJcM4KXPUAltAd2BSfabmFN70ffz+QracEkgdDu1JXaHDy7XSziRQXEyRL7WoxCOxGX8ngUYTDY
GJWusK8+DxoPPurnWrpR+NnGzaKrcb/0/Bb6nizElna6y5s89NS24Et3MJerXgSWa3scnLlFEpZx
UxdyJ4upHuaxOMDYpqpnIvh1pNZyS8BB/W1qtFjGRabfRdOnO+xLy3fX+IZ46hFbjZ6Tm+UfgtBi
FPTEfpSuX7QcVQiKnntG0OTf2vmtdKuwnkO+tb8Ij0EiQuZMVys07LrAq789aq/RM5YZZN9eSQRX
WUILaT18vTqOmiX85Z1ozTbggCJ0CnApMHGUUB+Elg7uWxmiAl7oAo9os42XkYxauTYjKcne7Sqa
SNq9XZf3m61go6ipRCYdKFd8chlspIctUVhSk4H/zxAiMiI33If+o/yEljFfEx/wRw1GW2EgTR8p
yXhBjJh3lDyxvQbowtLKi+BzG1h/VAWf6tQLYfF+K0DrNWJCD06OfZv7/mSSVB2JtUsBVuchmNWM
O97xrDYTj6M1w30Kb+t4Ul3aTzBB6CDYeBb+ztMt3H/pOXO/FhNjhlyo2zgttwa/cBvYuOaHmdFC
RcUIdJgWmG+nxSxj4W5MMaSSVvHTa6A71WwzJnXG4r/FkZC5K/WMsu//IEmZXugQiXJlZrS94cGN
4wZYXMoIas8Ei+IMGyCr5VScGpSE8Gv0jk9AEixGN/p1MJGMd4C8mpazf4s5D50Ghw6tbtFPhrbC
ks8lOb6pkI0kQep118CvNmiSZNf0S9rd3ZrfNjS1tK2Eg/ST2251YVmk0YzdqNBmNruUavb7NqU4
obu1TQrd7Elfjgdjg2jh7ot/a5Vw2xIGXp2DDCfXzQIyffSV6WMKk9ZEfNU5ZE+xQjQLZuRY85VT
G2bGi/1B5LvSuFNLU42Ngzxwus/AQES2k3MtXGDa+rDU5e2daJ9QJi+A8CT3JzuB/1CkEaOnkkd+
3meZoijVWp9uD304MPPyoYeR3rHkHshhsVUr5P5x7bFI4AnTvD/jX9pot0JPZPh3dO2Ru0xdY8ru
ayvmHNuWBxdUUCNk3Gx4KvkXTYmRouV/6cSWLjrAuvJaA3uFbKth74L1oFuYJPjHiX/cB6lZpxHF
jC0LfRleR7TIWLRrfU1sQDtZrusdvoroYPJQLn+iJDgG1N+iKasPLqPMWniFtHLWaxaLRmyaxg91
1vqdvle9IkIsGtR+p8hDeh4WzvlTCvcaAVc8caDjJ5kokRt0bf4BTj/X00uhgKiyBaW/SYnZml6v
iCKJ8PCrUh0OhhVwqq+m2jw3NABXAZp8w925jhZ0u7dCRHoPSnyhTUudOXZFJtPCvdK0ojzgTMMV
Rpe0xj1d4zaAL8NxoYhD2wsVz7MHokops/+IRjXqk/k5m0Sc7xQhKzj45Za3eOI5kXvrj9CuHFe7
33gbT/rfWw9HPqEOO3xYqm7mSXlGJIkLzM2FKplkmvaRKZgCrVtmaku/fg/66odFP5rldL4p+QfG
hyV5J+6QD49SO6GkoGq24dw2MYgUQVvv0HFAajs/ahISXLq1PpzzrXD6u1SXWuQBOkY78WrNprHR
GHzGgIhTnmmWDF+PGnP/POfRGxrpf7wxeltVMGSEFpfDvo0Wd2yt4ufIAvGBZ6Yydk1xoTIS5U3v
XUbhpmddg9C8DDqyk5x0fXTej19SP8kAVU7NkJ4XDjuYJlOfCLzBESq7NmZbbsD9SfexeEwg9Dup
woL1fvGMcEBFKhHJiGPaILujk8NKwlmUGHjtP1fof/k7XgTuqQh/pZKIXfBbbXbfH2sCO0uKlxfa
N+ZjCNpsqDccujXXQhf7bTvJLwp7HiTIslg1lJeMowI5uyDC5FYA3ByS81bgRxJpzoYTtikcAXc1
4IpB59Ga34C+A24px8xLHp+o0d79B93k8m4+Cnd1oh3fOAGNV6PyUzOPAVg17COo7Dxpnf2hh/uU
DFSu4UnJNLov5mj6JfE4uSxGjqsmwv0lLA78ryJ4d/RlezuWPuFLV0VA1Bm6HOdy00tkskAsScCx
0Zcgpz9qPzlan7uDjsbH+6f9szaiGcO6zaTcvf/kQNJyWr62m0a4IjXkfufdVBcpfXj7P43vvBtD
9MdYszFr3otFzMAfqdMcYITJ+JwEZFWCKsgLzwR0MEqMWXjkzx/yG/yXjcBNOdmhSxt62EjwX1Z1
1JK7wBbYC/Zkf8fAqC2KLvNajdqSg99/Rsi6x7lvZQ64udOzFtGJPDnes+IqlrdsGQtU5WvwNAC/
TV47XHcyYWg8Pa/rRtDCKww+3EYGIEizjtlqWpjKmUqt9fu64PbVNkfQk5/RI9I6iku1OWFQcYF8
WGtjkccuCmIAD6IJDB1sJvdA9DPP8wDVlDaqzXnWX92Z3uJf0NoO5QfTzwb0Hp6E7wBEQ1onoXKn
jHyjRe7PYcc5eGqyNuotoJNxn0w3PS50zKNnA2BAq2sKAwgFwd8l+beQVWgDn4XEePBtsv/n5fX3
Kf+4NXtZXsC2YRUikL99lE9LLnglsDy9SGw84wDKTYnNOsoU6FrHs3JFTsPF0sesQ65UwS92rC9f
MgyeiuUXaUxvxeBZB3SLjvUrS7jD3JkfiduWKc18zOhprlgjFO7cv2Uc/wVMwPVCg30nKeBpK9ca
rEsBokJX722y1nz0lFRuaLchs1ihq60TVUCSAGXT4PcSSMiw/ycSqSTfrnB9QCtJXzudvqiFbTdH
/LChxTu1drZ1VngoJpldj4KgtNv0oKAM/y6ip2Aa/ajt/7a+qAKSLdWUoy5DPjE6aGg2mddTPTZT
la68192G4p909khFwP0XXSKv0GYbaqcl4jqe0m98+hNKs8saexf6B7dDWK/z4TMycZMDODorReVx
W/pRsjQsNVF7a6UKBob5qeFQdR0enOsuHV8w6WE/h6Mt6g/Id4c4hb+PMtvpVdL191g+2kGC3iNX
KWiYETqFcR0SzDuAzjtkxNTTg1qoLl1Y9Py7MlPX2H3367EFCWGMRx2ttI10tx/pJfv0x9n5eJrA
QEIGTFDt5fkJS5OKYqLiHmVINvlmgYF6H7BeB6PvuKUdVJ057DYsrAkA1X0GHgsmPygjT/ilcXLp
lXmDs13TTwoTIx+vcp4m+g1psvUkRN9m8nEiwV0eeLpY9FachpXbsbhff+MKwzERf9Jnir1WSsHd
y6I5nJIl87i4qBhmbkjiiH4ufZjuPY66AZclfUS8/3epMb+9W/yiLXDeLf4gU0awlzBDnBIE1KFz
4xToW8rxOze7Zww/+Qm0fwxODa3gOJoz5orWZB4QXv/PoQr+bbR1KGIbdEYKH0OM90MA+szFDawA
Pcga7Pr6LXWobAoxvqELjhu/WfpSSmAYaE8zYj+KAXNKM/poA5RHjvgqE7E76MM4arXHIy0LnxXq
dzg0+VNjJEHM8V/vGcObwupCYtrjbL52CgH30dB9PBcts3IQBwxkD3829oDn7VoLdp4V259efQlO
jFJxqAowfY2hdzNTFRhIaKw7Ojep9zI8JrFXQ9ytArNYD/O+8u0Fk0gqZCfxxp5HuJ8J1IbHeJxa
cAJzA0VGtimppAqU8bo6HLWbGV+fhY+5ALO5QHo/RN5DI7LklNYyACZMvP25zAZQ6YUH73DbukBP
V4Uc7q469P7rmJ+huCztfnIUfEIFiJ0DeqOvEsx9nFi1L5QXx8+PGWJFGDopraCt+5O7kirXCTo6
hNFfqqdxKlAUsJZ0+BtiZaQzKGIQ6zjYUsVIDwEfe0yPFPytvnctUyWdLHv8EQCxXKd+TAr+Rmxk
FaxTrPlzz/cR3eocCo7VC/cUJs9Cz/POArnGkC0yphfsv42uG1XzKHwQa8+cE5t5b12+uCwfCOUZ
1svpyNb/bGW8GzbL9PMWKdnkG9UGkYWG6zsrrfxM4gDg3hRXbBH8IC5lhLKyI1fVhnR6NT3sEFMb
zHdGTqOaASS/zEKul19eis6yGSCz/UJOG0OgkITX/mTjX3LKWagmS1r3JyENER9RAuNEcPqpDSMj
MdKCZb3FzdtkqxtnqkIN7gyGVV8utQSxTaDmrlMH35lDoWYWX71PVYOEtm6EVwGqS1dZA6l9Ercy
n7IhLOJ4hfAcYHRwjZSLWboMEx91K03oBSObynt6TC1T3tynRR+zgM6tWUE7Tv/M7M4A6a/hNX1O
t99Eb92vznfhfAYTmBMMOf5Xpdua3yeh+05q0dNif9H27/DoelPpL8v6xFfhW8NOZIUN/kxpvTlS
amD/HmANXRNFybcWDrpYgMd9/SghTk6u4gpJbaKSuw7U4YpXzkJfIQWfVU+lslL+Wr9jnHLf2o/H
ft8Q9GfScRQx/GCTAfGr51/jMRta6kx2JNRkLM2O1yIThpaNqApkgLP4cIPhp/Kn4VaxnBigXcET
RzPwnxXCTW+x9kufHMJj8ixcB5aZqcroP5g2bQXRdk/O78NtvKtKVbgmTNoHrSYVbzio2r1QnXx8
xvGUIPKp/eUzACqpMY1AUkJsMMiU9w/Z8J7cYvd4CuTavDrDT0wvYIzlMyYLCGVv5C56rErjDr0x
DXhh6A/8wLedwnFPc8MS9l1jRhhpPWeEGWo7TYCRtD1zluDh87DTlapTBd96ZOXoLrBQrQAZY9Re
sbTUTYlDa1/vwMNayPRsX5IXpWESwTE3m1Bp8TG7r9YwPwjO252hFUitJySiLirxfMsq72erxMzI
hpfvcfJzx7rBRHyGzcu6Tt/R/Jfor/AV2+vj74IaIB4MeMVCA0PbIQBwepEK8j5OLeEpJ+IzVtoF
5Ub6k1QI3J2iUuXb6o0OJVEdVJBhfKRk2VKGsTizE+oGYGdi5rPBDR3twaH/m0wCWryCV5j/ixEq
h8CXRPxkD0hN+BxTVrB78agF/p0+0mLDwfDcMgNLGMxHCjLlyi8ampNx83swnxuxk46rW4feNZeE
tCQ2/d+ZJFyBZfwPnzGo8Xt3lEyHu2sqDIHZFah7+5QBKbTsBdUjd3N9g07IDY0JeiA3I5MtMQxz
TQBFB7XykixGWatK8SrK5G1F7ljqhduEms/qAiAvDa7idp8SnOrn4oHRpAV2YZOXb6F9ku3lMBBf
z3PYi9QNOEQvOJcH1lyPqhnKAUh0TjlRCtkbkwDlDd+ddkLXy2q+gVnjMxWrKQKkCThq6Pd2ZWYa
vkLdf6WBdNRFdciWhBNkFrzGeElyKoZp/TjaROrCigHqzzRKe84iOav0RaMgOXUvfmIEWWY2bTY1
yKp8kYDJ8bCoH1gOYeaLMzu/C62k2T+GHggmEvq4qqe1mxaViInBxx3PFj1U3u+R5i63KcP82rnY
DfKI5WkD4xjUEE1AKnpDrlYdKvQPfIwUmBgMTQkqxw1PWTFaO2PA4ZvMSZT6vDJk5wbbxzXiKdN5
Iu0hj3LEyAl+Mk0Gp7OzhDr2bKHWicNDCWyK1iy5ONpIyKdVb1/+MAfZvqcIJaKxq4T7vVtSOYwT
mugfduSN/IQCryD5jLOtwnTutpphbPZATKzxSnY/xnpp//ThDTjYw23K+GKmzDcZChcp29v/oO8X
pJN0cRYbhknGM23g72fpCS25Yac1w75i6/63x3x1i8fF+qby1nEYQqY+y3kQpDGfO2sF5LigZSCc
FXp3LGGq5Y04EEnqLnx/+jmgI+SkvqglLepqxbALzJ0kRuZV0TdUBLDp6Daa1awdxoOOdP/ofBJN
uQ7OIbH3VJ4nEGwMgmKRk4fIeKKNc6ZRjtsa+kn6+ctIAoCxUUUPP9F1/lbD4/vIkxLEwJkWQ0dm
GNQfa3U5UINrWcNqiuA2IHEWiSvTUCxO2vP3SEjOXFWqW+dyPLKBPFvAhBCRHcwV500SozjPyZ+H
oxXITZ3kPAvoTU2z1GaBBnlHpGYlIDbhOuazV214+Es3cg+i+hqAz5RnR5Kp3AfIGcaxXqiYpi2i
BmLaEG8Vo3mxdXUz9mIHosSzgCOLR2fv3ZKkVOtJhg7G/rrmhsxklouj7o2Sfg/n8ZhHIaLZ8bF8
brq0EetS4QZc/cyMTgfZgQzVbcxJlMu+XW50J8LDAOCPwDbvKQDzHIG7tKCdLnNn3pVCLK25bjab
oPAiLPyb6KTNIkWd79HV1lPuUJ4G6oNbObpjR006PXILa7X2/uaV62uIhJ5N55D+RKsAxK5k/cWG
tGlsCzRkSeigGm9YCfSV4OYgN9H+JqlXs85tuP09u1p2PFGLJh48PZJRM3lllELDJ1pzE8baJMG2
AGsMsiohT5Q/2KX1pVJx3lK8LEQk9n+B9Qe4KU1r14YwKE2IThrzI3XLeKWKVV4TZ5bmj/9/4X67
ouN1TV67/wHrkKNGIkBm6ydy/J/1kAjxIzKWAgUi77o/C03X6xzkmghPKnAM3vIKcOQYFcmfW6QH
F3uunyWpXl/PiGfgZH1tHbwpUMiwMdQUexzRn0TmzSsAt18Euvhfl6oNI0ItQfKL+BNObtdYXlh4
gayKjORPIrwjgZbBQkQfBMLuk43xfNpqagjQ3eW+V/L/zZBfLuMo7vnq6i2frwQjYxapJDQBg2hm
BjKpgYq81aXgLe5vtC5XXOu6EoHJ6HAQtngw5fx5EANo+wQxlHcYAPes8KWZORfknfeCQTzLA/0G
9qnrIvwmAXEDoCH/btcjppJAmwoJUutjmTG9PWsVH6g0oJEoZ3JzCTuUEmmdYTKT2hKut4vScxqv
mLtbG6g2FfxchU1TJcgUUOY8gbLF9vHHPOu42q6+VNopT84N3Iuuh6TWezD4bdz4eGZf0OMoTB8C
/+spstHPrVI6KgMmHbQ/iLZ9ktX1NTmEJUjPfvMq11pepH+Y3d3ndqXyo1h/8xOE5ZEUQWsPScLN
jwRdbLxzHJLbeo8FUZ9qHNXHa3qTOX3Wb9/crcLOp3fEQ7JOWiVr4R09aiDxOPm106By1ZJ5i4GC
W5QNrDdUuGPyEBKY77LwPMhX7UKGUy/OLWMhLgW29Yvvg0dWmzPuNl78udsJms3TjGM9b9mP6YaI
2if+QcsRpKdwxtGonHOXVoG0sYq4kLuyrtz+RpVybf3f3WjPGGOGcQ50ImQ77NzFMfhcj9sHNGNo
JzxOcWPa9KjGIXWBgQe5Z5Ei/JWdXtnnIRaYM/3uk+kbBYwivbBCxbCi0+pQe5krzvkKCHMJF4lp
gGUrsJPdq7tR+Oyn7YPMvavOqGEYHA8dWVx9emM8cbZzTM7aaIwDuio6Tscv0J5eaOzPzNQIYVQ3
TwM9d4Wl0rf5NiayiZIIFI9HtXldiEbbz6/LyBG1otVtwTJNrFTAeWH0GIkkxLLUfMh1mNSlH55/
XmjrDZ250sUNVjQcVJy+YZ/AxE7C+lwxA1QK9PcvOsdjW1j9bcIfsa/lp2/A/I0vvdDH1gBB/t2O
sixKh7D52kRpW+hUrQCe36Ry0TLi6d0T+4STJ9/Nwrvc+3pLVQrJQp469uemqwujNOsKvfZBY+3k
QdPiekBrcS0GmY9gDFDeGcTZH30nqOneWOSgmbiOGx5tuDutSEwtI7cz5ipLleoo+hWkU0yWtlzj
gvGwZ2mg5E1f3vaqkJTRFBrIwIFAxQthHiXhMU0HJeaRvfzEoEmhQi2wptgePCpadno/dOF4K9JU
4xTzKrNs+vK2jXJ+hLpZUmYZZXRbyk5cRdE925D28iWGwM2yN+vjJJ/MZ82HakRd73ZOU8vIECME
Qq7sIRk+MbXa5BVkWfA6owoTJAlrnUuWMPyDtn/Uu+PvzRoxd7uQF3xjHaKdPJx/eiDZ+43Eb/WX
eVHDKn6RWdWMB2qiqFipeYJQu7UlSu43F+nP6vh0KV2PL+0H0iM0D6wQhRJ+vE/4wTa8fvuWa306
2JgsbtNI1CQOmTDSariMB/Ic1Jzv3z1bFXeplmpxlZic/MZFgZE/DAHxedWeOIFGcfjIK5ovAwTQ
wa/YGeD7VTgtUyfO4z8GxWkryu/lqsDPPZOZAoUNx/a/L5L6RQ8nVzj/RQGHR/L1pug3B5OHTp6l
wRz9bze5GO++RtHDXdPJB8x21f+1LnicF2uzM9IOBlLCl6YEh4q9byRSpXqtxD7kn1gh+G2l3EtU
/aOQs1CPvcyTkznbWYQbHL/AR2rgGIgJ0Uiv6dxatgBQOU7oXdWpL8f0JRhnUM7Dlm1lcMJxH7RC
yj+iaw7xehguJJIvguTcrlbVs4AfrFiqQFFD+Dz43d+QfmIhv7hBTOVHnUXKk1fmwmJ5rE2jPBUc
B65+ricDQGG0s/66tu9ShjLoNYLRw1+CIIVYxBzZFR4hP2oWxmdT4t+zRnZZZt+U9EXN2J0J4KLY
i8Mz//mIvPjvE3Hl7vo8NfF4aNWftnHzk/gggn4c6Pk0gfZy9chhzL1fxG+9d1xY38qrxgWnK8LD
ePk+FFf54zPtTANEY4TKyY78bK3TccSIhfAyxleScPlhWPg8hDc/T3lWzszz28TUCYnmNGpz4h2Y
oNhoLqxbCKDQHUZ0Sl1/gEtmo5JNDjyNmIcIJ+Leltr3M4Zw306b414eJAVfPPvCwQD7Co/z52C0
PLaqdxrKFcuZFg3+AnHT1TkisiwjDvKJ9jSed6aVIePx5BgVWCOWIFyz2iU77VgDNhfeq6s/Ene6
nIcr4EXY3td4LoadbQPdp+u8fUIB1dajWX3rL+mAdmb3UEkB8Twwe/4QsMM7NU6FHva4kdgH097j
dR4/anJZadZSYzKcanTa57gBcre7RZBi8qYWzMjak3sSEuawle6CGjAQOZ3t4XEwbVk7YELCgAyy
3oKW3SRa99syzhtCI20jCc7aXecbV1/wECCw4OjZQIMC3IyPSqShUHEjDh/kqfytWidQJ6vbYgZz
NPdY6x6xPyG+OP5vjqW7LyNXHfSghbPlOR+bMpDBwKDg7uwUcx/KsxysR65TaWnMn5ollIBdzjrP
zi2QTwzfBEJQyNEb7Ht8xjz+KI+NyGjukTMHegjD2ArIHkmE53v4ysGtTTkJh4Qy6JYjp1pP3AQy
53a+59Xsa4Yxi7C9u0uzhusyBh4sPzn3aoCB2ss3svr1eSaMyWzKaRUmwsOT28kxXBmn8i9NCtXM
W6jeSzHR8mgEANYZrARlyxM3kvA7trS6hgF1YI5q1kqNG2HKCsIYFBG9NUs09dHCaUjon0+73dTH
kl87UJN6gxBOHZrz7lkDwIpXAPVhgixjV8ElSle3FUgT35aHfdE58tvzvbANkx9dUujOOsGE+flo
uhj9aKfbaAlcWCqIijJDjnGBS+LnriSjfnTodoKOwLyOzIVJ2kEfg4OaJ+DTdYJw/EDATWiolOw4
Nec4O2MP67lMuo/p9FnRwxUmDJz5AqPPM/FH3JdZNAGLQqzYWnOPkAqAsneauLsZ5FKU+JDK1Oeh
+ap9C1ainTLDK6JP3erw4jLGobp85YWkjBaSCrZL2oqf5gwEIIJjJ/Tm0Rqu2mQkN+KoYdC99Ku7
s/Gjqa57V+6BX+6MmpQ/1jyYWGUgvHsZK4jaldGRjvVJQZRA9OGVv2//mMOj2QL2gx4UAvikgyER
oDW+4TNueyJ8dGghGw4KtaAuTml5zS3nnLHRusBnRJ5+XdtfE6HxAPjnJlGjAxlLrfxI9jXpKB8w
vYc2aYzO/XXJX5o7+y1pveGW+a79+yImCK5j/M+gFYH17Ug3SDDog8UXa9fmaUjgQwwQYWJrYmoz
6AqNFn14Wu/JzWqAVpvasxEwZNgusx/+CUdnQ65udttXU3DgKZ8OKG1zbNbHh7HzK9EPDls7wOmv
gJVId0QGXHsFAIOSEkkV5TlHAcgffzDp3GmEiiHv/IG9Oii2rNwK/EMXBw8igHlEFxR6pvPKN2mS
eXGxtgAgDbf/23ujhEpTKS6Ux7APOFE+rUxKko21EvJaym/ZpKNpW2LtrAZOacuu+IG7IdYiimF5
fXa83Z5m1JgMG4myAAKcL4bUC9sn834fSQE7Qwqwm2UvXpE8zADPkHknaUMpEks17CeLXFB4NI+j
WAAeWIdpvn7uboMMMYMEN2TxDaSzSz6YdIZPzfbOtQta4VKIX0PdE6A511D5TPXmBzbkwbOro0b5
9vk4hhlFbiVZCLHyaGP7wbVXLlEwrzzpmtxJK7wQi//C0Qe/N9m6tsy9VVN0w9pp0hxi1s90L/RG
E96pzn5sF5HiBf4X01O9G0mb7rQvxhYxSiWjKmM7/WjGN8TJlskn/nzpMyFcta2VVnGgNyU7GI9V
80mF5rcfmsoZkaKIXY1NM1+TKZ95hBB0TM8cA1ilZMR7kr8h3KmvT67e4jVe88J1bBK0gDE3m+PE
Wd3wA25lE3IuydDfO8RqxA9AWi2bc8wMrDqQTjSUqtUsiB26UFgluBUzpHcs/s8+0QjpzS0ADOUX
mO3hO9KRgQhMWNqjShN8o1vyydf+dzlarFRYQ9qlQpMPyZo0Crm9hOFbOJ9Gi4hu3IrB5dKu/zYR
zkJRJOKHVPLYsZTByBgjJgQSd+q7ED+mZ1U1HSIzHEibYgf6Ky7xQZeas+R3QRb+mBFWgTgGnZvU
btJxphTdyO7b1Cn2w6IlCL20MCmrDV4/9YgC7Boo97OksoYeXtwB0R3A9GqY4yJP7DvohZFe4P5w
LytbQw0i/xhpmz0tm0elfmplhrhwVprFZZ2+NgUk+q7WAd3+sDBhxVAUf8J9IysaSLes7hccvfny
kswk+HnX5vyZrGCNY8SgEKwMT0bjR5TSzmKT9NevUD2/+NI1l8b2TYnM0CSSKw+z/mbF0bV/0BEI
sfibwVSQQxxqv6uF0HsnkelQQ9ckxlnbrYpJ1aSMgaeUdGc0+9wo0MhAlCNUhsJBzwncZRPf0Vyh
SLgyfpbsDnSRnJf/DDf2NkU72aqUWeEGPhHd9RIyCZvM+mCXhJXSZht+lLXAjdl31bpw236H3/BW
T23l25/TDdR68EtfwNXyH8+A9nfaBYxnFuVq4R3PFfhDTF9YXamxOv0LQ+8E4KmEFaYXbf02tw6i
m5nQAhoMMgHfKPvzWGk0wfd0QVQUVk1xsFEbmaDoslGsEitAzrqnUDhY5jN1R+fQXxd+SeuWWG6C
XQOFYWX9028LMUOVjJ8a0P6YKtVnKLlN4y16yBM14VGVaQtqgnbgzvqssdZG0hiRbf5xaWG9m7i8
NkpwjbC/OxVf/Ti4l8CJZky5puR7AKeiYl+jrAn6ZbeHUwpZNOz4hpJayitleL/fjS25dB4QvJuA
5VzcZHeL1tMs/DDuUWkgYZ1hbh9bpIuZY6jfshLq/fkUZjnVUHLpk8we54T0b6+peffXaunzTBzU
jVH3ULw1QY72GpMODVB+8XeFIoCa0HA6HCsP/Pzl+PFs2UM0Ji5U9VUfsHzDEe4tiyTmrxbMPwkg
ebNg8JC/e8+7NDP9tTLBTcdDvPSezYNlAHybBT2A8WR2chVGAvirsEuqLURdCfsPUgixvBt2b1vM
odrzJch/UeWdQdZAZ+vIybIe3hyU9zdqjIKajw2pPCf7n7SixwTtSpOyqllWoj1TRS5N1WJp7G9G
nEKYo7ySseOR77W081npWa0+PTfUaHR7U9LCT2JQjVv23NjS7l2W/aXtjTUUn+43iSRTDc8nyx2X
LcDxox2ovJ3p8NTa4K3YW/AiZUvn28aZezkGq1VTJYfbFEOxwNp3RhMoSNtM21YQagaypyLkVvis
E5jPO11mV0lOFkddmZRalc9hJy0ME9NTBMKWGRUxn39QJKrC8k6SV93SoNoLLyQfTnKvk0LHrVL0
rVLR9/xiFp7aTSV+Qsn++2WMZPQFo6U75yBiwB+/v8t1qWLZZMpmdjdL8yRemiZIzvSiRv/vxiF+
Ilr7TlT5336Rw561OjOioEpPz/qxr4qhX5aFxpdFKDn2dMVvuZh7t/5wWQ52EdORicQp9Y5OMhzH
qx5BD0ghN4u7yt14Fhs+1GHGnlruV4kXYAaqF8FwbtmJFaHqzHc8/QZRYd46wHCT2OeBwDRDUXLK
E+epl5wPYkaMzB3h90M6orx517pfGE07x4iZA38n7qtmMIplRaYW7drZweKYTdddSrNx/Huo23t7
mLJ42CTAzMYgxsIAJSG6Yk0KU14hdhNzPRWFVkmVfllIGH6bTsXlPlIGSllePEUiYFPYZ52mNJCr
V4i1p0GI/ZkFK+jDPC9J0Y+6e3k7lv897fKql4BvRgTHCVsvjULnmuVXwypobdHlSPaUcgwlE3ly
pUV3Cz1tEfP6HILdzGYh4mZxiNRHQv+7SGYwKgiAdDxaND/9PoxVVI7cZnFUX88GVuULQMfE4ntp
O+bv2R6FbpXKu/19969m3WZJmQrXUf3sus4IOBbW3rhYXaUaWbIDKdUrByTLgv3/gqcHOZSndxd7
byD+0lmheHr3dAArhoJqCn6n2sfKzWD4iOSkv1b0QGxsxE8vsdqI9/xF63U2TgfAsK2UJ8BSQlbw
PItBd2ncwf4aPb9Mpx9/FFkJJYfY8dIOtC5Q7G7njVfdo9p6yALW0g1AeTSwCZmYgNaPmYTMS+zx
2RWULR4LtK5WcLI0V+VsZbA0kKLZgdUVHOi3hHOaqQKix4iA6iHkU9ENduqSJ9MvG9feOOEDnrgO
xRi1yOHC6tDGboSU+pzKIqVYk5oEZXb3rDBbeN/VP+iIVhqKbvZeOoJjIj4//bDLCqsY6oKLs0Nz
tnUJJkd6246giP1rVs3U8XBAdIcT/Uj8d/vWqn5bP6HGMIAq9DSXu8lD1hGERhMcbv9wVhxI9+qA
dooBesicsE+xkWTwcmep0A7W5iEfaa2h3ksVgsQau/obkgu3Tf1v5M8LVJmK/xCy0dGawYM3O4F5
I/rRthxafY7O/gbikAys0NuVpygDBFB5QRrBV6Z50Bdhpmhwx8zVJtcRCMCrbRTYURShJ8Y8L7aW
Qn5lzSstDnMLvXBdqoR8ZNOsau5x4DYaqPaafFh/OYLkIuk7nx14yKhFEYO1ZyinMNzvMtGf0pLV
OWiYHbltCYzjfGoBxtb0EFTJwMjKChezXSP/4hStB7hMOq9nMQ56KC7e5asuNqN1mmoASCt1iZM/
KcW+jVXXHp7J9LOws4S5qmFms8VlFqSjDHWEpYjKuvt6x/v/4EVfQp+nYSL+WUxq+uDKk+KrQoUO
6SYg7GJP+gIgJ5AkvmZ496qbk79KhnjKUiVr6K+zauI0wgig8qSMKnDmtzkkgNqLozkCYdc59t9z
qIEHXMYpQm9FgKYbyI6Q8vZfxOX9bPeLC/IDcLvvadUuDuwpk7rYsK1WPuKeQnPe+Yufjbtv3dXz
ecmq7KZ8zfmBso8M8UCYfu+vWrDG6bP4mabLwv5WvrB8KbbknOWoBlYZxTN9gkhvaCZ0MEjx3IVB
S0whazlcT5DSEd+ItRApENjwfuush0zgRAhiYXQk3gTPChg8H/EnNiK1dEQIeSGjCTIF2MuQADXX
3R08/5HOAJJP0F2wvXC5GRx4sq6JzgrL83xU7rDLbbY22PUJx3/T7P7Ovf2rjfiOKyUg5/B2zJl7
LcpvlhqVkLQImZu4NtvMf+DCUkEm1XJpQV9lR3wSRBvObdppZDvv3CUPn2DBAwBpiZuU8xi+iLD0
N0DN0gaQIVbF1Nb1uLXH+HlimYYnt+knwTgi4D8kq1IOHRxIWdY+rZg58TXG8jkpd6pBvgb+TdSS
O6DqSygXufyLfrqHgqYmy9mE2hS5PwJQfIr4zcqFgWmWzfuKHocq/1Dc/RlFpyTOlEC9tpMQ5mtg
VCn4bUkzskNIiRJ3TP4oK9ixaQ1mdrp6dCrGsFKIWKZt7X9MpGNFFhVnT85q9KnKYrzT5EIb+0zR
kI2BH2/7AFq8YFRKNSbtQLbbDlphwl7SZbdq2qJB8OllmzhZbX5f7Vjm1dSmtkbIkeCdW754uJ9t
lIhu2FNg5oZq7wNCH9ifJuKZqLpQCyAnikMYErbLh8jzD5nXoiOII8qVp67w0T/K6jhNB1o1/RiA
VCJOren6it/zwh9exQovM7cCCzEbfZxIkeKltl2saIX3ppXuAnYSERhxKsLbQZ6AAZYyfpJzgpAw
nHjxybSrBZy5Ue8x5FnjBlVFHLtvedGxES0wwKCrJhi3jH02Mx+gipdjdgp+T0CsAZREuuCZt5mM
Oi4CaJvsM0x8m53UUbFrelsgDS9h3mHHo09t9cC7pDY1Tf9YdTrptfJAutiK0mcG0s0XN4AAt8UE
hy01vSSI2wmzcHXpFNK4P/LgvdQ1lZn8zMdFk9AIuoEoycVgr8FdECUMQpx0+E17Dk4kHnaGWAG7
KFdH047nsLEwQrRFHXEclEj2kUpawE0QK20BdE/hbER02j/fN1VJh7ABFRLH9r56wlxV9bgfNtQ6
+bgM/4dM74XDTNW0utIguwhb1gNcIY3Af5VbtndiEla9DOumI+C/xKA1tLwWi4r/Zqin8rSVgkLj
T425gUqrWMRFDyPPKKKGevAAoRYrnznAAs/MaAIh0/bS71dmbQ1pDyLjkGbGoIGILInsuGfzjuHp
/6nbl8uJ7yGtb0acAd6EZ+kgW10cNvmg1NKC0pPVQEMxm5oWqghiZXksMDCDbCbEPohjwrkDQfHp
lVr47wJ2tBYViMGa3gMz6SQIsixAmP+EfRt4E6GP2UZo8KZrm7iK60HNIuOXjYSFho1DiOCGDSOx
bV4vsbR5HWRKdIL1+uxvxNYyrHJWs74LnbDkVGGGGeRNrNpXEZC4rOKULjmk5+uy65zJS8weKBe8
fZIfkGz3XY7REuh/mPBgIuge/bxxgtS3fTKijzipeRvAVIfg0Dduct5EXRV6Tpa6QfxYDH+2fgB9
lYPge7ElV4xIQNuSB/jfmyMJh+86uQ5QobemE+2jINPeQZUcQwlQ3nSlsE3TXLpKcqdQLibE4iG2
Yk8/vfmPysOyIOMLoqySaE6axXshpYOE76hfeGoXbQ9k93MacnU9dHPDUhZTs2m4BXPvYJam+mUL
GcL736Wkspd7FjRYP6afthbWW278TaeTsLiv+IOv+c8FFkrWy9Bdwv46jyWx2Nv90nenQZgaOWbQ
65yVQLjD6GoA1YawrK11Yf3Manjse1QqJqW7HvcE1UxFwyCddC4iaOzFTmNgGjvXY23y0qKADcLt
IcMrBNoD3gLrbSWSI7OoDaCHN5SjZouJc6IDu7YDZhmiobrUXIuv98G44KNjQbtEH7MbwIZTkB5i
M34tXN+rTiA8+kKN9BcbUCn3qjFKbRzcXRXy10WgOMwjVoCBMQjVIW2ERtWShDffjkoRMTSob7w2
sFQt6vV9E/3spUsQWFm20YVb2sLeUfqbevuhhPPtWpysCInUYWWFP+Zy1IYuQFFdVSOBaCXBgDEz
eF8wh9/2OXVz45uhhYP7u1KsWP3nme5K/T9oYuaCIt40oUtqzmzR5pV4uDzl8Vr4dhoRXZfEmu7e
aWpi/Z3D8qRmVeaw1Qa5qz6QowICRLFa4iYWvYtfccZl/D0JCTqvQaqs7mQ9r2dURit2mZorI9UP
WA4djp3c2NKcZZAzLqoA1bnBODbnMLQ7INP67Iq9gDX8abgdFniAv91QtdkZgvWr4/z65/v1obFQ
ncyfO6IGeLYCeFCGcz+UbHEuX6yij3lz6eF+UMGTp7XDu5Yva4/5RLcPzUSvYXTXlWLuSlkySuTd
siYJqd8M2okqzvSKeeBcIYYd7FnKawcGP6MQeGzU/XdYivfzsFwgTOgMVcg1CqOyp2BeVcSd4M5z
p4GdZWx4c6LrBG9R3FgfQbO1EnuBrDR6NjWN0NMpmPPPSXJBrJNb81DhZ+tPPpxkd32+K8cTXDPG
cPLuLJOyo47R4sdb6mbK9yLwy8vp72F+UWYstaYKmSGd/qnxdnqdFIvoRwtq181SStYZxo1bTAWb
NBWKB/PqJ0LDxtzDvOLS6kHS4n0ySyw2PdnBOB0cHV6TvwwNJupkv26+ics42LkwhWZ8sUtZO6jj
lUJxBNuq1TE/eKdAD3TQ+dybJ8pnG8+wdwqp0VhL89fUS+6wO1qJrXnUGNvU6pHIL7BBEUZAOrwN
hQbKTZmvWwjxOHuawnFw+ArBrExPXRwGr5T6XWWFhs9nIzTLDBbEzV0ziijwRX2YS/VxRBLk34Oz
VfTeIlpgKXd8VdvuRUnvl3uzulozfe9aqbbrnFSYNDFebhpYGB32OSwLez4b2zS7PXEPX/zCze1S
cgoMoNF6IoP4CqFUWdrb+4RGqMerrN/PgN3ZSN8RgRyqDIjVdY9IK6+t9zftcRqZGrTnkN1it2w2
9iGW6bJd9Tklv5xS8zG7S9qKVw6P2rcClh2AK41MELdJuQq3x89D7Xroxnk3N9GLg++6URGj69Ba
5aKWzKQMw1YzSyEzhtsVlLQjfe+3ooIBrma/Zx0939MfivcPN722QOtd65IXRn6NZ1NIqXS/gXIh
Kha+97TuUNo0g3+qzQYuKstXPaV1/yjLmB3wPiKY2KMolt6u9smTJvXGY2rNk6pZjywjFfMKIwoP
DD0woV43o4RrI0XxwOjr+Jv/UKK31YsdMtQs6wiMb1mTgKU0M5lW13kRtYShowoLW9u0mAbtVB7p
c5TVTTBc2X/3crgYxhiEakvvN4P4YjViJENA/U8FfR26rdo/trySLq4/lxtXpzg3B39yhWMRvte7
CF0wojWOxdGxTJB5QUWyGiCes/Wfno4Gv4X3S+KgI3sX6qDxJQU01wVhpKNGBFkzNJkuf/IBwqxl
+yWf5tslVheg0HOczwKlU14osh/GyU/HUCU0EUm7LpPiK0lNrtTJ0l55oeOUUh0MtWBfjHKW2TnD
ytsfn2xlRVoh/+UX5Jr0G45WWIAIpApZ2BlfCauOvgrpVNNnMKaelDb+eBP3mfARe52mAAgGC1A7
lOvCJ7fFXljYjmnuGYfrJKBGyHu6lhWKs1YuXG5qXIUsPvvCkhcnao9Xz3YX9Xsi3+o5Vdb5FxKJ
vjXAGYkcxTNLA+DAtDZ4zehtzNdPu5vxvhGsLA10Ix24+QImlwTogqsdgKDsXR5Rvj1cGg+pF1Cx
65Uphe+OrnSF6BES3E/BkyxawHW5RgB1OfhEhMX/BWWT6uKkt7n1WH0lvmbGlbS1/VmWGax3w1KF
DMs8p8vIBA2r/2A/WFHgszPV+T26EvcQCR1rZ9vf9fsK5nAWuhlFKdz0JpKozAzJoFNN7HEy3Y3j
TyKXXdo+n+9qjL0eyxbNyFtaP2U9lpsUiPeu7liRfK4eO/0GChwCyeg5z7zYpafOB+kiFEHKgZXu
OUUTxNbUxc71Uukx0kxvT1AOIXEOn+P/jPJtAUS/1uCYHI5GT4dxOBoTaaVvOnw7jzy+k9PDD2fr
8dMgyWAdMQ+6SspBUELxC1Qx2dZ9R7xYQ81Iwhg9ML7gMdBQ8hyPlrzSZ0iw6/nj347qFSmlxKp9
1WBPRVhQdAN53YEH2OSkVP4SkdAg0EWLBKfsZZKjg9sJxNvR1XcY/DfaDmRng52xUsT2T1SYxmXg
lhpSivLsvbd09RsCUvO+bXKSrGaYBtJX/13Nltaof8RD89pzd9slOaUfBsCP45f0jcwj9ERRS2bL
qteb14y2MVCMuXDYeafvd417xph9ZYsMcvH2kzf2XthZewlOjSmx+SSoqSo7baqkqc8qLITOvZhY
RJOB8oViGxtjstNVDqrcd2/ZyXjIi/ZzS3rESdFfqQGU/6WLJDVwB+vaVCeAJAIHrIxYeTOqFJNF
F8lylhoy82OPpev0hZdG6FKFbDgJ+A4M3H0rGMQ0XOIDNv3+HfQoaMjFDrKzc/Xzeza5QvIMTgao
rY5RK2OiEOteQsReALN68eYvXK8/ElaTDsKg908sEQVUNztyXKG8tifEMChPslc3Oj663zIIymTR
X6MakDoW+DArCAl+BuMniIW7uLTmW5wWxHJyUICazrYZyEHDPo1Etoiu+6QkxQ46acYzfpDZyiaA
/MSi/eQrxI7gkw+MbZ2ciIFX791qXbJZdlkyATrJmjK70wXYd2CT0F+agpsu8ypyu7+clLtuG4v+
tthpCG8hDyWkJqNoIu7Ng6IXs/lA2J+FhERAvWi4AXs7rRQnfxmttaDfBS/CA6G8YzZd3rRnNFew
aSgxJ59GVxqBQBG9jNEpIlpVcmZtYVzBmUGdBTLumVqeedconHdluxrSkHWl6tnJsgjMNxZINoua
QrtQhH5nMlS0uZ/n5orZERONsDIrutnFQbg2VWVdSvzlG8/Ex4kcIgFeFVUhB4H6SrAJ0+vui9AH
/vfWY41GKM07E24FsqS5tDlxE7VGXRefRcHmXK2bQ23Ck4fHJs1xN8zZWq67mpImGLiqQpfOIZ1D
3TFZeeRhVKjE04A4MKurTQl6zi6jRa4xvc32R/yM6T+YhbaQ5xdWZnvNq+Hnr3J3CnOxvC4mXCSt
BSp4D4FPHzJ88X726d7zMjRAQSQWmav8m7SwunzJszkKqrTkFWZ/FLbU6TOyIdgZjb0ugiMIXE2w
/5RBpmcIfnfMA0kq24nHjdPmW68//qIhCzaWY/Xj5fVE8IVqv8YPQBJeAGdFLCefZQZ5KsBl4tLH
ZKgWYrz9SY90x4dLktpg9m/VYDMItlTIYU3OTAhKZW2Gn7KIc9ILJnO3U8TZ6qygp3IxhyaoKpPN
A3Vfs1jojjk940hf4nbMGmOJEnTC7HKKGd9bBpTY0YmgpfKNZMTGrqgQBYWJAeNTimk2Sk/qshPk
uJYrkHgsonrkOCpPo5vVNMa2HR0MZ/Ea/AOwiMCAlNxfDUlv3FLzgXUd9/HxozjyURCHDdKQqSfp
uZqflZHZZWGsQuATE9v8IxAH3LnXI/1ntyl1+stPWnzJv8ArS8f9o/KLz0lq9+DvGN5+05VbrGHq
o58c5AG7tpEzMTLh5Wo9LgM9lnKfJ0Zpte4dE2HFrK1NrA5XNIUys2fnMzOtqpzNahrLLLKtnio5
bShHlpen40OT0rrIPr0p4xOQCubLZ+JHeIgd9DdzLZKIAE1MhOaleDPLdJG30rmvFufNfvfIvzS2
5q67ChfX76CVymKw1tpapgQbN2PQaNXMTsgDZYDup2OOf1L5BOPXni5o9+ccCneldUCoPuYXJtE2
DEGsWifcEqadnM9qJTQduyFv4J7fg1j3lttcJqf7u+X6+SsvWVD4M/crit2GArLk8wMdr7zcFqRt
hzbvaOAc6J2BFy5drvYxkSWWDEULJ2OTfDjOH+buP8jgxZCioTrdBc65BUO7eh/bXKSkTh2R79Dh
wxLwY5Xjz1RylVq/UGtloNqULJbEL90xQapIOerm6BxOyhMn0gJmM/x0oB0ySBHr5CE+olxo3LqN
P09iO9CdJGJ4Vsje8BMi4xHMTvPNO2nh9U4CBPfBHmWnRnRKzOI9wDj4e3rNhW9UUMkV7lGFXZSw
8VGrbXB9OoOAyWz4DuPxglkDO/uo47/ZpHT9BuH8FeMqC9R3y3YWd/icmnGfgpY2fUM+lFrteV4p
R4ff8GKqdpHAVKikBtz+YgMA0D5IM9z9DZF6Ax+Gm8LplnMAarNlFxAMhvMVeMuRgEcNbBvTbGYG
qjv5TXpw41un94NNRiVqeKnROh5EdeacjQmu8ooim3r3YIMDYwBXT20ydY8qAAPFTGKuC7Q9eiDx
t80Ha3IMIO6qu2C8VCgQk3wMliEB4gCGBeuKoPi0ONUtQKB5JnfEwvbN6jWGDZpcgw39G9pnsArg
vkJfwqQuEuB9AHKafMWg9hRFmr0e6CAD0hQymap8XefA5+TQeuVh4JaD6y0Xa29g4QDheKMydv92
C9X0ct2RM8PPHIEX+DDks+SSL4Kj1idPb+pLeaaMCr2rKveZ/UGFwjo4IbGqYb0tBvyr2cO8SgHY
+GhhzeWIcKI7Zn0wWdf3OBwyIH32C3UMIJ2v/yb9NXW0uMzA6jaj2LTQsaaX+QTjMYrR8TXEIQyE
SAF/1ybxjeJd1QkYmhw2yjpCxtgnfGuGWXQoTVH134VKvzAXx85FLhMDUmJ6qAq9C95oFI9Xr/nV
wRAu4L3m1m/q1PLFUkCQgeeBd4IqwvpJS5y2dGc/aNUoSHZ801umRotcjcmpR1KyY52a+hl0GGXi
XgD8myk5rEDLFhmamWBxmNQJ3m10zwIXDxzeYRh8s9BOQ5LuLFRvVwtYY1Eg7nV4wm0YrdD4k1U0
uD8Mm6W+1fJhHfDcKZ6Ko5d/4ovkvTFu35xQU7xyCjMMnYF6gnuobjMjkxShC6tQV3d2t+nhF8Pc
bcec6Lq1fNIBTd3+Rr2043Pz4uGE0PMyEC3PAGOqJ14Nuh3eUu635+nrDwjQmCmWHXlzbWcqidBl
DgseX+kSrIKiPQv0xZubt3/I0I6yeRMwX4oQmo6WfyX9l1hTnBtuy6SrlaqIhlAusd/V/QKH01ss
BPhMmQK6YisO+Dt8wzlRkgiqNl/shThH+KxAef7xjQVeS2Vb/cd8hQuLkibXbm853NrZmrAteT0c
79kvwSHWOo1RkcoHhczHq3iwq5R7LNtvgHFSFUXCInj1jVL6idC73b6UfwkKZUr1f+ukAQlDThwG
jp4nK8k0zt8EOjp33Us9n2zh3vs3JSDksONBt9+pke6/1WVWyS4xFP5HuToMizalnNwtT9kd1jJo
w2CPHcz3P9OfetU5BsxiuUyXatVaBH5ezFgBhKbZPzxZC3COrShoOTyZL5NZqx+H6wgzDaMuUdf+
7LsNF3blhNPhxNBf2KiS94BIKOO0sDbFYdvTF5nNS3tKyzoQWEHWAD60lhqWp2myFNFq6/+2DcoB
L5Fn8YZyyvy7zMWJ/BeMzvgYwyS39QiwBrw+ZMP5dKgGbJ392ugCRFQQZnGlv1McshASLJ/bEqHk
LCsZXE+AzE1Q4K/xFBfachyQwXpvnM4ZgBPU7KlpkXa1lAUk2v8BuyxceRTk0tPvGhK2qyzGPfND
hzO2V4EQ8fkKov4jjX214e6k8sG+L0HyRw4Wqdv1MugWiV6xfrtP/u+S+OS5TW4eX9zwYa6538GJ
p8G7seM63VkH06eam+hc5ikuqTobS+0f5HYt17ld5L96QFH642TTh478/kLFYB/Mq2gmb44SUReL
hYKk8b4F0yBRBfBTgCh7iFkH4YGMEWlq5uwyzhjlBREJGHMqKE/jxvjRVDISCJ8/yDvJyka31uhD
Wg75rhKuqRrUJUdlr554Df54W8UuaxkLQ8JEvAtcnoX1cwOw5iS6vLJZwP1w+FJ0201vBoQs1z6X
ggkXDSsCvq9Ea7KYHWrugm0RlOPcfjULnOzYBBnyDfWflLjj2hL14mrUqj4wDYkoVyAX8kL4rqgC
DaANy+eMfqqoY60ogQFcd1SbOp+it7QzcmzMSju1cFVzoJei6MrDqbIm3jglJPJ3j9OEkPo1/HNo
GWQ0wK9YPHs2SUwOOauBiXGuvzrLS4XA3WejkWzBZLmixSXw/0ghJfpOuT2AJIQ4j3K5h48LAal0
vEOHlGRk4JC8fuj83Nz9aiVmh9oN2Qg8pdV6CTaApojVE3aedQrSi+yW9vKS2Q4r8kbofc74G6Ja
wccQIxtLF99XC/SedSaFs25v50SKstpfX5PAtOkGXpb4dI/tKlgA5t3P7Up+kTx3hkItkVq6fg25
N6VOiZRhlbHJoc1YsLvkW3ejQ37Clt0YI51uNAfHg/ijLCyWfAkaXesy2pw947u9VHf5PZARg+ni
bHYClp97EtBgDIY7+emsNX9Nh7Wv1iCL21zAAMGmiF6GO7JzPMIUeFqMnRmKko6uzpU1fQXhNyGS
G4qsOS9CeTPaE4CF4SHKpW0QXZe6nWwxeOu375QW46QqMKGCiwo48O//gT0WlxW10JO+maRdzsgN
GADWC21JLVbWPmv5xfKgMwddzN0ZnW2PcakwA8M3gTG3zkoJVYI9LnG6ff4qOyE/q9dV9Pwx/bB8
XJwhrAUyoIhjdHzom/EoitgkO4aK+YB+mFGIajhyEXqbeXIEckqPfGhFsfYtRpnSgx2hbxC11vVa
EYM+flpr2gNVpkLi0uUEhejtnPhIzTmN8agC+wcD+qM/MhX2a31lvBOFOlYrD1XYqtlARFrsJ/Mj
UoGS2iv5QbivDBQtvmzaHYSJFhiiouBy/zUy+8COjT5X7ibKdWDaD6CMwgEDH8B/foy2JsuZ/nCd
6T2ziP4YcBnjvYnPabW+nHfhQjUJBkG8Q8ivx1VZQUe/HI9zDLxgL2Inwdel+jofVKfgjtPRtyWB
bji2ZY3Fvv6BN6FaZdnOexGdpVxQ/+V+t8ECTpsWhYLX++GPRohV9b5sDYf44YH3X1xqlt4uD4YB
4YAiSET+8tcq1QXls/qHB+Td+Q9v966BIZpkCnt+GWpclt39+YyQF1Imft6Fyzp0hAxVJbzYaa7u
XOlHFiAiwjzhblhjCpAFCqsnZNG+qu5+xa6Y6ZydISZ5nBmiCmwkZdmeNOQmaXbsf6IwTrQbLqAx
BPabaZ/BRSmBd3s6pjDGedsh7xSvtaK2K7YjJpOT2A7p/yHSMn/grn1LH7ZeGON42PZsOkfTnvts
2vSIOQ1GGoVabSghWPRO4DZU5kD7Mfh11oIgxJXmA8QHE1euhig8MZQ/ojPHuRTxYtdMqYvOotLh
wH+nOUSzXOAArs33gv0VRIic0Bul9kQSGDzzoSh7YT0GlU32YWgHTetBiJUDKNCivzhdv8aKookJ
gb3YjSNfJo/z/Rwhm6eqrlY5n4uNjnDH1tVRWqbxcCCyRLfpVDC2zcUOUsr/XEcmsVvEAlTkIwdM
2rumYoVu9YbSiQ5u0nPMc1t1BJ6NfBueR3dfLZas6zL5G/4H/kf6IjTZDvy7ZruPqdj48wuLiiqp
axi0qFusa9HSL8ajFOwWgFA3LOCdrTQy4dG6Ky8GcXNmkouAu7tcOEEbaS+R+Qg0RkpL9z3MIOfq
WZUVT4Rm66yx4QLRrLNx0Z86WPGrJQlyiE4JWQmHfMv6uAVLDVzXf8+nPmriHL4dOBOrSsZjR5kd
YgLV78XWE+zcXEsQwx6BSpuMjpT69N81Wra4bTm/4fsMnrcqwHSFOWio3P+Cw5aO9dhiRlbKp0mN
wOWVpPT3brI6EjTiRYn+ncc4K10Q+OLLZZo+GpaEo2OOXV9W35nYXqfCWpGZh33dT34kdSFTz7ms
xLYaZzyF4SNSlJCyOZRCciq8sDQNFMcMfbbhrnk2FHG59GMEfc8aqvyKe4oRjWQ3S6nUlejOcC7z
1QlidiuZE9193wQwfRflRMyEXdGn8BVhKTqPhIx+ffHCnX/fezdb/PTO4eSZ0BHKtZQh23h38iMH
wNlUDAyTevb5Ly/rXLn7+u/fGC52S9uAQzy9VYQxmk2aaG7o8cw5aPCDQEuvQ8D4hsO8Tof7S8ym
n92vmYSzwUUpiQQ7oFbcJ2fQRaOJZCNRxbId7QpBQM/YuG3UArk4VSL2Q6X08jY7/YCg/fSDcdja
UVrhE457c6kebChbHO5av7Yaas0+QnDoFuIGLvJINU1sydSpUqcPJ/IcpX0hryDQUXu+Mb/6puLE
v90AVKbXwRTrwUIOzIWJf1VIz+O9U01iqFQBgoYCSTlu1dLlfgOYqiFdRyIbLpwey2WpxvNadNN1
OTLv31jMisLShucSjhv7wm950//6+gDj5h+UQfdZ01gGTaSfPvmE85WpCDis4cxDBMUSqh+cMyHS
GaffQ6ieAqDIMwz9MNaXw/TaU708/JCfY3pBEA8lObA/YaF/uy63UR715i/DO2K+4f2cTezbq+Kb
SaREEW7c2vsep5Kv3pa9hVuvEaWKnzHeir6++Bv8+NzJ0gJ9M/MjRqfWI0LDEPLkV+oWFW0fWALN
IQlh6x5nANAVfcs7Uu5tPc+9JG1DzPkvWDcljS7MWKl6IfnP76iSi6s79EKOnOTjPHqBJDU60uEJ
urcALxb0VcoQDLOVMhih9TAaXE032SVWO3ONGe4M//6ecl3LT6BDvwsmywLaHLzOJmDpZvi68P//
HulsGLttCMBM1Tp2JuSrHMJVVMW36aFVckxQsbmybVrHzE83OP878KnHsBcUVufVUCKs4ch8IZxs
UYj0KGDLFrznInzlfceA6pCHuNTcb878dLs+v0KWIiPfEQAUneaLF/xShbXr8kDwUIJizTTexPgl
lrRmkNZGmmc3GAKw6Kgwq8Rq0/k1bKpTu4Y6pfqLX9Lf6bqV4Ez9jT+GXFPsvVBQQbPPOwyltDww
LkE6VAY6Ik6+vOPvkQmX8MZooN483KTVFIMNZIKyka0BcuGO4jQX7sMLW3ekItS6KxDVfPpkfRxh
TAZajBy7sMJvjw35wRI9u9waKIv1Ia42hWJ2i/wu/z1TLJQqgZ7sIiNnqaD7OHC88Mz7aLmhH1k+
KDVRDzLhscPOV6YWcCXmk2OYmzFo3dJXF7/+N9+icNL9o3CiMNBIoqOAkFGvgx6sVww2RnDGskuM
Z9WWq6rzM3fNtC3Fi2k7fmCHpQo1wIAPsjPes2X5vUDjDYRYXDb5XwLCvLZSfbmXSWX+MoIj76pj
k4c280EvE+xQKasbOeL2L9npEA9b3Lm6TUBaDMPI1Yn98tN4vTwHQELBRe2ZbO/kznn0jLolzhiH
6oJ9WkjZVykxsKUbmYmY39LfaV6/p+kALQxOuWhFx9A03m4BDoO8qNbqQgIIV+jLKtV00f3DdvYm
kaBuvqF6smCj/x2PjL4u7Ub+gpKwO3iAqVeSSCBF0ll/yb3RaGFAOoD5hk4D/f1A/o3dY4vP02n7
81Sih4+4dJ/1TqpbolzH4GkAWd7Z4Ug2gOx1HsGz5z6eDGzvVKYAOuug+L5FsJ78HUuOmisPUmUa
STra3vcf6d7qbB7SEWWZRfUm1TBGhsgYYEdh9L4SeL093Neu3KcpRik9cx8w71Mtrc6izx+Esli1
D/5CmmGFHbiFVpvESlfHBw8N+ejnO64H6DG6P5Z7mRme2hRwlqDnQb4AxQfG58IydRqQyYYrmflR
ut6ArcFeFhnH95xXVy73naEN/54D5Y74wm1Qyf/jeTqM1nCSB8Rq/i/B698r4P1idracuL1yWJKF
vMC9wVwqsDRETiEjU4uO1X7wVEwXumbDu3qm4NZ4N3CU9E08ZtYJS8GbXE2tzlSV1r24W5zV+rV1
FUGLuZ7UZZ5fHnIHEj5DSHYnx3a7N9EH6wgGyamzwF+jVn/KeZaH51WI2x/gJ/mPLGsJiy7ZN5u9
+kpLhpywBdAKCOQi3wt7sFSsE0+Fuouq5wer3K1XfcQFnWPmbdcmceNQeWF07OFf0ip0r1rVew00
ZjlxERL4hzHMeTP9w6espItQeFNEKf4kU2h+V0UmUeHT95TV/ak66ZfVdkOuPfSnriJRo9pCR5M2
Rrpq8HxhJhFDI/uHLp+Yg7pJkknYRBzZF3rvAnV7cP5SujM858W/y6j6tP+WJ4PGICil5amNtuAt
Z2kk5oHAcCvsrnqo0i2wDRZzlC7F+cICcBkPy5Tk8sw04gDak16ifekbcqR3YOuwSk2gPb0YctjB
ZKejGO5qysrtsFnzs53cjH5CMxhW8u8msschgMWXqMEbAgZst6PHqIiPNnZjaoh0onPFYpRUAL/s
l9eVjwzkFE6k9w9eHh2Kiheeo9YWGiROeZ14s27lsJyvV+WEEyVGwyJkRUT6aQeRXT43ybBhSZdH
VFVtaUWIlbio9bOeosHG9Jqdk7pVrJtGcVwSyZ0gnP2BgKbyAeb5p/Uvw0hsIo0HhEGHEBSE4vCA
bwMv3MaUFOIa8SzLT/kZegB8jdDfvdVK30cPreSVJxEWw4oVWSVg/pggWFrrmzSEu3Ra+9OKGtuG
FWmmJUje6Q1VYQBfcldXNy6Xr9tjVeCX4Ix57Km5bnaKd5yQ+gHPAejvX+JdpOFxjZLsiWh/UDpn
9reXNyPYEPh7nOOBfu+XHKInpZCcRVQJQS8xuBwC9NTl6eQqZVTbXIjV7uRL0/TJ17mRQX91ZCL5
U5Qw+3U7ejewoyIgpRdxcj/KiVYZMXqE4M0QKUMfz9FhDduczc/ZmJo5MwGs94ZG5CSEAKYSQYqf
neTnQRqrYp4cZfOJLp1RB8rGbN1zq9q4m4dWUg9TelvOFBCAFPU13K5OtljUK4ShZvRqjHoNQmJ1
Cv9Cd6Ja3TpXE+at/YLenB6hRk1j8oA63CXX4HCbLn19a/DiJDLgfYXv5xIb5dol9OwjRIwR8sbu
bqXpddj52cb6YRzI2xe+Xqdj+09shC/+H1IA6DvFIs7796hpmYoHfTQtCu+sPy1/8+hwGkmm+F6O
ZCOARg2kdkmaUVozWOSeCV1wWmAqt2MbsCQy+fo/VYf6i3qXlY3WN+5h/3YI8KPgNNbuhSbDB1od
FWYXkenr1bPQ0/iY/HOCp1mYNc40nqdgoWsZq7NKEhMC1c3YjHtWS3+F+YK3PI8BI7GNzSccTwHG
tJY3kaz2nh9NKVBgg3Mk1/CZfZygkYsBcc7KolM632OU5Y3vXz6Zuk3rssuaAQFKSVx3sErd2a4t
I5IDT0mQgj935isPU/qNS6evhhLZnvPoLU35y49d4uYRcrSa/xatvMknl2oUliEwDh5dweMmoqaW
jF26O7ER6qOEi0HVO3AnM5Op9CMi+51JkZWZT+5TO4cfA20O3HDwpfvoMTQSBKeBy/uyh1fgPFg5
aIYSVfD3c5u+W2NoEffcyfzJvc3PiVphaE7m1MdS12anYUggcahQIuCLMhC34rwPVdioezTEFIIq
Xl2jMuaoJKhOSvvIW6hptRrGD6DkGAWv2R40CTlUWhKJqfPLQE9qpKlQV5bQHsQVHUtad//91Czy
gdWbhE5jWJPp1xeBDSPaI0TW0oQPbqBlMgJwt4laFiXHbtxSkLSxg2cZDyuyC8Vn8VFOJwte7ezf
EN8Sa6mCeWjB7k+tCuuTJGTX7kLYCrKVIfCnjrWtjh2rEf7lg3aAGkJ3fvy0RJE5pSwBo+f7FCT9
EUb4zxFjd/izL++4NUITjOc4BCS6zEb/lKMwJnHK2ws+sdyYFZ43Fg3mELDVCwt0bXwh95j/Odzi
DVLgJEwrWRayOw59PDVhmznJEg5W/dfLU+MgdUvghxabsT7k+Z2oVJUou3ENlhc1mY5SRmXUzK14
GJheQHApdfD1ezYJhPXTP4miQ/imL1TcoUS1gDP4eYT+eTDwUP+ATU1wTFzFfHzsOi/pNedADU/c
+TC9h6E4q7UOUtlF2YigcIdzlYcoBBA+Au8ephG3R0kJCfQhjxYQcfCVAqTeTU6h1qe0QA2owi0m
HyJSgxGj1E8dVlz5RnZYccfJdUz4JbLed/1sxyBh/q0NY9i921aMJNGjLq1rXkzid3GI1NPJFTYc
JNKRlEoLwbdTiFrpqHOy6SPFQZqY12A8OihpHZSLWu6ZCx4H+GAFw5vnQMmv1+N0nO69xeoecYBk
O3pOf8zRMuDLS50LSnH2lC86x1YXVhdA7Qq9Xmyd5oRiaPIxWCP5ekftR+uPAj2A2jyTZIJd7ltQ
lO+8+pk652eHImI5lbuPwvN7q4dnR+GSP2Eeesb1wU/W1azUaPHC7xPOtMLDQ9Ls7/F0tBd8eSAs
tggfsplCwmUeN6aWrhvflbwhIOz/STyWSlXDRv2BLFg/zJF5IgK+pRS/5dEQ8J82ioR28X1PUcBJ
8LHSLJT6OCZhXd9De7S4vcWHZ9MmB8vP3Du54BQXmVmriW2kMLIaKFZZRfvIuO2Cwvu1cGAXZHrD
YhThv0UOKB1K1o0VjOTiCh7C0S0KA29UELfI/y1lpHXVZYdE24i+dc/AI3S+2aubnfVEUAGqBuqt
gVKJeAcGbsH6X/lTjRpsyvlU+jcpXlCH2rlqYUd3Hxy89CDh4zNWAubr4W+SmeaMpnPsAMJxDa03
D9rEnREYyt7mfNFlJhxyjK+hgVBPwO73O4fop+es02CAmcQ8YaY/AHBSKufw7wBFR7VqcfEn1Tcy
eLkxHpi2QAjVf9QuJWhVDyWkpOjDWMf6Fqguztf1r0Dg4oFfNNi43mzVAI2ACbtxhdiZonCd8auT
yZf2TgS2EUw0aoIq/v2o49Z9zM70buwT/VPCxvxkuE8wAkCAZcZXUz/kkN+h2EslvwiMrKDy00iX
WgfuRda0S9q+CleNSSDTF5TQKleuneSVnoQ2v5tLUf44ypnrvXffrfcgv0vhjwGvrcwOVhPhAqKf
PZahfHrp93qkhqLXFOVFBDAnXylkTWwMsCZkNw/2ic2J9V/NCua1DcMOLQmIqGLNXF38qHVkSe+n
BJaLMRuyHWOCorj/yBAOQv/Grru6tmHPpILWtTPN3K6ctKjdkHEY8RLDJQ+W2DLohA2qwCa+/Gtf
AcNKiD0fxxyhE7F1fUDFZ1WWoBQXqDK7cB4leNGZNhn2GMfYrX2Rf2FL5x2ROTd9yYqtFRv9fd81
lODeHbuEkyWCeO+ZnR/wr5w7bcUbPTwjoDUGWwsvrChoUqfpohxbX3PFleacSVJXodTd7FOREW9C
pxifFatmhkXfoOhdTQO71fsy4hgVAyWBhthKh+4rqw3CoIxr6nomASl72aTl98/gWSlqZCtAQvCJ
oEMU8JBUoEVRQaBhWwT+ut1ffwxKUxqVByFkKyVYdur6cMsGxH+xFMGGq1wZlqvEWaj9B2p5vT9U
AnlM8yFdWekSRQ0LHDKQ3y0H1JBVyMAp774Pu+fIfEZbdAJbKkuDVVYbXZiiphXT4znR+o4FElt+
9Jrl6iGO0gFESdjHn4yfSo+rvxo04anL+Yvko839dVa9lfuZ7xXuxyge4Io3TNlXhL27A/h79+h2
KbpCJMaKqdPDETYVe3n6s4oUhm92elQHa+C44c8xrSLJQskPI9LO7gvhfY73/hnlAlCoFWl453MD
mqhqiJiuGI8J4n1PB2bk4LtdWpCFqUjkagU2TyqSpX5ajyfO2zSkt8EeZgJdpr2kMbbdycFZvQ2L
9W7zNd+QdYQ7fejTn737GptbmUNVVWRAJl++J4GkWZAKWQf0ehyOqINlHXuB9MlxC8suqFlTt5W5
XD8+QSfCUjo5zLRfvb7EluZ+jk9c3dhfD0KGK5jfG2wZ2sSMg73mKIX4Ye5D+giE29cQ5dc12KAQ
dU5IaPhGE+pdvjv2tPDULEaGieavWCNzZgF94JTlMdmWlGUf4ppf4I6ICWVAEn4OBz5iq/AqkpL9
JRPCX4ah0S15ivY9NHIbOcGEzk7PxUOFgXciikGg7f41ihl020Rn0JP4PgzkTzlQnLcbjYGzNton
wVV66h/czY6379NeaGxWD3/sFYSZa5D2mvDAoooXx3bAjQP9oQFHQgpzQvLAnO6g1MVPX/UoZ+vN
q2E66OHGu+jY5fAsJorLIhph8RHerb0al43qGgq6x4gSJvt+uAHn4UOVEK0ujt1v6+Q/Je4J+WoR
QxBQHd5N1g92AEhWk5Ygwm8Dzce6/8MAGZDeN07GmmEqf4pD+I+f9nJ14l4wGWuJH85L9kTV1tn7
EGlqeR8wAgNH/jZJDZONBEa39RnelAWFYWlqGNwjDFLtwAmrJ0PwJram9B9pcpkw+e4yXLabHPQM
13dPMWUhsW2Te8yb787Ph2oyWfYPGTvdI61o1hUPNxeCsfehWNxH1WJt8O9lkFexfI9gxox7i+TN
e9kA2S6HGlEW6sU+b1dF/v7qmFNM9lcyis3TTsOBkndJYh3WYiJ1hvJSCmIoCXshelccpKXvGYB6
dzeBCqm1OVJNMpmL5wwc/Svm0fWiE17hBDA02oNU3lg0RrgwKd4G4W1CHwaGQU0bLrH5FHvsapNT
U8c4DkwBVT5NU0QBEDhnA1ktL1rXS+/OenrkG4RRQxaRfmlaw6sZiUw6xgxJI5x3IcAJ9/fI8yIh
bQHzmICh71mF35BjrwMmLnHPBnce7WHGp1XfCF7AmU1AxZN1FNLdQApMyw6nYfCUfy+DDsodBLTr
I14bt329CxXGzA/9uIsT6bnIxlDsVTY7R+81wxJdWKf0BU3bvKSTZ0apFWInwK7oupuK3jQ8/csD
t0BjSEHCWXs+kvxtZXgyXJRTzIaxmVIkwxV4av9aFOSv9Jf4MehDEVVYRpDdXJJpfGR90982Iiz/
JQFGk969EO91NMOjuce0VKcE/FLSB+A40sV5fE/eX3wRQjZRAw9/X5Ca2HgArYrvV0vj+z1CyF8P
SWt3aa8MxpZn4tWeX9GzTHTo9ZEmYRfn+6wcita/gCEoCEvYjeMoV9BKHnk1uFlyBPs9ZAMcpdgA
7l+USlwS2Ut0aTMlSZn0okpRio7/yd6peEO+iaiA4zgVjfNjL4y5LY8aC2uUHTYFADnNHLN5k3C1
e8MHym8HOYsr9ug86r7SLcm4FaYw2yC2fq8hHHIXzPD+I05ypLHes2KzGaSDfFhNPzTZC22s8WV2
C4/EQlpOl13t+ycP6GTMu5wf9x6d9WgHS2mA+6XZtEsZ1VptzjSHUXp5yJSbGXDaaOsTlprb2/4R
JpmbfRVj3dcxWS4mp8f6ReDH0yfNxzF5nvOiM4w54C/CAQd44TXQoe7JBOsTEKfZeYMrdv1cl74f
xEByc5fpikivmHjZ9xDbpATocWF0qMiLGw4pjLxw4LRpqJ28CFzWBsmym0q3/gd02+wolgejD6pU
TN9yXsFoqnI4kDiUxZwqgYYeAvVGM5LPxScOWN2jO4VX8vrOXwIkjjImSsDoXwHY1kbICK2eTnAH
7u7Hkoa8FEatR0XIyLCcfXqv9nK4u/MCz6MKkXxZ7vakL/9MBaQwo/4svk115Zq4ivxa+BHR7JjI
mGSOYxK/ZXeGqVqBqWqa9IQh/FQdax5rzIZVXvLlhBrG1mQRHsu2oSmRJm3t7RLFIPAC91LMYwpz
MG5GndyMBPGI0BtpCA8jcbAOPX4/1DRbVc/6IPcPWh3+4k6bd4Xs8LcTJ4DpE7M6hWi13fiO6KMQ
99oavWbei9R5tOHudD8j89xDYli5eDZmQGIRdrYXYC6mR76Tuw1pFpHV+1QHzpFZD/qqGLUrzTTj
w18dTKVfc1vGtBcQJ8rMNj0aQb/63grWUAo8RPZ15pCyTHiiCBR8kn2MHyfMa/DmzR2DAMYY4QVg
RL+/xN4CE95CNxwiCm8hesqVUpSS55z5FTpBLmbQVPJAAjPUKl1Ahmrr/R7X+UQh0m2KkrRcPP8K
8A6Zx8p9b7i/4PyCmT5IYBsFhCO0srkJac+/PtHyf2rH58si3s95ocfTtGDFkgt8lo0U618lIPdU
F1qqVV86UmwEkdjfeD2PI71lY/P783dF3+gDPfyuT+WibbN3qlBPhByWgR4gVPCz2QvTPEPZNFh/
+oqi2vrDFXbdJY6pyUVvfuCBd2rNvzhZMAJGUN33sNBe3JxAoDIf9jPiMz9LYchiXVUNE27j/lxJ
RN7f4ZHiCVi9JLj57+91/evijeM2bzFi/U59JgDMavp1H+vdG/0ftsLhCTE7e3Pf5NiYcvYGBrT7
153mtGq3wZhDdbCmgX99sSjmtm3ufLbGU5ie+FZv9x8rug/NcXXzFTgOJ/2R4T6APGZK19HX6v7h
BrN19yFZPAnuQJL6otZ4ct6b1vF8kn9tzMezhtJuOhNr63KMZlt/tmFP6afoPENY4quc4gY51hE9
IuH5TgCJEcCJcLwrP3PL50cujzzD3Lniqg8W/lnwVcR7TOv8s5jNwu6oKVfQ8bBqwbVVXc1DKHL+
sURZrIB1C6kANxEuARvmuwyXBHMFHkgXgm3hEkZ/OFjE2LgMczgOsG1zQjlcAuNJftfvixo2LnV6
VNpdwFgvCBikwEtzdrMJIBt8Z1LsE09n+g16K9P01Yo2ZTP0Ht+C2TapPaAuAzf8IBbyL7pzqmgb
rHiLab5ecX66lURuw8cqUi/1laO7ndJcBOjbDSdnYm+4e99NRoEpNRImhCf5SSHrHEhCsDeDSMqC
BQeRwImehDaQDInYbNgqixiU8Xd+f60uKAZgc/bqluysGMBfnCDyGiBXbTKcJgcnttj0g/D+HYLW
q4q/E9a9tk1mQBmouydRcm7iidZ+mHQXzHI/5JKei3MTbMhQl14LKc8BMsVGevMiYpe/Z1s0vnST
BUish4pQJgH/dxyIkbXCKy8w9XJ6cyUH+uIlg92N/uNZze5WeKpKhFXDQskTsEwNofl7P41ciKfn
F0gxGFxs1/NwuJjU8DGI1T45xUPX420lrjtbOeGoarvKzCDLEZ2+SUEUoFTPbYsGU+BnmCXUJ98P
btELOpAmrAHHBL0RustMD6CXBnxPZqhuD6v1pwafkkoxFTS8HDvo/zcHuMHLWA9qY5hOh/dVx4kK
WOKr9MVsfVnLSc1wAPAiG++4ezGzuipTFeChmoGFkfj/nWjm5cwekFhgCsmeJHphM7s/FGC9ggaQ
XBUel0KZHrZaPVKQkDQDli3l0n32GB7p58i1KUzF4GRlzjNhguh3wUhOSjKvnB7TsQE4TRrhA5Gu
x3qkfaXPYE2yUlv8UtxSg1uOd4OUSHnfLG0BIB8waadleKe/PN0BdQicwBCPWi9gZHtmMuGB3MCu
kM9h68D8fmeWeqmYURn4AEZttKA+j6hqVRfNKNRy3/if84wk3rj8pbsLL/x56IeqEYKH3cnjcslm
djf4KgDyLCnVn7U4380nlJmePNWkFXJGTXrWwjMMvt9TMOQoa3hOpiFIPZDSwTV71qiJQr3TPq6h
3v6EFyb+HnIufZq2V03v3Om6MBPC1QHjGk6dh0LgrXhJmy+pWna8zva34JfWu8/TmSnFwi0xEcWP
IfnuFCUS1e/a7cGtY2lEPH2U2YEC20tEoNJJLFUWFDzuzxofIYqjy+maf0cmE+5KhdEo7OJxjpM+
2CL2bHnMIl7aOyWlYytVrgL18WkPY9bs96mGuvcH/CFryy6RC8S9Csyl5UP82HJ7rTU3/0JFz6ZW
lioRZSsQPRgQRUKF96SC4kDqUVIqfW0Wn4wHFdRh/PGgIGIBUC+YKnl7BskA463uAFmg3a5RVNia
gMkYjzZSnQ3OkSn2eqWGxcKe8OGDxXp2OfYI76e5+pDPkCDKaUvsiqXfO28HWN+pKDpf83NV0zo7
1T3HMCBmDJHUg6Sr1/rwFPEBj+EgZRE5TzPN0N7XAdIRs5NPcVRP1lkrptIxIzXotfjXw3aXIVRq
chHIg818Pw4b93I7N5Hsa3WjU5u46mGkjoR38IZeMKONkXDKrEvsy/Vnjjgqd8OieisfYrGFT3Vn
xgBSmgQcTPKX/dqaNUYumpgWEFdHUIgF7zndPDGTln0lnaZ04xAyfTvn4bHx/rsGO3Sm0isNC5Za
TaWFOwIpdvTEUHDxi+s8vbZrpjviWiVkT3FnP9bSqy13Vm7kN7sSM2NcdMtHrW17ZapbkPLAF/aN
o7ArYO1/mGmLKxFL9nrH0sx8Y5R+U0bRnUEEi9qKdppQGBvb/TNMo14cGx5lV6ggusTW4A1nHabv
Ug6C1Ik9yqDAFu/e89lfQ/8fz52TOGvHeD3m1+EW5Ytmj1lnW5aVT80+vrSU3mMlaSrC8Xu+Rv2N
Lv6U40ak8rxcGWIDpe9PbSuYcQAybOC1OoTRN58FvqH2Doq4HqGChkfSDc6EjVroBP3ROt64FVxB
PBNyyNCBe3fqsa1kb95qWRjd5gCCxv8RoaUArDpHCdTs/PHlwAWl7gfm8SQe5Lg52EhDLhoXOGXL
dgTwCyBRjQ3tCZ2NHf7vD9y9QyNzwC2m3S55GYK2n17NIyzorRW65X1XWI2WoOzEorzDa0y5qBmm
vj4wF3nYDLru0kn8kAnZsZbvdEbUBLLkHsTgeB3GvLDVFBgDDbNJATNG/AG53EkijAYzjwgZP0g/
ayNMAzU5FOd9ngK+02Rv8XHkVZAkxIAFFC0SWBPilyEWAvqXEZKKVTvbkk8rmg0YTqrCdpYMjUkN
b1yV/b5rYgNoYFFfjNjQfnf+sCHa4cZvQhtr9MLNTMRJBlYJD1f4C0T6Jwy0faluJhLeBVEemO4q
hAahZJsd5aMMagEmYaTqLqLYV1GksI8KRcMJMjlYRD3jV4+BKUeBY2rjmsE0/XMFYIk4mEXwJKIn
UvLawHwqZjci4n0Fx41j8Wfzz9nXmKTi8TFzMRUEP+OJUTwJeZdnIfXqp1BcCbLac50cPr/Rly9l
Ok10EBAHAKk6EeMWhF1Gw5b9MVwC0cXg0C7Xsrvv6VGg8oE0xHyLZE+KLHw+VZqBtxKWkxVUXwFo
WDhRweZNIw0VSEoDB7S5F8M6WR4xjMixa9KqvqCsb9mnmBRty+LRmzFIxup+UimYr9ULFwMjOlgL
Q/boGtsERQDWOp6/9asXNfYTiNHtcA6itVPgagEijgtJYPpN0VzUrHDQLtgNINKAWkZc1aH+9nwe
CIQIzh23bniZMLtaEZmy3sMTUtHQuFSQxj9PJuBtz3zoaAM3l5+uO92iXo2w+Pi2BzGENK1r8KBx
b340fD2/jFYrteFsEnxCXEttvT+899MOrDHYXHJouQpGfV8Zo+QV4vVwiayuU43HTQMbfBY1Zd7E
N+pweDjy8jkKK8hA5+TY5meIAhKKMS+/m84AGC4BzLIMGrvupTqZERTrTj+SqIiUWroNykHkFEOO
21zVPLg4J1THR/BoH8mACU0GqrnMiIKXAdfW23wZNiF8cO4hyCP9fxkDEtyaKRILdbtzTD/nItip
nXeY5zRX/zl2BttPCFbSLwBUhNUorxxw0/K63JGCyE0/9zZkWqKaFUjAOB59qDeW8qFLXjTefMhN
pOxP0jQjx/AKM6mCHHm0Fcg45Kd60Gj6IYD1HLTFC65vYF1P0GkO3WkhpCc6WHgAg+ue3yrOgq4U
5D/GW/xk1TLilNdlFggQ5N8+RkoMWMqjt0ABP9xJtOapY6sofmrVcMNikfKMflST6XM4BRpQ7ULl
1gdpmMCu7XB7Zic1Ppel362ptLuKx5wwevhGbE7+3xWFIpBnpxq+HRMM2vU7qbe++XfcHq67lsd0
dz9UFGCmr2chTuJhgxvoFLEMPlgQXo9WNzTU6grQEBjIw4mjG0APMk6w/VHdCm+joEpTzAT7AvAA
hR1/NFwX8BfL42FpkO5cek1EZsF2EIEfRDSVcnZA1bPWjcw9UcViYvjuXFUAAV43mf1/RUpvPPOE
qN2G7Kqn3FBgjyQmfJ0wFG7D2P+FAEM5MO2DczjJBhL8SVCdBvzG41DesrFLpmpOxI91Lhef5mmQ
ALPCok+Q/9M9diisKvnbyDY0SyMV86EakuMpgmilZWhXWQfj00u9Wtf3i/O2yViJEBrt176ewbF4
/6AGxFpInJq2YhSW9WNuU6qt4u7FRPadjXAYLuZugCoR9lw1t1W0b+wmLw+kifxrQ1xIc8nMEUpF
6XEYIfMZEfZNwWPhujwDSsTshYJ307gPmdfO3vQ3aZvZzFTssq8uf2gLWiJUU64L3reOt3NkkgNn
lXOPA5nRDe2iRKHwco1vVS1O+94FBDWF+cFzU/+JteycO+bryHeEtzGZIi6rIvMWqCaFfL9XGzuf
x3Gb5MbIYtsUCdKVYkX0yL4AXREsSf3l59Ky4bEZungIMMJpG0VMcFzDjd5ywyfa5COafBAYXZC6
gPAv2JUPIq4KwxHnOa3eprdxGaxx+WwCAjWIAKllUqRZJBqWzq1MQxtjMEvq6mxQC85ntk4OqLI2
kySh51t+mjgFc8UEFpfNa7/9OzgbB4hKgVo+9V4GrD7xLEm35BEwCPVp/Sa99z6byP6MEMQkNREi
28zuHa3azIXZF+ON+4WOx6vRHGBXk5gew2QAgXAonMAb7yoj6ZAU+kcSgOhE+IlMNNJEJXdXadhQ
ZrUiujqZRiNhRfvex/rhBoPPXZkyPW/E2fvEhmNa70E+YFeWEMoUMhB2gS1SzCN4NJhBliwMszBz
Vf8JpXAbilan0SqTKieYkMmHDjkOoPebgZKfXJtxQE/35lBHd+DjFQARSHwmCoV6gO0oU7EG5SAG
NeIjC4xKftDxhbQ5jxAwkVAjB73IpOBgCRemNctBOoVloojyZgb+mCBgkJJh1+1Ivo91RQV1iN4L
35AySYEBYpxhre4qqUWk+ywZAO4m7mrmZDR6P78C0svX1E5iDjDR/0MzPCdLln78Gy3Bnq0UNMjd
xMgoXwEqt/tishtoR2vfPS0dcD9BH22iezm2RJtNsFYUcXI6cIJlyS8EeAssNEg9bzvwYUtaNkTQ
y726hyOWFk+x5IIgB0GIHAe4BBlYS8KzfZdSYfOp2PCGbYQpTB2Ecny7G9F9IbkzyIUVyq0i+EgZ
jcpEWjs/Fc3kvNBlIZgsLQGTpDe9RM7csX8yLwJzD6b4Z+pL8vE8sfahFXBEFp+dkQGi5/VEI0Sh
YW1n5aXnrnqRXkw2KiSYklJGBOnKvxL+ZVhnp8PYIuNHE4ntXpxJnAFnJtY2Mcaoew+c1VUxpT4t
4osnBSE5gjORVyMcD5Wo+TvkMs7o3GL9gLnSt+5d1PSsPtAblqLmFmzmvZyJ02u7IbaSpgSqFUy+
gCXRvPj98NIjAmW8MWfTsxiRleXXxcw9IVGIHCKGdk1LLHPwAl/YyNuSQy6apA7PwgaRxY1vEbzR
KEBkwsSeS/ieD8wn6ih8zRY5xy7niD+uNssS9cWKz/a5SnY1KXfyZr0zmx7G+bAaTzqDDg01xCEX
Jss8PBDq/OlEL2ECFoX6WVGeu84uql3628JOxVDZlg6asSIf2GEr/3f9CHNbOGhKb1AYFLXVyLbr
orsvcBDXcC2lz8HBJqUsIRkvllzKQidTv4YTgDBwseZjesTkV6GHVebTekBfladEAFitOxWxGttf
SlILlv+EkoRg4/aZRRdMkJ65Qyrq8J4ELye4QOfyvjxNVoY5fwk+ptaALPd+cOdOt7kM9MDxRJiq
v34X8xEMxJNF6qToDcidDeAlKuMZBwL1Y0FVgKVK7gI7+IJwWBt96DwOy2lO6ggwzH1ooKdXtygG
rYVVABQkMHEN9fuqAFU9mYRzoq7Ct2f5AOmofFw7ffMufwyVFk2LnGImZoWcBlEeQkW0ra01GKBc
d9fe4JN0ifXVzXiT1lCp70f2q4h7AtfoxzLU0qTfX1FK0enYo6MWT9ZfyE+lx0kCTFR0w9spVPwy
7yR7cU7/gvpHferMuPTqZfF28x+Cr51uAXtef283GSzw6DuybosYmdRcXQjBwWKlbn/PnJz1mw0w
OHmjmbKT+BvD1E95kB5VxtlxX6TtWfsUfV04tRpvd/4/Q+nqWuRmT1FeWe3IrjETSw+OTbMK5vJ1
52kE4j6m+URjJomNXDlGeZO6jbRbxHVtFCY79ucLJ8uzFEc87z65LFCuEmWWKiKZewItLqb9x0S0
TjThnNgYsZaGDdpebIeWXxRqxxoAWZKajUwbjguO/A7tTW6eHxr/rDLK/TEvtfeKxxsOYGolg0Tf
fkJCp66DZ96Ui6fncDv5Nbash0rV62AK3le8sMBR6ln8hp9MAEYKPANq6Kdr38aqlXlOKnhpufXj
TeXL2gxR8IOYInlRDq/zvb8yPK+vQ8gmSbim1elmOv1rDZfX/NDXn8tb1XT5bo5SmJ0Eax0HKBOk
UN3piuL8+60QTW30mP+IimvVvI0RD83XEjwn5ppq7QGiIcQubBVhyKWy/CSJ188GUxdTea4/vXfD
w/bgMKS5dpaqtzR6L4NZBSKN2875QtkKx+Av02D2Yqv2eN32YlaRufT/zFv9dGYZFwwmHBcpoDfK
yqow7wR5b64aeFiaL+AIiTHpBW0RB+cnJ0BrLFSpZJK0ucqQWN+Y4P/Sa/DXRbjDXID8KhSCRW1T
wTskG+MVsO0lnCEKdzovMI8t8PWjriJPh/yMCKiO1F4RqwE5qruyGGmccIyeEYqFwmdJiALvVjcx
RjRvY/cGZVnojdHzLEFO/DRxjc9vTx2IVco5TLYk7weGWjjTFf4j6LEqx99zaUabZiCFcmRkus8E
DZmI2NgChIFZf6A+SD2sjPl8uooMIEnMc7IPffkGWGFCK8dkjlCmtjAtvfVRk7MLqYKZMVA8Erq2
O/Bus5kUGrN7EftcY1WVgcCK3QBGDHxWcRZdmUCtsdpzK/qXwQRLmB0XUfddA0/7g9sZ381tUVVO
krjN9UldeVfzTdOlwYpYjtq9ceDWFsgtSK4A9BAMHzxLsis9kihlKurFuVsqmWhfUXYLrdLQbPWd
awizM2LtOHJHIe9G3hofmtd1DOMmYFsmxykZjSZNUwU7IM21dYAOEg8IobSUKxH6JKY0xvZidlSj
3nFIkuX3bGQXO7c2yIwNWQ8we/V7lqs5pM9RLaQwqddspEWGqJhLlPip+kxfbiXp5qxysMXCysw8
JKGoMZMdFt8uLCjVYEV2B8NO1Z76moMwQnMyiS858rkN1V/EmlZl1+CyuuVDH+VqbjqcWGzUnfE2
zd4GJu2CijQQLOoy/LNjhsTIyJrBX1w+cEGuL4vXBLLqiq1qS4ZXzpSr/rCkw80UhHlsvrWODwRn
0WJIuVUjh7f7daHLsaaAfYM7XIJ8uI2TRx9jCLlmIB7Il8/9ROk3nQmIG4AzxsZ4Y2AURPQZn0La
xkj3rtB8dYba8nddXMP4Wu2RFgaVerPzFspWgF3pWhedPA8Krh6uwrRyINHUR6BFZnttfCem56XL
XATeXlFHknKHOqtHVSgJURTjTL6r4oFo+C8ngVYEyWFAXKNGx9WyoDx6zZiuoS/skPfNCngw27KB
KLQsLdX4T7if0k1MzRwkamFAIHfmukj50OR+3QvKtIOfuSOxMT2Uk752f7+5zpAZyTfR7kLF/who
JS3WU4iDnezgPyypSXp8FUBnvcSi8zwgJVHSrN+ndwrkSKTMBxJwGkpPXyWxW+NIvYF9Plqq7d6H
d2Ry/qeHZVZrxqHgHu92ERuKPiC+wSAZw6m/lZkmvlmHeSzgvv+wv50NWDPgg3pqlp8zyWzGc2EZ
BcIHzh45YQilOV53lrC8OAIjhf28Z7kPdTHsi6+5X8bY6x8TTgOhszedDuz8pdJpIpGPgwjDv0bl
vKU01Xk8gC+ssSNDDqhm71gfMBCoGbvHA4O82Mh7ZywvHMRGkUUEe5j1iHtjP5hbYw/PrMGvSbEb
Fca6ZJ9B4z9QdIZaq74QOOXxiz58pKXg4brn7geKJLMVge7YenQFfVS4XCP0BTLoTb1aRgvSNArJ
6rctRYw5+Y8DhX4B95VJjxufS3X+F6BZL6FdJfY/gpp/F/OTbTCFKLmwFkjVdzIZgpoOZigcvyOT
GNQ0igz8O/UIXWee8x4RScp+lP2cOX59UqmyQYFFSLZO5l2rYEECdyy/5SxZ/mYEIkvkaYsbByDK
PdwWquqBFbtM2RHN6fdWiPWVwnslb6oeL+p9bZWMNPCUxTAUdnzNTVhW2Y3HIyDmCfGlewsIlErG
L9cLjZI4IquAXDzpjowZP76w7jtTxkVg94DmZq1l5pJF1C0DcD0EfLisGapNHUj30BmxJA/UnyE0
fjh/zVFPWyNAV2kPKzVI/5LYI1zpp2/5FBYhM/XwFJU5dS2l6ourI3SW1xomAIO5zYBVRlpAdvKM
hGuYIcbOa0wf0KkeQt1j8vxBgI7H90Jdc4NkLRtvaGP1toCrtpDUOLY4nohX0nEDvXjt+pa/GHL9
8DpXIWG7PA91xkYymK5yyWJbBA7mWypBvFHmDHQriU9HO2QiQaDvZ8kLC3OTsiZhBGYeHowaUrtR
KFyN4JzHrSVdKtP1u/wCfIDMwICBqFodUGL2LwqDLeG29oGSJsaC6DxnwspZsh3qWnlCv6zZ8DRF
wpq7E7M4+7mJbR8c++i2GUBvaVS7DbaAS7wHoAKz2HP/JQwmw6G4lQzk7Ghv5/uVW16wfJ3ApH0k
JkF1BcCa5IpSGxrNfXiPoAaRZKBhQsoAbPii6jGCSFvt0clbcaGWhU9qz2GpNaLG0FtTVZuSeiaZ
HekeEdyfcpThxXIVKjdT6IndNiOLciRYDIVrfxfrMCHGiMorgZEGZh0LzusoZYWa32sffXFp/gcO
gPgV3sqbaAU4LlCKBdZnsOdEmlDJa+o92HOrv11gik5WpyAqbZ1j3weqw1HNz0vZGzlcbGGC0lg5
qPhPOa45F3qKy+YIaVBm/ZuvfBzHAgOGm0tLMFuXqWzp19Ikr7QnXXpWmOvdAwtrpi8DAhbS9ScN
TbZ2uZ2PNLNZQj3JJFyQtajeRebqgSVw6G7b5HzYKwqhj/4xnW7xljVtmpRYTgpqEOQNz6UvgmHN
6k0ClU0hgI63kunRKdJjs7xdJ2kTvgtWrIEMmrGuYoJTe8xB3AFfpmBiXMwbmCwbCEM1d31HhUxG
9+od64hoDrp497NWEhsKrKwsUyrzH+o32dL4cJN8Svh+YVl94pgJ0xaoZBzYifhxae58ANFXUXrk
YabBXhlwVDR/7Zfp+prgKeZxHyXsxLM8n0j6Jm8hsEOrMNpT9na5D1SiwM1I7koY+f3Cuf8ONu9Q
nHjrrspjw2VsH0Udc+ijvihT4w+PnoCDpaRNhmvJ/j3Q+VLfu5MfgOx7okkqQIsNiFdalNL/yfQg
amCag8P16Zh/MJqnYiahk2avpg2BiygSODSrpBrETHx7cv3+Th0cf7f7RR86OYOH7HEqQTFgXyDF
up2bXC4fnq3G5JIOIkIvk63L/fMRSg5VQXg/H8ji1vf8kLOAZ8Z/50JZYpw53pxlC0S+PkeTvfJ+
1kQW6HGslg5SoOszXnOenc4m8DGPFe/8lPW2M12lQv0aH1Oo/3hbxTE2J3r51cAnHW0ivyvNvj1m
tbPHns9kV4YzaMrmOgVi6qWdMjAoUD8bXSsJSkD2elpIIl8HOhH76EW4RBoSvlbAo42X2/KDvUfY
oFLSdfzHCDQt0S5uxzKrUiN6ezk/ooeKbiTjUl0CkcAHP9qEm98QcjwSZj41HirD2CDOWepJSt1x
g+USgMnkeW2j/rUz9CZQopAyBYsPK2TmX3MsqUz3dNDKNrOGDxf4yJDaXaV5jkPG1fYQkFexNqwn
FAT4fN+Zw8kUE7Qx3RIrDh08T6B5A770EoM9lI2MFXfPwNgJ+EzWvDC3jnVG7Tkuf6rAzSguMSzO
jhzbWfOzkPQR/ObTbTxGCEZA6AwbXbvbJwMUPBSuho7koE3qE/QTE76Swcwk/351cfCRQWj/ny2s
Uqjkz9n/49+6qLA7VS//hyoZhbWpj4WTBU22Ff70QNG6pfyWTGwvhhlIXUWbYY8djDuj1Silmh1M
H+vqSrfQPY7iaYS6VuSJSZ6w1Nz13vW/X0c0rfQmdRAnHwem4K2tmpQNijtUw3iXQL5ZaPn+9Fd/
ozh3sT0WklHWnG5EoQ/Yo55LoT1INYNUA4YRPvNG41dWKpoM4omJNR5Xlsp5ZV4GlKfLROyy5MAd
PxQQ131Mo35RNOFaY7u7xiyNdK1WwnTirT7nXTYMfKl5Zvuow8416r4W59kkk84sFULm67medeK2
69HFqtXVhwaabh9yezlUdRz+tcyPL2Dxu12ePvko8WfM0Q40oF1SjEmABh4WiuT+0ZqZDnQUK5BD
tCeBYDxANPC6ynRkENw+ayByVCP/PAryodojJRPtBkaOUyTKTYQQmVzX/XDOZow9zYrVf+S4S4An
0zuyz8o2FxA159VbmA62VaHwE66OcvXys9miRt0M/wB9RSXhnAt54prKxeeOCgz0Cny1YUjHmwX1
uMsEstnoD/NnToZDwnscF6DqM8W6DEEvfzBQpzMjHeSFZ/R+ldW751l/D30TD43Ffml22zNWR4yT
rLvR5iq57HTGyQaO+6Tf7I7rxurfMkHj53eFd24K/Zy9p0w6nP0AGzjTxpf4SeS6mekf2eunf7g9
vuJDSTKknsZXUurod7vGzta4AhMLHWyovAzpacuWA7OAicMYZQwSf3H9aw/VOC2bW3ypaog7tO8v
7fRGCmUNCWtNJeFyzbEBPJSOgBqhu23XAhPcCJG/02PNlQ4dWgZEpyAs08e/tYUkPm9RGHzX375R
OUfrcY4KADjz/JPAboh4LCFJQYdoksPcRpz/wADquYiDOZI8hGm5i4Te+E6QCerMUnqFl7aCTzX2
AzBN7SyiG6/sF/1SYdYxcwp1N0IpVk4R4iYzPRNzYhBhX6JKEDvemii6bhnIcdNHEMns38mAq8du
6sK9JyTx9R99JmWYniz/TJMlxiyxIpBUGALT3KcU/0WrcYf7gVoJv6Pt3pooDJL8p9Sz3yww831F
pMB3oVSJL+5J2CGpPHf9lxGdghquan58RvH7N/gqxcGJA+QEcWPkyEbHc8K1JFqDIFotYPP4rE4l
cyHMePxYq0p/43b5U1DLO7XdXITUuc3DFw54yYsnU/wqpr664viQ+iV6V3lWCkrmq1vBDoVC4UF2
Vri7VzPYFIkoDKCvr4n4sHW7CDDIdPr80whr6vAXizjuu2/TifEe3D48J1azC7TIXZCatu884XzI
Gu1cy7otmhT61TXNjz23rEDgYdSawIbGnHHlTyPdKPXm/ANCenLxMhNWrHROiOn8DVuw3QK8eAn6
+CM/esuhBb0xfG2mQPon4tCsg2A8cJ0y7nb+JvENv6JvB4EN03sk+amQ3rC1LsbygJGAsRiUVzXU
g/ti5n0IluLiMVlvw9tWAS76uWV+CViBsThRZ+DFlpN6hveq0g2e8hh8FWYsgc5en6ipYP56ttpH
yXLp3A94vjxyu+mezcO/xVz6M7WLam5JJ/SQRrjAl3UzEVZplaX4pVcE6i/j9B8jr0ODNF/pFZpE
6sClK79GEH7uJOUp8S46f+sCM5hTTvOdXLG9QALXCI/bTenXoMj0Bd+lMru4bpG2x+oN5h/PND4Q
y197jVM32A1lVAiKLM3N76CqkyWntjV2tuArMgF7G59HO4d7KZnS1Gl5Qu+PUvEFJwKFZP0ym35g
a7OOz1HMRTXO05MPRC6wZ0zkWVIWavJjQuNl6AHJEmA6qEMq6JXXDtF872BaF4nUL8zAnYavNTye
6XxTJhvBnLcmjV9OiZFJEJijcKo6XWHG9V6QdKJID4qGpHBysaPHNM4b6Tf+BPWDGObRWbNczpzF
DhNu8aZJKY1+jy2jDFSZXlgrik3P3XzJcpM/kCXqMH/oBbJdjzyOmVTNpBnmJ0hyCi2IDbRnrQ+Z
7lP+mHdf3IBqg3C0yCWiiJOUa8g+d+wW0A/HLUgOEs99oyXbBz0DF3MImquGXEpTE7aF5cGUoZhQ
644BOKl4hIYNR4LD8GWCPGX4nQhqDfxrbq9Q3C4EnjIwql2DroRgGq/lhdFm/TYAGTlq1f3erfdE
9FZaxomvset9I9wiLpnLGc4gars0HflCq3ka34eneV3Rjbp5418UcWnau4uTj8KC2NcMX6EogwkL
gXqiFMd6jizADOF/IirDFAD9elXKKc9OUjdqASR+ZlUJd3EjRS6MFfaiF04pWO0JhO9qiarxbA6a
aUiq6UyFmj/WaoI0xI519XO3qb/5hTI6pe71P5Iiepovq6nFVhOonUvru/n/blLqZrDAWUHh6k1h
T0C53w+xfzjrCIWQPY4G43TRQQ4rVrpLn16Ht0Od18+0u4oQytNHAMjMoOp1p565Ebz7xhx6jToU
aaPrr0368qfTctobHV2bQVomwsfca0/2FRt4x+g5X1bv8Gm7DzBdp2k97q95NqHw9akYJv64QneO
frApATFOPNTa/wX62hLWqfOMwJlJSyCd9hIGBGeJAeRUe4Egny3QEbUBkYhF0ufePib6FQONcKKM
rrIWLE7qv7UqFu1OB/WAEgaCHBvS+vw2/ZWVzqd/W2nScOrmA4JWNAgA06sys6EidUyR42ZDJkdP
PZFUHz0wuvRmSTmae27iNeywfDtHw3U2vB7rJVc4uTElfuG71bJtksMxPCB7rljGw/V2E97tokWg
xErBkb2W9KLxcs1Q4hOl3X3TS1hkmLUd5nUpFYDk+zk/8L+6WA9/dyka19NgFEf347C2wdgETe8v
2z+Yqp6LHkGElTh5pJTH2Q1NvHXKkzCdPLX4hkgM2Ql/opijdBS6b8uhxJ5OI2C9A3hnrV+yqXiH
D/ilxNOiiT/zniT0IB0KHDSAmFwDITJHgLZUgy2Xtx6LPY3zCOyEflcYa5Mqar8JGAXUOnq2NCVn
gTBpjIykduwrDSr5LE5smQt1gwiJWBV7U/DbYcaJcF+qN136fcyizhEI9p8OVPko25JTcemWrXXY
m3mnVE7vChzThUazy6TQZ0UUUx9FgXTc+azvWldmRlJnRw6uIG/ThwBLYHAq0Ggu3L1piGcjacFP
DD4ubskq8D04oCIiBaUw/euCy9i9m5lDbf3QdHnNObwVtgqZZmcqN63tBktSp5ny266TRSwBUEsC
C1yIgjy9l2hKoeeRCxJwkXS3ax2rN+WGDs1BsN8U2kvk9wLnDlEDGduw+1r6VPF3C7TkfwykoXHn
nM/FfIpj5LtqoxBInWr+DzJaqTfOxptsRVkPfWZvxgqXOj+jLNqTI1X9WkEJtRYMiQwiQXcP9VSf
jfOzPDfr5qx0YiIRRPmban85goVuA9Rl0g/aEeHthycCbfD4v7x0rGpSN72ozfRMTmlTKl+LR6gM
gxzWw5aRunT3bfBn9RUDdVmwlUXGaxI1hraHigsQ/r0i0+hPqlb0R5GJYg00AfvB5A/6NpRCDoeE
MgoqnS1b0/Q6VWwEeWz7wJUKTHc71M4WiT8CqjqFy1mFD0lf2U/5xEZ0B4/lHDTFHCxOJXIjfVfc
2v1REnBZcscJ0w8HHe+4vMxp4KVcWX3rjh8/NaHj63zzdhmOFoqzKb5bdZr2/VrGDginZHIYO9uZ
99P9tAQG0qEIydWM6DhahuPFNBVoH4udsiFjM8S6LL6F/ymfyBR0ffVjd3diJPV33Uro1yupmduv
tPl9mjanHHMIY+SSVG1bu7C2c+IBFRWjT3oZB6qXVv9HlaB2nM+otNN0Q83xoKsMe1uXFyOTUdGs
IjxeiB/SFjIKVC5zxmBF02SnHEhRLDmtBvLaT/ZEmbAcIg/CRwRn8mGj8d93A7/Y/s3GTYrF6D5Y
NSTs/WILNgxB3K7j+GVYvCPNiRrtdAfkeVTQyBWByvu9tjB+FICG74tdl2JMJZL4WFd2UdkkF1zM
lZl0AVxYUhJpVYABWM2IC7Op7q3YnAwCU8qVW9pDJLQ8wIizf9dADZAEYJCQ4Au9T3ZPJy6zyyWZ
a+Ah1pLH+iEllJ/+XzSnQaRY44kUiUPIbizbquV7nYoBXMBUIYYu4TM4P1s75tXY4Qxti/9gVcCo
F4ePJFWiivLMihVYjFHm95G6RpiNWGZ386E5dRGakvVL3krdFimxTxmmP5QorkHbkRqFCRzG4OG7
DlSrsLHOAkRkdelWbhrOEua7iaU8SOju5VQJ6yiCU4xgGnwHqrPUngaTphC92GgtKPPKk7l7AbjW
6EkGQFOw6CiuTXyHVEhDJt99U/Vj8bFRRAfUfGaPw+7YEWUZEwaXzKiSsZ2ikmRBtUwgB8o859mR
D8oFKMVqg9aONik1iI+/2mzeW3aUAOafUI7IkfezC/e6CnmwwdFhUSNLB+HdrApfToglNHR3zqhs
Du8pESP7/tvQRL+54PBmOCvFzsm19Gi37BNsUWQ61lUA0+Raz1oSycXaYfLV+spSCa755+1C+8QL
aThRZqM2YMpbZVGRwONrbnat4dtc6fRWqPruqOKogM/2it2/okpiE0EJ8YTl74unWMKxXGK3hrvL
BN24Hc0mp+gNUkrKMjFTFURjp7SXlvHVve9ARCZKCJs/7ymE1PhUYBeWLV7RGVwCFwU/BVcQehuv
iMqovg2/is5Y/KAZNJDZ6tqusGBZjNLpN4L1raSMvXiuUtZU65Ohp3VizNSXbPicSOHAhkYZAhg1
ZO0t9JIdvU7xgXhXbl4gEL3XDB6NKRu5+9C3SfVp7RFzqENranuaOcMttswRnwAl6bgscbeJ+75j
0NhY53z1GtGL/VU83qcF6O1dM0HNeHWeo06sxY+aK+a/shYJ8pqlglHAycgFmXcl3EUiSWANulcF
/+KXnzZFdHTpqs7yThstenbwAlclL+M89p+bucC88O3OaZWAghT72zk+CX/G8jqCmx7LAyuPV5jd
BuPiA9demketdzqw9MQofWnzU3jIMNnbiLdP9vC0QTUKt977PfaIt8V/TtWoXLROdH7UGhYwiZDJ
Fhdrv4ynzybZqawQU/qzIuIL3FR3pxH+RbfVDZF0L5+KnJffXyQKmMarih24fxm581JtwDcAk0ym
DOSD/qghNRl0qF2RoigE8ny0l37ItgSVWWTr2lYJs/iVAXrCazcSm4Gq1u12bd6hBVH3Z0XJlUPc
8nbOD1damAMuWLSF2H5g2flzW5jgGPheO57PLRsg0IQWWBRFI+kcPhsb3UWCdUhiVjQIStHBlNRk
17uo7SZkkhG5J4jeXJi39mMkdafnhUeAP1elVq+AejDhZ5phxRQAFCTQkwmV67h5PNBc1qAyMkgR
swVvFJvnFaAmS8hOqFhL4HV7xR5bM2fEg+ladQiNYTszwde46bfr98ff1J8XTAW8OwaEOZECxCgM
uE3uer6ajNJ455ts0utn+KcXR+NZkqmsAKxjnMZaNhNw/A8F0sxWFB5tGeTH3f3/UqUCnAQZZ6mT
VS14sVKdY5ysO9ScNwr1GKlx7guLnbzCxpBcrAa94iw4Q/s766wn3V3VklUEwJqUy3i/eibVkmai
TNAR+tW7zWxjjt6UFM2FzbRt3kNQmtyPYcBGPWSzsSoUz2mqMFX4BBtZYKNVuYEhHc6wII9ZGvPv
hu9pbhkVxHaVFMALG0wGCb9/MXzKaO3KFI5NGTo75m/L/Kt2INDqvHWf3GBmgeGMsW/BSQyMB8DG
inaO1+mEcyNJa6l7qhJj1wugMS5w+ZmTNdTpZ6wBrCl4ZpvIqevmvxIzut8rPDTvq5GHKRH1rmOP
Bbx+tnwExl0RC4481eLow7/BM4zp9Xmf2go1qnhpMRTn6JlRQ83nryRtyPSJnYxpOkubIsAE7Beb
kkoqpwyJF/KXoWjvPlBxZhPi7fG9ciu6PWKEBZxOmoOVeCWnHSZlV0m8n3nUfLrIX7t/za4YxH3b
PibPLur6wnbbR5ZaFzI/0g9xVScGIGXr0ktph7E6jSOMjj2oJi/xXgrVpJJatxCdui+onfLPwu2P
FryomcP9nEV8AHmcj0JasAMvljTSX4eNH0OTt+B8ZahFE+gAxH8wgy23wvvs/FZsh3LcVVzoAidj
5CZzjXwAs3iRCUgLt5X3rgZv97uZJW6KvVrVmGAx+K4hI5+4Dv91iBHHQrNU84wkCWpdaEkx64gF
0lTVL5twAy6/VRFgYHM3W406CBmWihBMFrArppO4NO9EI1XkgA0fILlEgzWsFcXzgTe9b1T0ZP8m
WXAbKL69OEdNJC14ynGuSbhaT15eFg3N+oL2cI0R6PHt4WHjGc3rMNFdbZFXkhyhUjkljSMSckCW
b/dMHmpaNSLf/6ARanac1bm+wa3Jf5p+rDDh3Ec/MM9d9VMeQmU0U0VwK67koUhL8oXSvXCS12Ek
oa8EYQj86almfE0e1RLNYRL4+20x85IfahvdCVV6SiVcPj12gPrAZiRJiRDgHra/kk9VHUXPG5N6
O61pX0qMnV/MZO4Q4tvhvlLT8qUOANiMSdwc9OeJi89aeEUw/4KVQ4b3W/DyztQlgQDP2EzzEUwe
I4OT8RVErzvDfWphRZZpYs1qQ/X+uZpUiCDhA2Z0Z+N/P913BECdnCXG0JZJeibrza8BhtKuu5wx
5l2uWRTXMBtOf3X7CXvXvH26XNj39aw9S6yFEpFLbKK8IVYnWGi2Gkc5VU8jxYAnU1zZJpbkYHQV
anO3M8NYx39mJyOyTTE1SPpOXEtPJ6q5AThhcpHNIkmF5hSxK6oXjETZwNjnA8EBIHGFF/NZgIsQ
2mEo0qA9lwzmJOdjBAOGAgs0HYeP2QNr5qbcm1040O/15g92MTsMhPUFKVL0RJKaFadf/wBDRwVs
Ph3IrRjWiVzNVJBjX3fotA0zQvpntgF3UUtApFMMqOG9fbjT9TtmR24RuHCkiDkJKw8mzzaVfIg+
qseep2in9hq3+V1w+y8FOkRnKfLFowuu4POfvcO50+nIqxGd7IFI/IHVkU0I+lRFz9dIB38VNuWK
B4Rbjb3Nnqrg1vy2aLrfrW3WP1FMaNHL5adMKaQpTQJ9YgHsFWgorfiXqFLbLTTYrfEJUDJhl1Us
bc9FchA5W/3+odT47IwQW3wqnan6n66evEqi8iYXhO6Mgr18AdNmUtHeRza5wxuBqrclBvVMscxR
lJkTDSvJbbX5zlbl0cMesITnSzakqyYK4wfgoPWl0+QwfF/HM4yX++oQz6oFcxaZV/L+l+n5lJL9
YQNBpsBOg1qI0BOR25K9FDL5zg5LjbruEzPGrvUJTx9ttcwff6eXgxn6K2rub2p8veeckxZ89Fi4
vix1zr6nUpYYFkUQ37tY9Q/4p9bk3gXMoK2SUDOKd3WcBYu6oGTHXo3GSfUoJUZxY1MvG1+pszV0
nxGqaCEo2TL+7YoVeBqxF0u0lijt/2CQIjER3VNGZHNdYkpWNY9KF+GX9UV/ExqGGH4WCPBvRFNU
LscLwDEAZPHjsX8bQIl9Q0OOl0Q7cRgrytCp8jyuYtKkYKYwQDKcXMm+13W2NAsbqA4qWlLE3xe/
zv49ZwELI+T9J6dPoyJ7LrwDMPXZMjscqEcG79vgrDzAaukKfwfd19rLYQU4uRNzcLw7898jFKjF
9Ct2TLkpf3nQ2KdQliM696+pke4ADeP9xiuZrct+JjTjwya2NATnHQuHz8w+Zxh5eaxKBBALttTj
Ac/R3F4z/UIGyZyXQ3KSAH5COr0ry4VdPe2Dbu1Qtbwtue8ZPAGPbHb19QUlewxbu/jP2C7ysF5a
AH2tAoaxbthuWP98JZ0UbOGpPmCDVUkYzM0G8ZZTGjp3W3Lnz/Gn/F23IKcuO4TZQsD6GUDyk6Dy
XAVb+RFkRbxNefp1oaox/7SkKPy8mjSiVbi8awHoyW9zZtV6LalZ5xozshCKcFQypUywEwBU617u
SKMLRtfrZYbzcXTudqgw0diazvXRRA1Rw8HYNWurdL43rmh+BnC9OcH6LHXV0cJCkmgaZvb160Jf
GvXDcN6mpykY7TQd/C3AvblBBw3znjf0AkvFPphrp/fjg3WXGb6vqrVv4u803Jej94yU5kkmy4GA
etR/mwterv69ct2WGCn0r2T8AROuJW0BjNIkmDOBvdsxL5Fpyy7k+o8HlszpBV/vLARNZQoxLq1h
p5ZT16QlKp7svL0VJ2E5564Si6IYEcIt/Gso6c4+mcHSXOB0la+dtsYEsqMme0Zamz0I+2vDt7Op
6QGGln3hrcWEJFC2lJztuUIlQA46KQ09Pb227HzAxgYTV8GJdqqaUZKmfCxSDVgGpF7J2KOH+WlB
TK75sAEL2Ho7wvFtjthWjnfA1bIfNJHjt9DFSF2FLzJX/JjCfagd/S8LEVhPn1daA0LuZhWXInjZ
oxlFlzCESvWdKFjm5QLHqNfQ7yKwFfph8BalrylescOwss+AFN9OIu4sGWkFCna2kO7Sz2bOom/F
SRvmha2tixlXus9tffyHdQo6+YTkyYzqQmbScXpu7uIqXVynPAGx17+6wPz74RskVslQr2aPJL++
n0A0Z6x7u9aW4NuYGDxTm31Ge2KY1uHThUQMxhAbU1imLUKe54AdDBgYJgUr6rhJRNVRBNguRwF7
oGcdq4zQPw26DoDcj0WWUAn5szCvdAvYGIrsjbBj5ULZnf5bdGLuCKhdjLYdCWPUiOI3xxa+V2m2
NbMcJmelBJm1uP/IR+rxCRiQXXrgOTod/Mca4PqwIi1clR0Ara9Z111rmBXeBZ8H19aRvNv2Pp67
ZxLblxXYsNM3jhp7B+h4/5ngkwpgS3M7XeyU5ARXb2YIy87CEGvaAvMuyYFiKIkCOU7vtZCaMb1Z
nPTdPjtjEr99lK116sHZW4tqFtYX8oEOYPXBFiKA3O/WRMLluKpPwg663TYjsLlzr2CAo8XRhel6
JG3oE2iIfn3dvqZJxg3Sj/So8D5qNrNQiEd1LfeN6l8WIDY8bFwjJ/S7axLLJn+2hbB9N+J5mjj/
TL1xkWL0OnKv2e0QI9hwr0ifHmRjZEMjW69fvdzEE2TKwV5ATCW8Xfj7hBy1AT6I9DDVikOcAL7o
sYE8hkvZTS2mdWt0Oos3QPMSEkdxPW85wCQt0wtq2tZ+v0Lfif0eUrN0cLxW2OoC5ikf6VOXfSPD
XJ0Y8BZk9ta1cAx/DZ0iic/j/6zHlSyGbWr8Vp69Fsw5iq3soh8K3f8MRKceAmw99E+XLEN8OalH
/kYnqLNoLQ/GXMKH+fm7zZ0PleDj7WUyVP1doIkBStZwmM14cx8GlHsm/kvoz9zbMJjNfIyw7qX0
iyDVEPP+gwplo8Pu7z16/7jGftTTrCe9h3UtjzJBQlaUjzgBxgGuvX4sSC1Mv0IzjBGRP6E7M2BC
WSxizrmET3BBBs30rr1W7bE6Ox0Cr5Pulabemoqj9y95CzFaE58DL7SDBBBjwVcXwtsbNeXdrFnD
kK2PIxAmPesAxGs1MQpfrBua1cTjVnXyTIxdhbqfZ+5KuflrdtL1pHzvpQdN6Rmaal5MfK/rihDe
1B1vKgC38Bw2ZWTyukAg0TDIF9bvt8JFK7KEPkiC+uo4Fe8lrY4r+Udvhl8zED1KWQ5Iwwde3GMD
KudDiaa+uOgY1ELZc08D3yd2cOTJBX5DaY+7x2UzNRm7HaRih7bkyqI3uZi9UChmn5MLFwNtv4iW
fswYoMMWMqaITQMdoG3pI3ibaLztvu16BFcqGRuMwsfwg3Kv9A2Svd5QlwgsBPtXy/tLy3P+xDhe
VgBUD/UVXi41yQWz9yZN1pLVMO5+LWwFb6cHjqeA6uuEMY4Xf8Bg3RsZ2FAJ/T9PtvhBJFkj/8Bz
+YqpxOegvVcBaHXrmO03V0jTitQEnVQbQbRDBIt8f72cI39he4WIGkx7p14cWIMtkYpOjmxTtONN
QLxbHSZEoswsD++dlJRdC97Rq8GWAX/588sN8Ta39zcO3Kgd2Fy5cULNQXN2PNmw06LhDZE1aazz
854QnlMR6ML4YRcOEvuxYXcrosSiG8VC5gdfGeOyx7rBjyBu09tmaGPukq2LHGKEP+piyu7fMnb5
eSKHDXgr6qybYhTy8zUCRAJUYAfJlhkAzBo1yjU+jiryO5nD0qZLPHF+2z0WwtvWYAl2K7FZUa5K
WaorLykAhzGNsQaw5DfFQjl7vOoiGOr7ZAGTovm9L7aCduN9q01qe+j3ublBX7YM1Oh5p4G3A3p+
Sfci5hAonbxFrw4qLIFWiX37Qxu23vHCOLhMefytLl/cimrvRVPAeQ==
`protect end_protected
