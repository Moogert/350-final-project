��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h}�iH��ẃ��>��8p��T��O{*f	���I�Q#a��09Pm9`����D��=���vJ������f��jb�_Gb��b�NX�J�H,3��S\h�;��R��ר��=�diZ�3$����IKf��Vu����ŀd5e*��og��t��!�n�w����V��Q�u�Tڮp�*>\_@�W��VRN��x\3�l�A6Ss�&���p�+�a�Kr���0s�/:'OqN�/Κ���ڸcQ��^O�ܖ#>�f5��|i6p��r1���tV��YZ ���ΰ������਑�&�8���L��zI�����iP3�p,Y�����ތ�^I���l^׬�FҤ�$D���Ѫ�ç����N�Oi6ա�\3$f�t��&���ʲ,��"ҩ�N�'��pF�ĺ+�����eA8C�����aՍ��7�\�{S������S>��f�Tk
�yQ|�o�.g�>�����Xy^U�I�	Kp<��}z�1��};t�4O��%\=?��H��P_^�?�3i�d���k*ȓ���9�֜,�yKfyp$�X>jD��qk��N
��J2��/b��7nچ���eEħ���?`�H�H$��v�֮�;r o�T^�E<���qH�$m-cj��&�+�����_���"��x)ܛk%�P��C�x[xݚ�����#�O{A�_ٙ$i�?w1#R�n�N&�/��'ô���W6�K� �	5��O�]��>x6(i(�T0t�<�P�z	a��hq�9w5��y���
��5�~�7"��.V_��֝�VI+�@c�(qm�y�U8�@�O9�&Ye]msl�q��!R^b���[�^b�E$Ƚ�����=2����s�Z��tQ7��d���b{��r�0Ѿ�:��~լ��$�lP�A)@ۉ�����
��2����/������&��dr}��{Y�+���cp2�R�?>�<�2����$���%=�?�$��q��_M;"X_D�_G�]/�J�fVJJ�ܹ�~���B����߂�!�Ȳ�u����ɝ]�BG �dK�������/?G^���S�;y]�,-�c�v0�6\���*�\mCHK���~>S���wf>7�xw|OR�`S��>��c���>�-�:b�5�|1axvChSO&���X�&���^�l�iZ�g��l�X-E�|�xX�����J�7df���R��B� ��b���^r�X�6!��֣�sx]v5�w��D�Q¨��z�K�<۹^��ťj���C�|��3E��g�f��x�\em�u|����d� �SD��S�V1Z������r����i%��gʉ*'̝q>wbv���y+�i��2B�{A��W�:�DL�d%���<�;�̙�|�X�"���^l4 �hȶ,���~�u�,���ǹQ��W�bb�fM''��8e�

�Y����:`�n<��6ZJ��7D�lE)�c뺑�M?���RF�V �U���i��u��u\���G����ygߙx�z)�,}����ɾ?�:�Y��{-|�D%�A�Ѵ~.-�o.��tm(�`t�xwh>�B�NE��Qh��A�^�0��������8�8�#s"�q����³rx͠0=�>��l�';����k����6:'�!�3N��vѵ
^A�|�.җ�*����Rsl [�w�% ~����Wp/�vcl�I�c�(�����+4�����F��6[������2�L����|`�� -X�yh]=�9'�ۆ�|0V�hv3��B��\Y����Q"���먱b���Va�j[?�~���]��0F��ߖ�opQ9�	L	ã�m���\�za��wVk>��#��P�a,{�S/�Gi��G|�	��xZ�a��ə\�5�`����7�m$�z�(N��Yg���Ft^�EVG����>�!������Ҡ�d-��	?Nq�{���8e��f�+`�oۆ�w�ᐮ��S¹ņ�}�4Zn�\L��l`̅���h7|܂EC����:4�W�"��C!n�+iEpA�������ϐ��dO\��=��_0�wK�]�w������|u��amoC�3#�CB�b8=\�aWc�Z��2@��z^���j������4�D�k��p��f8����b)�ʈ�����EUc���/� '��˯��8���	eW�{�T����.Δ��"62�%�ɱ*#;8gOMv�k���v7&���E�=�<��LY�h�/M�X���r�����se�pPJ)�6�͓��&(gamȡ�\~ٟAQ{6a]�&"| 4Y�e�^�/	�ؿV�ά��>
tj92����(���KEx$(n��0kF����vP�j�
�D���" �V��[D�k���?]k�n!�p0�nsQ��\�z�Y`Q��G���]��c��'�AfW��S���Q�r�`C��3����=��W���GT�5�A�ǚ0�/!����ξl�s��%����T�O��{�{ܚ�Oc"���O��G���"k�E &�p�����?hqw�u	��+5����1�.�NK<-��/�L<1�3�F���fC �Y�c�&����S9��hR���['��c4G�;T@�KH�"��@ܰl'��_�~BP!mN�i�S��A�P�gI���ӷo�z��}��=@a�K�6v&WH��qy���]g��`���=I�ѐ�@���t,�c�Y�&���H,�O;>�t�ֻ�Х3���D�ag@2z.�A����c�u�?g����,�a��<H�>����*bo<�(2�B�ޓE�:u�snW$�LF��� ��Fd��MCܘ2��5��Ce�+Ͳ �T:h߯M�[�t�>Ң�(B�v�*>O^�=;,%�l,��7�dD��v�Aײf���\�L�� �=G�2����o��O���v���I����i�1��G�0�&��[j��;4�����	t��^�CT��Mgm�U�E,8r0Ʌ�Wh&�垉���1�>j ��)|1��Q�V����O��2�j�vɣ�~ÿ�Awa����	���e�fy��f����[E�P�Kи�˕:1:�`���kO��7�/"�(c��5��b2���9���{�X�Ntg���Wx<1�]4wr�81���f��V�̋�m��PH��ð���F�I�AT3��Z�@u��D�4�`5�	��`�c�ݞ��Z}�=V�!�������������?�Y}�0o�[�����:���:#���|��I.�)�����sf|�x)L�M����C�MW�hb2ڛx.��5�x�p�Ԋj�a��
������'�#n���Yqg:�K�8n'/��2�c�ꏎ?&U���%�	��:q�A��\�j��i1�1�bm��aj�H�;J@!A���$�+5S��b2K�����_d��?ۻ�d�?,�����E�����d#_���E�=ϼ(S㟕?T�5Q��G3��mp2VE�A?k�O�?��.o�+Czڝ7L�I+�ZB�'ot�Faa�v�f�$��i���q�'����ٱ��N7�uk0�P5���(	b�JQ%�A�gF�Ϯ{��r}@�g ��A,! �lП�z�5�̀�V8*���\�cq!�X�#	�����<|~�[E���bz��e�5�/p��LQw{Q9�;L�Y����i�Z��7�ܖ�G6����V��պ����ڴ�KH�d]�-�~a�W
���ݧ����c�O�Zۯ�P�<y��;������n/-=*B�]�W� ���]�b_'��@"�aW /7��(�dN�| Y�����3T��h��
F�[OJ�Y2dM�@�Y�����A���v��;k!K��p���M�T�E��i��G����3U�׆:յ��9d5e�MbG��|�xU"����M�[fw]�t&�� ��'�e��3�/7�h�T�����#�U���mA��f0�~?LB��p&(>9w�7�������|�Ymj� \���~	�A�_2��T0�Y`kD�SX̀6�i4�����^�7Ș��oq�Y���F�Ʃv�	�S���'�7���\��f���Ϥs8�Mĳ�h�7/Iv�H��b˝<s�|uW�눢I�1��eR�$/��Yq�^7�4����(��7=Ou"-�r���P�`F�8���y4���0���@��F��<�ܲ�*����kogX��y!�-�$�?�E���}	>\��8z�L�8��!�z� oՊOS"����%f�k����z�i?��J����]f�B��F��;�
����������S����c/�rs�V<a�T�d���EQ|�m�g}��#��x�;�R����6���v��@�͉ᾩ���Fz ��j%�qa�Se��+�IP�/���?��(p��
�<��!��*���^�7�M:k�?e�ҿb$a���ӹyȱn̥��}�.�ۇ�nU�U7�ےa^������� �.[���9GN��ݛ����(�K���t�C>�`�������7C���
Ѵ+���6�d(/��
�y�<)�O�~g�����u@zOG�X�XW�Q+�Ⳍ$n��]W��n[�V���n����Aԑ���4y_���ø�1'�]�	ե�v�(�u��QK	����" A�7��SWC�X��<e8`y�e�C6߄ hzf�8��
���3}���r�	�+@��ΈX��?[��w���R
����yi�|��"
���q`?�uG⷗����,���A�~��d�����c���?����F�o�f蒚��y���_�Ov�3�=_z a[v��O^�V-5̀:>m�QD��U��C�r�D"��$j����l��6:i!X*����ڤ��j���h���{,+a��3a�O��L�o9�HJ)�`v��=�����%�f��.ھ�[_�Q}ׁ~���s+�b�D��t%��!=�UR5l�G��ʫ���٧d��I����s�wS\ʁ��z;��u����~z��d��#�+)�bB"4�e��á��'Wv�����)V7�.�e������X{�z��������hT"�J�+�1L|��4Ax��yɆ�Bc��mȯE���h��Ƕ'�^�_�ULdBY�k����1ղ��#���Q��[��|�_�P�P!���˅� ���L�Au�<-�����i��M'/]��Ϭ��ڻy�W����ݞI]F/[@+���Ƭ���8�[
C���[���<jl�Y���%�049o.2w1+L�:I�m���zf���I��Mc�(��L�t����Į/����Ͼ�)����{�(K��l:\;�61^ֲOZHh���s�Zh�*⥔���mƖʾ��󻗟��z�@t�#�����ts��b��^b��Kt��>�r���:۱�T�(�S�� w���Y�}�hB
^[���jK@�NB�|������Q��2�Y(��J�Xr��G\�s�(�:,�N��C�&�&��I�.��l<�?(����"�8[Q���-l�89p��a bE#A��SZ���h�-7�N�A f�_q����&�?$���&����9���  ���t����4�!��7��Lf��%�S��a�SE2�W��FN��ZKO��UV�s��6��x-��X��mJt�]�qP|�'�R�־�%���@!;����[D#�Ʀ�x�S5��=x��c�k
f�.�`�7,~�؆��U#�U�(տ��5���U�<4n� ��`�e�&�r�ʤ�'2��>p~��^N��Y.�]BFkm ��z���ϨN>�V��]ūU�
�h*�L;!(G�ux�w[i