-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IDC+xBaFnQ6HoKAYb5I+ZMRE02fnNQf9YqPsDcXkP76L+01yUiPQPNHafnazkB+CCyfGf4zYylHe
e3GqZyMDa1TwJct7129bJgdqh1ocGcw8dzcvt6sCYudu7yuXMYNh88QRUqnmbAlfUq1MbESZcLBM
IzI8jbXWqHsH7UWjpo399iDsOrAMnCYYHDN0GGzSk+/SJzgCzOeweIlcxugVT2UbB4MQUlub/G2G
zZOCpwuOfZbvq4B3zBw3dpKH8O/UXF+XuCnU/iGp4SfhZSiHsm8s8PwledOBYadGVrlXrIg9wXJy
hgUzoi8Wqto6XigsKLK5oysWCqytRYn13oqyWQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
2DmT0cp7liuDrty1ASDh2aRtZ6PCKtTDtXkeHkSsTYXKfTEncbyzANwblHaNswjLXWOvUxUYIAG8
c1k7txeUgVIHHbqfWDiJt4MqnC2DVnBbYZbS1xBi3nWNJqN/7EG9tNK1GMJbNivvycNmajBqtF+N
Vez5AFNbHxAvFhUosXVswhRD6/D9HXsctm2pJI+KcoRPXxepI2biVfaAzN7RiChNdEOX3BNZdJGc
iFU8KOAN7lEYOGHD6f2cj6dWJ1SIZ+9C0vhmyuC/SGmFmjCVGt8dngp3T0lEgq2P8E19e5xn+i15
eiw2JLCodMb4sV8eIJCNA+xujMOntstD+3tIb34a+RQZd8l3bStQ7mAP5McXB+YSv1dhc1Kl97Qb
ftrtk9OcRIZ7ZuIMv2W3khDl2i0LE/gNjNGrCU3n7STO1Y81JvomPW/2VXmTP6jUWXGjlfcrZaT8
A1FnjRJ0XNoNAADmqzScOCflKCNT9OvURVELr9hAdnosOSU53VXDAOS89cfHJmCQ59dJISSi0853
8dNfB278NswgtqoZmZ2eGo87Jgho7u4hkpLnKS/+zUMgQja3/geZs7ClRySLVkYgUC5S/LoW4moS
pdUcXHnRxFSG+2L4Ow7dAHCfwLxZZYjK4dmIlygBEDq6+B13lAVO9YRsyYgPIukzkfc8mqVaeXf3
R4CpR2+7WcFtCj+c9CVA5ds5qXSkj0rU2bXvE0dUikUdG3ol8v/q6GCj6TkieDZBqxE0RcLuDAaD
lC7wTeg6aO24G5woYlwD+UxC60BTt+hgVOIDHNzTn/tHIfPRvZhP0Xm1dDulxY3DNOJZYw/NhgMQ
mb76ofX6WhYADHUXM0ks9pJbfioofaEdwDGH+QrUg7q0on1QbgOdib4sHPZ9sv+dIeOztRTPRoxS
2dw/fU6h7VNf5SFeWOitC8DqP+UxHCzKw3MyZaIk3rEVh0ube6Odv/5MORFNen7FPU1FQSyQ7WLw
l9ZMNeJ25lBdbABDG4SbtGdN0naaEjc9O8J2BTnvNaYGrmPbSPIOD66hlWhqXN5IUaW/bbUy1JOP
HJnnwGrQaBMMgOikkyjtDr/D+VDfGjA6aCzk1Sw8DnuQZvloY05WQWPg0qdMf5HSCGLEx8V3bxf0
4MXbNTJFS2O9J/wcBix7ewtEHZvx2gDSS4Mh5nzj+UXkmlxs3I61NFDhcNwzODH6wnIIatCXf1M0
/1UQIJEUd4c1V7iHaq+qJewpgfBj5B4RR9alQokOJiP+ruIDesvZROYRh2MeuBJHjoUeYFUdOkne
T70Btrf06Q+4nV3SdmFw4DxO/6b8l/eR0oYcsA8QC1yv0ZDZ5rFsx2U5f8UnaGb7/k2akkW6vwdr
ZFsanyMava5gcQjnVFRqvLUFxNlhux7Si9SSYrTpGS24b+EcxXIiOwe46V9HfXjO2zx6U87TFRvx
6EI2VffnsfNjuvTc1hIUFThmD+vx6kN8NDb3yDcvV4XjFrmE1tfuZRZeaOBovWPFapet6eiB5zwd
ojWMj9GX9LXHw4nM1OSJarQNisBMnbB2TXEr+zx3ozoRglqKnA57SRxRVE2yElEe9b+GL+tpWWH7
VZ65cqi4omXQgJA7NtHJZz9YB+zcEfHfe/qND/Ll4YO4I2C+5R1I4AZlw4p0I5ojZWE92DlXYYhU
XX790wAL+fscvS5gzV0MOByu2bRn2nUy+Iv9IKNu+YnsrYqSnnNom36jibSgEdtoRbvFjcnSA1VR
jguAXMlhZMqJMcxsyjT6ipPbhVx4R7ZtHJewRK/o/3hHOI7Z6TF0Sb1NFqzNg5xnHH1oZFK43o4X
ybpG1Zm0Q8zQLZTaD8JWj1knTfh9c78+1TYtHeCDiPcJ0q3/H3eNw0MH34/a+PxWna59wvzgalo/
iK5E1hB5dKtwY+WbOVc5ComS4XEGU5CAoaOWU3TlXpnlhyd3+HPGZiVSqBv2F1z7DTCHe9H1D5gF
XS0hCTV4Iadww1HTepDluI2nVAgZFqoAEXp3+K0Vompyfkh2zSrBPnfPJGj+mNvnmpU0fc4O9Cyn
+XIJzGGhR3rCfhV5FOM2jStWG4oShFq+MmmH7mAyTKi0ROamlfm48snOEdjtTcQCAaMfpWckbE7t
kyOuAnoNDN8mEQZvNrQIu77ZbTJkmplU8cxiJMW97VAyDtgoeQi4jDU7J0siRB/aLp+OLWync2UT
ozW0Gr3gIOdwG1+zXropCzbIZYmEsAMh3EjJJwP+JJNWwmamycbXUDBwZ20tkH9ncQ4uqc+eHL1l
QhzGGQ0IQObLbPNpY3n2UX6nDPaR65WGjcOq4/zTi6VoLhfd0Q/AuIS5jAe1Fxewp9DbgMc7R+UH
33CQvWDYxxcnxf2ZqaeKSM6sPll8fy8l4dKJypq/Z5OnuDKgoQPF2RWGWL7NvT6blBRjzBavv+EW
Qhn45LBUC5ppWXiGJfEl4YRCyjKfmdIm2IsLfT6WIQAE9aX5KZIq6X6fEhsb/3LMfiBHGj2HZBvv
H2gF4hQyBUVvd8hi5w+xwHQFGQ2uxeMJqVjLnOR0cR+CQ26k/HZRJv5CscKzHVF8HBP9UFwjmY7f
4/QBgjiVQsKumIcRh7EPleZAaUncAfd5jVyTJDPtO11nMDJd4KUbaaCHFUh1UwtedENCqv8iVPnP
Av8GI11OZoFYCpGFcV0mSLF9427fHqPbHfNLCrsnS2QUNupz4zfjE0hHNp3etTu3DJ+2KO2im4p8
W/oOHkt37Kc8Zjc/MUJetP2Hewj4ghPN5CEh5+fIsdWZOVO95WGN7BYMlD4qFOGQtWyGMAD2Zz4d
NpT/8CY3EJvpFoQUob/SOEiPrwOLtDe9c41QDe/0om2qF4puzQj6nztxa6zk4+9t7L7rFzSDOspb
eN4S7j74lbs1pIk7xxKAb86/RdGgb/H4n9ft9xhLRS2R99wdLp2HjadzIqRcEgJY5jouXkBHpmtv
wbE88wDeHDVbYMLwg4w0b4jXOWDkacgjK+rBAbSqhH4iL9N4NsiaC9gl6ebtl3EBVOJG48v40Tfu
/UMx9Eh/AGf3DvRx4ZcERZaC67VxGm+r3X45Zrr17fZ268rGFWf6xAT4ciq5dOr85vy/BuI2611A
NXgF4w721HHzjFyunzJVwC+Bas9izh7UbrHaGlKDQZPdK4tCbZuPAGPANlCTmH0ABihr59laYPi8
BVvQEvaINTjxLLQH+t+vPkfKkdUt6mwDgCgbD3LHb5iFWTtcZjgGJ1MIgkOxpniuLfqQkw3LGZ5o
GuY4f/iD8ifsnVEwLbDuLFVRavgx3NjE+FIxXEe2YHAwfhVuf12MQQRSAOkN17hnvoArWOi5Gbwe
E6YgcgMrndV5hZv3marDRGCSqpBrL9a+U1KY89WGf4sd6FvW5xeOAvn3Thrrxgolh0Wp5nBSdygZ
h5PH7e40cYiivYGtP+WcimEKIty18q8ZCG865NDacwzEtb6bDcop+7LGGrX8+mW2+SDkyH2x3IbC
b4T1ANccyhJfdQswSo2QkGedUlwwiCXWK8YB0Ypi9MiFol2iZFGbCoHSq0DWKhZsMXtUtnInXTmt
PBEkU2924cI3G9+KqmrzcWpHtWDSK6BLA18w3ChNPTE9V0eYxandXpwpijkEBNuXbbdlvr5hEmxE
3UqSfx4TYu4/Vlx+5GToFjJ99ViH9/OPRzEnGnUh66CwE5fb2JkFlnE9ADGnSyFZ9eO+/dGio5WM
nO+2cgERC+DjaEV+pYEvszmnx3bC4zmYdryTISzlLyfthissFemqIbXG7km/FTtG26OL8U6qJq9D
ABWR1iCIE3hYsIILmq9vmAU4qFoP4egSUVqy4BYhkeUBBBl1WaXoyDrXUCCmOLOw+PIbM7Bb0DqW
j9zeC490Wj4ia4nx/XXuxr7qhO6AQad3B3roruLRgTRcoWjxXrKAD1HH5HDH2AkmeyK4VzWEPCpD
czm9zUM3u1+scggWT5n1WKByvvsj2cFVZtcIOy+60q9hvmLkQIH+Htj8QmRQ9n35XdS28l4Ecv9F
7h+5b3emAK5m6zPlhG71+ukSxvKuJMH1eEG3/Vq3HjjHzH/0P5NPx0hf9ycTUc5oeTvM8kJDabgh
EJXIqGAmmrqrdKMAMoJbHV+u2V69O533CFXZS8+pyWDyAufEYopC5Q1/+MnVBVSLynqStMUeVjJz
ebVhihXn68W11lqzZrffDq01iaRQgWtsUHADx4Di0ZlRItLkOipLDJQQJejt5gpmdhXKXvJR0cwm
mRFgDsy92vGdUfh3iSWVjVLGZDFW27XkjypsoTNkXoeqCJluybhkfeC0W/jFGQST8fSCNl1l4GSI
Qftqe9VcJW8WD7hLYLb/P6jRrCONOcMJDB79JED5dlhT1K38qY+SJQOeSP7FAd7XLSFxLgucnTmR
0EsR1uVA6R01X5SX3qV/9wIGeMR0No2qhLB8w7b5dXchMly1lI90ZnPkmC+oKlnDHKU4kP/nkTMy
weIVggC8K5xWcAhA46pHhG96/W7AaTBBcv7zBMgjI5YQ9uiAboLj230ibEX4S3IDmEOuAStNgV9I
N8CNKKQ7MaahU7IGgCYHr+oavzBoHgnCNvtzYVNUm5PdCXbv8WqGwD8BuDk2krWI/cQIhHSR3ZY/
GMfhaSOolbNXHLS4AtmrYjWgjp9FSLk1N99U9oBxx8t3QsonC0LpyWDV+HrRJ/a14o3pA9d+qgL7
OcfiIu4aVkUFcp54sHLYoHDKR7F+o5Hnx5b6ULbHIH/T6olY9RWzFOsRm2i4PbW/uaQ1mRFX2wOJ
UTipd8SYi3HWjMlWV1DbmIu5A2A7nVlDx0wYTCVCf3IjzoP6D+vPhw6UIUPgdLprOILGyg5zlvzR
6QPvWQUc4RVlG88Nw8derR2syn5813GaanCu3xwhdXOognP6riuuyyCv8Ke5k52ADgq7bv/0qxph
YrBBod61fMoFYTkh6eOGqZWWF/KXNh5tkltJujtuCNENd/IHHn5RNZTBHuF3CiZo49vXmSDMOzJx
qG0hPQAziWf9z+MYptdkZE8rGIA+bGREyV4JZsLyP4YwxFCyqmEw9XbEhg/muASCEE0STdRz2IKH
HG4XtqF/VNyurQLQeu7B8EyQXmu0CqE/FncnpvkjXsJfAcjRTdoeZ6Sxvm892EtbY5YeufQjqf75
R4GoRU8cU+oG6d7/IgC/hjfVyXI3jHKeBk5QIqA4ynQ9cemH0rZ2ESZ9Xmc7tRJ8jHu3oI0q0+Z6
IVLFtOnhScmm8psoC0LPvkiFzZaYn8GsWRPGT0lSY6lnShE6MgsXb0TWaJ7lutxITrv9bLlmlWUj
ha4nTWPyJdn0Q4aRByVvQWUo08hm0gHpv++d5juaW2Zdce0AnROQI5rQ6ErwEWm4XDoU1E3RClLC
uDTh6OpjlcBMJJjRk0Wne5vMHTc55vFQi0Er+RAT0iL3V+68Bl8uxJSaoV88VUMLAWI2APzADPKW
R4NFuq0QzHp4TpKprN5h0xrEQvuCjzHyaZdhyieGzTZ0Fi/UpnvBSEAze5HKyPWRvmKAIA3njbI1
vQ2QwU9hS7suLa+oLsHLLMcM9hJP0NaHiAJrytIlEz/ZhYm9MrM4PZbd8ory04SGX3dmueh2pUkm
Q01ghi+ERfccCN43cO8z82wd9m5c2eKvdcI+56jqhpwreMF9nMGaxLGwSGrIwFkck8kk0u6TvueB
yJYAfa+0K2b3rJ2uMrsitdjjf6porVdxvyq/EdoSEgqLEzibFH+CgT1Eid0ANGyxvsdpIr9ujd6K
vyK4pjji5WpZCYpEryikZVlkV0Kf1+A02U0heHHLMWTp3xq391Vo9Krx/7yOVDKOdC3dgslaSAAR
+o+y8m2Ts/KceqVN3wBlFFZugvsCOmp4Ne1HApsBx5MKUD8uVHs14LtBEESzMr/gEfIlUaq99uM+
5LI6ir8YaxGUvIXN+5CV+0uBoC9I15AL38XcNPxo2GpIS+uY+IfZjePcqJQGA8EHlcKiOMbBIYAM
izIwAGjyQNnVJzcx8VcxD6y3YxOR/4JniPz1S+Ee2feOffKbHOjO2CdcItOIS0PctpsJ+4QiKGQq
k7rc/NCdux+V2EfSnQ/TjqJXUenyUqsF26L6u8rJhrLIHp7Fah4+rKktFwAgU4iHXLQYD/Rh37sO
zJJokDcLsE5yoErCURduIsQjciAvekGeTfPZRUnv6+sTktEdRZcgBCZufRQC3QhTfHvpL9fdE7Xc
F+VX6yOOOS3WIRlxla2voB/+JphkWQCHGuSTHTh10cJsdLDyH1d+c3NMLo+4HSs5xhk6xZEfUWr6
HbKc+yZwv4A0sl8xb+HjFhpg7TnT0Hd9nGkVX5G0MJjI+Jz9ZSpHoEfXGnpWHBUxwCZhJoVUfO7U
jzFnkT5auhns4oPd83w1IIal/pz9039wN7Tfi3Q8FeAiT66CpSDR0mbT+GZPcWJ0816T71EQ+NEb
kafTqB77dDVIdOUJ5WnLZsYyf1e6bTEQocuRGhe1gGmtg2xzJJG4qgMv1KicrmD6KkyOoWw/KfWP
6zkTuEm43eNtiyDltX7r3TmI6LSZJOkmOrH9SBOamYNqam7rH1/scGn1xGyjCs3T71XhcDXkdShg
WslqT0Ikgi19SAZBoPGokvCISXBP3ss3M6OTlPFICpAuLnS78/yoL3tr3eOiUKnxs4FPB1gV2VZn
5oLGNfx1W2Anm+aHuyiBl2zzCzFkp4a3RCUzalw+IDmaAtsJtgQG/bx/Y3vjPYUT85REkmRvHYNe
qtdD89cGv1MGSJWKu8g/tNp2x08qFwbGp8cspVghd/3ksPafSQbSBoLdHsNYUtgBqKz17oihk02m
GJ21S41ZjmYmpTpTcj1g4wVGm8ku5A1lUgBEJYsQz65NvSGY0Y4LOA8WLDI5n4rYdOnO+wG+j6ad
B7rXhTGGwtR098+ooUj067l+jAgMLvsq9nRQQSdzpVKlp0ZpgFdCLeF2Y0VzAKCdKoJbg+a0vVia
infcBTEn9KXIT5p9ymyhx0FFwD1v5O4L3n9f4Rw4th1gv7Rt4YKR0lJ1ucVQZmbMx3n21cpIReDP
aQxm6HItOAy+dt75pjJHSV1SSb33HUdENQgYJToQq3bnDff/6zhIXUpo7X2RAFLWAZFhio6YKVw0
qxSA38ZtxRTGhO/pYm8iQdmxsXItfFcvPXvI/0EFCLgbrZyDJUlmuVEzB7G+QBd0XnKOHB1RBBg/
Y1/cVwJcU2voXJUGIrOolN3iA1MQpP+UVaUr0RfscfGv/DbfsYbAtv1Tpisr1SiXRFFTuf+TvKGo
iflVxUelG77pCHZI7xxtnqD44nnzwullumyMvoVwDdvnl52qJkE0j2X/fnyZqOpHaHIddcsYlV/N
Y3LM6RR/3CZ3HBt9H7WHqrFl7lxjL++xC0BG5+7UqIwFuFvDnuAjdjSG0TUTn9ds5TMl43x0tNWS
KR2B772zuEaInaQQ3nLvKFFpkMQkDmzqC/LEL6rmH0FMG5iOAttwRI9tUh5TbBR2u1bksXJphlf/
JHLYYTEwjHY7nos2Bsid95SobQVTRbG3TTPYSJtwlMU+JsQCnpBoyQb87F0Jw3/lGKl/sklk3hOE
0pI3raapIo80b/pmzTUZqVn7ir5Zk1pRNioIVj/bWqoPT1bN+SxLRsFVBSPsq93iN1ZC6mj7Kr6U
Hu59WnNKTEl45ZbX5Lbjba8FTXKhwSGnuETPE2BIrr1fkgvyy72WtqVTQh0WVxSYuwEFRDwhSpCh
j3sQCswGDUYHNX/+mwJKtl4ORqVVZmvLIpXSsWo7uMzgmW5p+Gk8h+zzO06UDneb1/Ut8iaZL0da
MYBG2Wk/nx+Tx25gZyd/K5cpEqbSb6K6nACcSHaKlt3j4+DWfcDkW7CNCWIs9jTtnV/+MTd8pd/H
LwKKN/P+hgmPm86dpzKDYiTsbHnwdAKlY5ehfTum3PeKXYg9FBcyTLQdkGxCdde4ptoGPGywiK8Y
4K3l0XNefs3sMB0gHqOvvXVR9htbEisoTkjp8exBvrW/sGnzYoB+9DhhKcwM7tax5N5X4dOvFd3K
xiaz+a8/jmWKaP1BIF6zcufQr43sjygVesc0/IAqEMWdpTUCFsKWAgBsI+nWHcAiQ7Z1F3tezN1g
lg5kgkDFHCzK/BuilHr+zBIEcTsFUDtRy1AlTPfXBPscT742b+f9GREFos27t8yy5KH7mov3zP8T
jUu+e9/LRsKRUyGpWWclCU5Ae3GHaxFa/QrndoJW12/uLnP1J3O2lVmZ+T5gJ8s9nKlhy0d+Ha1f
wliEmebHRyiMCvPd6P2Q81aTZ9o6kNnXzRbIXaSlA7cjb1JTA2m1ltvDaUHk2luQlAYWcDVMtcNs
E0fJ/fgYh2mVPhlYAzakGdW3CRlLvBS+sV2BYpHiTn5ox+gX6PK6ft9VWfssown/n1hpnpP0su9M
MWr8qS4Cmu36mhW+GAdDKG3CoSfIXvnl4G13FyYlZ2empr2/6WGiSkpNBEYS1E69rEr/XSleKd4H
Abqi11DOlhDIaq7NMaeEghwttKnGq90c7pvgK7h1Rx50SYYXkkwnI1cyaftyZ4WrP29CLq6fAzDa
0rHfT+siSZA2Dy108EWNpsVrkjZV2VzOrmP6umjMm6SHkbbr2W8y9MnUguquS57gldi/YFGEfavF
UL7e8HNO7mUIJXEK+h//rRJ13mDgSvq9SqaaiEGeQ39t//FJWZS3Unb8RfKCc0SZvczyyUcbgnbW
L9KDI19uWbip7TXnb59TAzCtpj/zM9/TOMCn5ELKghx0DUSI/W2j3oCmWXFJOJ9n1Ld2kEAf1AMx
iADLS1+Ct3180zimRx6vwk8jYYbKUfSRqGVu9NkY0i9FdKGAV3jybeSAz3YTSP3LRneXb1PWe461
hi9BXbuXK4olhBF3HSfarEiBLCUnoepiil6Y0seOMJje2ywOH2RHoxMTufffDdY6uNmVLvj84Iws
AXYZrV9KSkB4ag8dFt0k5H2zt79zCjY0NGkopevZprJWSgyjkauO+FMXLXZ7bi54tT1Zh8X8Vp2h
MILbjR05oiPn1f8vCYPU1AAt1x0I9zTRYe/xHtI37NT7VLsIHTtzlbU5eN4iTwIjafSxQHQUI8KV
f6IqykcNIrbxL1qNYqc+hKa7g7Pcc6Kn9gZ1gl30IS3hmzarQnMtkolLkLS0w2S7Aud4YZWe+w7w
Y8XQolA2tzjFa9n6ZkixXa/XOC/jrvYN/Gcd0MDaSczJpoOCcD32RG1x0iYgRoj3LsbjO5PEzII+
zOD0nZLAcMi8+s/HH6NFRdsQWdMecQD/aPCR+N0lfg3lrobwG3uwogYT1XGHzO4NvqWcPigOz+UL
Rn0cO/4KMf0ZXrpK0Lvq9jVnmiciwqH4BNYlR4IZAvfFgb8Bxnf3X1+BEzg+9ZYYKaBQsrzyr/4d
yYNIlrFAgsxeGhBTwHSIA0x+G9ElnFQ3wghgguzyDW1ye8T6dujKr2924jT+UMkGwnsjsTdo/91h
nJvUdf0z5qU0KVI0QnTQc2gL+DOxBFIOdfv8kugr/pQ6GqFWxG7I/qLhsQ1dBwZpjMBF/Nu2sLVb
GdlCJ2X/lafsiOjwsHYwL9ndulrUyVTTGV45+R22DlGAtMhRrChN3fwrN+0iq32lvk/N/ySNj76/
XBgYmGb60ipyCaWym2pWOM5+RfaVhNjVkDRriPiwAW0x4maKjjfB1uRL/cJGJcjpFXhSGocBZXE2
qZLoLOwSIMy+cqyXVq9NVyEsSNZTWjKkbA1Ptf1Cl7mXQ2t+qpJ1Mgks45Vo86Wx7XIqAFhr1EGJ
h46WXyvHMI6e8HVYrWmWeQFYiCeRRF3UVVSHrunuF+9I2MFLD1XCEJ4lZJ9bL1tF+72mJTa5ug2U
c59yLPM8a86+hT8a+Cses44ilQooF4WoiNJUnrMZJ/e+xjENmucxS1UjYCR7EGTIznJOdDiP6x+d
6hQZU6dPRk8PmInqAqdkusNzkEWeBfvVO0X63eACNXDywAH7rxA6Bro5MSDd1X/pwNsPem1V9FSK
8X0OQ7Mc4+LH9VGNn+Zy1YOkQ1RvFiXE+GhhGFpnW0GCNHxU5tKRrhb9184CBFXUZL1Fvco6wfdt
Rvfi19+sEnWZQgdJcX4+ItS423WXX98Epc7G41rBkD3yH9LXDh0DooLZ0p6l0YOSGsWuGpsgeyjS
VUriIYZg8e551zpwjzErzZIWWU8pmnz7TrzwHMyMDjSggBTwquBNs+ec1Hrk0U5gs8n7hdZk3TZr
wJ1cZeK8WusrmnwOxq1RFGdwdxcAJib+bNeG8xu2vtn07tHYRKxn6nWc88HRJgMqUS3o6xT03msi
l5oAJ2DzL2OVDPnAD9kjLEInoaBqKhbipirslTYt6DUqUsfUUuBWZDPjeeD5mnqvP/Hti/LMyJh5
P0029jZWCNx6uQhksBxLvsGjv/R2HK9sCvRJFzmAK96MsTvnEwm1RdyaZlgpiuplT+WvsXlbuxFo
tPUGtM7aJNzIxvH2F/O4xxnHbXE8FU8DKiFe7SWIhHwHYOaYQH2pyfroxuWl0stX19Z73kfTvFbH
lcM4lgy12X0PjXsIYhNpJzVIatB7zxxbHqurhwEr/SE6JujmSL9ZmLOSypsFHIVcmXx+eJ2zz7HA
FDgXyMNwbUXn/pfUggjdJVIrFfFZz4srI6EHx2soL6dsUsQXWS2emsTE8x/BhaHJSjVjSeW+dVTU
RZzMGJsfkvMkxR/Hdvpu0HjQFl/XK2KvCNYagNdOqKFFOalUCHjc5wDAlBOq0bwKSs4odeTci7Mv
kL0Qlw+TaDGBEabbgx+EmnqE6MwknviWcTd4ev20lPbxVbnseBS4WwJz7yu++Nj482ElxnZcZ8mt
rq8uCnd2DH/QQVPN1HyabIsTL2fIjIVCQ0Pz+NiwTJQHPtoWFJYCp1h8tyoH6kuqURV23urWY65n
Vc64JEawtAR4xPqGn747taUfK8kyi6aj4L6G3yfgOXwrnHMUpgoY85leqkZRfJczb38Za4u276Ik
+JDii0n/bOPOyfFQFkMZLOg5GERAY1kLzkrRFIn1rtJMOTp67Ygz1LjlKXA0xPv2V3O5yXXC4NkR
Hrga1no74FypqjeD2OIqM1LiEzw7jzDxtPTxl920sXhPvBd6Ebj+4A9EKQkwkDIAy0dJcilYRdmZ
LEUG4BRXAQS+FcWDa7KbFfifWsNQ7RjlBnF8InBalknJ2udXW2UPJ56900uuNIaayeKCZDcAAYMb
7WxH7P70+VVemZD3IPv8tlMOEUeelbE3ACel0efh1R87droHRYWxGjfobNiIBkdkgeluPDnMmw2d
Ydy6jkmXaK9VX8QQiDYX+v9rPRl3vmSzxkKmwoEpRbj6oxzE6IUJM8JpjMKzim0LOxSIGkeTqoip
xV2IJp3oKxYgNYgNMD0yeBXrZPSVBQAtL+lWnQvOtK0ZiXVqUfjMR6gikqvYnMnUTI8GHtxXS4Ec
YxpSqg9z2guB2wXIlL6Fe08QTy1aZYPGdceNVN9aKO+Nqp9AKYx7RM/Fdd0gKiHBl8ZZGvkrbWrG
Jp/1qfYpDmQoVr4VPLMbrW60xbVke40EYtZV04GWmFaFJFUQ8vpoNaZE5Wv3mSAhkcqNExCFNsma
27OnNLN0OQ/afGBiGL2XqJ06etfJsOpAWHt7wQZ5ZLk0/SKouf7Gnqu7Pfb38G90PYqiBv/+M3ni
c2CJ5brem1aqTls520RAHWf01FOAtER8XjkoP21+KmUqTr4obbQR9cyw4B9sJE7n8ukz8BrYbUcw
6qZlrAAcFz5si08e3jBhqAVv9rXJuLSbWCbI72FKeVjlJfJWK2T2Fr+JjTXzwPCsUpCUZO1r9BeI
3kwJG1NnOWpeTSNL6p4z5P+yeLSe/gmSjztD0cJfPv7j2bFw5NfICsXXUhbq2RyjSsz4hZTcdcEj
GbqtvkvFg9ZgUfEp+UQNK5X9g3cYHRIgXgZ6eML0cXK37kJOWwJqINYyEHLyn0wMqWLWEuh9hPsj
jlWcBdtIOd7dHjM6WIPytVdyHVfqgvLtnH4K/36yI4PwDFJE51fbhJVdK+meSWszp73IVeVibGJQ
sDnEWhD+BFPieKe7qGUX4ZrpgL7ZpDArgLQlF27xGwpca4EwDM9A7O+t/AWUKYA5nuI2spH8ssNg
VZU897omkidlZj7bpd9XmxuFga8k22UHqb7zaQrbpG7BpHUGgJwrSjZru68lfF739XK5ecwL+LTa
MXZW24QdO6g+uDxZCa4DNj5CCIgjUV7ijRywez+ysI4V3EKci+5fT2aLcuEDvd/u1Px9h6h48yRh
t/NlF+aCeBNXDskVtPJ5b2MH+F/iWAnDbb96xnJtroaqVFe+mfApBKKfMZ3Om0zzOd8dfjErVVeg
kglsz9UxpnjfMxMHdckoYW8azi3X1i586ls1yNPs4EgmBt3Qnb/K7Hi+e5arzgWP7DsaAIi5qeMb
QBXWcJuER/+5S0j7p0TOGNxhcUVNUxZfkkRUBszUoEaXOxK5mZPZj6KrUH54eO7KtLoDHWhRuu2x
vq4l3uxwKdO1AqJ/qiQJIQVeqmCO+mGq93dYDMpMPm+R2y2jRhc9DqlpN9AVq4RKb0pForD6K7Ua
A+m1TvEWGANFx44XoDqR5QbJ/e/lcbpumzF9hoPCvU9bQGssrRF6BaduTcVJHD92snkk9TvBJ2gw
dIkzgus1g1+KtXj3jKGXbOy7SlXqUsbvL8+hNyHSJJi0sdMAPebtaT1SAFzqDML8fevg0BMuCsqG
tO8EFUcTkLmlv6eGYNtORLtrUH9kxstHxInfuoLiWFJw+W+g4H94Gj742nenptk40ivWitIEHIiB
cw8klZDs5u6F62rc17ZF3lKCnq/zm1j2+kKoPYN42zQq8CauJrzzJBMnqe4dsLc0aQS+eAZcpnOD
EuWr1Kxs7sEI3MlF9tvROQMGu+Vi/J+auCgjFtQf/YODl0S8T8OczOnROv20biyV8ym7vsn1yeg5
dryHou1KljRFnYfX8JeQxoQ0/13FTNGHIWFR6OPiIXJ/W9dDALj4LVZjdopOAhXl6t4l7iMPtfZZ
r1kZWxBIlwAC6fxxHKeZqO76d+ilR8EZYtLnmTe3pWBkbT1oqJnMlHb7nDxCzFHvzlKL9PgCZb8S
M6ifU3/d4LbuOcH+h0seTueyQiHq7kBR0JFf4QN0xXRv6g/MS2V3LRKGXLC4AXidd+oW4MHY2WZp
YMN1SBmN92RErK6Hx4kkubZYQ38HYMg6KCjapnoW5z1uvN8bE4IE8uolhEOhvkSyK7VN0bJGFDEE
IOnQUJ0YNvS0iUSPJWQzXKO+45wDFGgMz+k2kCj50AJ+i7msH9puGHpS3OXz4cvSLDQjgpf79yi8
JCEs7LICWfG6QohD4uiZdRPEr9oCpSqL92io97K5v/pQMFV6XQT0ivJNdr5g6Zhj2aFKe72Q3oAS
Pi/gvLV2fRK1gUXN5RwQ5ex2q0DJeDhTziPe1a4plt+bGdfdl67RrdXL9D0UocTuQdC8+V4NoGdk
jHz7wuC/9rmSLddhtkoxXoamfKyCgcvhj975zFWqDgGF6nga/YTjiMy0ZoU7KXYhdayxXfxeM6q6
Wl7w1FPlKNLhIVscwk+4MgrOcZXxA4Jny0Jma45JxaCwo/9CURZNCWfdBa0a/35OeHptR8gw3+Oq
WgRsFRBdftkQm0oyYFfcM2LcTbQAY6kYnV7W63O/3gES+oQkaluhpwr2pCvizSdVHA5eOyF/khz6
nU6/u6Gm2UCmax9G81hTVdr56yhO82lAkcTwjS9Uy6/OjIdGtif8N2J2e1hLWva+CdaGkt2Fl5IW
7QYs0MbfU8TNN9SWF0WS+NRj/7bWwTQ1h7CLoMgje1eRxN/z8UZt5Z+iPOGBvA/OVxrgUuY7v7PR
XqNm+yMzud0DT8gs+TeMg7H26UIVoPVghspOclS5dmspKSHl1M9hT2Pm13iJScAXUr7qZBpj1zFO
fWkDns5xUI7473m1Bp+s4n65eWHUrMsDxV5MTAys1Qb6YsZrOjDVLYZh4Anf4jRDFA9BEZej7lEB
pp4I0cOWlAhmR4FiyChOJKWJOFB/NADMe5E5BOzCNiimBP88UMjEdw7QYAVnAFWMcilw7+m0DfN8
FbAluY5JvzPEVsGv/UpizxFMBUXpAgAB1JsEUEdVvxN9YxRmaYL3D3Q5IkYjy/VVBeFcXem8haFR
V3EuyVqI048gjB8UyfpFOyVZkir0j/0mFda+/KjQGOoD7cuDp9pfcT9ALmXYbo9r5Ur0rOMB05cN
lkXOE0Rutoa3Dq1NC70AlEpdh7cMCvJRZ66u9A7NjTH/XbLI3ecHeA9PhgGp0ytyP4xuUuIpH+fx
4JJ6IsgJJbq45P2VroCgjcSqAiKvDOiPKUTJayCW4bzZad8cER96nfV43ZSeQsmePd4I0ssDlOLv
XlWDmK1TdirQ/n0eNaY7TNJ/XK439Y1F+PfYR22vVx0YUbKE9d79BsWWFID5KPNChBhxFkH3Ps4r
cPAuFrTV2N0ORe+jTMb/PFS2mZ6dMc3AskssNdACs1vRYKnOrZ4Sl11P7wZMgCXR9e9993wHle7h
WUn3nF57MLl/3vrEdTIylGShj9ZWKMYfuYR/sIi0y/3X+i8zzX9+E9Ov85CnZUm1CLCKPx8yEHZX
P407yjt/QOzCpzGet0pSRvZYWjUQwbcxxHxCi4AX04RpB4d8I8qf1xJZ7QdNNZkSLF8aP139XK9W
1LHSa5vFNmvh+H5D9bMSSE24ejZEc2YHkJyJjI6sN4fI3KKIresALcGT+9j5RPH9Ig4kybnxedEL
7H5BW0ZpzCLxSczivdbtUasdkGZVXNsc58njMaawVPDV1k1j1iWarC7IHsNtIWkejGSu7s7fFM/A
/pfQB2qewgBtLRI90jKcaY99W7uM8taf14z+OndaloV7g2ptyaN7pI/A9JqStVUL8YqWsQ/3oeQ8
0mhLnYkY3F/6xfzHN6JCm3JkJBK6VA9nVy1hIA3opOp3qlzOT8tFa5u6rP5kqfXpa5josORdiPYG
vbvkDTcIFmGUIX6jCflKDasUSl5XcFvOii2SFbFOTMUVaRV6CsxL0dzGYr2829LCSmxNF1qGdjCQ
8fQJLRFso5AoIdUhcIaWvFUEHwbyBxiAuFG4dHneM8utw95vSUN7u4StlYf7T4l1wft9P6NWFs9b
vYjT8DPgHRPJg0rfCt6SzmB2jAm4LXE7m1eE1B8iVHobLX6GJTLV6wSGiytswN9djZMjd/sV1Y8z
rGYORrc2FvPZiLyrnJpOg9CrQ/c9MWlyOn7sTP8C1Uj8x3L9U8W2b1xKzG+J5S/gMou95T+p+N9D
3J+CmSeqxMV6sytTi70zLuvwggxx2/CpqlBty1WP6UBLoB8RSewuJtYkEqTSt6l9O6cyfL21FbHg
/jmFYrqce2IBXjqMx9yZWzLBlFzF2Nh2spvzF/5Zs3Q8KUA66b9K7F7Xge4+/zwwIwJ+AzJvUrkT
MLNMtTZ7vXosbH4Xm54GBvXRl5gnSH+/K5qtCdQTfwfRpcH7DqSx8ggTUrQru/xTipr/XMjWeSVI
Ro2pxY+QgSAy35po2v28om+u9vXpF7xe0zS73u/a8rg9yGjAveRGlUF2fxb1xAzf9feCj/diSnod
Y2Y69co3lXFUI5OHIyAJC9/2d91EZgBH1rZKBi1Z7858Tt7epiRZO6ZjTh21MByd7jDQiblWObb3
yADImFeWkhZglDrZTn2c7+qLkIlkm9myQ6ito5iOXhCe+KEiZrCxM8eE8+yLkUJQjOg8P+NsTTm0
+9Y4WqxeT0MsCxls9NUZXareUPBaXca3sNOuK51vcLaFJklKUWmZ5+vulUf23apNoRaZUkpI/moD
b08A9lf3o53Q7fJWNMvAVLzCkplD5SWJGmSLTtIY6Fbmo4BmIvDM9WapP8kzii50Y7bOjGEXk24l
qI0sGTlaCUzLep5E64HFtJcZjfMAz4s2T5ZxNhKcr0lm+b/BlTT7ICSq0zy4TSYLFyP2zof+QzzJ
ZR+9gW+kY22EZMLB+kXP3YxrAQNfmHwVWThFcU0zqf0zsHPHeW5tQLZfgiEzN0saIT2U6RAe1W/9
t6ZAxUwBG9a93AVVAQk1f9tO6W95xRYs67eH5l5Y03oaBR9MlSSRZox16phSYsrh5l0OGBPiQuI/
iI/R3Qt+r33Zmhn/HYxTQkz3vsHEZdadSjoinsXnGCami59J4ie5LepFd0NUAFXOkEiNoeN3GrSK
0jO5G+UoXSxskmSHXZX4xNR4HbImuYxWrfUzuG0VQGE8cGsUlV7WnrvwQiLwJ8Xu49DZdgnpSoiW
4YrrOPB2YG9EaG5k0PX2MiI839KF2OxInxWf/DLagqE05zYHBoi6upMSQkNrCp/fAhPspuPaxDdO
kMW35ynVENDV8SpGSpbTeRJ2VZG4Hltdf20NnyQ3t2UsQiv4fyxOhx9+7/VMb7Tzh2sHRD4XR0mJ
PO3xpFA4QVCvfzVIDOGvQbsDGvxnlRCgZs8Cebq5OI69jir22ej2Er14PVSrFzAtamFIGT+EYHoY
9OsF7n1nukRJesqdI1OhFqbw4seCChn7Pfqs0mzYO5AUDqBx5X6WoKO+rC0+4wOn98vrAKe5YeZQ
Fy4Bgb7AatIexMcWF7/FpwC6VEaYCR7mAJauCZ9CgLY1Y84qcGrpW22f3mMx2cat09iaeq/DC7Fm
L1Eh8NWOB4QfKHDGfp6tN/xQxUoaei4qiL3ssIMjg6+ufI8Q/8wfLDUpv22bG+zgj3rRD1j3Ne8X
yD35WEQfuRFxnmiIj8UuHpX5a16CSzd0ORaCZPIAnVzLhI0uftduH36/msIKhzQN5qRsiydx4t0B
W4d8B4FRqMqyeDhOZ7JLwz/4R5FBuXWwAAeKRl614dS0iAjt90TYXHtySgp6iOW/NQa/MFEdNggP
aw1UoIZQ8yTRGFjj+xTe1F8A8I39yd4WelnqjjmuBwWfmc7e+80Yi49Bsx7e6eBVc24aBTkqYLdK
LaNaeuGkNYzuRjVBS/YxTl0uyoj71z1eA+MfWN4vY7pUgK2i1ZPUucEYbcbAdi0fBz90YsKIMWnd
n0FScSFbywWEyKDmE/XxAwBFyxAP5IribQN+0PWRCeGl71mHQ8N7S7VKiDBbe5IwgzKlg3kieQjP
yYFsjWrzpfRnMM9LC4O+ZXSuMDbvEsAnTv0nhRHTyvaAorIN7wNRbI0Y+CKVB9ID7MylcskZzANm
5CPkAzcjE1XwqmpnjNvS6lK+aw3I4Tdr8a+qVGbmw3p2mUI/k+u32FYA3wfAHqj68c84W1ktR8VN
FfJMpb1Pyx7LYtXk6dWjr5077RzZF+ZWzQJTzHklZU/pnn9fZBxdsXrNhIigH1RtF/ejzUHTzm6x
IrV0RoCelM3uOJrLvrkLuJ5hAk3FYjODnOaqGyaZqS5zrvjMY2gBCYkyFr+U7QEXeiBO+NWZCdjw
NwCfzxCcoDBtpadhuwnYReANj0aqsdYPCGoZPd4yBVACV2TBl/sVEm6vu2vFI8AwIBFHtxzn3h5i
C9oi0Ewale1scApAXQhaPnHOIloBB1MVbA1LO3pL2f2bTC/E/4eL/S1tJ0ExzX1e+0zK4Ih38gcX
NSOWDMpJUsfCRYxJR8BvA6rxTeopL2RoXlpu2JQ5N7ldjtwSC6u4v1a+gDBBbct3VtcfpmZovksZ
T6hcuSL4GxSXjlBSJAB+sN59rna85MuHIM6PBI2rFc0xQNPf0Fj8p8+va7vstDLng8aiGypiPPK/
NsywdNT3DKlVzQcNXewnNRWkcLLpIFGviHZEgo+YZy4/S/d0RlbKmqVoopUnAEE9pYMeCktN4JAy
Gk6rWOEFeamriYx5loBBKSu3qIAhwc0tcLNM+4hTARdAOUmS2GJuxlFcwNFEB0EPIGTIINkabP/P
MsD8Yp0yMleR5tdX1I+z3UXTBFm9JLMHHoa4OQeOo1oQJ+17WIiMUGivatvWhmca0aeQ7v0+kdZU
JRVhl5QEg1sf9c/lHKqigrhFAyFV/d0DtA6XGkwavKZCK1dRKKKvKf73kcQ2byYS+otwjsmvoeVV
I9/h4Ig6MbZUj27RpV3+ljBkPMhgiP99JLbe7sNq89VQC9vcwAefpwAmRXtGthNhRcTyZIXXODBI
Bd26phmcfdpQTd28fPaUwRcWnhYlIFdmUHj/P0xgmafpFcNDrW2gvZaz/RvDsT4xjSmUnARtGDEz
xp8pStCdygo7baW13bizJny7bjXyvFM+cxFmUBq5VhIxoKM2MYHpKG5im8sHyIHNMLyv8cQgpzek
UFm9Y+gtLsj2uZbpfJtwZFMuaEnymOtKFN+4KgE/DKMrLkOv0zeA/fYyNghjOOynwG1GkVjSc6t7
CRzTzMNJvKY5lV0ual6rDhpqArq7C2n+wfW7mXq2gURPHgezysNvlbd2ZWp+FGaXWkxCZ9LZFs/S
JgxRFkh6bk+DS/SyT1+Rv1OKGoEQmQ29gjyfBnu7H59sNTkmlz3X344P1NlAz9bWN2V28lWRf/yI
yermSI/gwqNjHa2iWRmiTqxOY4nAQVGIJwOxY8mR0Ubl17T39G8zzOxHIOrpGsEkCknus3UN+H9b
1yiXZbHrrFcjruq8cqOW0Xr7XuERORuokBgR5pe5PVBJOFQ+UTsjic4n/2cn+0WHg5Z0M36B8U2x
Gprzjqh8IzF95UdBorXMUdFLC/Q4xnTE/e1GcP4OBWA5R+0OTkX1HS/Lgk1GXE40KFrRYniNgkJb
e3FLh+2FKl0aT8lnRAt4AJa934l1F/bbGvyxh9rU7FstvG1c5PSRAydND8DcX5rLKlSmzdJbE+7j
8XqKeWpUEe0ssjX1cBMg+c9WkSm88Nsi5TPTyZLXe8mflD5D2FYt9/SUu7sl2FgJKWD6KKnE0yVb
DdrXu4TIBSVpsNcEB4DF1RBvBz3AcSUgmGMfW9T8QDCGcJhaGLaElWGX4wqBoQU7nGr/jehvlU1I
gunu7KLmVzcgBvps2miY74897PH88R1HBgS49M68+ELBI+pEWz4HD8MWp9m4SvPB8rIXVhxZKzXD
CV2j/thGM8S+gbxyBN+SGQ6uhIXyqPvDVr8VG/cIQqFy3bNreWRwYhfsRVxgLFnHtMyRTgLynjVK
57CUtZ/h/80mxwnZ4jKNAVwdQZWrgUXKCvfQXNODCETj6m+LwYe5+os25bqZEbbfiKL0u90ed4ya
gvUa2cYcPa4Yf13zmRVOkwHX+orTp31UCVNtxktmW9MZ1uoVuLGSsWAhyGW1mqpBgttQeeWp8ZnJ
9MxxLG5F9lLkW9Uh4frvLwPF8+65E7P2NjbQ5EC1PbaujJ2djygMsd4iI8CKUAZ/pvTshnGZfJCT
61HP/NSaMqmcAW64Itu3ONpTfXCov16nY/egQSfq2Yws7zQlPN2+8HO2NRw+L8L3A+vTNU3Q2EVc
3gz4IescEElSaCTiqEg8e6qPjjjc3AOaZChQ+Olbqh3gQPnNjzRFUzTxQCXzMKXuwtfWFQx9Cp46
6M+UnvI0I95gjl5p3iAjU+o98MZLI3rMTjlT4AZ66pwAsWihYDOWMKmBYg1DAeypVf0r2BC7sNV2
wjwjJqqcGSgqFnkpUfUV6oQXm9F9I14KWbSyhORbnY4D7octoLE3sJqiOU+2WvYMnwOVdE0PwC9f
f5BFP/bBIAya8JB9sI0dv+T1JPtCNDZdKickRIKA4FIh8O25XlNGlpRLEKJsP09aKMgZaAplsmL0
GibobSml8/obabgXKAA6M6SfANFPS6c3GT6fLcSqVQwP4/sesOQbf0mrmOAK2l0BfFXyFSDdUKtL
aL/59ShsnwL6pX6e2lzz/gRZrq9NWRgvgEnl6GmfTnSUHPVrM4v4Ocvgc5A1C/YMgF5rdDslKbix
LdTcQORQjcAm9tTJrS3r0WFT641VuL3piKHM0QjOxAA0Ku6GsyMQWnu5JC40DKngM5KpqwIbHnGw
GIY5y3UTyRlIltpJjTg+EFRV2n8p0xcHpTsyvBe2Hmt32TEJymuseog7ohbdajaKDP59uiWMb8/x
RBdmdm548Qgj5E3IrQMY5QisW40EMNP1lXj6HNsreSLndJhTg4sIN8U8ImKzk9sF4395HVwoPz5Q
A0eVZaXQuWQ+wLQQgYsFpDCc5d/KH0RxY/DCkzi/eXnhgry5qbzwQI4doKi3oxBhg+ACBIEjjGK3
0SM7XJyjhwu+Y6RKPxZPjNfnZKkX7QhwGUTKu7llXUePBw8YK2vIK9r6QXBjoZ4brXtuHiNXvopt
i8/wlvHPkg8YQbt4SBzyojDsF1RUOKVhmQqbdX4ngzhpFVh7G1Wkh/WcD6+OxAStnW2GUSG3XP6g
sNeobd8LDdulGjrt+y8r+LVT5/9s6F76lyd1AZSUBY8Gsp0jdl3r0KIFTprKvex6zdN0u3KBtrkg
bg71HkVkp5ditpXnOdywEBgBNC6g/4YFiMCdpajkuCqaAlVTGANmznUT8eRccwEtNvGX8YoH3tUm
5ujrrPWmxZCGHXSoAyLGr2TqLm34Zruuzf18strUu3k+WP0k+WZbRsPPJTJ3lPsV7I/o97L0HODQ
GEdv1ozk5FfS0bsVmGBInUkbnx2eGsll1zzNTVurH40TccZnjYxp7OsvthQglXubWuGIeJakGggj
9rcLfPzRjegDrag2WNo28bIus1VqVpvKd12SctEqGX1V0VAKiVYxqSUctguZUGaOyNm6jMi6XX1u
wN0MzNWzD1PSdiQ916RbjF5r28PvmXyBpBqwJ1d1QASXQ2Dg6HASbZqZY0zEIcSSouXC4wnWmmd+
kOGSd1jxWe1wJ5oMDKFn+gFYKu+5ouq0IFPsG1VmaXKE5L65pQupraPwIIXErWw/B33ODTsgkdBy
4q6YnsxuWx49DOuhemeCV0JRa+ftjVsT0vFr4y148bp7AqPPdA+hh6mhGEGWnZ5Q3DQM4FqDFQyN
fymWql0RIcBZNVskDNERlDMWdViSMhy/Xy7iwo5bQpCOrhjW051JGc+rwKme4La4aH/Ke4FrqOpc
ucD6yZFMtK63OGnINito7nWIrpr5WpWe8Qss/EDRtIy8AxhNyYg4DXQxAqzvd0YA3RZaH8w8CwVQ
tGjp/xST2ZZwnSOAS8AhMdQRfKsO1EO8CgCUPQzGZgzTad2B5gIIhCz1XlyVg/Ujcs2IsGIrsRFZ
L5oKgeWVamgAKvTLmVnj3GNVEsCtkW8mZ5M6Qmry2Crocu405S+6rsMJ4uJ5lJpwWd4fTq01AIfM
IvLuzIbTtIXLzBhWdEl+T6ChGGwrX/Y/Q468/ADqp5X+ScExonlsJP01854lKXzpF/v93X7pMdT+
Ud4o2pTYZyJ19J8yDosRbDDmgryFZPR4d4gvxEHhq+u3vfcjvcHeW1M1quRTXdfh+YOEOCANkAfs
r8irgELTKEzzr7HyoSc7ldSbHBuxYbDSkBiB2zj6jPLOpIAqNlfk9DyiZnO5+MjcwsMXNMUweUcn
SHre4xnaqVFlPf/+0mlqzrMlWLb1obW+V1sb3hSsmo+ubDeYXj8wMz6aCaAMVSSIsNRfK8u2D6bO
NeY53WtlEmIJOh8iJTzvcJudGSTPG7hAlPCpLJN2ee6ifbsOnml+ZWge/noESLvJ9t8t4AM5zhiC
+YbVCgL7XQiWVolCa4LIKLQz+om/J3gdDdvWvMou7VapWmdjdQxKeYyxrFsfwFhgO/AVb1maJZ1B
yWoysiGhCd9uHp4vTTHgnmTmbiD012slPjRUkOk3OaW5CzxFYetsqDQnCly8z1/ovAOxnyGBcVWO
PW+kkxdxifjgL1uYuOd5hh5zWIQWyvolm1Fnq3WFSxNWuBuPZxOSWx5JnNR3JZ9nEc13198KcA+w
WHV2/xUDAZ+h1POn2QJH3lw8rL27mcmTJGCyLxuf3unJCOfq2hCajmH/ibQa5AKBXIjtiVPxw6Xb
0/djIjvKT/jw8Qfn40hLuNKac1/4/ElLtlys+uV+AVM1fygxRxe/3WQN3LvQYzqEDhfuno0Zb6pt
wpCFLHYt/0FNcs6He/CqIZBiBTu5Wa8acuLSILKZcN6zSneF4quuCFJiE926b5ywOZBRvDmT0vil
znJJSz37G2TqzZDXm+X+ZTBQ2yjNLbd9TjphURierzx24v9bktE3VtZywhHmwN+qMWiLRnfwvJaT
We/MWuM4SI7vb6s2jN4caWboxtfFTlPQC4NORHyCLuaS7nQPjjRtlkiYZo7VGyzlK/4HCaN2Vc6F
dOtUT2cscbdDrn0ONO5QWQ6CwrfMYQ8Y+YMfiXgEaZLiuOYN7Bvsq37Ip6oN7k/U0SpPTgfzXeK1
W06XF3OWqkdNj1DtQo7WVYB5Zw/Q+NfKlTVQGGzL8Kf+04J60iNsojQdSB3RnV15yYZobjCZWGtq
4Fvm6PXIyc0osbFCgQJxLmf5r2dJJaNyS9S1agWU6bi4WetnpmoduhYoKK0s5l4wEBVI71XaVWQO
LV6wOlw9PNQEWB26os0M0sWPY/453N9fLnlk92ley/CJXs6olFNhQBIMdCopF3kxAwZTEXxdZvhJ
oPaNW8EOn6lkgWZe0Nrax6npJIrwnR+DIve4QRvsinyxeXh9n0UcxRujLNbbwRvngubWkEObE0vh
kEjz/Dd/iDA2h1nYPNs/kpZ0V2rCdKko0VcBazH6KU4In0kDssW4nbC/6Bzfs5DRbpzMW8iwPDew
kpb0CNj0PRpe9sUiIokR5eb27hIAP97ZTtnDjxmOz80WmYwnhwgxGcosMnbsH4RJoJh3RHpDyYOD
FjzlQDUZHUPixQQQsTVrwdV12yEbZ4rtasEAliRiJUuzwfXn/IZrwOtymN1YNbQVtT7FK2D58Mg5
Zb/izajiHzK4687Up2S7EYkYUaJASloGfs1Kov+30ga26305fgBcesDBtkn0w3ewkSHyLcWDLUz2
/ko+ceQJtJ601MmYmY+vi7o6r1YbxurSNK6E68+b4ab5uiWp6bEQlbnAusjGunHUy2cieCUrLg/h
WjhE9un4/6KcjVZ9DF3rqQRg4HP7l17OJ4ZiQJxcSv+HLsqpQX6qeWqlIWo9ntj8ZJ0TKiwJS2OB
Tk7f1OnZFQDqNqz8M1GNAa36U7X2jfydsdq38uCNht347xMFJdrO1raFD/oG1somytXM/9I6EI1c
4bIql7R3c2ILfTmcVb4Z3vlyTlon/fvxj4PLofyAhACcNaY1KNUBr78v2II+OUg5/nr1Ry+JJlCj
M55Qt9SPySi8dWmM3Wf3pK2jhoyFFVjyFgzYJ88w2qyOZQ62Ty6wN5BokkiHslB80DTnBX6isazs
65l3+jRUCIP4eJOMtasM8bjvP4IY//tEtGgi+plMxZjKxq8gpTFpT17uNYzSsKK7NAEtIwuChYCm
fmoLQRTjeLimEqnCC1afMH3WsvyIjivwMDTAffWsmXNSZMk33JytDznAN/brJAtSzZfCjQKKOmuC
VFkvDtQAF03eQiamrPfI4ibVamjzppVMo8mIEtPZPfgDzktD87CY3D52PwXKmK5Q/MMtrP3MSmzz
gAt9Im4w8JcZ/ABoZTv/y8CY3tcPu5v/BCsY7LuHQtNvbUt5Qq03irlfgoGd/Qj1cn+e0fNtuD5q
L6AdQW16W+q4WAP2e1lylxUYWoPsdcG7EwDFN/za5fAKxKJrhZEr/Jraeo/qNb2YJaNQjOHDk+Sa
QxQxB9DhJGIyVtBF+oqTziaDwXz5aI+SapmnOcCb5tP+1GZaBndqmG4LoX6UIhsVOKi+ZclG1W8P
tG+MGqY5fZZppEgPoI1/Me/h4QYUKEcdNvmyqO+lMF8PplK5gTbb6a/10hMXby7EnICVtjiKsVFq
l7w0N1KtW3tjFO/gngAbZXXXnEFHAWZ94dWmEEoMB+uPcNGXY8tKe9hSWGtU8fP1j0oualO5gFrN
2MwXU8zQNfaNG0DB0bZ7Tmwb5gbbnq7lXCSWZPbPrjXPjdRe4AMHXyyibSU+hnBjeoAy3HIPGZEc
1QrWxknYkkkCsH2QBFvW6s9VEAD+YVPsSef2xmRBeDMWpqWclxSMvqMMo4XNhzCWLEY0YQ9otpEz
lG/3bHoVnmBrLmh01y7eVTsolko92G+HkaCOlJZDmwqB3JgH2bUrXLeAJunMVVh85u7gR40uP3X2
1ISXa7O/NTg4CKEdgStMFYb1eUya4YysIJN6JGwpNH9l9DWJe7khvBZW1RAXL9kA1RiPxnTmVS+8
haOzZEmcSbBN4VLQVPMOEjshCtI5uy2gRJjTwXVECYhG8266g3Pa9rcvW6BF+5yIoMWOvV60bOK6
wU5jGHcvH4f8FtI84+Ofe3gQrhSX4RYOAtXOq9ycV31SWh1EQdgB3T0nbs44YTQuILICPrenxoxW
tZ/K0kFloHSfAuO1EdvIRwh8b3j+SZsKE0O7wZZ9RkceL/ezo7L2//uYt5RqlfOIqefXXMNQteGQ
m9uYYz9IuiwhsmlLvnwaAX2UN2YUGtc9v8Dqb29frnmIRBwKc1pAW2HbgXBzRMqqNxe64Pjn3B7e
l7NfDgtYKA2L2QyGd46gpt+NggF7RqDeJjjqCVlreQS97GuXuSfRbNlvG/y41D58M6VRTf//n9zW
YmnPr++yr+k3sahVOHJ7/CrlXFvmql4v3c501WK1UoqTZ0w428GI0zvyrAYIUYa2LhM3xsOFlprI
SPJ116VGdbJ1rtXOOXHHJVQvYJGvXOqTVhcTeClrM7/aivDGubarY5WW9k7EE3U5+oJXIxMoH2Gt
CY034SeVp2MO3uEOfi9XRyp9kjbZh/i4y4MaK6q5vcw+xMc2IHh/PjEkT1Nv6i370auKETghCJYP
/rbaDV0sFsJr9/f1UKHsQ/r5IpXP5CvaWomHcBc8NmP559yShzIN6uEFJxm/ujRJ3U/6yTXUeUfg
4zdRro+JIORMIVmifQ1gZyvQgTnNynd43Zgk309suEVgm2SDYnuskr5fXL8UlJ60gX5K+PXGlxGI
7DC8WyWXlt1rH9Btd2q8A4ZOw41AAKX80HaHZG+QpU4+dPtBXl43W3j9JdDBQkocPUk8yM7u34Sf
Ovt9z6UjbC2Rlvn/lsZRYp+krSewaf1oVx3G6rpnMriXuJXYNRHWV/+MeFtpR85DZHUWfJAmqRKZ
0wxFNm6gBWXXAI4Lv7mrgSVZbxM6KMDEX1bO+Oe5pS45ReQGsPjTVa8UdVFyKc4hER0TTZTayv7k
GOyYSfikhqJwpuvb7qoUM0DvMNlJNlfZhlvoVgHdNp4Ev4m0eyGE5uLueO+QaSED7cBHH3I6G26c
MYoflT2V6QBL6IHDA20TPPC9j+rNWCaXiYkMSqUh4O0Ose3Ny9ookCsV5wWk7Ny3b5gBo6PfZnbA
zaEgiqaxDF/jcXtjdsH7w3YJaSQ1EjS8fvxs6OUsK/yQhy4NFh+mozc+5rKmA+uYX3qMqI2uvaf5
ub+wWyTdOLPwNci3VKxWorhTmzZ5Fcl04c4ivqwRuMRnKHo3fAOX4GEn/IKjacKbcTFR/lM7Oh3p
YM5VEK87H4hJIgdnDshQcleAVK/w5zSSIYRJ+r+W/PrGkMnM3Nu4eGP/fYt68Wvc6VZ2xBb/9pGg
gHhrgbbPZj2RroouCU8odyehOi56YPUN0MWm/U77NeP1lsbhaVw/3hdZV+S3ga9kxEM1YHQbJxuE
YpCipKrNehbM19aKwAqVBgtCvNEfqkCZkJV6lTJtyPn9qF49oeHKQpKlNyd4fTmI/Ri7UizkAewY
DcVO+w2zlvTYlDrDhNOCHgx4y8U17Ktf8KLyPNQM24/GeQDstisvnAQmex386VDryfxQk/wFnRea
gPExRZs/BN79+7XSpLm5DPki9iiRinhuJUrKw6oKPgTiIFwTCoLq5VEbsNq5LqyW/5lkHBgvMgyp
YboidSCkjsm28lrMloyZH1prWBnLtPTdAZjKzOJ22B7EVero7DhMpMsEEo3hF2dKDfYEmo5RWssz
akq4CpyQfN6RZHfhBjiSzsfP6aPGUEb2iYj4mKVQJtg3ZKmQflAwlV9U0P3enezSY5gvKpW3NoG8
CNHsocWZdsoxjM8tUAEDy7l6rIxFFFKDYfx51ZNLwcgEuqeYfc4gYJOxwqZNkfRiHfGyb10Q2HJW
i7ZMxVjSXwwzZ6qX59bDnVfY5SBllWiKjuD84vqgehBBmu0X7BebXTEZbN1bpQSNFBTtxY3gCxg9
PMHj+hafsgmO5+vIFzG8MK6kmFO8mVUbXr82beCHyhY9yWGv6OdF8qjHH/H2rbpsjWkS/4QQ7RoY
htgl0DSzhI0KrHL91Dgl6JgDQAFdJVymIAsk+PeU4CJIr7mgDShkvKkox1K3oL2effSduHRohVDh
DiCsmfwiHSvLplGcfASxrB66Nscul2O1kY5qp1YcbmjnEMIawNAlZdneKxn3pWdkbAnwzeqbKBKN
qaD2RUUMXmA5sORqXLOHU/UwTagpm0bpAhit6s3zVSKWwkQntUREi8LSWPR8LUGooIGyzuL2Xlpk
+tw0t6SZsevy1PKJTXULYXTEqfvWMNpxOte6fxhDioOKwjCGRM9gwTit89xSEzjzVBmob4TQLqCW
/9nshyXTcZGWLJgmEYAJ7LK+hzU+q34Is6h5BmpbKfoIwQqUS16O+fGQsANPehL0Uk3J8zwR8dmv
wb51+c/jTh89/42Z07ZbwuIpuEj4CDpcRlVJWU6irInmYXqS8k1uqR+gbfm+UHox7tdVqHYw4aOB
f4K73HxZZ03iUZh52EHggXjBdFh4s4czPEWJ+TY2huwbplSI9BsXHRUeV2ypNL+byHl+sknkgapl
GpbN6e6jXQEPAYDYH7DcJ73qMRK3jrqPGze2Pd4DqRdp7YMiOKAvTU8LaouxOq/blWpzPOIPTA3b
rGeqGm4Ei2wTGklPQRerRf4YZGlt5mX3EmpIWb14nIOTz4oG9YxoM6RHfM6h9wDHAyVI5zvhJR93
DipWKDtfYjHC2sWgSSrrXiSTN7sxgpDiZols4mROGOldbDB+7NDHkx//tc3iBecUqYV35ysQh1yL
KrtuRfxqOps+pabPgKyL6vXPJyP4KPiWocnlVI7k/+6suw7S0qEVN7MXLR4ifnCUYO1autZIOtku
OlRpnXQTdJBiVxUlTgJ2rc7k2eflgRfMMjdGr7xB7WS/J9ofpCORU+8WuYkYH0qLkgrOjORdz85m
gEFaIQYlyClUqzqN+SBALcYn6Zgw10hgoL4Gg3gzKQ8CZls4aDoCNmloomQXVKV1BZMl0efqmjPz
FYtfoj76eQWRmrazn/nmSWhF1Kd2CRSe3NklWKyfvouhureFAXVt6PQPYVi0zpzjU4gvOX8NxjSg
h7PCvDFvqtwUv40mFr1vwDEZ7XOnhHYTanyLAXcN4oJVJLfz1ND2emOyy/BSIxY0jLZ0x4I+KJJK
svuiiN0t+KLdCzWJf56xMyjHuJvITa65dNsLHUOasiDkH8EltBxHynuTPULn1L7Xuc4Zh3z0vFPt
Lz4y+HuVVjum58Ln7PgP605SzwkoCgK5OzGhnSIMIwTtEnhZ2OE6T6o0FdQPSjqQKvKlNPZSexMT
FwurIwCWvOYQN1zYmqkkaGRZU/Il99e+gCgbQhn7JfdqYxMCXSP2+f3pb3YxNjToPynUyItmtk5m
NA8MoyjZeoAMcjRxvipOiv3okRNeavcQ0CJJrmmXAZ+72i/dqiYd4BRDWCO3KJTVkCXOblSSYB2c
jvhvKb4ga8OnpP4AhJ3ICRXuAgQ3YzN4zIfGQRYHmuJEur1XTWqGGf2IKMiATqfB3J1+CWb/A+M5
sES6o7u5NVBbdt1q60gc7MkqFgVLtOZjaZM4Eu6lQwQrBysqMejZKoG1gFNEn+LWv56YysWKGfKG
2/f3YDBDlLG3PF4Ig/5VjH3s4sXhwg8HFcy604q3GhQisoztdQINcPs/MWJuz7Gq2nx2XM/ppHeU
zO6xcI0acZjas8zi7alycGgsMtFTCzml+Vz9OpkCKll2xCtmEFqGDzz4B6eah5sasD/b3WBzNMIu
BJ2fCJ3eyFf1b/8byKtzD0jMNPWXy8xWu951jg4MRU5Qr/ptvIhfvhSQDHeoq2ECTgbp8D3XorpV
5r0GLJ0P56WqrTEBsUq7FIUKwqd7+DbAv+6pUcpep4nNfXeJejNqzRrHFdHDj8wpS/acFEsRF8av
30LA6CTtOaJNantmrPflDY5ceU7koniA/PHkEqiPn4XTUqFMVc4+kXwOHb9+TR0RyejcHVKASQ7d
D6X4VHEFSEI9FDc3PWRZSUL+WX4mBIT3OTaeFnaxfW66LpXiSw6vms9B7xJ1yguEM0iMTsB6iVsJ
gJpq0+ueWl2TwQ14XHYGACkfSwzH7FrG8gTZ15ueKnG6IbymrnssqiQJ5zm1X+MPny9jFOhuGm4P
1n44H55Ob7a5SONLWM3agSoXuBgDkEuwWL9wBD0xuCXB7RigXIpRDVsLQHahLux3x7f4yRyz7vtT
yGAZiVtbJ45YB7AAc4Ld6RIU4pONTGr5lbRYBd69PK8r/V3fzCBuTZlNpOqVsgCEpmb6qBl6jlWF
7enCMYI1fMV47PsZVH/C5hpQO+GZRS6cN0LCE8FOUm4qYMULqdBbBVhGdKuV2ADstX95/1YZSqDZ
n3cxj78RmdKYXAUgMOgACL9bgXICCPP7ZWtgqzK50kEWs+h975jPRiblG4getGlzalXVJfbZBEQ0
l94eRYsYaDkj8K+8YPaw+JbHhUnP0065A85moj3jnh5BS8StA7K+GZKc5mzTBEmMpNa7YfUEIa2q
0TYCq2L+OD7WQQO8+aQLkQQf9CXwW0TIrCpVkH/PtoJ5Vn6BhDU0aAmmvOrNz8IEfBgvCqKE7liR
tiqDH3UxOLGafWEqnpzLfw93ny0e6jIcpbG9siFwKn/h0xHzmTYnrrmPUgbbcFLC7E9jHuaPHkZS
s1VIfPAdIel5xPzgpQoA5kR9wOWmty1qELAPr6wR9FbdXKSynyfcJcrVDj0trbd2p3l77R4YUIjp
ww06Epk33AFMHvAfixvS9kDCvaS8KnhAPR3u7wHQUV1oLTMJJLCDye3vtw7/5yhUEaSfshTJEuyJ
7vQWZwq4Vg0VdyjjOCE8ZVZW8LQgDVFs0+pTpGsMkkCaq3BmHvFFJdu3Fu/esyW6PFLQAzlxIFV3
hmTMGYbXForLN/q3pl7s0WUD9eLLGHccejNBEC6ouqDlTxWdAjIz0PUkfFhFfn5P0cwqh+Pi5WL9
cu/36w1QdaFCo44uyjmHOZ8QYTOZF+QI3nYopUTZe7cxXem1DyDL/rDIjTm7lfKLCWiUEp2qJzFj
Kg27DrAqZ/ADiDnAEASqGJ93lGJ9oM/G1VVtqUdrQpDsImBrDOIlmddeHIWh7WtB6bbBj9IOGiMl
7/XQOPKUTRB+cp1seoWp7HtXL4w3hnQLFTQDEmcYfmJYTz/4YrWAJsdrQtYrBLc9Ne7ao4w6eilZ
bkyRYBiXnIXV73DViE8lPax4Y0Xv2LOdW78F8sJ2+NlcTaZgGHWtLPc7Y+lSGgr/veHEkIe/Tx6Y
QtAkTo1Z8p3dwCP6vOqP8FbMjOUY/iiZpB3fBbeRK8FKm3RZlhPFTBlJkN+6A0lY2pQjR4q4iwvL
fRaO0qd4UHAdAo6cqLTKKzjPmuVIfta+DYQ1M75//3KLm/cBQZxuSmM/kMwYkmRRf/9lVJg+BHbp
qyC3Ea+qozX+/czUTwHg2zhfMYavILFeGOCVv9FP0791EkRfYRDwuuVw7oKQpaov0AA84EuQVwb5
d8ZHITKqbStmYQ5UCZlPAxOKCXV7IYE6YTafjRe+PCPaOIU7DUxHYT4CyZ5+/ciwYXRbRskhiFX9
58lxp2kX2H1ilhKivS/l8np7/VhfqVR6EX1Z4FgFunksa+8Vsl+SCf762fMW01EpeFQc71T2+qTX
sOph5f5Izofpq4/iY1j3/Wmx1rGDVNAMBXau3cpjT4GSAkSMND7DbFFenlxaEFKBCmrvBsnAt8fX
7qFe59Uw6d/glkoyn8Gbp204caeDhIhQJcSOUVxYC7ewVbMgoO0OTmKvqClGFWtpcxaUb6r+paZ9
Cp7eHHRbVoyiRDAEECr99tgfE6FJoqSAeQbxzPLHTnORJG7MAVcr45ijqZ5JPjX7YgS84nN61WLB
D6BgSLGdiL+FhyWviZcME2QmeQira7liJE9Vr3CH0beJfa4+8cgtlVa/JajHFdZ/Y9phsYxgbXaL
vhtZP8HwHvp5DiFw6LFWW8FV3lO3mkGmu9iKjXd+wJcTAxc8KcRFvbI0cSj4WhyH0EQE+77Pj71i
n/Zyzz4Kj7H0w9loB8L4TA6AdmrToCVa3EWJfZyE62MqzG4pBs4uRw2QzLWATGb1M5qqqG4OMcjH
PDatzILwBF0qbVbmX+HL2OUllBOvTtrGwYG9hjwjaUMXEesTzIChNt1f6EfpwZFSjx3Ys9Q6M+1S
19RH6sfRiEmozweeHu4IP87MLgCy1rwA3+hDTHGlRGw2p2kcR6bkmlHN1CXs7JLAYXafHoYERoJz
FGffeUsggzC96tT+Z9QZ5qCQl5G6ZvsrVnEKzY/YEbgi6+2I8LSLHpTqLojTV2hmwC2OwDETlG2k
jic022O7jz2YuYzVJsXCqq7PY2MzdNzDfYSPOcficgkBZMqAOlxCWffvS4KywivCQYv0MKcljMxj
98JCTCAzU9gaqnGbYwhXsTd5lmeIQdOlR0v/BZGeaNf6FH33YhOIJkSoKWFa6uOj9C1NUfGYvRAQ
+MTBWbVh4vBoQ2d+jmpIDvtmYnTIOSsAGvs3GqEfLhq7du8uiCq3glAO9Bw28G6mtNS36H9bFa4O
TvsUsKdWRWbnTWWGxIM3ZMfF85bicQCtkcuSn/Cvmcr5aTjrnPjnUEKrqVLpzdFqDMk+5NWJ9obd
nXEjutjdc40pTCq+HxuE+tMO0gXLBqCHYygjLPGusK4iQYcP6CSP7Osyyxm/lcxqbT1SXHchLaZE
f/4qVYdTGo4C/Ca4mFWMOs7aJ7/ICun38tecrfrqlbYwPOrRCjGfGEqt6UQa8XqCe9eRnUmOsiuu
kAbvnBQo14tiLP9t/0ZbqoVqlCuiVBgwFRS3nms+erW1bPlERH0j3gU83CsVn8VgwnutDaQ8F3bj
yLGGaG+Uv7R3lz3Nj+Vn4ocW1OHTyMvjRCnA3QMFOOg1HjPPSDCDoZUqJVhnRU7hEWeYnOdEt8gA
d11uzWOnRNEpzcXAO/G0t1xtQba1dEF7kDNkM8XYhHBVMmW/sbUGtByIuw+83rrL50f7xl6j8NtZ
jvXUE+vM2hXQKZ7XJu8CfahqwDJFRH08g0Fp7bAsXU5sGKWajQOkR2zbEzV+iv7b4+9ImkpSzrIV
e9u2K/Z9IeM+gaxl6EUvboXTdVY4apl5NXvfnJ2cGe1S85UJrNy6EO9skNQkXFMDsI6wm+NVlxiu
WR6mY2n06l1d47btpUP9BkFvM6xkX+TJPwfAvBsYJTOK33dAG3uVTOlOY5L0KSCBhdVQvYGtcDhT
f1M6thTucVC/fxWA9D2g3zqg97PmhfWt4tPlhr9ezyMS2a0IY+BoDfb1CwqVoAbYIKK3nIEflrtp
7uwh8Wx+NoqNfmcUgNB4dadFkjejfAps8okcj78tMMOWhHxYOIJd3brqo5UuCwvhV5YkDWJkriL0
MPw1XNBfWVmL0RVwkHE22buvrNWlyHXAU7WuBk2hLdQe/styxge2qVJ7uDqj1lWJdYMRzF3h8Ymr
jqw1xYklnqnLUSncXX7CIje9Vyb1IQ+1RwfUQ6o2odneAfApI6l9aJNoOXM8r9D7mw0ssKZe8ZRT
Eu+ZThZzsrzxAhSVv4IXm53HNB8SA8flqqKX11pJuqoRBUpTo1i2zqdTYBvpwt8W2i2HdfynGRrs
+SKieQbxpNQk35i145QBVxZQHyDdZpiER2MMApDBSuTnY3VtYKob8bjmrc5kSNzDSJex0X36ys2B
hxor3KrLW/6EO2sJQcPBBaBWQZUrqbqjnHSCeR16AGgXX0eezpqYQWyWGwf1uNmKyviY9A/WKO4/
VVASfbCOZYFiYKgxpljtjCpSdtK0T7bYEZsbA4bOqPmwvhmTAaQvojlWCIVUhRgWg2otoLBZSecm
xxNeYa6AvTuZ1hzLHZ+vbSx9pIOnkMDOAMKYfaK+lcluyqGJwgxTU76V1n81PeAS22IdQxBMe961
l3XiEMZ8B5nHihwPZpjYDCs2Mv7rpjyQDYMZMAmxH7mu9bwEdrGSmUKDJzVPbcTSjXKr3AeTH5W0
jRE7O70NnYLhxvCuCDiTgb+XHm+0fUFGJc5pMo07GCdJIA+xfpSq56fsyv1VjFC++I5pPCXnIOPh
e1lZxNGConJHIk/zKOf63z9PY8eQ0zKGVa+sHxW0/ZrNMi2M4wJBL9/bdDUv42m1AzlotB+hPgGa
Tk6qkhwzD3ANi0esTpgTVQ+erj26TwkAm9O34r2iY337B8KndgDbeG8Yu0oqAcKBHDra71AvUThR
L8tKSkSsPXNjDZtrDVeG4RENM/FWfyV4I+UW5b0Y5MG7NG/cgYWjX7sigAbxq6szRbpg2IJf4qR0
z0JgOm5fWBMnveE/F0lLxU5GO0AyaElODwOSuXaDOQ8KoVeWGS6G73mhAA85rbJaczUKATi/m2cH
bm0/m2TP9wWK0qDyEYPKg11lmb8MmtljMeA6f0Im8fz0ONe8nl1xKsubzrInBCLGSnORKCBLuWzp
HGUud3OEdvXur51ln+jeu/NcSpFpopMGr/gboZDboEvwtAS8QwojhnxbWTq9ESn1XgCoiWI1q6bb
tf+uGjcSD78B/H1oUv9iT9xXC7W80x6wZFEBiv9ejbMokiyGQ5o/KBfxNUaPTnKYjUa+aHnUJrqQ
wcieOcidP4SR1ogLOef1WotVoJjfCMA8tHyWGKxVsAtOON5QCe8kaBC+lPBk9HeMKeaLIM5Ns2QN
MH5bmjHUqV5csjedadWXKn3nAYcU5/quV8Wl1myzSGRY3QO5XMOrmcGE+11YQ5FIXFJBmUmv2v/b
GJ9BxbLKR/LsxKlaFOvQdBav+0XYpKzu5d4U6AqRUQYQxT7kC5+HDZ+1nmF9IZjsSu+iQTeExonf
lDssui1+idA5LCLwJsBYrj7ex2oNIIX1uKpwtyWTXqfQSPMNZ+ks+zy7npVQ+HIJ3pVbUsfIDMeg
tRHw1xhb6qqqTJbrXc+gYyyK2hFNlyc+GYaxq3B9jS1v6Mp5HZCqpCXvNPAC58BHlIHTEr+ZhCF5
EOCQH6+6I2OLlKl6VElSzywYb3oxVqB/9DiUILlB0ldbNwL17++ofnFXa8wxaL7/kV7CIX8wxlZD
VICxo4o84t1oPaWjOhNDetBFnUE/tMlvTc818e1WPXdysqpU3yr4QqqrRhLsfprZlT3Myw54/7cZ
6HFleUnURFkdpNoiHNxb5r3MdSVOk0dmD2ZiY7ozqNWyY+tMagyiHkWypDj37B0mZuXgcLD20OUz
vVu1K3hMJSMNdd6CwsIAU1AvmIpSUz2mkV3muyllYhtrKe+zRShVC9WG1s9NV7RyiAwfkQE7y4S2
fp79w2c0E8XvQbYf9DaT8RUbvhpiUwYRI/3+gcpSeRfFFgGfd7qA10g7fcH6oxYxGhV9i0nXgD/f
Cmld4yQt50a6uo5SMaIP3COfwZBnm0gZGWs1m8uumxkwYAe9XTYf2xMRYXFwj+vGyHN0zwO1YfBk
zYxFRHjwpFIM3SkpE5s6CZ0DD3ICn43BETpCLalehkIC5ELr1clBKULNT0Nh2mQsr4ju6K+Md404
pCLXwDN/6Iiz1z12hoZ+RwQ6Xdtq7R0GN6Eu+6ddWAMuGnaG0nUZAe596w420lNhBJokA122Yxrf
ckD2AZ0ITED6uE7MEiujKfgt8bCic2boeW+5uKx+d1KgZErqnC7IJ7nXq/3F27gor6QaWR5tLVHP
gTOQY/ooq94EBSkBgDFXjg+bNvZ4+1pdvFikrdJRHBkeSGD9wWiEKwdRtmqmMggO0a3rD491kGF3
Q+Fv4vigMvEZD8neRNkM58zZrjn6wyfDo6Qyk/35CYqq5fL2hdqAI2lsh465SQ1iWlDcsZ5qcFar
AeaS+9UwRCyydc3czjPifCtaFCrkaZ3ht219TiUs8YyDeqmmbDnfDMTmVwDK+Lk52PZAWRisRQbx
l356pDO0Ivq4GkbUKmAnZDdgph9z++xSnFhZiOcNHkagozFC7tJMX9KfkG2Ngd+PM9szI9y3PLKx
RXcebfnznd/fB9Dv8UNCuYfniwowNPjSE8eUOVHmZJ0V+BtzcDODu0gU6VyqWPFou/IBJOpJxGtf
xg/9zhtpfiGKpQTqDfC9gvh+Puo559PtVU6Rik9/RBuELIfmIceWHp9skIgu/sWU8ByTGG/B8Zb3
eZ96bes73Xzdpyn6bxnjaUESiSkMMtECOcZXaRWV17y712MIpAZ+hlkIttJJfqxHHP5CfxUR3hjt
fXg7XkFjd26uvrH73Cm9O4UXjYhQTxyTnngBYA5fR7XTvLVjAj346GhBv4+x1Lvr1Bshfh6DrSil
Hqij27onIycB2xWmBeWzSQ51zskpvEeoXQQTuo/ddbpxU9pau1hbl9kwXIgxidVlyuoqKOp8GoIb
OOfIUz/VCDx828hU7tJIq3NQuARynBKvkYiqUF8NzrgmcfJ1ry5f+ZeRtaZt6WlYH8nX9QeqSt7m
vfzirajLGw1o1pjKrsaiLo7jf6tpqA4iHe9TUhXkJm/RX0AssWnHvtLDVt2AYXafsED++PcGwTVn
/M4tM0ZTEaa16bwHQegICBMeoptf88ym8gCx7rzawE2SiaERJS+UiHWN0r67qaRCCAYrh7gwRYv9
py1Zcv+KNE26Eg8/+QfkzMF2zrPDLYT3G666Jc48ufez46qmixOtkeS9lrN95BtaD42grZIq4iEi
Q4n5r6FZK3AfN95fSYtcjA9QJb+tD7Ui8oBNnw3IVFUuru60Yw0X53ZRF5lMyeXhOUWINVOW9J52
4DKUokx1vT5g4LIq24fGEobNJ7eMJMIpR6Sv5jukt3gK7xGPPdy7rGCun8NTOMFbwUmzIzf/MCxx
D7Yav7QR80MOY9FgjLNQX7SRZ/U+PJz0T+Xgbl1fT2rWlmEpQ2kzJwJTzv8MXW4Eb/fEgw6rOMI/
A7kjuUE3O/oh6ZBOcdkRkuvFNBAHvQwAj0ljahETiVNfkl6L0mqRybVCEiPvncaNhCb+8BUFqC7D
e+C3VojYxaI+FgI7FjtIeTzSG5mlgAUy+CB0V6NACErYmq6KcV5Ec/LgKe3F4twOtdJoZk1hYemp
eGIOeUth8JDB43umbB22UU2Raklhd2e1W0oK5P5B2Tz5zU2hrn+GS/5ncpguagTA0pEuA9GqA0HD
gCV0vdRToP9X19CUaYecJzbjXf0PWmZcJiurkcQVKmBg0aHSFyDN4GKgkvlYr0BeT8JZj78gf/ah
eilwRHYWueUdoyy2IzvN1tHQSBci6LQPd+sAyfWi/8I+JCjcocF38OaGANgF/ndahKWojTAi6zJE
oQ5lbuORBMtt+HIISNqxwAbjJYoes/0QDpNMw9Ezeafh/nbVRSS5b23iCZ6BadFmttHCfcmpzNKk
qRYPIb4yz8cFsHMDAhYBlpCjhsfctbPQloBvJV/O5SruUa+hvL1zo7j38Xt1pJpKeaMJZqoQqkvk
wvxa1qSnX5qyA7P8I1Hq0YdKe5DiVJsY4P5iq7NmeYXGlQAFfrb3XYwAu2eA29CSyKTfYHbfDlNH
FuDFiENnZ8t7Z57aTrcl0wV4ByeyGZ2aO+okvi/rpf+0s3TMdWNBWPBuUFIiI5ND1HeP3Uk+czZi
nlZ59rEaxG/xFsqqrknCNIBQt8C/7bCkV10nMuI2SJNqqEMa75Ok6rjkkOfgTt19BfxXlDjWx+5a
oYgS4H56rHsXTJDhyJcEPveYqPn9qKarZiHlrbEgfuT3gwJ09o8A4Br001zYnmb0hydHxelPExiX
BN7G3KMHjp7ly9mGtAGAIwVK/t67JaZmcnIB1Pda5BBOJFa0eCDn9WzDTy4+EK4ZnOO91k2g4PFy
ez9DbDvfo/dOOxZ157firKft4cOJ0WWdvzAEz2jOdpymaUV8m2xr+0mtmLtGAdsJW/y8sjxKgxBL
7OONdjIGmpBQf6VpDc2Jx/5HGMBZ28kGiN6twdvNi7UT3cjaB/RhGq0O5DO58a7wy9qVhXrUN0Re
W84JpuBJHKb5EEQmdpOv3rMfuQ8emrrRQ3AvLrktqOFTKfEjRGdDl8d3UUcGygwtgISJi3EiFdOg
sB9sGKZQ0wSG//s/LYbZ1FO96JOctm/nExjgEuuarFxs+pEwUZ2oYyLNUy9M74D/42mk5IBRimOX
+WToohV4wHVenGY7DYKosFgORpUd2DJLLbqkXsc8WJRpKTEDsWYuIEXY0GcBqAxUnSzFtFY8R+LF
Ea4J8jOw0IYAKJmiC81uxpAJsxV5ANKBm4jNdS8a8jwRY5WmX7CekFH7h3I5KXGbKKoQUUIiu+zQ
aRUpwTZ4yT0VE6jrMK5qoaRF/XSB8Hxn/J9Rk9cR6r0Jd995kuB+03JGs6OuKncu4Rgx4ygsKEOc
eybRkEXSurjYpOrCWkyxH++t8Grr46iEeZNz+9O4yTMr82c6xO1CKFeGmbq26o+z+t9zYk9Q/Cp9
bZUQXvQgyPgpFK/ukmCksCE3Z80WKkA4+S94LVor05gw3iBOmHrgStbsoz/44G623Sbumb3BFwSp
pPGQZ2uT6pWQG1POENWfKtUvfIaeQynVXuKXzmL3q7jwtYF+Z7FOv+jwo69HptGi3mrf8RA8Ip1R
+6JS4JPqj/pb5Kt/ruWKGA5Y0aN1ek+LAasCemO/7ecf1MZjAGMrsGna9Mjaa4iUQE3PK2zUvP7O
BLKMIXbU74T1hODpihMomeQc96ZJZgQx/FmO8hblnfsi4UwNAzeqAjjrVCmlJKLyJeCQJlRp7DG+
AnfSzLxihTO/6UxrVKuHvU877nmcvOXa2r4R7+riG4QoJIwiaEc8ZyGiyGh5fh1VbKX2klTylHts
T7/JNHl+J/u/+EH2J33tx9XUOoY3gy4Ln9izdlu1WjtwC96878WPJqtU2dW6To26f4daVbn1UPM/
nXpJJ74G7sGJdwvQPya58BBbSnGHJ/VdZRWGV0osG8iji6BstQK8Ph9tftd0QVwehUpm2vvPhiCE
Bs1usmyXzmCtX15nEQ8DhVOBdLR0olA66WCNhciuA0g8F7amaOe2X2S2RJLNvVTb6lccxA/oIhZs
oXyrMNSAyAyoX1Ze2c4diQ7Z6w4R6joP9nRCoeqgCF3zjjV7PNACcInU9RCZn8ugebMeL34dNpFs
DCCxThci5WfarOV3ovHN48cyUfCRRviFEn/uGVT8dNNWG3PXVusE5fTv0oSBDEiorwdi9x/6ZcH3
bqWYQnD0y4K7cnUZgAetW/EO4vPlqe73QNxQfp/HDuIaspVBK+Y1R+GBW1BkhX4dWKrYGYEv9P9d
nfdCMu6v6WklFiPvzg+o7qwLYrW2pVmoCptduHzvPA+DXb9eFKntt+3jMjFm+Sj934o5JRAQp5oJ
EJW5foBkqDzSwWDWpA9j6qdxbpuLpQFPQgeLylR58/SW2YE9ctYdCqW4X7js5bNvafisM3rgdqbO
U3TNBNmvHGhSrWJE6sXOLfxv0Bqropm6yFwT1ySgL2d7z5mdabz14XX2Z3BJJpUt4tv/o8Eo46YT
ZeV+FSf0zL+/9LQqrAXlT5AUsxJFJcSjM3vbTZ9da1oVH1m8OdjVlsTZxS4kg5Q7s20weN1cbQPg
U660XvSpA26d0XgKRcitmgxANgTiJi/CVsDuOLDdjpw9NxQjHkcNjY6xtTW2EJIw5xj3Cgbe2ujt
lDvKgJ+RdtiomqUughF1kLvgC8E5/zJy9a+7+vWh5NeC91vMtkI16qxRub49Z3liFdIH2oKkGraB
URHfgSHbY1tJtxlAeAHEZLexSsdvw8V4f+uRo/Xy5kkgHgzcWlJyvAMGLhEtCGUnVFOYzoPywhH/
H+QwKk+VtuU7s7L7rpYpZW0d+XNZ7/A/M91s3RNUSL9JNy/lFl205znVPDuTBICKCMIAItaiqkMZ
YfaNgSx1grmyVzl+ljFFVVavXucdMDk7pxw+Sqpu8jUaKqH49XzPOrImgalpVJhmAjhc5exYEqpi
b6KcM40P73dD3+3deR500/Sw4nAELohnV8wl9v65A+kZkPLnQeDh9Ss5bXAUQXBKjk1ev2GRp0Nx
iWYcWm9uFQA9vojQy0nnO/5LHkH7oVgYOCPnCKcT+VWESZ4lk3lS4VdQWHcNxgEWLdjNs3AFgUqZ
3TAc3ywjGJ2DM0z4ORqfnCF8iLa2fWuORhKdnnsFSK+MrPmNzuDfhZ85PuLSJtUGKPeCjtpB6QQ9
mXNT0LSjP8ciz2En+XcqRWsZLPEDL7RxJgZhavhEEf90vrY7qpfaggbAxz4ZMkyCzIVFgwqOb8If
AMlHHUiHPbH8mDqTdjVU7weYi2hIImq/SmVroyffwpRrR31laG3pQ1u3CLoWXQBQAloJPhI/fzs6
3Ge/xITVeXz3KH1jkuu5urFTG8q/QG9dx/92ywa3o2dX7NpwnLOWfRQXS9ZAtccoTp5J1Vuw26+2
eNBT/2n8AIYJxE4ftGIKnIgJe0UhuC5CpDY0XlV6ncNDruihfmtupp5WzXvmcwslaSH4xBYtwoGC
RK/5y7o1PwjtH0g5qKpvFk4maeyYOga2xezjpHF125r0DEzegP97//Q4nExCCVZ+y4ms8aCCSm/Z
K1Gd7AhOY0C8EfOLY4bO2ZFQ2+q/XatbCCT0Wvs3DPtEiLoGwp+dUlnA6fJdckoBYsPLwXiceMqH
yvR81sWES2Xqxh/2WLu4NP38el1jJTDa6zqJC5yU7MPn+LnoLKF4QExuEaiVgEVACn0MGBspl3VB
ZmFji7wvAgTB43vebdV3cnm2tAIbH1K/MDN+NKpWxno6Ac/1upMIaIQlHIE4fDvjQ8fND9vqs+Er
bGj3flSkpH2jZjYwKJn01Dl3zzP2+7jFkszsZRImftUvEDXX5jvg91lngHxz/Wam12QTmAFioWfd
n+ka4KDlAzHAFQXzKMfOJ+nAVHM/BJVENvH5NK0teiW2Rx7qm5rXBeAFo97rejA6wgKGRJhopy3g
alW3kuLXb9vC4RFO74tR9mkYzIwJUWNYiR/AH565ct4LoGvPjSH9kFqTAenZvToLOybiHNkVTvpZ
kagGDv0o6SqCg2GKPIHR3F8mQfCApsiDMRs7Gaic/oGCxsyfRVUVxRI8ay0Z2N4+BMqxBuiQAIpl
5/+UveYfsu+Shtz+hdfN1UQ8D3/H22uV30uvYpKTrTFzLnXmVDvVyNKjafAgaWsjURlU2f8AD8uz
BQCQqR4txrv5NDv1ARDJ5AwcEN71dZwSexVTfMaQ0SVKSI+casJ46rq7ia4f/oIzk+Aqq/XMkgPv
mzcArxlMsCyKn53vV5gILGHtKglCWWt1FbswkMs9brTPS5fLTijb867eFNY8HKSzc5rsizLgzrbR
7DiGptjYe5Y6LAqavp1yHy+XXj/HVtQGZR8ucBc3mQTaqE18c2n1/MR71urQYWzbgauWcV+O0A+N
2dpaciEzUv4SITTE5zatQb4oAGiFD8BN0CJZMa8ymP5fJp+ByjtMlR3dCrA4CqyNBzkVw78caXlL
q9gKgTwOVJFOVwiyYj5LcA8eTHWDUG97Cum3TkAdKeMb1l+pN5XKULiViT09vRIhZYXGgnAg7zGe
qbSOC3/dUw+GXKyB0pC6Yf0xsfV9zcQrd67kcKpvMkgOYWMeF6eAvKK6ItXZT+yUqJFZLAekMhug
dvMkTo96h8CLqGl+8UG4CXCsZVqgd03ha3AdBKqQ3imPmr16BLWZsA5MmbeHG2C83vyHPaZ8Pcup
8AKGu4biEreCwDKd9XwWiZD/cICpWCUBZeVENZjjrYSzBDCzex+ySEcVakV0zZg3WnK03JSlbDMM
3zGQiRtBMeu2mlMpP3BF4HXRn8TSH6VgVg+l9/HoGYZ2/77vHtPM3p9+r6hchLQS9FJWWgbeA2Z6
HbSxuAfx6GbQKs5ODDRTdYF2eWfNQZP3cfdhlEXjbkMst+bKdsgkYlVE0UrYBKH8mN+7EEGm8A8U
T7rZNU0qF/CzG0GVlYguFEj5ik15X5mCCSOg8vbc+gkdjtNdkTbbVIs0OxLRO35Xcbb9wmxYADbH
mniIgAkPuevPbf9t4u5ZYo9hvwb5od1qixtDn9lOwfF0gAU5R/RWHZ8XmsPBRy7bo1S3BrvXmaG/
WViq6lAeesI4VmjmDfnt2qdON80gA90GOvFDFJvcn/elXWSU70I4Mf9Z/cmVzdZxORl1caN9dmJD
cVc+gkvZiwa+48CSePAkckoaq28Nli8jlb0GnjGncR3WJPIoZwdQUt2VwfGo1RVXmStdo+MX09QH
DUbATFGRNRIEpDpe8+hgY0TplZghKh8ECe+35wYV9LeJmrnTJcLI7rMjbxE8lxkjG5rY6B5RWOk3
lNpugPI23mkhVvXPfVscoxABqZDiwhx8nzJ2B23rf3noyq7UNGZMROpmiZnZfrMHD/ykmqDN/gNn
B/9A+V6wwcKSbUm38+GSCLA6JATbMPcMif+Cogx2fFzenomMP2Lr8HN+ziZSDWxJmnA31P3DUxRr
SmziTZl+Ni7eX753MktzKJHXdBfT0Cdn3hAJ4pp36QHRhpdqrQSqRcmHdUkIKdCNAlb0vtGXKXCO
3Ids4SfP4l0g4OY7W1M6FE7k4p+3T/OWgJbK2WuOqRM4yIIGm7vwax4a58fN8Cux3QKfK+8ystYs
Y61ibE7a4l12wobT7hYu+VZOjk/Gwvqb4QN3aNDcWtb2HNuGY6H+gCsk/5pKDEpz+cLyssktc3wg
Va9Y0Ksv++5IZBjE0tQv6SNI1LE39IyEQU6inuDNKws6Zu5mb/qYKgnRibzDhg3/4t123dJAV34/
6ZIlRgB/lOAttWDQrpne8PRHCh5ydZC4AHlJKmAFcQXAOOUhDGwfJeN4MrQtf3ty73rY0wHkTy70
r9Lw029R7GSyPW/c89+BKzNdzqBj8zaOo2yJg0Ev19mx7eStftUpv8FL/es/RvbkdDkSl1mu/taa
9TVfa4MdjsrKTlioq+/KNkvgUaD/ux4YJQnqBtpt+3/sbJ21dw32tNo06ye3F9sIMNuzyf6qqzvW
b6ggKzKomhoglnLHQFsaJXnQmhPMw1JgKuSiBQ35ozeEc4wsEl0yKGTiOasLJJPAZcSIIQ90I+FS
eFq7uUXCClDTxTjctdk+CGaAaNdgmXsTLgVoniEQZgjl9DPac40xXhbzcuUHe9t84/bQfyZyS6FT
4FEl+aHTKDpFworbU2iVHXpMjzWx3f4RQORDFHMCjPahYXP68cuvlAW0duGbt2g7WCHBs/BH37bk
Dbqj9mroigI3kKp4StHBwEoLTlQ4vQRB4CmppqIpXqXlGKE4ZeXRQSzMPe7TiNeFRTzi7TuFotn2
6d0Zysk25pUX2cEpINdNgnxTKvIezOu1yVAGrtiDopfI37FefRsV7SENtoluNUJ2FyPIpL1hk/YY
Jlb1puNMJ2kTNsqlfl+6DrHILz4CFXMSsiZ/fDSWINkg1Pzjc5seqpJR7qhtsxKuwQnyGJva2XUZ
fHblKtmzPncYr4eHLpcU84Lkyy5RpiptSiwL37EpVT0NXBrSfR6SDrxqw+O/F/oVzCyvCZGiE3Rt
rVo+zeTSmq3GpZJT2oXDarzv7c5INaAzkAVWYfZ1GFhKydTjjiamJucvzL7xs6g69GU7VFuMmRDZ
AK9Xt1EO4r8GyOIT5LF9oLfPRKg/KToz3Wa05OrECSVcjHIuar2/A1GXD7/zPgfo7DJxMXKFoZVL
+OUJkP8ELUMoq9DkVF9AR0NaOd7ApSTz8J0HpAN55eC+griyNSmXlLZlTilJv7k8KIpdmZao74+T
LaquNI0KMx7y69l4OlgFRMinS0VN+J8Pl0iHj1mFU0LwSD2hhZaQ4XIe7BZ65zUfr6SwcVEP8VZL
rEBmQYtL6T3aLneEKQSS9BPpOv3YGHB8pCEjh+Zh+Ml1ZmQVwBKGXmN4jo3d6EMvPW4IXrysA/ow
W1JZKiXusVWDlpUfaljTgYD3eoN1MPVNxVKql5rbbgm8YkxPPz8qRtKB3Ounjw7DeN3g+IL52egA
wUCwncjP8Ls2YwBdGkzeN5o+bQgbeD1X/4cNTBrop8u850jIBs0W75Ooox2/LsqJ+x2qW7yz0vy2
tYgm0b6vUEqoZo6Kqkq8e5TpawW5RYmE/R1xy4YaRpS5W5ykMTlo3MHF+pID6hP0lq3+uGJMH3Vh
lFf5KUYzcpltBLbjWAf/iyTA/Bbkuq4yeF5EQRxir+tnP86y/jqRqyyTQJCkEW8p8jyB1oxRQhB6
oxbwbfXndp37OJTj/wLTPiDOTyWZVenEBvVBTXbARU30pJQJ6sJ3F4WOcj8pg1XIiVlvCN0pBF38
gTpMQ2mmWVIrBU4rW0FhIidZmHbOiLvhftg1d25zI5u+VqYTYelXCRmRtTj6WglRN5UMW/on9gFn
iTFPtOhZBS/kYep1H0QVFI82NFEx5lRxnpFxctvisJPYeUZFImFOQOPMcUj/e2DhEJGSwIB92J3F
d48M9mrrX67Ij5KNq7mYAw0SkAmWAUe8Ri3KY9hVNng1qhdGwBDVr3iEGRvbgQ2onKpAdcivfuIP
UBstOAkNgFl8afff9nXXYuBwU8PCCKnOE0z6FaK6KgkV3aV90ddnwlYj+Q743PuPygcPZgRB6ckn
wooLs1ZZxGTrHMcgXRNm+Gu/otQuD8Py3mrD5I8IbtCUfVoonjS74L6Zxel4GHtwSrcBfOj/g0/8
EFBa8x4WS5puxxc7GTHDiPOovQzuX4UKmJJcYk/tIeQIVdyEGYWvKFLlNOgT4+tdGOdyYiZdVvwn
wLDgtqdef/HaHKCJmW6DTdoOJmBwGD7E+yeIrkcItx2tHPJAJ18g12QC9tTtA9WdlCxuWQrLUWb5
Gzc04m5+aAWZfvHYXEhKIaISGFpywTs1D4neOoGsoEq1j0cuOn41/385NrKwvKfY+7wX6iSKAFq5
eYt81918s+our+Xp6IsnDZdNZRQmsn88D+i2mrcOrRj7ozDPmcZBOY6nR8+7KvrehAcm/JreWxu4
gOUIYIRkEPCsry6gu4dCCraxVn5sjR3EQbqgmpBLBdmtMh9e6FHew4DYmNJhXXB8lWKr0R5QIQoV
YQZNt72IgKi+kg9v68hfQu/dID7T7kCdnNRr6LYlcme2RxRI0L0Tf3HYJRSQPbqjsjTqZvrdteTl
ns+Z3mykwMz/rMoKyhBtFhhqxGEYpsLyH02QspT220yNKKwlnyQ8C6qWbD6dsrhtgNhp/eo25yLT
/ZBoHLii8ofiSh3R38lwxo5N+JNJ96Mdeqz8Z3NyoVD6SsVJk4UmUPtZLzm+D1AFvTNR3FFJNCsQ
mANU8qqH3xdww58L9+tQZrnjAd5LqvMkYUwC/gIHsTqiBVONB2PkymyW1EYgwntZXALij2i4Z8Pf
R65cI28Wu1mQFVvvTpWCSmbYW1stTT3m5TDsE/5gs4paRn64/0uU2eJrfXYsQrVZKPJ4bx0e0K8A
emqAso67lLkI9w3/0Ka1eAl+iQIW4LT01s/8sYIGb0oZF/5uDN3n6Nyy4V5BBNjHd7vqAyrQBA3e
07U0QFg6uQSIHkPZUeR882aLkCVqd3j3wtCLhm18Kr42k6d+CxUIZ951Nr7RWhEWfEPUw8dLTu1m
3/SrLZ3CZp6849z16tP87yG5ytrAawYAGCX8WFcWkZZxXgJh+NkJeMZFCt316GhuOyR6L9DMstbk
8zdNBoFB3WiBDcSkIP/Tsh252OtYy33F2jXpj98vxah1JzUA5cLdRlMu+oBpGlmcfsf7VLHE8J/L
yKXNwKgezBoZo4Q4g8QsjuTOxsntJuEus2d50q5BcZkoftty2CuWNbsOWysU0AzDXlX/kvZi/Lsv
PrhCSfDziDJjrGt0oTC1gfuvIO1+Q5IBp4zZj6FxM/72iowvFWKNnRNYzDs2VQOTGR6WBAT1TjUZ
XqGGYkHXZbehepussfgVKrG8UaDKknTvNf3llUlZ/uIY6UUj0vaXd/Km7wmEVeY+NcyKp3to1WpV
dy99OOI1O+jvV9nWTq7XYx5tGz/1xTjoOV43tpHofVXsLT99KTce/JfsMeFz2N9idTZ/ibAfNsqj
DXpA5Gub2uvKDkhhoNS4DUQ0vSOCPObaM3CqZaCYGTRJh4O776vsJdX+6DfO5YK/1Ydre//ImIQE
MRjfd0bpC3mBHrTewDnwNjw0IKlK9/+ZAH0RuIC2fEEuRh3TIg16Cq5xxI1nrteJCYBhVrhaUSEj
81Y4wSR0A+FjOfXKfnWvSsr6ivJImCqZVBFrY9NYR+qqHkUpLk2WcSVNV8r/lAXda98YzLdl0X5v
tkm1Yxln6WtPdrkG9cbDZ2EBwtDa8kJUyD6zzZ3HTTBxYJu9slm2RD1uzLUd48EQjcG5RNM23iYz
j7NZte56+9LaEm1zTfK/e2StvIr4WMTOL3nfKbxIfgaUCS9kJ9W4FwBWhgLK6FALJIJbHD9WxHNR
/QblpSTlhhYQ7uC8t2H6QPy1q281raGiN29yGgAMczEmKsCaBcOK10TkQhDIpFLeT/lKgztQb4Qh
7OrCjErCUGUAPjqEnGs054CukVMyfnufzHkeMup1mtMu9HRQL7def9TPvYqTHdsoSxQU5asyjB/R
Ugupv0rsJsk+gT6HjRN0DR1xdnvg6yTiZJCy/YvC8mfbMrWSAuyJcbwZInH+QRD+5T9KGwiS/nho
S42fipW2c4ga/8Jjm3J7tdRpz3AzWpXj9S1Fltnz2bLOiHDd/dsduMxs+1C0zpMYqE8h+bXOwDE+
zF0iPQaxUFogbTgilmIOz89OR1ihkDXZhK1w98njFIeCyhNfbN0ttfC4ZPTOVy5gT4hwTH0xflBp
4xXvz9etpbZ3yrKWhcS5WeiHA+8d5C+YhsljG0X9gQZxhJpYZTfQb4n3hX9IV02x8YvxSdNOR/WJ
SC5zVpOURCvcTrE8I0xUhYQhgUpcfsjLAqz3KTzkFvKZKCEIQXWuxaYoU9fA6wtoH01hlM0Zi6tO
mR+dFVNkrs99vEBLHy4Hr35cLpKTuUaZcAf/IEvBeOoPoCP18+3R2CvXmg7WfUgmt42arL4OobK1
T+yMRogAzKqolkK7ikEYa2FZ2zsWgGva0/ObHlz3cJXNmk/sSDLcfgbRnCIaWudDVaPFAwgQzHzm
+MTD5s1gK9X2vOR1Kxq4wwKk50dXPaB08dvn2uZbGHx7fTTOKLTZA/bYJlgT42+FyFZIja9SCOAD
Q1iHqgBYEtNGhc/aZ5bjsgdIcPGfH+4iX5xQb7aKd8FXxrV6wBuCfsU6h0sbT318o9s3WEr3UkRX
NvO5vwHt0uD5vSHp3+IbVg4+H2O7Qey5mhtjVBoCXx/koKOFq/7/obdz09fk+NPTmt8Yp/0x6etk
0Z1yOGHQef9gi1VEz+KW/CIxdUKMIdsbycM2QWvvDb8t4Zbjl//3viEmzz+QgRzX4JfJJh6oqjr0
6iPqRV315nVEwJIolm5zibO/a/V/cLRZEgnQTPrPEZVlFidg4kbA8mIMT+1IukNgvjT9Wti3ybDo
M9jkC2sZ1rG5iXJPG39tY7egrf70eyIl4I4VNQotTCb5lwO9OlhRuj0MDKoY254jezcn2jrPu3YX
pZyixwV0zAXlwJB0rGArjq0g+8+8yNKdzGrcJlluNTWwIGJGAdrVDKLFAxrwTK9SEhk1tU9iO0SL
3DHwAhcKTZP964FkA1eFLnPJmRB9uXKifLyfi3JX4RlG9F+OB802KwF/pMh8/LyUZzLKzVpUM6Oa
9mTAPnT41gRPc47ut3l06voBIKQK9dMNJPBojtOpnvBogEJMCc+hlfrKvWmbxRIhe2bjmR4glHBm
Shl5YH3hLBxCPgC1OfA3tW5Qj9TAzJKRAhjTXjS0ekxI0LfztHm329uT5HVutXdDqYlRBpUrPbhK
DV0/p/56WukSKzSfxB/R+0tXSI1hxYhiIOboW9B5rrGIC820maruDsKQzghbSAYs2ODZQ3aVcHuM
vR0jstKJ9exAx2L1hnk8YcOIfBNUxStcL3850NuAeRcbOmR4uwPMOSwhca/O4wnDrYezwDAN8tpR
XXB7wOex5Q1fmNfZZ0vI+wnbmda4KG4ATzhtfp/S19FJToIxtj/C84H6AsyynfLowRESn535RUYf
EQKQkiL7bWcF70rG2bDZZ+RWvxhR2iHFTR60U/6suLWyjiEgz4yym+xv8QmtQa1346hQ/hjFUvKc
QgsQcvgWUpWr54BrA4W56yYpG+72P+DtLrXkw1Ug1zNA+K+7Kkkl1JhR0aeA2i/8IbCeN0DlFRG0
h6QjCXn2Wl9RcLI2RsNqATOOpoe/IO965hTuAdg2hdkePjgAGDVqdsGsDXU8Jppgh8pszS4rQ48z
LhskWQy7Ckp0cGLQ5F7JCkR4LFdv7FQEzPVtkKJqge04ma8NnhAMupLWJYSwa8erywAWRUl1/kcM
So0TgZ7gMMM0ZV8RSqh8zCdBe2fXtuSkXZA5jq7MgOjGo6B+4XJtlYyPTdTkqCwfBMhM6+p/EsOq
GPfgQeBLD0kY+iq2cL9lwNufX7xNkQpm5STXH/AgL70+rqgEy5+fd1dTglI3OmNGOeZWPfJ3eqAI
UKybCxi+rhSNBtqoK0enLQVf5anc/auNJCQ9Jxby2NrMGqFZffZ0nh5I4W5T/4+HsNbO55yXSk9P
NKeEj8T2Pd50kUSbd68F+63caKQlCWdZ40QXeQ/SKp87ghvv4y0xhc/OdH1uqIEZ6cTAXpYLYnhk
SD5+R0bHxsVj7u1WHpSCifuNY+J6x6H/9zA31pkYcIqcDjHa3EqmQH/ZD8/VP+33OQp//b7i9UjX
bZ6xLmfM+zDoqMzRO6wm9dlYSXJcSR0JJH6ZZUd3ABQOzgfJ+frS/VkvisdxU5Kl5C6w1fkLBpXT
zXEggrc2MyWQQQHYqHneiprCqy0HdudqVj36MK3mD+g0AFtPOnwSG69MSMFMpcYfy8UaTYDkHmsJ
EzVSNjaq79kL+5caPzAawzQ5E0clfvNSMwF8tPdDzmnxUUUEzr5j1sLZfia0/9rRFbtI/ipZsMiL
igHxG5RwPpHToOk1h4cwMSulZPiLm35dd2ltDb1HMFJ2yEIkK9XFpyNIb8qFUFsShvpaIw6AkQsH
DKo1ekOJc90+iT6pVA9MrT/4Bo4F5MSo/2RWyTRnYePRs5I2c8U6FU9xGloLwUZytJUbZwBKvom4
inW2OTq9nGV+tP/x1LUmEHkKGevrWPheiVHLzDtHCVcXuulURzunp3I+U/OhW27LWAywuNh2bUI1
DVCQeD+r/kL6zgo/UpYhQ5N/rI0Y24PjNeng55aFn7/z45QiM243307b36t/I48/qefMFrZi8wzx
O4tDocxr1hkpvI5Uvv3/x7ItGhzh5r5unJm11bsg3w+AKQIWuul5Wg3xTzmKxdNFFiopxdBhFDdv
/jMXbVPqAHbUWRnOInlTwlQYeu2mYJzDT5QIB7JKN1ofM+Bz/sXN3AU8nwKE4+cHosUlnSzJe2Xd
t9DT4K0ey8sCJKiGll9iO8WNDhQ6FZG9JDnfGVAb/NQZnJUtu21PS1wvE1sBalwIggmyZqh/ADsx
0O3ZZyx/RqiocaurNycBfDUmQSHtAmV011s8xDv9qQdvI5lA4t4Haqiwu420NqZax0xj0nz5lz9k
m2S9vGJNmf7s31ADxTxoH4BM+iF7cvyy63QyI3ELov8pgAUE4HJFguhLA+m01PRxbi0bVXaTmcKv
DpS4pLTBl/VdjUlFVCIyQPHxdmMom9Z2aqnykXoP4oamF7LAa11Bo5BTgwWWt3llFDC9nfd7dBzG
0G51x/rABaQ7M0Rby6h4XgWwMLv0ECgcVwsqq1ubGi5LexAxFeWW24sGMbcRG8ci+OzzLae2RvH8
4RotBQD29/dbV89nztmhm2tHJVOX8NNghcVbBBBhwzPeu/4KUjHXdeZ7LakbWUMtq2JJRGBfs/xP
X0z7X2oZDkhXNXgZuWKjdxOJt6EBNuwODDzL03XiwuLt2s7ja5uKh2+QF6agXqFmOqqbOoxahYTR
Oc3iVqyNb8nYXbhrTXOG8QWm1D13MfMXwkrDBiHnSLhzpYkGTno5ueN9FPBx8tYIAiCsbvzJj7Es
i12Iyvf3j3/xi3T2/Y7pyD94Ah0cTmbHQ2LjwYqlszKJU+ykVUoJ9e2uov2IEOYJQOEtdX6lWv4S
iGTNhBUoiX8VmFMxF5/1syA9ExHKmx1ipcd6122t1SSSLnmsgOy0h4lnuRY83hLEbOOiqazq47Lk
3x3X2sy7iTd3RZU8Je8eSLzg858ued2G8rJPirQAqxzwfaNqJTilEfXEEk5XO8lXhPQGQO11MnZA
+/Ue+HGBzgHTYfkrTAehfSCtBJONw1YERmeD9a9nHcWVRLlbvE1CTrsqO0WgSUCAs6nEfB+BBh7z
ycPn/J8kulyDtWfPB5yBByXS/E+KbnW7IU+Hn4qaJahUOAaNOxDoPM7XrvowWPQ3cF/e7W+Yid3d
MKQnNkmoCvVKzuTYY6vbIKlDjfZJj16PfyluIWPPrJbUY+KTAiDqqxMNqy8vHeuN0d9l+waRN5nF
5Rui07rCM0rrHnp3UxxZLYYm6UPXSKmlsrGVzlYQR9cNS6q6aAZSb/PQK2KilWnl/Tj67BIvO8T9
sjHcl8MXvYqSSncmb27kkHPAhtYAPI05xGUrOVv99uhoHquRlmYZLFoiF0/TIE9HaI9shd2qV0Eh
J0C7hR68ndmHiU+5zBGI6yV7hBvw9nzP/h427/uS67JcvLjIMkMCJhoMcVROsQ8dV9RBLS9hjSr+
mh2dHPVAp+g5QoK7LUV/43cMwy9xhvd2x1EqR0ilNRYnWIF1IRYp90XAOkmJpAQgM55IEjJV0zDQ
4mfP3lHZHsTQCRpGx20Tu0LIJmubyyZ6LAkznz5Kq+/BqpPFwglDcX9WRSGTE82MygK1RcLtxMki
GnRNDdxcGikOxUWpkGIOOZqlTfUgOXmkmXxRcUDeIOILbIz5HNPENPgkuZgOWxquBGqndE7LPYzJ
n0U2Cl7/uQzsRAmPO1fiXku2THdIT1JpjDEQnLvMfw+RwX7qiZ2e5PVSktQvcXkLI4035Iy8+Y4b
zPa32ytIzcqjS97roKRv6nCJxxBxEnYaWh5Y0fG4gHezJ0qqwOsC20oVk7fBuob3NBAqbo76QGvH
czmKuQKtnEckuh6zWFYQkdE/hfJ94IuvIDoqj62+C1mbjSCnrwU7mObKMyItkB4pOFdkyr1JqEoZ
+f2wkDDaLB2AuVFLqFBLbMWqvegCXt4NkgaEMLd+Tqkig6bk9DDDbZRewuSxrjlBzIQ+lAzgIqQx
tClunqkhZDnhgjZiCGCKO1RRATY3GfyRMfqRo0oIwR03lPtX2SHdWRf4kCrVqrPj1b2dkwdbF24U
/feW98IMGsmzbejry2MAI+wqn4SCNTp/WQ3t+GsZQ+IegVxu3lZX5m8AfxLeKGhTxcPYDvbxBsTZ
cN6lB1UFsJ6xibSiw2dF+iqaiB5evxUXwpR6fkktoG3L6q9yT85IxDlQRPRg6NhtsvbmU6GScdE8
urlAYNx2elhiFQnydgcuBAAw96i/fatu/bRrqU5qAXdoKuzXzqh9N3/EgUx4d1Z4Mf620OMK5lbJ
tgJ0mInf82Lw77e1uAatpfIvGgtchfO3dHWTAKsQwSigojA/hV0Vs3Fr5KdTN34G6cJGcOqvChUf
R4HV5beZz1lJGKUiI0fJm3gpJk9XRpH/qcSWaOScx1g404rlwn1d76aQMlZb6qAlL2BO4VdHSmww
TxD5I+yPkkUDu6Ps+nuNDt1XxdniQ4txs0yPET6ivUT0IGRCdSlOWHS9vyuGUWl5dg0vmlMnOhNI
Tb/ZHSdjYew+4XzrrI2vWpb0Sisv/cS0ID04YwhALoioSWl50z5auj4uDvFOO0JI6yI/6J5fvBGs
6FmFs8wsRJeTfXeKHJsMppS49qMf6D6Tk8YIV2Uh9ymgqhreLOhKBZ508fnUR6/yNZ1kaeMv8Bfv
q1IaHo2wHlziBioMQhz3L2BlDHg0AbVaefercKaCz/7aWqnkOGhqa7xaDYAANf8mt37c6aE4pdvi
vsUdB1ItwIl5vnSxgijRcnxQrtLnOVe3fjtqiCVlFVKEE/mPVdEzA9XXkTHaTxsE/0o4GERHtbBS
PX6ExUr+nr/x3u4SAAQhR9CZBEveSM/HkpYcY1tAtBx1BQi5yICD5kYtGvcWzHITVcfsfJRV0wh4
21FvUezTljBaRH4gukP8Etf6iK4mDE9ygX0aCmxYZ1QKKYVTdwMNO9PfoWjNflp3HZBmvlZph51l
8ZaHot6+VEP43UZAGankQV9Ao2KupwYFZEdLoHmUpRyYgLCvVx6rDaKNbSaPq4gl3pR7346Yew6n
iUcwVYSwcaI1zej3jTlZsPhIeKfl4s5srsGNeK1V7J1e1C8sUP43mgvmrRhAOmbTjm5Ul/d5lcop
Uj5hfqFnzKxBNS0DID1EOVbntbS9emDO6F30MZUHZ27gS8nHbiH3+KHoEH8x8Vkkm5xYvjHNzTm2
d+eTj/35F8ri3BX8LQQx88UDcxSDRfEaHgvcA5kxa21tE6J4sLTMExNEHvYD81SRvuDAlew7ggno
dKcHJBEx+mby5NzBLkAYppBw51X0zX0bkFS9b4ALrmdnWbpOjqXDzc7z9t4YI4S4iuGFd2x3H7P7
nejA5T/sPMqQW7Mqo+JmSJdh4Od2rvkFR+6nmFpZNSH58H71Bd4GpiATDo/Al9y5WjE8YnJ+GmOn
fZZKbglv0M1BoUfRpml2e5SK9yvtRFLItyTZ/nOhDBCQCWDYDaBVOK6k389Pkkj0RzEJGn/mfzpN
tq2WLMdkJWIQhhnjROJFW2fly9C5NzFDQYtcGMHPUtG/Mk3tbo8yX0zVo5+JM+2KhTESGpO5j7kT
Ug5N7pUczCW9eBO4FdpNvKsTPn8+VzRDGwsX6w0ozba5NXyZmqlk73rdx8ptd20jWwtERdNoPk07
FA0trntDgNosOtS1rX0gYSDwqFmI/VtqI+bktw6atDihPBJ24pl+puFkGgYqRXmUt4OlPUt5bJ+K
FpLYhN3EhF3E4Y3d5gdbseG2Tyh9KLx1wPR6J2L+2MDwGDii2YwzuPJji65EEuYJNqllA2P5xEqd
iAR0Nqv4dixv7lFftqNaGYL0u+pjprMbTSImEJIrN8ngAdEHGfogUvLJrmXbS9OYWZUlTKe9nKIz
CUUXVAWK4Zmy1jgwavZ0u0q9IvLyeU6c3HyHTXmoDsZIOFd2ThEL0K8Pw3T6aCBVIU4LW0jy69qd
nWT4ANmBSCFK1Fx80VfTVE9dljm6525E3N0ENpvllCiMmH8ur05pOFv0TjAl97/RLJvfiiLpeYp5
Q74xZgaDVTVNsXbeDMc72ZwxaTqE8342D9BF58hd0MocK0WNaGfyEIxwKveZ2hheUVASbZYllF6T
a+xpuqIL5Sl6O//9V7ltQZIMAYrMf0WYvWGZOb03YeOGwtF3qnEepmG5HpUN70JgknIFXKxBIgIH
6+ODuzhyuzr/4vTBfOYfnUcbw6V9q480fy5YUoZgni2eVpZNItDHQYEx0qVVEx1D9Xsr1P3ie8Tn
TJbtiaLVHap3CYfoB7DOu9UKimfbRIIRdfRWaFwZHIhfRRCTfCTAwxkqApGrJxPh3557++wA2Q+i
K9PrJoFtYbHstR1q8nKEhaO4LLFj2x0GfNdoaUfPzbAvKHGrMuPpo2qpFwrXvYZ8s6E29z6176W7
bG6+wIYh5OPZfnqLyq86Gzxh79jHZ24At2+mIEhwkSzwoVqRpQd+lBmFRphn2tcidqhm7pZULrwZ
P6gOZwSKz6bDxQbyHMr4ai7KEqxWcNOy9rqn+9m6q3Wa/EaTICEik34B65K4ZZsV58YRkKRNfhHQ
CcmtnLrkIqZab0nyZwbyU9r9Ir0gQZCz8uFJ8TQQg0/9wbXBegz/WIMFm15giSx4I7tRXLe7lRF4
mbty2DeZ9A8fnvqF1YGuQMaAY03D43cGa3mUXnNpOhtJtejPki7E1V2ekiPRjodc7e+1836mL4jZ
QBm35XhH6ijPrw35AYbJzAXvi9cP3PSyuFdx+2OGUvqpP+O1bYbVlHlTJ3RHGcSb3lsqrHDtX1ba
0kb6ET1XIHzWDmwkPybzcB7jBEDBJ9br+3BD7BgL0f2e3cDCivdyOEOG+7IHRei/ZKAKW0MK0yya
FHAKO1W+5Ae3KuZHRy0mROBROu6LXhJac7v4TKWJBu5rKaOBrpK8o2RV80F7Pb/Y/61GSL1OBGfi
5UBtL3vFh5F8q2ECOWAs3ebc8VMv9cJz4rGBi6KyYxGvfncAAJfVkBSKrdQ/Utfq3vLRGV08h8UV
5som37vhlxF5kak2nRTvqgxQxA5Kk05o8B64YqXMybK+gkFCn9Y1HkA/NL64FwxN23TXpx0OeBYR
5Z9rslBJm6GvN/5dbfeRpMSuYJvm2anp9sSd4qXNCqA/7KJMBiJT1jc/Z9WBaiJyTNKrGm5s0o5j
vJZGhjEH8CCcDwuSHWmXscflTFeMoybSPqqvMyJedwqRA1bQSL95TUt0EtgRG2OW2XJE5tEjNK+G
6VrMZ+EKJ3uNqvZqScoxyQBksFr50eBoJDb1v4yRWZ5WT76itNHrPP/GvT4diTKT4HfzcDe3U/g9
hl6et3+0GdKWjnZnTwEl2mS4l2acar5iNI8qxRWNGI+0RRHo0E9DmJcnLHd9EgW8hqHYe1waaPEH
HfjJT807N8zLFac9eQ2FBN1DliZKlS/fUdwx5LIAtIuuRhKzsKxNQ+1aaHYScD1re4TJou6xsA/H
5TT7q10sNliHkL2a0LuYf6YT03DDVRRRIyrNJY6iRSj700WH6eUp9B4VYFAf0/i/3o9JS8ZXrD+Y
cyXckN95aGwvUOimGI/hLa1FfE9WLPq+z/STOtVdHFyggqkT7adrzPLij/yf6BQgclSBQaBq7wFz
cHFd32Uad3cqArSjrH+Uh3U9Mx4XIx72+VaUpgv2AEPdCdc77DN8shAEkxxLOQCjIv1sD4dgGBwe
qVyz9Re9L5KZZHJVdaIEhgnN7RIRXRN4BCVS1KUFWt7UH05KGmpzRMbWEyVgbJFRkmQedPZa+l8O
ilThO+PQ8JOjHBRgf91k/W3khw9L1wATt6kGcsIWzDsWq3qoFZKCtXMD+SByXxvCIaBk4Ml3qe9B
5GIyZh6DeKjI8nPXmfE8blh0HbJ5H5DX6maHzZyYxygjxiiEaROlSPa0C1Jr5+9VqMBHsa9mRbqP
NR8sA3EG3KAFCukc1psCnutopf/LMEY/aCp4u6la0qvlyhcVjfoKyO2ZByV+SQGwbbZLHK61Dxcg
sN9gj31CVGHvN1BunI+9GYqYHo8TqKFj3ktNbsHfvo2Dx1pwhCB2f4ZmgvugcvJ+UzCCp2yNcDEb
x0s5PVIPXeXKh9BGIEspmQabFN3biqYABxSKIJondxBScmWWrxhDEvRkrnmyzOiMw8VXnQQvt/kg
mupATOoRW4rZ6kcm3eRSm38PYzfQi9HbbVC43A/Eoot5rw5H9AvpCRT9Gh23PVoPuTcPQx+SCAFa
ux3coJS2PZqs8LMemuQWl5OX1tGwLEmIhykA+IoTpWrr4obZEH8rbRAs2VxWIjY8NAkfJoVSTh7S
m+7a4kJKG1893UqHJgWh4gEf3Slv826vQeUGjNLL0UWS0HYMg9G0LukhVQWCJbXBkV8ODiVJGPZQ
jURWMEXnhaOAyWTlA1+P3th4nwo+puPcmYJ8ygrdhhgYoNO1QSzukLgjiZj/1wu9aCb9qNI89RUt
1Ycoe+eeek2Sn1h0Fn4/dGG6OBoAsNfDbpKzT3c3QDTxr8xdqh/9AUQ9gPmzFYgcMws/vVWrBgpu
RS/skgct14fJkOy7OJj6gEktHsTUX0yLnJDPHzJ9adxwL50fF5cgC8YVVo4oTz5YxQZUaRjEoGOs
g2/rWesVIzpFJPrvxU+dFccd3Yy6LSVwM83xYSh2yjv4+cgt7lHAJZovSPYTaXpLO5R3S9tEFWJd
s3kNTtQVzFt9MgIxQmjxJxx8Q6D9DpL8EIGidRFoiE2GruPRkyIaRu14U5bwCEct0YEMz+hTI5z0
WnvEV45xjQ3OcGhKhyj3U+nJn/i6jrnH53IrH8jh+u2LKAt6cRAOGmeAW8rAoRLpUsRxPp4PCqMO
7K+DBpS9hiKjFt9av3f4eNufn5A/cxUigkjyaAiXZADxjf/NPxgb6574AclyTIAv4vgQqEGL7XDf
THA68va9XR4MXouVco+v9hJN/T/KOvFNA9Wnu0XCV6Doc60PMAJClk3rJ1MG78Eiyh3W2Btuipqk
v8PdPpbuS0Lz6sF7W2a7k7sQ5hbNF7W4ZJHHDJAZZah+zcOOpBChHERx6TJBIpY+QHbE1DSqojNo
UypHopO5GH76Ht5bOEp6qOtvFFD2EQgcFnf0MwUZ9wuoGZpkZNU4BU8KXQXij5XPbtHOrfq7lci/
PnddnxqcHeWsnC8dgxVXO4QLKgObt8F9fhxG5w61/d2uHiAylpJTxKuPl6CP3vKus9u8GMjxJgAU
UEwYb3XKIfyDlw9d2+b13aGjjIClcNqDoF1v6BJthb8K6qlDUBMgmdDcCOBcGL5uv4Et5RuqB1c1
0LeP6aeeWmQ8BNeQtHKsaPysxbI0m2TRivNthn3n8fcAE/KbXPtlb+etT+GNBJaih5MhuPSDdaJ4
MAONlrt3av+c71nKI9cMwDSJjSH81fh6SSxrPOwqgind1oKocn+1w0UnMxz87kVX0yt1Jl9kRL8r
x7LYpoGJBkqAuv+qw3ZHQbEHywiR70TLcCFu+aoJdSSsIZr3/zQPbiKhK2JaPhVmHyOjjDWtGKX4
eks/c8zUlbnfCeUUJuxjPuTgLmphTFpAPQUQ52PspISDcg8+9dR0t5rLe8L/ayuF77AKvJePlteW
srKf1rtJTjmvaLSFpQlWVgIJMLd6JXHlEXX4rSwONDh47aetD+jKvu9hFOvhSLGstoDZ6UYCOwWA
JDR4OdUTxjpJtM8i8Kz4uy3Wmib8GI0/vQfBZJs7k8fNg21F59A+rP8tw+doHTEDR3wS8B5peERS
MBfte3hUrvKxzeDU1yeWafCBYEB6LQ7Tsed4FT7pfAuAsmqZaLu59RMp2Lxmvu3ry6Gvfu7vXNJF
0icSPOeQEJRKQc9IU2yFZUjfLT1ZLpiKTShF2sZPocfDJUOzIqe9+JCcC4AEx3mEAqoRFJ+QTk8V
TJ3k0jAQrSWMk/+CyId9Q3UNIIYm8rHDhaFmOfj4mgEgOo8ItSTVbO9L+AI1VROfdS22QLEIQANR
obBcQNgM5zdpSbVagbSm70y7g+ZQ4K1JTxQve9QSy+R2dM0VM9Vj6KH5n/9ZdO9lXbJzfKiqYkWC
XwpM0xbBB6uwRf2WkIoT8DYKOHp+Q7skGRdxO08kR24AH5ckZTH13U0u8RhQYVKz7VEDUf1Rtt2e
KeVHDZIyyTRTU7F/r1KwqwuQJElYBkhIVBZF2mFPEyMJO4x6w6Oaequu5qXao/SfyVyRSbir5owW
Lgy9uK8asnouSQf9Ld8wGfPnvnl5mjeDIZ1uqwIMBHBcH0rLlrd1Wp940JhTcUVLHUmXyzP83P98
3PHhJmfmykaZLTyv4iwBrQb4NRjbwSL7Gv5630Pyu2RVmWiAueZGqy1RY6hLC6Xqyv3vouXJwgL+
DsDF56vq9U8PvSkZGdI16WNnGDJmaQEytgwvkQCfFh8RR/EBVMZXj9oaYZD6K16WWIvEweWE4ZsD
AHpxo7yikk7y3z8AFhXZnfWzciVi8RVkZML/5xUzlQMHoMbKkBgWJPARYYxbkuvnXV4po5JSQ3wC
DjNeqcoXNIig7wWPkq80qBx6CZMkj3tyFKyk+3fOsk2TRwPyHY/3yMc7Uxg9AYiPpoLNECl2Jtn3
CD0xtizRLZxC6omVVv3Dem6FpFDdSL5FDmsrqqfYaeAKod+4QgYUFBS7K4khX+5bygdIM/gjAE/0
0i6Q2X5MplXnD0Ucez5iF7HPhwJPNMRLgnfOJ1tUwkAxgrBWUqK6iUs5v4Wwlwe+kwaG8VrGoUBO
XMr2hTMd284GKUB0IBhGdCpRCT8qdfprHbIgmjXPg/cckfBhz2RfVaxKHOd6+TPgNlmc024yRl/X
TmpgAkgExgpXtJgjF0DmPaHmgt6AG/yMEsFYQSHSddfqQb/Yq5QgyaZXNnFBnfDMxyP9rcRnnKDY
KGH+wSNKJiyhkGhlDi5o7ANcG3neccqAPbyerBUqMV8hHFYW/gscpM0o8Q8IzUIMcBJ7waKG4qL2
hZgbIEUd8I76Pqw1qBtY0C5o9Gf7WjHFFZmE+BxinP760PlGMniF3Z2oViCL23RqdfOMGssvuVPy
2BpJQTyQ5CmPmlcBtv1zDNoO8ducyrv8VzfYJphFOKDXivJ8yoX8CGM6lDSbIlSc5JxlDcNqfQtN
DAlQ0Uhb1cRtsM8uozz3V5gCbYdZQv16Vb2d8E612GZA4/l8YlbyXgKqVoyk3vtv+7bZEbdOG7T8
RaPFdzgHbH2nWtSy/B/oisurswM8jGyzsQ+YW/oFTcJ/pJn15laHxMnfl0nhDR4gSJ8yx0Yx0BfS
fT05Rwlc/sPnobFwz0OsmMrhOcUCEVfQf2EvZHD7fnXRHhGbGATBVhHeOCMyVxPpzZd0vUwyMs82
BAsVogehwByovRJ/XoLpUNo3/+7+DI95xdX12t0hKDLwrjtw4QxOS91xTZ3nPaWQU0pTGlnIIhYl
0PCrZu9sQu7jkGUoUbCNRwFS5o4gTmaRI89hqmn7rSHxf0gP8ID7U6t5NRyCH5GOmkI119WvFsW6
3VlbgpN8lASvU5GBSOM8VaD8fWdYtEzm029CcGhyFTCDKuthknzo1qTR2VIiSswIFFpl2Vtu9alg
/4JGN4jHNieHm5y+Ubf/hxtmlzi6r7Ij0V6K7//DviMziPM40IF4ozKsdsiCHRFePKs9apAiKHqO
Iv+UQ9MPPyAJoBPETkIabu7RajO4kh64HYfTG5VFwXYCMGK+OOcoeNeSw1Y4q9ltxd7jVph45ku4
ThMZk/TQJAZak7CIqWo9tkj3ano3KuUEEfTSQ3qjdJZ8QOwGfzk2VUKgDfNkzPkSq849bZvv047s
KZJpJ5mJT27mobuUlhMeHBNTWYIzIwia8q6TJKexCoDQiLvx/MgHBvKB8aVUhqRejjYhkZmv9dNR
kkcPwr+MkZr4BgrkjrZhTmzpfKE6KOXCIR5p54vowhPcsrhuq80Mtfsz/+aRM0oPjKU9OEMcPvk6
GwJtNmulxTVxcoeC2YRV3kz4BSKsDb6O6JfcO4Bw2OKdwru3skEaHTHh6m07j2RyezoqIXUY3Mfx
s4ItSJuVHYlIFEGdI7ErhxhX4exVMB8ybpmL1zZ0dU0zudwUGwFqqJWYA4wsspQ307a97StHBdoX
UWt7/DpCSpSVbv2LMzK7ohTwacWxBiY4pWcAmQftDKytfg/d3bjtE6Xc2B0xFWS4HYp78Bwa9Qsv
BP94t7FJ8pSVnZazdGw8ffWWZj+UQge5dzLQimtZPiC/lzf17LNn/t6+mRuosfJ10N2QOFzr7tM4
HppqqzJUHz5SDFJkOhKonpCDtLhj1BX8gFFa6ahNNSIy+RfroawLi3jKi8JAsEp//dHQbYkl7OyY
1Lzh74qeFrD+vCwqV2JsRqV7dCPKD4pPwmBE4E26zvLLV1YwzTZUmt7L+hkWqYdVZfrIDnOku3mU
x9RWinw6FChmXXJP5cENCYb9r11Dq35Hb7gE59xrk7tQhMRbBv89UaUgUIGYWLuZouDlYE1zixZL
TQOTDjpm0B9C2YAZf4lAdYeuiARaYjoIpJu73p52n+VonCB4Gn2kmR/DMKBmBm2fMAeizaJ7hfr3
FgaZiCn+ZDEFql8jACTt19vvQaQW7/t98NFLdv+TgNvYHWz8QZisBcs/3A9DJXf2PWRPm67GpUNd
IhzwYSL1/BENZGb+ZwDVm2fl7ExwFPxDZxpqmJ+yWUqCZL1K3QQPXou1buXEhRa6jSuD/+I+A+gm
QEKmXGB2cxuwBTw98o/msJMYZDi3eovSfy1pW4j/DvCaZ2WGU9rVKKuiCZQ6MI/1tR/KRp1t3H3J
neE5n4J/EsmC4FlHo+BH/hqpU8u9oylCQpWxgbdhz+fcv+9JzQ73FzAkQx7Qz9mg/RPBeiQjgTpV
KXJIHPgTJofpi3NGzml0taLtlXjpUBRwqdVEjPbLFsHOuc72+PRIWQxAzHBcTWQgIZpNq+Kq1dpQ
8IzFAMPdEeKjAKT44U1fV7v1oHzllospxwIzXUZZYk9x0BLiCglV5uCOiZeuSi6OTA2qc6A1G5ww
kcvyPbLNpzWaIBCXLEJkLCgsHvU3BBifuYbevPyO3/OHC152vWG/QyrL6BpKRJtkcMbg0PXEnzAr
tORikZMQN1/HIEiiADfeoPBT5Fk2vXkkfMh7sSte7wVthuSph0wh3ho4662mw3oomu6m/xfXw6dV
c8pBPO7erS+Dj87tNHrUgbw0GVqCsOoapApHGPzwJwJdwoSFQs9FTgdzf49PkOvllhcIu+OsOSxg
bsaLeDGwqWe8TkD0WQMFRsYe9GdkCHU4kNpgSVxpQ5mEx1FWlnu4GzyjnV1QBBa1pDdldDGlB3kM
aC6awpjCkMm9lHR6htIztXMSYNH7kNn/YDMIhzuiLTbqffIEG3cwWD1O/X1IG3bI9/qawG6PjtWE
jZRXvVv2uCgu85ebt8IWaxQzpnPNC72Pshhcq0uqPcx957D7tm346lBhuN1gziyR5xynlMEZ4+bt
nhPdhUeGCEK8JwjWiEH4Rt5ypd3iExNgpoQaHdv3HuQM2dnGTnykJ91ZPjzAZp0AbDWQpdh290xi
S0A3s6G+ZeQW9kbV78Bec4LIVaCKu84rlLJX7+t3jZjB82Qf9tMukZcXKKEdx8CkTvDAa+VisgKU
YREIdKoHLB5WXdsdPfTmx6jbL7By5P/iSBNVSedIv1V3a5LXdnqPsPpw7U3WjQvTNn53OPFko3qc
W9ZjwZdAoxGSYqxT10Cwx/SN1+cIfu+xv1JVVc9e76sOXuDBD8BK3u23TkIPM+mo7fx48uwJRTiu
LCstUmaN9+Wdy4tWs1LmXBWdZ7GhxOnwkdDCTAmQim6UGaL77dapfDevjkXVrwvibp7iRhYpoV42
/14dpzVplrUexGSCsH0dGEOQFg/yOMMejIq1gPJiGN1W73vWkfJ5w9BJNgnQykybG2Z6wcg3VeH0
YR79P4xy8tJcVoThidQqJrhN17FYFKkRcZGfjtlmV2mN6JIECxFVj2WCov3yLvgQiLtOhGXrmDHl
/2rJqHPJHWDQwg6B7pd1X+i/22m9ow2ofepaeAk3ionzwwar2MW70+Zm5lx18qB8dAkFtC04RN9G
sHSAtivvxfIxVJZYoqkjH9Zi9ANC9YFGslnbpY5qJRBsChqoQtF9fsORKD5XcLYrM839fSEWcVsI
+hgNY+jciQAHSCBBaci/RtjZRJjhPOkZ5ciuGZCRqYA8tfuuh+0zZlk41++ExkHc12aTfKPOFZwz
oiFenrAbxieZDZa6GJVnXXWpLo8CCoIPmBDf0oXl2d++CfRt1Tkh2yrOCjDK+qeY713NES98BZjv
FKggXEQVqCGw4alEby3TqLrgjcf34jw3pCucMpQkoXTmMNBp9mMFAWeTaoEHptXFfZQZw2okFsVV
gxqChYlofHWaaUO2YWotPsT7ohCoMqoFGK+SK04iIfo2VQlHZg7BEw2+IHVwP1BIJl5RiAPLR2So
Vyzpr98HlSA533K9XQOP5O8asoPEQK01rz8ad6LjuFd082+AUF4vsBeaUZohGuWlisGOb1cLUtjP
RfcKmR/lgozkd/+6LnSwGxitQuOnzv0O9GfizvViuCN8MSzVSJG2QWROz4zKMCE+gjDTXAE+lzKP
/RxjxkgS1BpmlVFWlv1QZQwQFdCz/XFvOVRhJMVOeBYFuFNYg57A0Oo546jWADTPtWNhJ/ltKzFb
EtokEkWpQDQy/KbXhMGAKzC0U8BZ/yUD4BDg1tefzrLifv5ntUen+d2ruBiyGfImQaTp8C0vXqkt
KaJ+Irp0dNWBsvzxVUb7XJLRiUJqNi0MNV+GDoBOaaSjU9qp5qscFypznU+Exzz2+/cIgi3gUymV
n19ZbIN5dxa74SLK0FtitR3eejBg9lyLxo+fjahMhskIuVbl6N2yBQDidtbFwVXC3Ck+6hQvsrXX
9ia+PGgqlmaeRZwni8N8ofBFRJEbxUGn1w7SX8fX3kafCESMaRAbFjU+TRCPBwCbWNGqING2eaS0
++sS1MHqVTL5PBxl2R6Zub2m4lAuEYWvL7miqyvaxpYALGRp0DW1aB2kVRC2YIuR+k+r7nUCVWNb
ABPG7INr1DPnAIjLACyebWV07NYvHd2aZpk6Q7nNSBS/SGM6xTRRgRpC+Bx1dC751RD5/7QtFEPZ
VdgRwrtedMNgjdZGP5s9MoJDXOvFTYqfg3J8MP0v+DPEskgtr3vjAU1Q2KK6zXWa7QRqlpgkGFgJ
CriGBi4PL10dp1XQF2o/Qj1zJuk/8w4BCc9Jl3Xpunj7vDu53FNkRec4YV2L0ru+GDwo3NBouDak
Dp+xLEnU3NZAmmAI2IhYd+YPJCoqB7cti223h7ne98lQPuZ6KEK5j/9GeX+yyIKVXcLAUhz6744+
QBVNwdBpbHq5a8TQ9F3NF79ef+vGBL9iihqUQgJHNZOfZXYJ1Q/KfewnMZuY0i28idTBWGbHd2b/
oIEJ0XOKSEmSqX/L6ALmzfH9IAfMQjpmxI8FIXYr2tOmPOaXpyNFnjoRXxC8sgZqs0W6v33mb09N
a5jWJpIWeBAaPJ8N2EqTFnFMjlRhO/ye5dlVLSB3AOWE252BZBksoMN/V6WIofdqNatoYSu8Ek6+
tnYfDXSvgKq7HOY2vdgulDf08Wt6Q7NfY4tVTRTw+DaSTk7IrwYOni8PS1fkEfGr8d+9lTtsnNJJ
0GnU2LgMPXLAGIlzXci91c4+k7fpRbeYu7mrRD5IPfFn0tJYutqqbeYGK53ka9wKpaQHnmL2xvY2
IRjpKNRMkyPLT0zxP03V/GFYjJtgk31i0hc/9M8ZkGeUDmkEmbbZiRANRnPL4EUOfnoliBmgtQac
bAHxUSESlDeNZGLOp8P0jpHjYpR+5Yb7tOCAlOt8r+NLQGUNFHhRLRe39D2bQwbNv8OQl0Q9Fafo
0FiaIgs5158u7CgXhNYBQPoYTwBypAhcvxdTOE2dgZ0X0CTyyl8HHas9HN8JdAlXWOJpLXSWYsaX
qzb+O0nYEVa4miU0B8vK89lWmdxSLLuvAPDZQFtCm8gifhWbV18KtW4sog0PJ4KagmXAH2x6COpV
T1B7jx1srNB6JTCaXmStw9p6GHckk0LdWI9pvJ22D76Y0zgrYzqKiJBlffnMBvtmYfJ54QD4zavZ
DXXsshJGygBieX0V0Zy2MMylt1DexgLQfPUZRalEJOkaxCufYvxmaGMSu9WNG1IP+IoTYuWyQMYe
bLrk3Wvylr0poIXPL589e4BgTlRRXSiGXIOSG3f/V2Ng16MbNgJS35QakDxWGEF2wROUImuyuoY9
i7hkwckbb1RcgkbTt2U7zHNkyAR5DyyFl0kIeQx4go7rmOtSLCVnS123jFXZuPFH/ZZrLPaKu02q
7fD2yGRwAlXQpO8Xi11vSkMuovP6iL8SpNHRFjHA5jVujEyW1Z0XaqPpJxdaBxEAx65EruW5igoy
DCvbuuAV9Er8J6oaxcZ7yhB7+JczxPzNRctng3A2VLRyOzoR/YZp1OeDJUL1Nzu7QFCdYefzxaFI
57/d+z1xwngPng4PV0MHxtvru6tC6qL+zGqsJPqLiRSms0Im2cOj9iOC2D1ZQ697D6BURmf2s9Lo
DrYtgvzQuR6z/lSmBhhj2J7ionzgWe/MVTufMNit0Y/vKgAgO1v+ExHye6LGgVTB7LvaBZNYxFab
cX2nvAEsmsSFhhA27JXYjt9XpDvhslH99RZ08ZQB0OJqJKm3j56+/FRwgXBKq6qHg1dEDCL8oWkN
YWf1JJhy9pdQxCMNv+ED55IhxE7s3PR55ieucSC+LRJt7Vad/Tcw324slLWSFm0gce4ca5ejwf8U
YJWMiJraEKm97W1m9ki1jyAXc22V+PDJyx+hOfQfPWIv+BVsKY3ryGffTB36QISw18FUFyqJ4vsV
j8/zswuNc11V0HzKt+cWKP3OIgZVp+3mM52UU180WLcWx+OWJ9kC8pOsJcRwEWwhijcnv25QV9Sd
muY57CCKvbLFXEhhe0//lDJYEp48fVhUw73WOM896dPgFwiLhOCf+TQJa8/4kqETszD65gVrWKjv
pRm/d/RSYZ5C78hmRRlhsfpXX/id05n2/eFxc5b+ul1zUAsaITsQEmgltqN22mzUwFpY9421eKBD
RBy+FXNR9/4m1q0UJqybsMN/eq5ryRdCOxew5zownYfJ6Vu5uEDhj5/xa8XYYBAKPwsZLS2Ew7p3
d2m26fd+rcKzyhe+X1/wqwN885uoQJOtveczlT3g4DlKaLHoHSH9QWc722Hd26Iyz3kfKC59bBxL
QZi5NE1sxZh0Q54SguGm/daohoj1nltTrZMFvc/mP2kPCB/QYbyuDvejoAIAAXtoXBK3SmyVm3Z2
GYmgmTqaJ5+oMt+4kf787R9tWs1m4M0yipTvNHG1sVfiHCcmGrIp3BxDfhFCMU33/1F7oN3UXGSC
Y8hCro6+TwpT82Pwzi11z0poB2G69a+NNihZ1YWY32TOVQYILm4hW1EnEspKyro1matliHXPogus
vTv6j/yCIDfz1/cD7TENmT7wyj0BA/4Dj8g/IrosI+IKysVONFmT3mWtAq/kRFoRY20NKE3vjDkV
DnU+L0T2Ll0sI6axp+AY8L4LaQdIGnPZb0GQfqt+hd/HyWHW8sJakbcunq6gXM1HzwuRj1kndqs9
qMwkrH+D6w5YV4clNnm/KQQFL6Uf85qIoQj+qS81Kz99xX++RHondn68/Bzxh51Mws40Sk3hQzJz
ya/+7S1ENVUjXOmR9UVK7gN4fkm/eCnQsh+Vgz2NXMDVv/sbR7FAEhD1jtS3OQK0M92Fu25swThL
iTmGAnc0UAF7L7H87K2hDxu3L90KwxXvpHYXHDqldtCaT+EcP29nHFCQuM09IGuXcMHIN0bGlRTj
14V1ENRosrqFj2uIPXLVAxDPilvauBOgcOD171a4CzjBXrwZWszC3sPGLYzsrFVUCEtcELd7BSQw
WkOdAfLnJhzNu39pVo6eZA9VqH3ZQXW6lxzDCUcaMq5aijEeOfDj5b6LcKSDFhVofka+u8jgLxF8
SOAwlIHS4BOF0TDm4jK+xgTCB8OorgQXvsodJNQI+QDyvy+goKDk2jjzfsfNKl5LhDu7dt+zuex/
UL0hs5SRprWe+LjaDQLAc0+7UPahVdMnfQwWPEMfv1ewFElhxfSWNpNoUB/NgMORTWQi22F8akIb
qccQSchwjYY3399e3hVhUZFWGZAFDhMSTAU2bhf4A6IdC59jvINv2t/IX0hil9FrHe5rnw40B3BE
1ePPof0+uNdDZ2Umo4jejyvXTwpkgQyJwO7LODMBl99RwZ+1Zrr8L3+DqdGKcQZwIliOEoge2ppW
jdl3rWHfOfNrTwB4YToN/r1/51Nr60c0riEnupP51t7HEmxZpoYvuTlot6ghFuY+QUgYu/8e41qp
BFuCy3Xce5inciSFXx/bL9gciBNGnTDRqYifLYxoiRBr6I0lihAz3Axdp/RxVmIQUqkeBHRkMXE1
eu6FBgJ74zM2PY1HgV8fLMNMlFUax9PSaGFTpCSVyhLZYI4wVm186OgAr0rZNJV1nDoUkFkDmuCG
rmJlBBxiormT7zKn/cELB92rwsrbfy+me13cRcfLs93PIQS1lH+G2lwxgj2xl6WE3Qy16DQRpo9u
mmHJGfwOBw5HcTq1dQCPoeH/1hF9RpKvy23gp4ryG83WGygfAZTXbjVbtgku2U8F7L8lbAmFo63K
PRKWZduubYr8Ibw+MU197nnTQ0Yk5VKVkm+3KiVkovlrKmfbnF77CNQ10V+on3sRkkp4LkYHYV7+
urTSXi+eN8eVm+56A7t3gtOEzPgQU4HWSX0OjAkhJDiioeSva2E4p2HoXW3ZZvRMrQOiNzdQNiiB
8IODpKmmPnW8tyUoNOP6/2iZM5FeeRhmIdLKKuMvK6dlNtMMWsO1rmC1jyhXafxNgEw26OZSQUdC
MKqoLGVLmyldKYEf4++OwiNLesZm22TgBRDiEUrkNBL8AGCmshsoXKou1Di++xqrXDDB+/4D7q3t
nJbI844988BcUp2HurBOHsdOtHjKROe/eR0arZZTuNdIhIGgCvAYu8acndF5j4/UEIgv6VdVgupA
bjxJMtalzAPAoeUEAs3Fd48DBlW8yT3lNwkJp8RJKs6W+grRDwOHMAAa45XLLqeTY3F9cSyZfOIt
WAbHFKWKJpeNF/dx8W8YvucBbekvYO6sXrAJ4NNVYInOUKL3lj1jab3lxoN7CKvWyy4oScK5F7ya
V9R9+D6vYO0FsBL7Z2X75JTzqD2MtmVlHIvo3slDwtt++QCaFEPIyan8zTFMTowx8D8chRbP3mnc
sO4VKK426IPDvvlwiw+LcT5E4Coi4oMGB+DQSGz+kl9z8Qg7dhQCILJ5aooIU3LVaiA0MGh3vhn4
Pq5qNmZe+ChwYXZv8n+HDA/SxphRW1cmR0sh6MnjtAcwn7pClzP81DxJ2PQVs7IEa6JXS0D7a8iV
AoBYy1oOTbTw1vdPPdUapn5iPNSHsG33sRnzDUsHRUz2H9bZjFf5anZRSVNbW5fyR3MYKsoSU/sf
NF5PhmAeiCwgi9R6BLYhB6X5twUvDOJQQ+ej/imo613z2UP8+xX/iPzWOMCyx6t6YM1eLS1uBFeg
VTTM03FqVrY6n9fPd8CjZW9t/WAa8JjtuBlYzTTNQAYB0qYunySH3PYUcbDBty6d8GImHmbDaSlD
9muDJIlug5llHoGri9tbgw8M6F7c2/JqozRds/aD5SFUIxx2dkQuuKwCoRCHlgrBbxytW/YZkxMo
UPGqPL4/Mr3uD8MiArjToqfpAEYsQsp3ac3zZY6gDR8SPWBZfTFRjXGHZ7SqnjL/V4LjvzvoqJE9
nesfAWizV3BKATenhC/X5HfyoCVwrtmpa1ZtQjXzbNivG2j4S8fdIt8Phq9CI4TvS3/epaAg61S9
0NLUDBWQxl7uw3MtfKNc9xqxit7Fo98sXwDhdfWYC+QzHR7QWCMRgL0cNPODJzqnjvJF6JiLSiwX
5OmG+kDJLgstED17IMtQPZidUIzni8dUcVeLT9wgz+47cZsEBMM4mqudNlck5YmwKdRrgd3wSeea
kwfgRunKkfMPseJZtHvOpKrto1edaVtYwRPlDucL3Xp6L9LYI8hGkwxP8EJeR5HZ7r6+hz/g4x5C
pUhubYr/SrYjldWRbLlAsQl9yf+Ow0QrSjJ6Zae95oh34wcj1UH+c3BaFaj7edi6fwgQzXDVUQ7H
CCjB+mF9PSeMX647phJsqryAZf3XsZIz4iLhL6Z/KrAZhdt4L4R/SY6OeVMGOnEWh5pZ+I2hZBFs
/kau6bjNWdIkxt0ySX2s5GMyushXOKl5jHleTuVcv4MEiXyi6M1GTXhHhWgvTPytpJzxOdZzGxbO
odm62GMTOnXIQ3BSMN2wb0KPy6XQc7FTZLqJzwaVXOKdPvJ2/IB7l7ib1vDprRebqt7GFcI9T8gH
EKTdClfcBKlsOwULm2nz8oIMgS0MAqUg9ae3JITShHHm7ElDfok/859rC1uoTFmPhvxv1uxN5qHP
0GadT9Y+B1rBisYqm7PnSJEECDjJ55c/653FqU9ueS4OQu9TFc0LWBmYcyZv68lj1lOMJ4oIJPwq
StbyL50KrM/+vJspyIgj23JyV5YP0IDu8Ul9P2ZHX54DH0y/SIpjlPwxKkOKMRLIRHgOOJhSy+Rp
RvNSF7gLe0XVSSVoDFcH6ZSFpFBaWCSS2VNNFA1RbIBSrN2qvsuywm3K2+5qhQTeGjs6MWktMEcD
SL7WTOlp/g9E+7+Gi3/FbC2WAupk7t2EJfhTXmsYcWR3eJR8G2E3BiGVzGEcfjx/Ssw9O53SA4dk
jkImNvzarVA/vQH5gFlIB7lj9PljSRWkTsIBJ9WP3+JI2+GmyPLIq9P8uBr6EjtYtdY2Auny1G1p
CY/YB7s/d0muJUliXADbFsv7feuKkJdQWRX4xJfZq7OxqHK6ARumFVXRLn7JLXy9+l0zYKqaresV
BqmyK+g3nWKXmlY0CQ4vjIbtgj8cDKVz3IMXNofTxtgtXb2Y55+Sm53p0qSJJ6xm1pjjKumuxnLT
QiNb4Dn0D+CaEQ6+cdryQKaFqKAxO66Esk1guyGnA/9rezG+/KULhjvmxJbXw3zs0r8CqQl31dlk
yS0ys2xLQZwDQe/ku3sQ1wt7P8UvAqhU2YzhiT0EHtJ/uwqLmprUw2wkyALG6QkpC84Z8m0Ax0A5
CJi/PfS/xaNMU9TULgUY2z9GisiHbluUPnqj1GkqIyEs/O8aaZX6DKYfM/Zhe+Bfu0i9HvmfKHkD
WdQcbuT///TBNROF1YjL4BAx1eeEqcDB/zL3XLsBkbLyg0fPTM1F7AS3F6rcO2EEpkznMQK+qpGm
QsLqS1ASmOMR9W1Mlt7GkDDmloLCj8ur5rjONzAiPU7tk923JuBVqrUjp2lwmuoiH4Wbk7oux80K
tHr+nFsly/Uu17/GBbYSBvNHcdWZbSJ3Ey+50yv0ZiNZ8dwHEmKbkWFLaLfokerm32nmqCwXT39j
TyncbEDrd+y00f1Y/kbQBBxIzrBoJj7mdACUmL02nE0lvcw6RfQbT4iqiVoOlNmrlPe9fxxZR194
tOyI8smDFkMpb1X6+XSIxCaJBu+rQCpBEraAlN1eYR82luFWcOTUzhTFXI8uFqzDSgmSIiG1cnpy
DU4dIJOZTBfQsiqm3XJ4NV9bKcSVmKcoH7M1IPDTfumOZwGph01uFwZT78sYP8OZZOy66OKClRu+
367nmOu8vXtIyzroIEhgUKWmJZdvr38/UEARg8mDe0vkNcwyyp2Q7lyX39qOc1rjaihzvlJtQX/I
EVHbvEa/p+nVZOD2W5wdNZogUIaZZ+dXUHfMFqSuMbE1yW+GhMg0ojTTNpDSlU3sd1Yrjp+KfOnu
3q5OlYSniNIPiaJG6OgqXMfp3o+yz0kFST3sb1n5LDA7yWNwMNWn+Im7Vo1T1l3oBkQ8Y1ZtnR14
Z8qWW7ABIWkgD7FYCkXE78oxzqWY5hyCvVdFxeSx22Ky0DSvBYZ6LTQ+6/uf5+visEthsJdMFgT+
5UjbrhdnmpFmd9QRhfwwe3iB2YlUj6OlCX1W7wpoaZ6dZqqq1h8gjXyczQ1shIPReUC6Do0GNAfH
c6hN/7N53Z2r3JZQ5+h4SgJ9haiQj4fdLFZyK1oKjtYD2gEMo7S7OVJTaj89853FNujFhQ+xnH8z
K+sicriWtCuFEOWxpWyyVkLfkNDkFYMoz0kqPnVQ274+KJhW01VmNKuFOETH/a+p9dJaZDPRQ4RQ
MIThIusMcob+HRhTCgMYmXu3f25ycILJXB+AgWB+ScqaPVh07PaoYsK54fCjLqY0GNjYDZAuptQs
N0BkBHFQxHH7/hHAM+vtu9vEztM91rzaim4uDahU9swy4laurr4LDqMOCVH04FSR0SGS5/qyTuJO
vNS77K0pEqolu1UOOBkIzgN19yZCDAUEst55YDV1TUKnpkvgQtA3pBhG49vqrwOa5Aw1Ude/GGs6
tnydjdkQbQo+fMJnJY0+vw==
`protect end_protected
