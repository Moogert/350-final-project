-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CDxMXndO2yRVxw25233fCWksK+VCrMuubKKin7dX+axe7JG+nZzAHu1QtJbyS/T4d3BKOip9mTCv
yINMvA6ejEZ82lvO3PRz/jy3MlKDM2W86E0wYg32HdI8xmD/MoU9s2K/zNGUdVRI3vo2IUhAYIbK
gDfBFJQY/CBx0U7SVuup797cMMIafC/9b7ZWZ80KIktWxnNkPQVBmEPGpCsq3xIfPSU9MNt3tfzn
19B9glYka6OHzTiZrINd17dq/fwkYb5BOzGuVuUXKFPrTnE657syDbOSU7zXVGwiP/YCrxoVRZc8
hibNfgPAKRHcCx+ResytHJLZEmsAZW78fhjrRQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8368)
`protect data_block
EIFH8kbGc1opoMPNKoe5dKXDyNKMEeO7yX2dWT4802PFzOiugRStNqnBQHrt6mzhL7YscX7VyGdU
/PtG34hVHKkC5BIb1DeQ0jSPw9Z8DR5dCxrrr17PBHcppdVIk+t1O7134g0kC9LAz1PbVQqHKdYT
viHoisWobb0wgPE5bRkV0zJnJdGlu/uMOqesrnA65V4U/L1d0f81qvegTcU7IbfFJyUEakA3LlUd
KE8+jy9m01gaLzNJQLKQGu9/3xcMWLB7U9xml8sjFFjA52ShVDOr1VPuECtdgDIyqU9Ke8kq2fcF
NRJQaX8I47vXMtOUjTkhfbferK97WaBUol5Rwo4ocZyodDxLimdmFDibOLDTwsIrHOU2ap0PPAKT
d6MnJKq2ibJAhInCmISEf3ObhNjN9gFKp7yoMrBSDzl8sf7T4c3RfZ94vVZRK2rhTSGNtyZ3dtwj
VUow0SxuCDItN9/mWR52ldYBiPifJrhDd8+BI46Ae7Z9OLSYXwE0AWKrOWowV18jSpmoP/6c/4QF
Zo/YHm9dF5gksF1VWBhHj6sA+hMQUMx/tXUiVCkDpyr9HHgqe+UHLxWoQ4FVFJ+qIXQTegRVopUk
2xaLMao6PjMTKvH0iHgHCsEL0PjerD4vbXqmpotxWhwm6krSDi2cEqYBMm90zZSTHzCUxOT94uIm
sV7c3MQxeZvNzBDrGhgJ9R3A/Fhp30ahydfsqUyo0aW7EeYJZNHM6mkvJHywH8RCaFKVU25616D3
M0+6u4cd34qHOymNf3Xpl8yjY5mkfJ+c/f/rmYjHyLS0CSU1NFZwNLyhfsIWFWDxPn5XzMdFrvkf
DFiyH0yyjT7d3ImGrqKpHrTiU/TNcaVKv+qYR4m925Qu+R1MHxztgmuOyKHN/7MeB5PVkByiJAfM
+mPXsKu5k00WaLLJZKtClJIwt9zIWDuzgS91OxTmyBgdS8PNUjmNbRulehvh5C5eKwlTGaiwO55K
Q0V9BNZJI1YD2TLTjrCyEkOwhavAwJRKri4stTt6MuknglGxDmCkMFQTFEqEleEbMZZhb0dZ+p39
XF4mrci0nfSSH+lRb8mTsBu5FGbj5UxZb4xIEuyukWPCT5C9amJJXLxgw8xBVdTld2NiC6axq1TJ
Ksw9hfW84HJ1mdXmDPfX/K5bgD3/LT8NbjFfIeL4p2tJ5mfJI4Fj8uPjRnAjFLGfXk6im6vneg4V
c6DG9UVJbuCqXrS9Rzx69Cq0HarPyZDG74QHkZ8w61di8DG5Y/+x+iw5GB+cKd2hEzVpZz/JH3Q1
oLgiSd5Zbn94D2JNmoIx9ZKnxvFR+LcA/m5Th6RcAFHDwYu9w8XemdgLwDl6jkN6qt+I5Bw+iT4Q
4pbZozrJjnad+L4kbfHfMgBbZlwqMT3Yr6RWba6NIeMVS/9X5y62mIgHjjUpTxLnI185g0vfBtZL
BR5uHNZxnpkNqlsHAxxG5T8zAoG55tSQQr3hCSzyNW0Ow2kLxq8IPmUeiCPmB3+r6fFM93/hghzS
XVPjLRE4xqumdh5C4D2s+hOvYK8jbvy6zC//NrkARVc3NlupHpbxRhldgsxf5TB0wF6nzaKfg4kX
YxZInPFfvt4fjBLTRVGq8u6dlRFReVMQMqnvYOfJk4j8/Fe2vnoVXGVLGHCwmXJfi4xvbPvTtjaX
RsC9aLXfzrUoK+8Taro0iFox9BlRMh7QVdf9HOrPGamnxn+sryYlWWd22AxDa3F9RIRZyQCfFxs0
WXtNb8Sjq67ft4gEN+2DG7sf1qwEyV7FdP9zPPNBYnjOdnEGX77KrZghnFuMR9s7Dci75rBDDCNn
G3T51hdOFEzfbpJXwP1PaPkhKsJkMuF+mTi56TC8bsfll5t4sBcQrWaaCWjpkGIXZoOXIh+aWlAG
ivw2pr4iLaIuOXT9wo+pXOiS8i3mcoFIvY80hlYIjq3iQmRNiSO+ETbaqZB7FWfJyfM2ok2i5fzy
n6MCRg2gEZZsJxbC4Uqj0s58qm9YHF3k2TtkrMKnKSdJ/MfQ39d1/05xVOUeiFZfUG9CclABDz8G
Aek6pfdOw/IaEYGv1IMCu61mRC/V66VLjcTj2PLjMA9Ep5s9bYmF/jSrG7iJm1uIvm4NHf7vkXmr
HeWuGnMHRM6i9cOXoxSdGA0JDz8dxQiZlFt43WoPf/GghweLmKz5gs9uq8QAhLidyINIuwRSw6pT
UXFXOuUVawIT01qtQW2B56n0obri87Yn7A/eAHCtMEQSjCS8zba599kuHCyDazINUPal8ZQFZZpk
g9kx/0yhkhZmXpZ8hQUh9gpfruS7AaBXDQqfR2vE34/LKOFzgSOyFUaMTgM/BVrkNtCmXS/3GzZk
w5Uuczr6e7/BcDbJLOT/Q8ta944liyg2JRALl9eji+iPD+QmgnDls2KCYLqa7sWh8ad2syiHJK19
XcVOJv6rxza8W8IOMPWFieb/y8CM8cuTtsvjmWAIpe4YGGZUA7f+CEPquv6k15dIxK2sa2OdAKKr
5hWHZ8TAmfop0opfXzecQE8zF1J1wZvDZW8F8w97++N/35902FRDBRP5f/jwEvSr2+4g8Mled1aZ
kb4n1oOBP5panE0R1gdbZfrhzYIAM3fVMWvnHwMN8OwR9k5T2DSyyaMQ3mgi6bpQIILZMqny5DtY
89YO8wuq7t4ujCQNnqSnEGGKQR1Cvn4VJajMKz4bo80AcAuX9zwvN29yEMeU+wk7Yk9pKTkrn32k
gZFpYuhGIgwmz9ULmNmUuw9+KxnAg2NmSCSXt7daZvQNrrOKn3GnI5matKC30H2h+4gwea39zXm2
1vZZUt86u7J1hbjyHJnVZwD2SwVP2HxtUF6luU5eos0Jp/DLSATFMC/XtVwSSHgWDOH9Et3lahZd
za35sHBwYEhg7cn8jTJj7ZAx+7vOdASqv65QGm5Dmmv2jJagm5J3Iu9E4PJE+ZByz3xPNj2L06R/
+FAkCFl/nfJJHP5WBwg/QMN+3xf6nYivSFvmJBbO67SZ9pbg5Kn1tvk7Bfa7ZvHU71Q3vaJRaTrx
xKEb6FO0nmRfqF2xed0fq0Q6EwJy3u3CXZO3CyzDbUsL41chPdClvAuKjQr7LQ6u/jv1V23nK4pj
0XyaNfGP1mkEzx8hxrLX61gxN9J6a5EEZ+9UFnIkmDtymRGPaxpDEBWnRd1OP3JS3SmmpPJz71oH
bwD7JYddWEvzoOkaCSFE4gpceTwyyQHJ2wlDwuD0KBJKaiv8wULh7/zxSPTJQ3Vf5PnhC/SIoZHY
nBXVdqJPQLMWL5b4Iqrt2aoUUGvpF9HiaQwfbf+elM07SJ3M0oaj79yUcZOYA0mvhaev7PpCRyXp
yruD/RWPctyCIQtB+LpJgcql1/MG9d+f6NrdWeKSa2FM13fmAvK6OUWV5x9jXte6kSv1heZl+3gA
T7H904Guk6gGuKDIGIY6avZnuaeKrDue2mTLG6E4YS7+B+9STqCP4Ij7aEtBEd0W2IDYrPHYP8gn
kEBYChY8ZW5HVH5Q/p498bbfY5YUrackyDSSOXyA0rXspZOpyffnIsY8rVjFzN9i+O4j0a3kiHCe
P18uuhXaJwm1bvZNxomKix9ohHc+XBKAJRiYihUQM579TntHwvZEoflSpy65ZM/+aiDKo1Aay1w4
7iAfVvRGQzUQFc5IVLFvWjuYU2W6++crvBVTeA2zknwOlzVekNw+aDM9vuVy+aqNI0CGlsbdcZaM
IDgKwpNaxq/Nlxm2NKZjfznDnz00/mZq10dC1il0H37K6mG0Vo+bEhTxWx8rl/nQovCxzNILqJde
F9BQJUURKe15HXHADfEuZ8WWRK9qrLYVGPVicQVhVzf+qbO9hIerd27JmaFMqlWLDzU2Q3wmp0Su
sfHi7gmyAw6Zr6siSMWy+r6RSWMK1V5D/FH3kvaP0UZqZzK/duoW7h7pUqUJMZ/tiiklddekCqCF
YNEOLDt/Ef/WfcQpjS3dCuIHWQuuy7lqmyb9xBz3C2oSfnlR5BRKUnwxi7eYQAAURABYRd9HiPvS
7WSK1YJAyBusstBJBQtu8jVZD+o5zX4Hsn8FWX7WdGvavMmLSfflevwBN10CBpay8c8Iwo+xwhHh
Payz1xBgkCQ+UiS8adWnwJIOkjfC23Bli64NgWisifIAPbSCpErXuvURmmgiUP3HrN5T3wNPXRP+
SgASCFHsTYklUO077lDDFHuDYJlf6nM8ydHaLzwx8vf4ejlzfZJAWGEcw5ZhSboeDiIvEL/k883t
wqIVGhNVWmXs5ufIghUzhJJfm2dTV1WCZ1c2wdvCtymV6Z9QvVsJwg6eTCrTz/w43y0zfMlBFWxm
ZwW4ELPcpkDvyfN/sGEXRFy/UOFwWy+lp0NKx2Z4B9m9ZTADaEGPZZmRar44V6Hd+VJBow6C/XQM
a5aHqHk6zLkMO6cazoRSwtNvBqMGS+lnzskEjFuIRxMX3QLdUgQ8zkt5PTCgN/wAsOt8Bp1WtEDR
Caq3vpnZvrWxRSKwoNP6qlVpEt4jcPYLXduAhxSHWnC5UZ9xx590Qx0o8YRRbyO5R/w3buO4Zv6N
HTkEoAsgeXir4778PXAtMqndgsscqG5Za/R+BmcG+coNDn6zoWFT4+OJ6zFg/WVHtkHd6LHI0hzU
Xe01PW6YpOAKOdxWKqAC8AQgSXnyAK49OfjQfmvmoqfw32JFC5zVe/xfJotO+8/z2Hnlq4oguB5M
uaWEyb61KYf7OYt4H5SteK76aE6j6ykLfTk/BxIRYdSRYzyIQbG5+3JfwHSUCNIcbhPM5nnf0Wao
PucBuVbt6A0mOFbhWAS287KyVpDSZba0KnaBRFmzozA8Lu10z1R9+io50LubPubNK35hujtCvNll
teXnpbGTgbtzGvjonejNQ29xl0Npycmqn+MUlbXDwaHy0i9g3X1H+fyPA2lfpl98AzOr0EUywNoA
6CkywTVg1fUzF2XLv0NfdNtLMP9J9R1a/DBrn01Rn84sUhAc/FGdnKmZjt1W3tyl3G1XIntcIIFY
nYwM6vrygP3aEN9xZ9ZeaxryO38mKdzswDtSK7IuTiChhISgW1vElNBu3Fk9nv4Y4c1wTPeFjKHS
dysyrYv5H5tHU2aHk5nzDUCQC/5hPfEwBb8zvfYhr/4BfXNC5VpTncAmD56npTfcX5atuiBioc45
Wta4RLxMWV14arEaDmt3arNWAc9Tbbq6SPH16K8eg+4MnuCoKgt4QYBRKznh6cRsmqAIV0olDNyW
E8etlgofYLhn7kqSZKR+/K8HbxGB8HJpVkG8JY6jzf9WJ5Onc02VtsnV8vQSbNqPR54l1TSuk+Zj
FNuafKXveAUwq0N3xE+zsTby/2zsIuDp10pi9MkTAeeKjQlz7Ea8bngod09DTByzIZM6mYKzF31M
FkqT/7Zt0v1qGQ2InY5lLwH0V97Pr2RwNwMxoogk01PZJ7qO75c4XgvS3XXhOn6zh7fid3p7W+Wn
aqdTqqd7pZ8gaRbrIRLYY94qN/qzaTIXkFumKvzwq2UuRyEk2yiLzKh3m5z/icjvDKpt25MX07e/
D/XLUDgGeIOGS2ywUQEzO50+gsZNuW8wuj/FfL863j79uUELVrkIgashUf1H8+WVO21ddyNETJ8e
1mW2jgi/fVd62YsF/hL9HwAcuYbB3kMYKj2pNj3m/vJp9kqAgfZAUVkOZP0gjgfLggeeSfPlehCk
+ZnpnJ/+z91jpR0TgUc7ybMSb9hoS3rmn1D76CpGNEkt8567rujbvxfZ9AxmH1bhO7LdOP0+SRQt
TigfzTCVIsAavNMGcbGI8xMEh1TzLmwjjvAUR/aUY5wVSLrqdLF+5TW6VKd69tL07bksw0RlIYAi
2n9D+VhXGuecnMseVVFi6Z0rUF/iJxUZwNc0qVI9xUjeCnggdtTo6HZHVataMhQbeuw/ALpe2Btz
G+DxbkRnhWXDgm3A6WlOIhk+86+RMXlimvmzt7jOtol85f1B26FMU73J7N6HpcMUKmCaAPljamdE
jiCBOoG2rGhsaAQaFkcfuMk/sk1pRQ2PYb+hP7bn/xddG/XJDahnXg0ydvkmV3oJ3iURQ3Zuz9in
ckEXjvI5IdwIEh58eukj1Qri3GyBnH+5MF3tdQmxhFYQbQspgiiOFee/AmuHGxKHT/4ulCab599y
HnnaN4j14Gb0GhNYAXuTGbxwU+eKXjdZsboZRu75h7KGJQZTtf0yAmQDjY+eb2iGWYCTwyIjg6GC
NkMwOFWOgMfbU3DLxTghS4XSGolktUTL/xcPTccq9IMkbpf6/HJJ2Ry4C4mYtsuCvqmE1NIuSYs2
j3URV2qrfgqTC8OWjt3rcXRXj6sl4+j91wY2b96c60MzLDollYwzuVjmnmL65I6rAHT2rp6EUtJL
Wi8RaxihsI4+gmkmUl3O3f3XFvA3PNFhswH7DqZEDg5nJNI50TVd8p6wd6zXmqRE8i5RUOYQdHxk
z6JlbxY0id532DQBonbRBQNPVpAjpUD1nUOUykUvgp/yq/v2Eq2o5jTs4Xxw4YH+nB00koA85dgg
QK/pG1A2gyvN2Kz/fpg+KXCeOwUku/47OWcAmvx3nsDxB4VClJS7BJ+SkVrTV38sUwxCVQIZXcRV
0QDVypiWM5WDa7QsSY5zRL5Vj5ue9eQKP0M48Fd3EsVq3W8in7mF13U4Jj6NEOjDk8kW/UXPryIs
nJNxdyPAp2xu97IuI8M+rJqkAeuTM7ORZxgy9l5mSsTXHtd25P6LpGc3CxbwNnv8VLRxRwAApB2z
nDgQhQp8Qj2HwNh9XMJtGwilafhKrxzBLs+U3/02qzs3SUtVuKOu9J1CdmwUmKa7cwj9ttC3p83M
jp49ORC6bedQZflTPiwcLA+2t62iLRg6O2q1faSxKtN3yJYUhUKj5RRJse5kbWj7D+3+s9GwWHed
r+QuAMWMH2Q08VSkhYS4QCdVL9BUpHAFk2iGYXvB7YEFRPxDFzVL9GH+mafiHxqmjcVsXpt1LNXz
+1l3bcoLII3mGVZufej7obAnh0d3bCFWpdhdTrmxDsMAGqKFb2x+3ne1IlFu/SnfijR0moCGHq8d
Fn+4ZRtqsGdqkhVaIP2a4WC+KA6XXV0HicR6Ni59nfDX//ov2dSjNJZx7k20wvO/IERzhB8JCWXw
lSntrTqh77nKPqCxA6NGkEVfajhecKnI29RP3NculmiXdqOGEFKlcG4mkPgd/4MF7Ei/afECYq6x
L7rghN9p2jJIhAmN/+8dtHTNl0lAAxUy3pdKQ1jV2gNshtEr0IDqxNyGwAFsT02uQ38CVLGk6MCP
OcQUohGdtfgqY8saOzdUh/uQkycOQLYgskixEfuZiLVgAbdZ3/92xQefNmr9pzMOikcgfi0LGRHQ
2Jg16CdwHqIy6lPNa7vc0/BjXHoKFWCW0FHGLzTHeTzldWmFVGzZaLuN0MoHR5YVRqIv+6WWPQIq
OMaqS5XdLK7nLXEMhXaWXGlkfoRKftpW9Ok5QiuCIQsN/pzdRNiy1AplRkUHirUreUqhcqDJ9ro9
yxlx+VYY2wbxi/sNaG8D6ZOjfPJG5rBVnsszxS1+rqOzPZ4DqnYRpeFTpvnGHLeYtclhKJiY/qP/
Y2WMc/KiBzMgCiFyXQCvRr4A7q6d5tGczXW1jd+E5cYDv4LHj87PJAgU469japTjX4mRAOAeRNBt
UsBTAG07OG59I4Rwgt8H0Zj5UonkE2sKtSUKOnG8FmSwNMo9GegRjy36WOlN3mPuzbZ6pUPpL+Tr
0+MkmxVwOsRI8FKO+mhpI/UhJaj3sXLyhjjaJUj9TiLVdRpTKgizAaLZS/MPgsmiyJNx2pYYVCt0
aOylyTcnsVuEGpEHEonRgVOcHPF9/Jn38PWdbSQ5ZiUUAMNFUo7dJ0iiIEiYx/nQl8W110J5v8sg
ZNSNrUITry/eloeY3SoOKqVVkV5lPbtPb8MT444/7UHMraiCFzvK5Qx0CF795YK8lXtCLG032+pA
ZtEPJ6a8PIVoFVFRP0yGNkxk8P854mEleWj+PatiKwDwUWjGMessrA00jB3cR34hQD6UZL0Z0m+n
/jgtGPBUQFruBMstGYGyHbyVMNIdfqpN9HRTyQgaRIuSbLTQJ/id02Vs/c0VFPbS65hl3bBdewnV
/JWwwP2jEMivVG9SgBjQ2tPxNsU4zdF2Rfp8MG0lvlHw4EVD3eP/3IXloYStIy17Flt2ujdZb4BL
SmfOCNLSYlWHwmxIQw14UgTOicIaF3rvHZnt1++lDoiST02EZQvhKiAABmKhKgHri/si3BYa9AB1
itekR7clGqDP3PK0eNsaAVz6TEkPrMOihaMKhfrP1v7BneH8mUPjojSJUB8D2ThSgr11KfeqQlsK
40C3qAfYP8ZdvIi6DopmFQn81MezZR8pQFiFcme46dksX3/k9dBPiWZAS6IaxU/Wh74BvtR+d1x3
8J5SXYt/BJ8vnw/YZB4VvWaxROLmgL7NuOFEs0lqYkEnTNgS8TO0oP8s3RZ4g40IVUHLBjnT+Uq3
hw5Q7S1u06HCnLuOjhqmuE/FHafviHLuu9RMy5/kDnHGHpA7MbqoCgjl3KfAAIDgIx3vU/2z3KSo
PVxX2twtQudrRbDrwCLPxUp+cs/94XJlaodsweugjripb3Ste7GvrdDFjzwa6IhlO1hoDNrHc0pG
jMrSfErQ6hDnBH/w/4mVFir+WkFlOXhjvecWNgATtaYEOAM7W4fbgDdkGV/g1Ft4aA7w2LDuvubR
czREDUe5SM4sHGuyp4HuXzqTr039+lVupTaxYHycxuKWH4wD5++EN/n9lK4s30bNDFjU9iMoon1Z
IMFCeI4k6PR37GiJMsq9IrJraGigDumP24Rs1tLrpi6+7FeCj9yfPnKuMnoXrOXoSAUQ3vSLjPSb
bO2SAwSZjF8R9oGoaE0y7SMXtGSN+gkMKgowtI//520i1dvbwSjIskgDH3LG+Hi237JQQIazRfRn
y3B5FD1THEQAP5+ymm0XIFFyr7y9mh5mNfLwgOcVvslAG5vDVGCCW4v8AtT4QXJrqOJomzOS1+Rk
XJR8dD+ltioipfahKE68Y+6nMrykUNWK0TKBRQQP+oZR1cCZhe8d+uiw9T49IrT0+oHwT7swHHmj
jcAltYIuG+BpjQbarqQhEIqsgB4o0V2pf9CXyPsZzzFbngs40nPThbJTdaNhMjn3THxLOclNgFzs
WN9FFZ9tIyNWReY7HfOEEhnpBdX08ovNdQz4uIgzUO43EiEdl/LkwH5AL4QldQxVN3hX/RCvITR+
WSbTqx/u1UlfCZu7AJLnK2uqb5fXFGJ+rqPswTLjnebCQYj2AqXO8JOIe8Imk1iNcI8yEBAl00tr
fUF8GR1i4Cq3CvAN5MZtUs+w/ZfzEjTRvHqANWAcZXbHe9dvhy2xukuhw0wdbmt7gEEmrwjyPCba
1HJRC7s8CbBdtf113/P3tb2y6bwGWCJfSp1l8lE3+71OlMBl9Wno19AxKVEVroMt620vp2ypVSRC
MKTz5fh1VWhXbXuroPsj/vMk4CezP66boxi3X4NbeYDzuLEjHAs3eeaRpHUTqIq892O2DJcXbVZx
zkY4xL74Jcu5w5RhnpcqVz4XfHtIXvx+Z+Iid0p1Qh0RZE7OdYVueoG2v4dfDrdxXbtUhRUrMVl9
Imt3HRQdV94QRGX2HC+SndLOL/W0A2kqlN/tj/8HAzHyo+Vnz7w2D/DOEbK6ZD8hkM16H4CFTa+m
faQnfWfDb/cJb6jGcnraJaO7ntiSPMVtcW9uw2X1upHVtQBABn/TKhrSDIixt/jsdwMMB6kcJf91
pveXjbPqcSAzRFGaWJNPAVYLh44PCEfeC+D2S6CNK1joNrw2pX+sCq9PwT7x95fy1MtCPamHfmVa
PgeaKLNJrGzZDIGYETo5DsADLlZFqgeJDp6jrv4Oto9poWwRgdKARmpBc1d2KsgDGRJ1Qo11X5nc
6F9KyelMwRkxuynI5HN6W9i1NSGFBvE80IWh8b5vb4RWGKgDO7fmVcqGN5PPHqmxTUSuzy4pvIgM
Lz9YX+ufHommuUcqKh2jAC2wpIvx6ETkm+YP5K6OmXiTDArmKIi6eseRsJpBFenDTaNTAq71aZdv
FIBXexrVtL1fhQDSUyupKxczA0scQToErlYRLRi50B8bv3c4etWdd5LsPq/XN11dR9A1wz4Y2HrA
RQPI1KX1IXGAoeNVMqaCf4f+y4AU/Xu+VFPYobFvVIzg64Y0wtdmkYSucbALojBvAMauZEITACIq
v5GSldnexpAs9K/sQDRAIsMOhzY40IjvMGzzbf4/A7ojIsReDs9Nhmj5NctJ6iZlS5Pjk2v50FG/
1glwUQFsRxOaFK6DDOWIIaqpK8hul4BIX7c41NMjCh3iZ2/djGb2mrVSK9u6xFGtJDbUxMK1K7gT
opLtvB/0WeXmNdyJjdIsnaL2JtRsCGPyqTgErUhcQElJUimeq++JCOchWsQpmX3mMYpis6RN2Ukq
yrHo7B6cMrnwKGcKZz4ep8TnIvv6prVPoY+O6mFPWKHLvNT2kq460/xy3BxsbLK75EDPuSmiuR2X
h+/olDdhieEc7QZDlaDf38UsXpfZHv/Nfb60tshfIAiUIPEAyHduBnokzdfPnwabHx2B4hKb/qdt
VSlLtAV+++zvNSw/g2NaEX9QoAN7k+QE1KLCYK5Qa3zEfOE/OzxQOyyx9Tb1fXYlwI4IYX//vtLT
NqO1N/iuep2eDQVn7o6Yen2eoP/YwljqriEKF6TsiHmrQmAlKLmuW2cLS2VXExHAUrfFbWoGyUZi
31cte5qkphdf6AJGdVjUU8ydTB6XJBbB+T0rSiZ9DiraDhIV/wwFk+0O3Mtn8Xs1cZRZR5DJ9O74
5TdqgZiuYAuFVpVDMmYRKE+fnYjrejjksBi/nAZGj5O0tBVNaAlED2tCb23m1ky/683NSMc/bHV6
G57btkkvTJCC1Pf/PHwYHLQMp+mjtuNkJRQV29GbfMGZXZE5Im8p4LE/Ad1wEedp+o1GFAgrqDt4
P3Qa98oDB+4MB4KloL+D0J06wiClfXt1ZsqDHSnVTjXNPhqE+yUuKmluRWf/2wzdL7KuaaSeoiLK
p73edN/7iidXVv0Z+OKdnLd/Vutl7hKNMWC3P+w/2gJz70CqX8PuWSNjAk0Cqg==
`protect end_protected
