-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Sd4pyN7JWuOZFQOc1sPO24A5b5XIFuF17TDZfz16KgPdrpdegXYVBAfbyCEQoMf7UuqP/+pW2KGB
xrLRWO/zhHv95dc/O+lr/JS0vaOCHWLy27kF/QTh0W3NWyRMgPpdUXRPdsINprZX1eWU3Ej6MWs6
C/O10ZndS+zm1epuNR2Szpq73ASWPDGoY7UIWV2MLca2wicXHazBMO/psQr7Iih6b00XvUcISZxJ
M1wkM6Zem+Dg764nWkD0Hms5sEEPjCs3UmPj1JdtA3ZRQ5LJGXzEur123NDZy6Eua+ju9dQtSAzw
8sIMFN6YrP0ra2VG3k7scFqTQIimpq70G8uLmQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10624)
`protect data_block
VYM2ThgCK15zLLDG+ZBYP8N4RzDJ3f+HBkTTKF7veMRqwmUN6VqdNbSUXwkHA/+VkTY9yZeUHSMc
wsCeZ2+5ygsOhP/ftefoZZblMnVliy9dL9Wj7xL6V7s3Bn69v/OWv3DySBKIrd/NnHaZeP0RMJ5i
23OyJ/ASzcQoMxzA1M5Odvx4s/7opzn2OBDVkdLuOExFkw/7qt8RJVErRjVqcD3Xqn8yv48eA9C6
Lt1St+YNjFob0Epy/4HinUK5E06OpFY/33CqmfJtbo8r6NMPoEtWjcjN4mftW712eB1/eRp4jkzC
EUao+3y3qmnPdB8Jy37wVrgfqJIFVlfI/qsE2YU3WRp13v8EYHnV8bhSJr1dBPt8nzOexOlEj94e
sF6tYTP+4XS3vgcLEH1sv/DZQho2o5eeldHJ4ac/N2Ngn14tr2Ig2bqmv50M8CYbVSbv+4v/dpMs
3yR2Qnl5E/ijapNv2Rzr8Cnlnwy9p4BpJLGOS7q2JCvzKZh4d8GV7B/VSmtQih63MmYga1+2zlLm
Z4kHbyON6PZTrqfZbzo73SrSKXKfqALkn6xHH/YW2o0bJezcEHljvBOwl3+hgA83lMkLnkST7OB6
3ITVg8wx6v79Q1fKoopkgzWJbhvUh1F6wjSeFtWsUlHoWC33UDr/jcQeVsG/0gFWu00jdEmX+h6/
mnsOtIcuEJWhuDWyl6qq14tgjeYvGep4bh+/Aqqq0vT8oBR5p+U9EBRMeogJFZrxZBRPbWM89fDu
EP45+1fg78vkrWzVqSMvhR8Mup6Y50/0WjF8T4IBebqH75KcUqyZYM4Va37VNW5EKxkQzCPAmqF4
Nyn5nibCfXLj/dtUtpu+nAjsaQm71B2sFbGq4tMKcZ9XgHiRAEZBboKVka8yEcGduBkN5vnUtSq/
lruus0QSsooJynyiU8KS5NLre5TpiWEn9xuXsiCcFZliJZpS78cxWXbebvwFZqFtEMgfsv3cOLCv
C5ZLr8NgsvVtM1LHgUQk85yKwm7bNJPeiA5aOPbB6cRA6diP9Sbvp9PPu07GDW7aS7pVeqgydQ7l
72N/HCGFK+895TSXgmw/X8IScY4p3L8hvu6D8gUEZb6jry3BteUMPfI4Y8v0hlDhFhdWNghvKXkp
vvx4un8so6E+/N5oGpwIe/Q4ShfoFYiyKJumw2fBQ4IHgz7TLeb0Zcy4tom37i3OQen8HSpFbUil
vBIADE0Oh9ixpEaJ9ipkS4eH7pBqPol6fns++x7U4V501xVEgdEb8YO3U+EhWkSR4cP+D5UnUJW4
+3KGDtqfCp3ILpB5ryrwblyR63fdm/H+Sq+SseFuLJq580RsPrkn658bN4YZbPrZ0Pc9ZOqLfF1B
374ey3+xvFgeJX1xJVFa7RR8OsC2H0ZVoxLHr+LTsnrzNI0P9RJl5ZNcg1dDezBPf/5H9pD0Gbu9
DbsXF9NiaG/zAmepsDxAmgepBOX8vtk6BLdOxTFKjitCimSY57oJMxjmROQ4WxZ7+AaWRflBUZKj
rMuM6YwdvPk/7KmclF5mmSfK5GPWH8TZ+ZnRGFML0LWT2xTaPLi0qyEEjoJUWwIfiyAOMNhK7Q+g
GwtgcTF1frZcl/CYYxCsl9hTOnigEXdrrERWLeKW7hd6GrIOuGyUPEr+qFZpMQcnqVqtxU++J1yU
DpSU1h6jGUkNqnUvfv8Nzv0gclx8vX7GJOnJPLWVJQKSJX9RQVK0R06g5dGw/7BFGgplNex9bVhm
dCKeZ/mIvHU5d1o3BzN8w9mASOPI2hxJF/e8oHE5bNAsFIAuqxjJHHlxdJuT/9vwfxP3yBYmyvDu
HUPzDQbAIHmhk7X5GHy2I94HqIUl48ukc4rNZwaAuICi13hCu4zUG+/Yk3+fAZdOtYGGmd62Dr5c
0fNi7ipVB48KJAz6hbSNgZqQzb1uq81VCO7lHdfWqbjpU9RdpdHEhBKea3hP+AUY/v4Twzfolrdk
0qFLd56xtvfEbZjJR3V8EZy6YLkvX/a3C7uJ1HqMQRwlDzGjbvRLPV0F5WOA51jNt4OKNrzLJPWQ
zHvMaVkN0dzbS71DVQ8W/yM/c5idrYoUdjgL/1HMK6O8GaQfRy3epi5BdbU5v34T7+qUracjdOfr
zGT9r6142zADcrZuJMJSff4KRiSgA9dbbaGGGZqLtRsFDlEAVKbb7fTQFFQK6YNy+f/RDqvZvuZ4
dh8pdbzQBFGaM7FMxGfi9so30y26+y0/OtvsxMU2OGhEUX0raRpl17q0tsmY271t9XRDpeAeqKIc
BpckDxkIwpmI/tGFGf69oVtXCkc5I48T/ec8zmZUdisnmtF81MCxMSwXlFPk+65G2X3TKMSBX145
JdXc0oXtHR+exP9c1tcb+ziIOisxs/3UU+mgNSRUdaHng41+3/FJOYP1anifRlUEZ7/6VL3yOVXZ
KAi9z3wJ5j9HBcubJzM2kbb7khQm9c0SM8yCl1RTbZ2Q8Z3V/5wMoZAeY1fATkz2xnDyLmZWF2GV
kPwBBt0+8QhDASwdr1CkTV5lJ5lI8mxcZXSyHoxnDVLDR+BMZXNtLOVxmUd/NKmvqNH+XQYOU/it
caB85Kl0QMJv6sAHswX1hLnGxb74yquJASVkn94TgEnfJbIc/rnRxKPUh6jcOahiWJ2Y/x/dmyPm
nQmBUZem8GcKK46h0Bkr7EXVppnQnobbhYdDMwPgyxnfSuu+pRGBAF9Y/MJXzUhsTk03xpK0QyLH
78pSRCKwohkJAvzEWk+6Kirhh904bNwE6RYZ66aWjud9H+ePUXVLY+u6eTwo1DahxX3NX6g7IA74
wkwy2G3/GdNhDXCDhXQXcyumc9af4XajbUKicG4BSyPx0tuNAupCz49tz8CkGXn3/ZKwCC9oYIMt
mohheaWeCehxH3L9pJ6VH2wmJ9vt/udzFwobO9rcpRalwLZBI9LZTYGtyRI6YhPlNG9nb1+vDtnc
9WzEF4xImceMZtlO9BJZ9hmNvbO+IY98CyrzKHyVuDVAWsjtsdTgNGV2j6e49C1DdAzCZu0SdMM5
L0Fq0qq1zzFB5oHjufj/eGFsoHr1kV/VSN4dUdljpGyv2OxcC0KBSH1AQP2hGD4fNYtjsBZruv1W
2MCDF2sOy97hDJYj9JoQ1P73DowADRJ8gben0STdF+P32s4qy3Pk3jrAHH38NMwuY/NufrYSPCrA
S9tUnMmOM5eRjTezcvFcAapOBU9dsSqOcXHO6HfP/0x9IUlFT6JSFUieXRxH9QuzAvSLJFaV7Ds9
oeOKH6MPuw8TalEtISmG5pofSBm8mDE3nkwkhYSFmh8vUWKgHK8HmlkCRZuN/jCWBpY/kBPbR+3g
GaopLmHkIQDka2LX4KvWjHT4hrOG5AfgnYNSR5yifA/QqFkFEQ3V+xRBQLva4HIRufxadQ4bk9oj
cEMQP7vo441D+k9sX+XiZdO9xkA89aFgw531jpZrSGXtvzGjq26oVc7pCtOjEGGjLYILpknh12WA
t3o2foqOYlN1HuXnBHORUM90VmFsys6HgUT9fnVwXMfhZMeSK71FJdjhm2NupIgxsvnk7oXiRsIs
aoDQgQzPsmfgePZhGd886Bm/6SQy6Bfmz7ezFnbaLQZbzNLpZHvrnQkNjAQYsGjmkYbgdCFHWpIm
CTaqsbiemkSt5YOD1RXagx9Hekw8yZ6tL55S7LsiqvWasBBfoRB37/jrQh038Yb6ubV2ufi3/mSq
wFzlba3ZraG02kG2OEknlYVaNFlcRKVU55xfl/cvwpG/u+PF4koRWDQRE5J5RxrI40wgZRM1AO9O
c3XXc2NpPTUy7aCyU1flyDLIoXVxspZ2ttKQ1prP3K4HfsMmaXr8c1R8JufKzecea9rgevJfSYMt
7geZWCfn3tn/5j2qU2V9LV2vBml4tZkZqxGf7QMWTQdWjqUrHuTDAfJxMyeqrX5arb3pYV4T+fj9
3YhZOCMDhVB3xeQDg4BKe31F6NSK+NVcJhfcrDhD/iOmR9C0a0EyNgmTnCuFnVEBQc1i4LVpaYKz
ya2ncLuQPlRZpd+NBrbUU2ZmlDH4NQllonWEIirzCfDrY6hZXKhkaeM7/DKyfyhpbHRzBRgARFN7
/j1XgD4XgtkyD4wv6khY/87D4U8akzqFvMUyisaCLQXo0L37FVTPmV1j5qirkWgHiP92UUGUEZ7p
kLZXjLnxN+UeI5gW9NaVl3Y6h4vdMLxBymUGTK3uVE/z6GmehR1GQWtuCkjHmPKGXejB/9rQFwtW
UALBi6kI1iI7k42hCRENiebC0nfmMt+CRo5+6OTyrZcKg3yg81L3SLQgKX4x8wa4HCuwnekzk6mr
IqabgbQIaBYU1N+/Msh+HihyBfhqv4Ny8ErWdjvn4TeGAwIil9mmxsgLkp+Mc+lbj2smb7alo+A2
m0CvVUgW6k+pQs1W2D9Hbxz8Xp+5fcDxgSiaBrDPVfcWbX/bwUf7T1aRG0CxXDOCsiRGJ/Ml3YxO
hSKBnoL/wJCSXDoq/mazVgI/riGu/i5oenO2Yp97Kj9D1nrGXhoh9fA3hx+lJw7XcH+dkMHSAzcV
CfE9X1C8bDPigNxbFVoi1q7TW72MgmJPRKX8vcaqz/q9sB1R4xyvtdvM6ivcW0yQ/5g83ZGcRapx
6/vEKCok+vtC3gMAZIKyWG58tbRRoO6F4lpuM0o/eczKoBEbg0hlzUcGl4nE0pDxr5sH+4/IzcFa
5wFzi2JNrp3HbOP82MJqCv0J+aPjngm6ApqjwKhg/qBV5vow+F1HLXSPJQLwRbRnHzCNc2W9qmLF
djsOhNlguItRKd5SQLgasQc+mUjUBcAi5oMHrrQj/WXh6RRFRWnBfwB42o3j4vvqvJJNBA66bA4y
VFIa7hhgq7zHVxnj+vVJLUtXbfsfTpXfIzSBDMfGLKuBdhJuTi0xAzI9l+CRpjkPfB+SCrklsAsT
r3PFMtt2llQ2iXDy1RecQASXH+neK4Q382jbLZG9DvnbzGRBfc8zwiBotvvx28efegc6BD8x0A88
oYJ24qNRk3NtUnpfE0RwTwNjC89EQuPTRy3c2Aib+IspOCLD/yjVpXBSwFpsfv1KqGmx92YlTrW9
1Aem3RlYhjrJBr1GjMivtY54CkpGS3OIin/XvnP72GANfT83S0yNtWlJqGvPGPLXdCyR5n1CmkXL
KlWWnDUq14KxDLXy0vVdmeMSg9ul7VuvNheh9LQ7Ac7ZxkQPzBBTwXaO1hR2c/8bv7gjT1gDlRX7
zGwsF4xx/50DbCqPqo80e4Bs1A0IPCU2I+E9WqRTk/3FErwM6FlIl99Z7ZK7VU3p3KGoyJdHznkG
TvuPw3y9m+bkXuU1+EUXNVK54AchwdSKNFm5EoH9WG8fqHdwpXNyMb3aK9h/HRYt2iMloyYuzHq9
tv53QmOL5IhaCyk0ydjsOahL5tKf0tB3f9o2O03paaWsxL+Z/DNz3xynX4cVHWZzfAOcJz6aU7u3
JIbpcg/qDRt6Kp+H5jKRN3RrIvMdsRCMipk9k8tqShbCOSd3R0FAcCPVKIQVO2Rxah6FP4/Q+p/z
att/0X/pN+0hYZrJ6j2+KBJIzasicRMJuBiTJoTEKhbmEF8qhLzH96Mez1gzsLWsSBWfVdVt0Xni
s+B4zVNMZrtt3Fo7iifZ+t6XRiVJSB6NL1YD6QLAuf7rVmUVEkUnbFWrTw4dyyUZw05F6/0QDkkm
iobxk3lBnaGFZbgI5MQLqilmEjiXPxai/hfwfUz8xthHZ6zDA/DCgZuU2UpoTWi6DoG6c5bZrT/6
z9fUtYXLtVl5H29Kj6IIz+nOV7SlAbEUUT3YTW905F/6dZ0E4i6gersD1E0xIn3sCge8UPW7QTVg
pBdlrPPH28CCZ4tMlKsKoBTrizAAFIbMskaTDlmhGEO5wGU2eTb72BsUmIU7p7fnKpKBphkj+ELN
ldcotA4BCgRtdj0QNz+QyT4swzPC48Wf49U9qAWaKR03BUyFuGG0J9jkVmENX9ruURZGvClIVhAz
eqwokAB5ZFCes5Tl2VKI69kAG7LMDpkBWZyYRtsSsRz4xuJgqS3RPzpG3Hw1n1HFGMQFEY7GqrFi
XcLqlow1UQEnpp91mOx6BIaaqEIfc+SqgpzzMlsnkFfGy77AYSfDLNGMPnXIw662oSmdCsfVqAJm
pIUOcQgLK7yvGgKjVdVx1FL0v+WZiE7whyjBhSqLHgrdpP4Qd8kEwfqGt8vfREd1xrLUAEI3Ksgj
I9Iye48s3Wf3Kb9WdQqsjfOdB7xzX8g3sgHAIYGBdY6Ki7d/TLEwY5PNT2lEyZUlavBapICrpsXk
tAtxlKZUJX0iyW1b0xuozO5QJzgh8bhjaaDvwinqL5eJexyhzknsNIc/W+cB+uyIcyb77XgdN7L4
Vu6XQMvxXUWnUOonGwIgH6Mg+aQLN4amPezkn6zEKb2Qduzx5adb1Gs6KpyH0lFqR5ltfhbln2zP
f6qdySnuM1l+orNNlrqxAkpDPOwS9sVXofyIG7AbXAYBcO52/aUZjleKQDRVmkRC+8UpeX1NuysN
mI7+D6g3WR6jAyqrQifQQoWEmmsHkGsvQGXlG/HB+/B+tOU20Ri1c+wci1T/V/lwIBVLsvefibGn
CMw59MwH3sg7tuz3L+bdWuhaZTSqIhZ79uPwtDC/dEvf/F7hZcwaX1mAXt0Dq99lETxlu1l7P+lg
gFE/phR0E5AHUmSLF6Dy5qMbrsQEqu0Jt5j/d24GR6BIYaLsTSC33g354DF51d5eIHpYhwo7hHHH
zxghinhMKsOm8HSMc1uYY/fLPO6/9SXKMJhD9+9pB1/u+L7+fqNZkjBzky9DMlZc30X8H973qRk9
Ncvg6X99RDjtp9zb2h3056UFlRpjqKIaInyvoIuvqer/Rq4cfuOhBJwGQAKQ2+DAO6uoGgOV63Wa
ECcynt76IohYM4vsQ/7O/uA9j2RU2pe5jTP8yGRM3z4HK6VZJ00/mempiIYEFyU8288W6n9lmM+Q
ZaT3E0icKMH+S/vysYBmmytRSTVel8G+Ydv3H7/LLmeVW40ZTm7SengBGs7Mpvs5wF1ttJd3aeWC
4WtsLXV112drU4J7rm6YUGM5B1brVUCxnBsaHpEsQiRyGKSz3DVhYD1tNIaMb4xj7VKnxH+YlWRH
BndbFIKEzTfl5OE6HZXtK9Q9TC9LvsWIXm+bCa7JPISgNyivtkB11SHRkJN+9WhOn/8HS9h79ONe
U4TFfc13ulPsjhjUdAir2Dn4vZ8CVKs3mqNjb+QuuHkUCNQiyHipMRWzI4jq1sIoNDjnueVlVIUf
7TOkXB/GcrHuXyzdD3Queg1Nq52ENcBYtBcEpnisN+U6lNajH6e1gnSdsWpPLm++pNTA8m0Cww6o
Cs7kFsB2UTAhdcm6wj3HyoWDN+LiGJ9HZk5ccPuvaYUWdzBakBFg+AN0tQ/niIn1vGdvBTenhLbv
YvwcmQhCxNFjfrMcUWk6INV3xceUAJUGj09fOqqHV95SSEcqeOEV9vCIVP5dyirUtBkWvRzClKAq
cLQc2HYrk7w/peMstr5UsEmB+FQLpZFugQWNEr9j2fWlD5viOf8NIn8Gjv58X39+aGilmN3KaIqI
FAHA8cg7OcCQD1Moc4c7l03L6sbSfcTyAwVsbbof1D5tck5ajuDmQX+JcQOKdct49KvZ9DgykKss
iSTPnYww8a0ZMtZG2CQK32HEw3yMluViWHm/bvvn2KBBJiXYFeS2/TE4boj+SxmpCWvxKDK6gM5H
vtxdCRryTjVLRer58DKKG+twqX27NJy7Xvqv0IrZaSxZbuunXsw3xIOZ+toVG96YeWx2ISslkdOE
MB2MhFo/+4DjAOi0cpq00N6VVJBxw28mJKAVh0LiTn3vHY0mdsNUZLfREN7YpMQO2kfvodUB5gRS
B5yI5nIqx85dh3QTDsQpvrtZ6QeHz5m8J1ScTmhitytCugyQtef2jZUvFZ8CJS6ytRP3ewoCNKTY
lc+5NJpmrVYzKa7+STXspC85jI9CJNjonwrhWWjWs99TYklGZywONtOsd9tBjZZ0VcNT1Mjsk5mn
1UECF1rLgCE1BjAPNmnHoaE2tX3s1Bz7YMOMMgsFMbHdBfDWWzmrg9y0IvBU4n3aUuiKGfAF359C
MjU1/xWGV/f8HRP0gBMzZ77/GQGF81OO3GfCSoKMIIT0793avWjNQoHMtSyXtlf2fPM6qJn2OVdT
R8VdNLKRUzemLRdg6pcKw2TEgI3Amj/Qp9LHrGc2CvifTLqs1I3hwifRpfF07gO2A+bI1TnFVWdX
PT+HiEnbmWpfcVo1XASN5Gtf1ng5gh14efnPriQQo1MM3RJjwAn6aQaKyvYcK80p48q+MecJLZWp
izdnCfKB33n5QpYRzGdIym2J15wB12XsktlXXkM4CtisUms/4qINjhHYRruJiCpT76Qmgj6BLF+p
mEjwOc4/XDf6kPSe3U4JQ9zd3wedNTE913C4yZZvclWkjOxJ9GR5Q02jgo8Y2vwZK2lMRoKSbEJy
aolcAioKZxh997oZO9VuzJh+OSg93OmywTrCwZ6wrzkUJp5JoL3ETKRR/3i/bpfGVzY6O860DY8+
dWGZJtGS6x3hCrpfl1pT87TxcC6XFRMwquO7TgEW0EFFVOjt2+F0qR0q8PkzATkL5YNMurtu1yP3
JujXxLMcv6gWLx4qlOIpcnmRux8ZEnHsAClLdemQcfSMKOBJu5DU8GhGJhEarrvOTdyIAEO+OIPK
6uJdbP54az7wlctsfzqo6rmahTGYuGOHEQncafkG8GrNR14Yc1jAiLHBqvpsm1wt689hejAiMgS8
WNF8Ms56bbVnUgR5WldSK1eZhK3UbFWa19NPJlsUequNcH4RYz6pjjAUqkI3ynrza+702AgcHuoG
L/+Zp6LA4XmL32VsuLJ9nRoTin+Dveu7Ms/+UlLy5Yt5IRa72NHYPa6p61t1zSPnU/VOiNWYgBUs
+L2rxsr5OC1a5Mj2SSZa6k8wgbTL4H+6T1m6tTMJfBPGUSj97TTRN+phsOaWD4PhPGQPaIN0xNPp
A3qEOb8cd44i8xCDSuOIdM4cgkTQdXjL36sEjnh1l24Qc7fuZgTujb1gZGyO2uLRdxYYyRoY47YV
dLCOj1D5C9vZ2Ndc4U7Z1IK9p0L+9AgUy89+pABFmig1ulSglRaPuo90cdXqiOfFuz0SPIiyfTWB
eXgmUniM0umZAUgaF5+lGVseNtZg8npEHvbUagse9F1Zlbdwlev3AoBS6cpK1ub8buL9uxUxKpAg
b/ImxwxLA1Y+jljxhMIW3G8y4zvryFkvMRbCWNKAhC5fKDNLjaZdWl+s6KJTA/UrkDY3jhbWQB7K
wRbVPiwoXLpUWd4PypzyDvz5x3HZLAE8PNpAPK5cw9kR8kgTDylLBnmtfNFSd/UDoD8giMAzoVon
7pahcVMFmS4bvQRbEhnfSnR9yW/EVE4tUXTYGWPavKoxwdqa5Cl5e5HWqxwIkjYMh50d3o6eimWo
azOb6Qu9N+1W/BgAIt3T06Bqx9mHsr/7rxjrShOT1I4FNnyo7WYcOTOe/Alxr7j4B+yZvspH09Hj
oyQgXL8lJCw2jNZ/XEiCnO7sz/coOVkNc3iTYVU4D57itSImIVRbFqzln2Ypae0vpQXpfmp8pU3I
5VpZHUTw0Vm9K8rc6EZkmvZx65W262Z9gMGpo95FmL3Tq5B+dCCnJVEisRyP0fG/l3pp/9vb0S/a
R4Q1caUtK0kGFtYc5PBkDO3I4sK/bDkHiiTW6r9YquzU/S1D0NX8aMyHtRwy/fh0g3EknbQhA5Gr
X8IEoo5ZYTc6YWm5FXBnfMKcEpzdyiygqsAvF1xPWsvRdZjZE5YI1CFwWdSR4Y9IAiVTZLrdjfwq
FoP2rH1xfXpqHz9mweX5UPLgkT+n8wUN0d+bTyBe6il6onSa9d/3va+xa/3VPbEXcaiLAJZhzPKI
t3vdcr4ge6R6JzJutWYdbANr4yaLBUUkDf3tLvbN1bLr1UboUfOknCvqLCLr3YbtEbQ5ibZLYpGC
TljODeotQ1YVNKrJveXAFRQseVoJxizBKsfl0X8uAWBN7Lfg88polZ5m/xJ51sFZmGh/HoK6GW92
yqip0R0KSaPVq8FOTNbLIUT/8tEZEMOLT/9carGU9LYO3tWrWAFTYnhbz2QrdI0EHAi1tGHv5J8o
ygoN9ZFmbAnQN1Gc92hH9HEDfdBO0809Fe3CgyOea97Aiqu6yGCe25d7DLKtcJz+0RbjEdd+6y9K
ZhBkftlXpW3R9Q1fsjI2HdZFj7curhcWWUPzU7LM2gfiwNzkCgxEf45+USaJyxj6a5sC3dksGpG1
vyH4gMKb9Q5bUtrYMX2qdOhlHuqIMYCSGqeElft5fuctxY8pV/08r0bkfnep9xfUGBbzRPJM2BqS
+1mFsnhb/sQPBTXS8EvDH9WswHR7C3h4RcPHnO3Fb5TV/zBnB0gDWzeAxZAivuAo7gzcJZfDTYre
s68vr5Qld4cHjeAhs7U+Qig8ElsahXP+Pkr3AE+N6iDpQ7moWeThWZ+KKS3CdebqnmBjOP36aoTT
lsdBd70trCOPyB3nuwesLrL7ElV7V4Xopaq4C6juilhOuTXcbMpLzkR0k5Z/xzLSlDDrW4T2XIgx
fKDeez7SNS7xlISrybZr6NkkNBC42eHEiCON0x/K9szB+AswbN1nrf2+YBFhEOl6GpjpCBG0PvzF
sfFEPDQ37iVI7SPjlJQr+Fatr9FeX6AbboOrwdo+u4drWrGcqPRoor/RpGtKk8m7dnt/nud7k5o6
mU1qp9aa/PRS8rSExXC9ps2NJob37rkf2EkfYK3EDrI5L/IXVXMh+D8EKJ9fwILEqS0TziUCTmmF
0fplQpLRuiDsGMBQyYZJeyWHRoN7yCodJXWxffKB216Q8dGKkIGyV92mqGMfDaX3GNzpnrglVyv1
JZScdl6W967aSD2d2KfFDuwYIaK0RRGtMhROAhquX57tCt+pI1o38KQX3XICadErF0eZd1pqguf0
fEemxh6LFkVoM9WeWh+oVP5KLe1UXE8wEuPdNtwkCTRvFir5k14LwAD+WFE/I/6rxU30VlS8L+Vl
qQmprDmcEKvyyctxoIFlAyjKR3/mTPbNWW7qhYLslF/XTFp/zjUFau1OyLQoGG8Rw+n43FkE6UiG
K2TCw/tCDSdNq3ybO0VjR/Hyjmzx/htBrjKsXKJ4PeY/AZ2M7GlLkcy+EZczRdDjnTWaRTloHEyO
wZQQQqTcA0EeakslfUh3afm/+JGezw8nObcwSTOs3Ix9o6uHX9qbjDF1WHuuzpmI9ysZmVN3MJd6
pD9rwI7zAPxMVttZu+1QqStNuLRkfTgeDamQ0aI8ZvcxjXi436MdHkb5/FSS/AEYNgjBiTOgBWiq
nfWx18hVOcEj5Pjk8vcGnaRqw1gf0IzzwV1LOW0w1w2B9I3qD+EbkSfyBgqZ5+yVJO+S1bc5PZqR
vUb37CfxkeHiJD4vsyFbGV0A0K4c7qGCdysNCmmpvtYAOMQFXnh38UXxEuR17xaYWk8KmWx8SdHo
oqwgMId4mxf+bbrS32rW9a4Qyzsp0hjwxpX4fCvm3cFFPffUa9l02aXSIEx7dzEJggSvw2s3e0dL
7Szq5US+oDsMTDp7n03uaoYkhXbEzVDAWMFD7E3OiU1TVNdc0Bp/Rzo5yARFzZx2HHhT+tkNtJen
ot22nGnRlR66prOPPhp6MVH05BvmE7oHHOLkaJ34njzaejZFT7+leknR/W2siQvfpSVPphJQ1B52
526Vy8wk1htc4v1shb2P22E81na9s4CaVrY9Do1QZS87EphXYdNUe2lJPMGCvG6b6sWLnpEZA25l
30p5+sG2H78xzclmGvYIGvyNyX1FIyPg6B1Wk6On1qNYvK8vnjkQRYYzrjTXCw5NVG/I0IpkVwGw
CO5INU0R3JGXhY87EcV6PF4/5xMyHUt1oXFzmz0/G1s78LySHr9z0OCZ3W4FfNVD6lz28s7kA1b+
0Ha0YzNGO0HhtRTdTxuUn3qutEmJC1j+ti6U91+1jb4sJ4LsAQICbCPxT19+dtK66y4eddO6YMgU
RM5zeJmFl+RiPNmqIIouapp5gmDRpaT0Yp0zySTBuAfJEoB1QSi9Chmk19jFM8+05x1FwmJ65mbn
ZRoDzosE5U+yrsrtnCBOPPfyXk+v1ilZHuqWS7q3gTBicIMAQGiEhaX/cUnnI30lMaH3piEThJPi
JLhjrn+viyOPOGqDks9Zzqfv4Bv8zka8ZiCVqaK+nGATogilX7nrlp8/uPSnPrP9usXE+PfO2EvC
F2pxGU/2q3NIeRi1gStF0AI5oMuo5rGLfDj50s0lyptLyt//YDPL0ikJghN8YNfcy0tougcgj+jD
r5lCPfjzmDPHodPntvXDOFUFEDadwCVXMcr0//by7KCcsLyINHKQeh5CicLDXwCjTiJkhCk+Mg/I
G3RYXhKjX+eyUGzsrXkL1O1PTl/Th7GguJt8dj8Eh7VBjJhaB59lD0U2fTWPuwocS3xT9An0Thlc
0nMkk49PeNOVi3DM4WLLtiquwypFZoMKWrBxjqdrmo/G1h1ti62qMo92HheTDYnK78s+sNhy3cm1
Rc0ftCmZiGpXNgDtql54rSJk1THrwXAgD65+FmIRxjF0OlIkma9xjCCxrrUBnwIWo8Obha/RSxKd
eftSqlcv5crOWrejBpS7UMT0sLCtJDD+7T2eeBQ5HYdNWHf8/ejasWE8CoBSpMbASfWjfMQKSv3e
pDItk1V7UBq/hChxe1yRgkip+jt6/gHqyqvEqWXhaRNlzjjxqeu2ADnycEmHyRWJXMhDHc7gBhnI
NXA3BAtyyHVpp4l1xaRJdt5M7AfSnmna+Rf3P4IAAQEdYfnx/WdNSd3DdUQ4QMg9agKLudPVYrkb
yYiWCL5Oe99PpR6qzJye5/MxJc3XvpXlTdWJI64la7gIs3eUUWuA6OmN85GlwpckaabfjWsGZv5P
/e1dVUAuIPpePIO38tKWw02Jtql/VSUDue9mX/idgqRRviuBE4ItwAU4xL1vjIarUGS8bre9zwfz
bxmF6ydjMItGsurxF4T2W/IHZSVSXgHWzTVbNoGWnBx56zreUMmVjY90Xwj2iu7Qoj/6ggURYVVu
0crW7HXd3KyC9HT92uDMkK7Sia2s2CeQugvZ/2u6VgIZa6VbTGsu7dwreeJMlyYtDrK7tY/OwlVL
qNHARjyPimzgtqaFp8tGMwfztEd2HjCyJc2crT24T2p0vdXIYYRmWJmNEV1SVDl/W+6bQgb3dOI7
1uBa0L+6n33sgjxHmwWylXwnf9oPqYosVHE/cd7SkBZCWenqfechiIPQTocJ8kZwWuK++tqHnd1O
3R8WySY06+9lHX2d5cjTSunsuNxMR9dZjHhXpHJJfHus7airPFsj0+OyNHiJUPtIaTfPY4x1fHrB
RJ5A5p99pCQ7xNpAhqb+nE6CSTdh8dFGBpJCAZwx0U0OlL1cG6GoUsNG1fYE759/PmnfEzI15uXP
HrwiUwuzKTbC5x55AXPUr/XajVXSqLkTGnEnkPbotj0un3UGmxQhUig0oSC7ne0Zk1sVdpT9yCgO
AE61qEi5f4Si21gAf8fZ5eUKxnMWnRsWq62Bwfn7QrJd+bO4+CKNzi0MxC/XU7lw76S+oc5ERjqh
HmsVUPQLXDWxDWoTGjzFYXFOllMHU6f04KZFwAsc5henod6P/G3/en01NutmOyFkWv7pg23+koCY
fgvfnmdATr2ZEEgUYXqOhmArwKBOeHsaHlZtLqxpujyO4Mo025w49BzZkzn/i3YEbdi91dodeSFQ
aN77Mi9HS1CBBcsYrDJxa8caGICJkI2Lbrhd11BPjt3mpdozBQd91t3OZaPvDE5bCq8OMZmCbaIP
7HTvmlmuED7yMjpQbAMq21mn4GII3TYFTYugqRSqJ8DniPs9OttaVDOj8l8vWHmirLJ9lcJKnrFB
7EkV84jaPjw5nOWxzZXwn6ZMRgQ+Fj/Gsfy9x1tyaZeKeDn/HBmpMZf+k2PZ7qphRktenYoy9h/m
YqLV1QYTaFjRyiTiaThewY7CE0BFxX2I/KsHaqMiBGaUVbEWsAeaXfjr27GSPg9zEfN9PdOleorP
Co0SsQZTHAX/yPOo8GzO/KXNjsI12A==
`protect end_protected
