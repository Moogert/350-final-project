��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g������*���Li�ĉ�3���R�\��0}��N��i�b�QO3s��N��㐝p�W ��Kl]���BI숹�(�a$����=ZA��Z��<e�TrRd���t�o#��K7�QX3��O���� eT�2j�Ŝ�5�| ҭ��\���I$��Ng��^�i�cۣ
,�P\��B:�CN� z���� ��hc��GB	:b�[�5Rf���il��.Q��</4X <�Z*�Zv[Sr�w�P�����˘��C��\&�η��zR��bA�AE�Y�w��\�7¿ȣ���p�A
 I�!�C�^�@��r�>���)�<˱2�H>P��.�2]D�$aj����t�2�^���ɥ�L��EW�~b�\P)s�`�0=&�؆5������	���5�K�<��_+
t�ᴬ]vM��{���ƨ��w�M�8��Oz���>��F�}g���c.t;#��⽄d�>7��?T��i��P�tsT��.Ổ��)粜P�:�{�(s�QZkq�R}1U�=�[o1V+�x9�q�3$�e�6(�Y C]b��}�F":���`Ml7�\טJ�n���I^(`������9E[�WԠ6��?��/��m���+NcKH�w��z�1K���V-���X'*���d(�|���I�e�E,uVw��f��v �
w���y��cj;y���5s^4"0���є|a?��O�)����##���^�Y�����Rz�<��ڱ;�Q�]�ʍD���ާ�x!]��'E1rb(��Ĥ�סk�L?^nb����~�R�2ꢭ�h�ַ>����.�5�N���Q��tV�|�+	!����+����yX.º˦���'~T��7��%��_0%���L��7�7p�k�L�@�q:>�X��&�Na��)��������;���nB���L&N�q��E�B7���~ޒCv"���N*�X�!���j�@�V3�0�U�����~�r�B��ې|���)��yw��������yD��	V~l����q���K�Tϭ�vo�P�Kks��X}���s�y��X/�g;5ޡ����IqDGCJ�d�erOv%N=��5��O�Y	�փ����_���������'�����=͊c�tX�W��M�`���#�4	�uCN^�Dy�4�N'}�N)Y<�~�ӽSx�?�#|��js����-��ivT嶻m�;(Jŭf��J)<?��'O�*�.zWb_�%���w��r���MU��\/��| �����"<�-�HH��L!��(G���ԝ�����ȞC���}M�v��R@I���e#X�]��)E�T������A����
V��aǇ��FO1a�MS�:4&b1�+-È_��19��Z�3K!��ļ���Tm�Le0�w��7K�`j6�G�Li��,	n�ݬ2�9Cjװ��5KEky����IS77=�����h�D��I��8�&Lr+��m�"*nCp��i��#��!k�a���vީ�×&�'Ic{HcWnT9�'�;ui�	r�oᓄUک1o�d���b�Ȟ@Ppü�0�l�e!b?T��m�
êEP�`�c�8"-��̵�� X#c�zŀ��j�[Gd��Y�Yݷ��~Y�ɗle'�W�.��������'�߳?�`ٴy��&��{w��(ށ�aV�q��O]@3#���ZB�!'#k��1?�f�"A;&�FA��.�����_~����h�M���("���lX�f4�0������$Yk7�;�����:`�^�I���j��.1aeD�,E�ٓž�]`�Lp��Y��=�l�Č��Ԅ�	���3.˩0s_�ea�h,��7MG�+zИ�3,:��
���@ޑA������9��v9'��(��c�LO������x2�\IO&�pN�UVe>��8�p�%�B�Q/[WvbzVٌk�h#�N����/��z���["4��i�gE�q6�r2���2���G��ӚoH�Hi����G� g���u��2n~~[�]������A$�u��gKy�p��� ,y�4e�������6Ef�Z�l/��V���������`�E�/T��<�S�H�`�D��z��T���J$��h���|d�_Kba�� �K�s�fQ�S%�����u
ﶂ���y{ayY���O����)nx�T��s��ى�e��J7����ǻZ�?*��M���bdqB��2����s)Q ��kY�s���\B	���̂��J>�T�vr����d^�5hG���&[�!w�}I􍖼���Q�V�Zb
��*��bM��6K��7����ՊD���h@�]^u;H�l��6��ȱ�'��!zfT�8xT!������%S�*���Tʴ�W�z�-1>d[g��HF?�� ��:�ox������v�3��e�E�:m 5�]�%����ev�`�bs5О���SQbcV@$�|�rL=oϩ��
Hݗ$糑��U���yݬ��%I��1@�}	zl1~�1����.��3;9uC]����
���Â�"H�����?�Q���2�����d]��:�.ڬ��dp�菄e0�����	�cp���>C5��8p5�"$wޞ3������^�;r�I����t&Z_��o,K��V�"�øl+-��$͙�,+�H�Z��,?N�D�3���zvb��u1�W?4��T�껻���c^����J1��w���w.���]%���S��-�e!���t��UP��E�3m��DB反�0��)��|,Q�)�����!(�]س�\���x�f��A@�F[w}�g}��<Ľ�o�/;~ ������(<�B�Lz�ʞ�Q��{\�}=��n&��-�d+�z��W4���R��5�rM>o:��O�k@�{���
�W�gd^�%/�1�-u��r������.��%��R6��ap��f:�"R�m�e�w&%�{���S��`�y2JG>����>*�L����B�����]f���-����8k�f��O�u����j�! �:ˋF�O�6e�d��J; �1�T�U��+��!=&\��A ձ��L��7�/m�1��� 5I�|f�;�}��Q�/V}�7S������h�Bé8l�a}C�]�dR��]��Ko��&VP�V�wL# ��W$�l��{PO�s9�ͤ=����� (o�(~���f��/�T@k�O���D�|�&c+���ĜL�K�ӰH�5�)�q��͡B�a�R��n2V>X������U��R�3ݗ���j��x���e�i�0 ��
KQ�\���މ�����t���3�@�y7�G���Ӑ�4�о�e�����`s���?Kon\X���)Qn!~��fsb@+t0��1��D �^[�гE����^�~�@�Z�_�\���<՜�B81	�?�@w�f0���{IX�2y �4��	m��v��z�j�%���j�� ��2��N��>�~�xh�~ҽ�?�+�p<�(�3ej�XW��CȮ��-�}f�����Y�E����k4Dz���x�Z�b"��[;�:9Kt�O���5.n0(p�����Q?X�0!#2C�ug��ͬ3�pSK���dz��V��ls�=�Y�^��� V!t�C�f*9S���PS�$*(ٿ��J;�0����:}J�ɻ�E�Re<����@��������sZ���t��؄�{Ě6���lR�hb/�b_�����7�ʠ��
�o��=����>g[����
2)�̇h�*�-��E�QR�F�#�n5)6na'�f�<�p�� ��8g��/�V��*m��ý0�W�)9��Ð)A�E	|��+�1�i���,���p�3<\GM�� ��I�_�x!�O��O/�b,0m��n�����۪Ӌ�h�S�M���`�}ǸVMH�
�G�1B��dF�6/��5	���Q�??��9}�3�K���(Ʌ��[�!d�+��gv�C�S���=$t�ƿ:���f�{�ʺ���;2k�w!���Ŷe雑�� HT�J��\5��B-O��J�y��⢵�;�&��QF��I�����,wy=�K�-huqʩ�M�	�̼��=�^jO �:�ƙWZoeY9W��e�î��V����cG�YBV|#�n��i 6�}�Z����%��;�@�2�w�E�X5��L1��WI�w!�*���9���;�(n�|��tU��%¡�R��`�Y���.|�2@b�M�C�]�첰яE�5�UX
�ur��\�W��@����I�)i���~|������h�ެ�����O՗Z�ߑh�N�!���D�mF��A�����JY<�?����9s%��V7<(YܔU�R�h��x���ތ�\o��V<�6agt<��3����b�q�';>1p|[�,d���:�W��4ѹX�BW��AhI���M�w!4	[J�y\�\]�O��vI+[ڇ&4d�,h�]�C8��K���)�N��=)�a�E�74[��?[�����]�kFշj3�<tW� <s{�JT���o�f+����p�݉Yt����h=	�߄5���%���J������9��w��ȴ�LOn����]�#*_�"ۻo�1k���^��"�$h����kv�m)�o	y&��=��H)�����۰I�+ȵ�Q69���!����OyZqV�	�<t`2=sG�����kAL��+�
�Xy1�Cl�� +Μ�%���]���2`�,Qy^��~	e��\�Y� ~q���j��tل�J��R���$�K`hZH{�{[aN�������tv:�Zr�&!�����6/�NB�7��D�^��ϻ�4��g�l"y������t̵X
�^���O��������HgS��H�ԈI�˯n���t�>w1��P�I�*P�SKM�
�O;�FDI{Pe���H�.�)��b_���w5!�x����qݜ�� PP�%��\� ��i;p�,n��R��z�ԕ5h{���XS3-��>��v��rL�7��0���'88��[99Y+��c0�U�{&D���7�Қ:�+����1���QB@)��6,#$5D+OG!{��*�:��;#4O���^ʈ�����de��r�%�O���)���͜�<��J��ԣ�W�oд6��ɉ���6�kͯ�g����%Q+���B�X�n�y��D�}R����:��6W�C3˽ĩ��B�rK/�V(��72�>=� c�uم`ͮ�����j�l���鸽^��^ŭ�����,���R�c����N���b-sz�s�|f\�����9ӽ)�� ��IZ_��+��A�w�K��p�3�P�P�F�}z��^�,=���R&~Mt�̃�-��%eRǏ��<礚Ke�s@��7�^�U`E����X�/;8j��RX��I���5�k/v+T�œ�t�G���ݿV�}��ȸ�R�A� Sr�#@���a%z���,�mT��(�<>�,�'�}{�#�����[��u�K	u�OK���5w�����'��o�C'���T��C`�!
��E�|Uq9��{�6�5Bz���2�3 k[!����]#Iﴻ=O�'���Q�SRq��i%�ό�J6ov���s�Q��g�R���1�_2��Q#8r�y��	������o֥
��R��>�V�jJ�V]D����V�~�>��.������Qgl=��ċ����"�ʌo�
x�/�P1��m,��:8W9(L�T�vUi��dF��U�Q�_�U<�����攥r#�J�Bb�v]���h�{D�
R�g�6��,���G�ο���i�����ٺ�lc	�O�伎�B�m����6+ɦ��0.\�g��4�)&n�c��-<;�#��P�9�V�l`x�+�ɫ���eFo��au�?v ��.�/�g{�/ж>B�rUN�F;u}Q��KK��<�SF��ѓ���N��LM:�2�1�Ұ_�DY |�=j���?9D����8s�˭�mGvz'	���q�������$ft�,և+�����5w�D�SX��u0��u�^��9J�Y���7��) �:����~
1�â�xf�|2\e�r��Ԏ���/����|�զ��D�M>תW��/�����9b6�R�$�LY�(��,�p�@:м�;���6"j�%��^eH|�(sǑM<ӺW�&#�5Z�㡞-��W[�@�w+���4�L��
xy\�:�X��ִyݤ��g����U�+�Õ�G��A\:;��! &g( �vT�ߥ�]��b�k��0�-���ke��3��ʧ���.4 =��o����7z���_�T�>~f-%)R�C%��D���(/�����P�͸u��R4L����P<ʻ��J8��	��J����:�͒x��Y��U��m�W)��$"�(Bj��<�E�����A`0v��vޮ��l�f���Xz����L:�fC0�Q�	t��u%��rX�(��5��H�]�F��oHt��@�x���}�$t�9�����21b4�B�� ŏ7�/\���\�E��;��c�GM� ��3R?4��ρZm�m�H�әn�b���sY��(RF ĝx�|�K����a��=���dsR	&D��!uK�p�'���E.1{�gY��P���K�W�v�|�d�w���X�q+Y�t���!/ŷ1���sp��dx�Ј뚈?ɵ��ӱ��0�G��������H�2��OM&q����~O\�laB�8R7+�|�sTjaɺ]1�1��x�i:eo�2�k�mŦ�@<�����ˣT��1��%4�/��w�=I��Z�(�Jq����|�O�lZL9��xh�}M���k]}���������}(��L�2�k��C�W;�b�ul��}��a�З�G&�&q����0˂��IiP&����2�5E�q�M��u/�Q��6γ�ZU���X8�ב����҇Te2����6"��h	uu�(�I�n઻�/8��u�GF�#O���H���0�Bx��@��B�j��4+�'$ah\\�����������`�@��WOE?{���}�Av�J�SZlOm��T]kq�d��ׇY��b�T,��a��ǧ�
�#K
�i��Z���D�߾��N���W�N�U�6:Hs�d;&g�$�6*����Ѿ��}{�ԆvԤ�\5+'�jw�rx�F	���Ӈ��^�y=���] ��·�<��ڋէ�q�9L��� �D�j��B��m�J�Bs������g$�o�(?Mw���PFn��������>�v[r���I(㐐\��
�q�S
0ޗ����4�@9-�&�qCM/����,�yD dp&l"�))"X���G�<��o!��l۹J g?1�����0/L��/�xx����+�z�z�|���:���S�pRE�G6 ����IL�O�0��v��"RI��h[)��^����Z\��w:��7Y�	0����3�C�d�p}�tӎe�CmKJ����5��qk�����ة�!X�v ����3���3]������&c0�LpV)�y� ms�hֵ�I����ù"����桢��׳'�,)����5�#ڑ1 h���B���^iZSܑL�9�?*)&H�b�z��V��x+��/�)c��m�K���@�[�o]9K�T)�ʷ�Ip�g>.�qu�V�E�֯`�4'�u�b�x�j����%3�z����]י�튍����b��W]܎���E�X��"z��ZL�A���f���~�BG���ä���L\����M��Bk�i���M�*U�b�S�Ą�����[�R\�������N�_�c�t�&�M��gx\���^P��3;���H���4cu��I�.�'���%� u{DU����㖓o��ra��X��.���C����n��0m,�8g�R�_���KZ"��c���B!��w�c+�f�2E����i��pA�KH�a���������P������T@���|4��	e4��LSI�3K�n=��r��Ʊ�8�+�|�T�x�4��pZ��*��Fü�������(�(	u�*�3�"2��A�_�\���a�+�8��ij}4��M������$ܝ��*���P�����ꂧL�7�a[�%�F��I�"����L�ըt����堿�����CQc��Ni2�Ì�r�B�cM.a����
��ϭ��<O��#�Z����4��O��z����p2�ǝ@��a�%�Y�K�B���M�����8�����t}\깱�޸����RE`T��Z�m��0��%��}X"T!��Z��YYu��#����}����M�WL��Y����o���)�B�ˋ?����.�
Zὓ�N��J-���~'`�w���Qj�X��l3�|+iQw�o�r�� E&R�[ԋ k�ȼJ��C� ���(�0�=y����bqN�RN��Y n�A=�]��(o�
��d����ldH���c+Sb���\�E�2���X���g���A$BJ���L�Ƹ�E�������[�&|���h�������S~s��;F�o��^/�8�Y�������f�ۻ�ӹ�
�bo%ᯌ�u�B�Ňf.c�̢`�6IS��כ�2�X�p���z8��A�<J�٘�z4�����_1y���T����
��L-��<��(L��geV�ZYw���ܬ�#��7��-�W~z��&���fhs��`��xV����sP���Y���a����!��z�r%�:�����Uy�ۄ�����%I��z��5�|_w�;�t�_Y���5�=ǧJ��>)�c�g&>�q'&l��]��	�(rφ�H~4H��|�~z�ob���b����YQ����\<u�e��}�n�I�S� ؇6#B�W�>��Z���z�D�*���	��+�l��i�PrZ5=W�"���zi����1@���b��cySR
�������X�vX�j/�X�N�4<3��V8�,�?@�@�E���/|���q�B�Z�&.�2f�9c�_���a�RK �i����S$�<���6�HO��
�&�Ҫhk0>���RH���N&�\T7م���	<1*�zl'Y�O��Ԑ��N�}��ߥ�# ݃�Ct3�+�L�(G/YM�,��Ӭwi����ݳ)h/�Q�b���2��
q����M������o������}���}u[Խ"店Fq�N7i�	3jWx*�qāP4R�C,��mZv�,׭����֭G�%�7Jt���� ����{�	v̚�m��,��v����u�M���]�����;�{ư��g���Jyy�3��Si1v��"��&"�-�D�ˮ9�5@���������v�t4�H��W�N��P��n��_���r{��T����g���3�T��i�I�;��K
�?g!A�f�B���`�/_�CWa �;M�K�q�����ū���Otm��3k���.	�m%�~�֣k��y�y����ٞ�w�̼��w(�Te>{�npܭ�,J��t�G<�S9���u O�]K�dUGZ{65[j�a:�cp2w��G!5�P;I�X�ڼP�{���r=Bb��n��MH�7��]0��,�����y����z���@��I&Cs 5�:��2�|�E�.��x�2���6!�J)��A|KV�[>{S��ܽM.m
�h�n����}�pn͕��j��(0��H�Q���n�Ưj�E����\{�/Q)O�琥�g��!�c���f�(���{3��]������T�}`����͈m`���}Ϗ*��Y�vŘ����:SlL�P�Bx_����(�`��o�9`I��S��`6�
�;�:�东���}0oi���d~� ��S�8���H��B����s�݅4�鐊����3�冋D�>FX0�t؈ �XG�i�~Jq�b�-��P�G��z=g�>ԕ��#�>�������k5f�0�F��s�܌_�9���m��jX�\�N���k�U���鷹}3s�JG�L=W���W�G�y��	M?p�x�}�&y8�(C;�c��g��F
��Iԏ ��G�����[N�AC��(�|X�}eX�D2Y���Gr�j\G���7��$��Bm
�ܬ�GDP[b�8��I�G-k<f�����e8�t�7!�t'���;;'�Z;�en�Q�V��u�CfF�4�-X����V��T��Y�����%y>[~{�� �}��Į�봫��(¿���m�;k����dg��yo���V곳d5O{����`N��|��G"�Ta�FƬ���ˡʓ��r^)P?�]�����]$r�wN~#Qc��E���0ǉ��ݥ�iq�E��R�5>���� _����x����(.Y��8�-��f2����'�����y fl�,c��E�ޝV�1�i���Ί�����;Q�HFT�9�u#;��鷿�d�]%���������}��d�M�_��8_��Zn੩�	�3���G��G�F�g?�ON��I�ð��}
���g���"��i�1+��;�������=�ʣn!��-��#��K=��,����A�������5�_�γ�Q��X�5Jcs$�o�N
	��#�0̩_g�z7���Ĕ�'s���=Ah���Y������5�.�\��E*H1 ������_�<�aC�Y4�՟�� N�d���vG��0�
&���J�8) ��|�DW�oJ�,;An���ޙ�%	ZͿ ��gܚ��t;�s\���j3�V�k��hn��
��5i��v6�Y�E��|�aE�E�qeH͡f��'c�ھ	@�A=w�oW�`S�+%���?��H!��lV������ʟjs����3P�+��������_�$�\�2a�P�4��'�x�?J�y�}���D��Bn��_~�)�'jkrc��$NS��?�̻W�]�>F4�ޥ��ݹ�W��aSG��X����vsVa��R���X�X絭+~�3��{��l��K�MU����S�뛙'FXzh8||�l
.�&_C��!��'���%�02��d2ԣ)�/O�	�c��G�AO���ۀ=sQ@"�+�� �3�����6׵<aͲ�3oǯ��}��F���K�P��s}Mw{��^�
�$�͓J Ng���6�w���:�����4�Q*��иW_�[mrO_��L�Л�����3s���M!*������X�Z�%�����5"^���`��ms'@OC,��c���5%�O�k�
#d����aQ���Rz9�;a�tތ��0��M�.���u�-j��	�t"Nm��n�Q"L�#tQy2�)����.�:7j���ۅ9��TX����p�<e������I�<h��W����ٽ��u|�O��^yt��M�Z�����~��"hƝ�+P�;38v̍Q�����te��(��Peec�Pz�-��>���>�x���l�-C���*���5�� ��Xi��������A���R�\�/^�)ڸ�5MT����M �u� z�I�Y�AM/
�Έ�F<�/�}� "����줫���/2[2��.t.oju�H��R�`�y�6�Ml����k��m�����fP�CW��6/�o@�����>���f/���Xo�QĴ�ْ���Ί?,j��~�9�g�[a}A�7ߊMr�#c����y��	��<iՏ��0c�T�I[��� 1챋�ǎs��M�([�:.��t�H"��w�H�93��i�5�[��|��2Y.�ɷ��햗S47�8E�];��?���\�[㘨6��?w&i�PZ�F����%I0��~��澩u�;8�I6^W�&E)�grH�'[��
/?�N^��w�A �x������f��R�,'�B�gD�s���j��/1?�n��B,�{"i�(����ibP-���D�bI�2|�G��>�TH�~�$�r�:6!�R>��\�;b�d�k���گ�J�O%H7йwZ'����sniQŧ7ዝ��4�e��;�c�<��� "RE�DwB҅�m;jf��}1��
g@0�x����Wr�����AD��q�a]��2�^0��P5
9~qz���<!���]��w�]d�#ړ�@�K���� �F��l��}.I��yHo��6�H������o�%:�Y���ku�Q��.����J=]�o/KO+�����`�^����.��ѕ.*锫�wA�M�Y+%t���yp=�eBe�3=��/�Wg���DB����	D�3���U��\(�i)N|'e�H��	܉����X�K[��l410Ǜ�'h:Vpi&�t����_l��nS�Y\Ͼ��_�FM�a����Ҵ$��0�ԉ ���'wY�0 ��h��pg<���4��o����Q(�y�?�p���*���/���Jճ纖[ �m%
`�e��+a&I��;z�!���iD�D������*;�w�M���,��` /�[�>sHm�ˈ�j<��)���襤��e`"���)�Q@�t�g$������ 
eG�.a/�X	j�/����$7�C���E��g��P����6LФ���փ��h��o/X֌qb�o��˶����u	2�r��Q�ƴ0��6�7w�WBoI���Y+��;�gzyƄ�����	��t0ޞ�ĸ. ���FQ�U���cX�ә�2�7��پ?��@�2�lj/_YV���e8�L����(�����Ib�&��� �����^��K�
��	d�P����	"����W5�dwm�8�_�bȹt�E*Rv�P���ɤՉ'QvN��S�ӹ�}����Jz��łe�EPv�4�dZ�X��^��@�ķ�*5d�2�X�ɉ���?)���Wi�IG��t����� ���3�����J��$(�[��M�["&{��/O�e](��Ӱ�� �r����;��\۩�ŗv���Ny��	q���*dsjR�y����V�oKXdc.s���&�!U�������RU���}��(���/�D48HG�l�y����[%��f\�D�_�ko'@�Fzg �ϓ��ۢ���v�)�03%1[tI������oԖS�K�PQ��St����ʢbHdM�����cI�$_�d魐�U�D_�{Q�!��k���c^kԊ��&��c��LX�jTJ����cȌ~�Fi���,?oS�+�H��m�k׾eӂk�����492����7o�:�c�ok�:{<��L<��׶⥶��"��M�~h����r���;c��I}n��IG��fh���"S>�I���޻�k��ŀ�ڰ��Z1�u��@��`�T�́s3��x�4û���\�wv4�7!����1?(y��|���:E������5��}[D�Ot햔vn�.1ի�#~
-���J�ֱ�~1�g��1����LZi����Ltw�8�ۧ�	�p�EY^z׻�J���چO��i�����&Z���v4����~l�Eߥk��!?d�4�������l1����b(�~�$����{�?u���
�
�z� �
=��� �Ib�_��b�#1	���h��?C����Z�;��հk�~B��3�4	�e��szN	H��/T2��'ܤy������g����K6�j�?ѓ���ܒ��/i=NX��'�h�F��H���2F\G����P���q����A+�R��
�p�6L�����q���璬(��_,�2� s*Ѵ���F>(|D6���G���x�٨M����yN��?�A�-<F�C]-��F�z�L���SM���k��wk�׵]���cCYX��xi
��>�h��[�ԖkC�p,L�X�H�u�gȈ�X�k�����枮Ue3���/�������7ei IZ؊H�����=<����:��&og�/^����`̻v:����Y�^�7�
�"��	�5�qt�)��`	ak�bO���oVj�� ��Ë��Bk�`����a"	�/r��H6�o��I�I�W���P���L�ϼ��M?��=���"���D*�X���PE���Zۚ�F�ʢ��P�Z��X�!�.,G�[C�ۙ���g�;t��.J�Nʳ°C�{����� +��/��c6�;��r�A���p;��#��8oP6�`�5��P�:�&��j���@�=���8�yƽڠ��RZ��R��T_��L]88�l�Xg(�-F�	�;s)I��%��)�1(��۫� #;��%.m#��E��TR�K�p3��K��zƯ	_7`J溧	�Ԇ�H(f�>��鼯����1] p�4I�.S"9�z!����z�I����\��sv+!O��l��ߴ�����M�i���Ou~Չ���n�q�6���Ֆ�P!��r8�};�`E�9Dz�+/�~o̤���`ƌ����m�D�>]u:̍:��C]'�k����Y|V��u�w8� ׾`�M���}�
�����_�oJ���F9�Z�>/���ÌĎ�g��N�TȌԼt22�eCE�;DT.]:���v�թc�6D����~;z�]�?!UMV��.��!W��βd]n_@x��9��5�!b�Upb�s�@���&&	.��P�>���
n�~eo:9�`S�(cTO^s9����pd��d~��p_e�#, ��UɎ`�֖�C�{)�u�V��1�]8ڪ��/��5*�Ƕ)��c�� �og/�G�t�-�"8rB�����w�+�^�LL�.��%�*�-Jg�>L�9�����Ԏ��T�h+�ӆր�>
��x?T=�t�7��~��7��D���m�-��L�"o�������HM��Ed���Xߢ!��h��Y��Кǫ�`��?���Ӑ��8�+������T#�e�8Ft�E��+h8k�T���� .��( v�v����Ȭ%r2aՙCt}���:�w���oN�]�1ׁ"�~H��Vj�j" D���.����- �	U�2�2��kG��~�>�p�X�!����m�}������ۛɂ�?�������*?Y�s��Z@R��V��	��V�]a�*��7Ŧ�㶯p;&�3j����$1f��#��bS�yD$DFڮ��tYJz���[��tZA�F�qo����Ay������̹/�O4�K]z"u�t�ӼX�^��>���枟��n������p#6v�֐��PV�,���/=0��6X���t�w�P��<���h����*ʖ����H��>��0��,CAӦ����)s$���C�=�_U�����[kS�7l8��,���\xb�A	Gn��L���)�'�,f��	���-��M�ݴ\��Z���T �Mt2n�@���D����>���dy�L��L��'ċ/���L͌�vf�+�<ZQ�J~b���Y���D��69$Y��au�d1��h|4�(4��1=�}�oȘR��pSjQ"I/0>Z�#� ��`��li�]�d��.7�����c�a�_���	0�0֢�x`���Lq#���JW�}�g!�J�Wl�'Z��ٷ�j��*d�A����q���,�W;�r ���Jz�c�!�n}�pl������<_�,�)'Ж� y�-?�J�� #�x��?��p}�/x	�����§��l�>Ue`W�5s�g��n�[������i���^�4�`��}v�	p�Yg*UaΪ�L	څ����W̿�{�R:���} Q�XC�~S��} � �\�'��q�$e}��XW��b�hot�ӛ�uQ�{p<:i9p��l�� VU]� :�t�jNz� �H7B�O �/:��*�D#ڟU��ڥ��&7@��&k[��<>�~$�����2�%b��:��(X�7�>+�J�}�_�܌U��VdD+�y�_6b����s p������Rjl��3�C#��UA��	U����,!��.Ub�3�عL�0Y,T�y�B�_o�_F
����6;ё�tY�J�s6����^�e�\N��)ښ]H�20V��NN6ZЖC]09bN�,%L�7jA\޹��]*���\���B�/"������f94t��Z�,�����p��J��|��x��L�"��J�7�.,�m'>~*�; ��ǈ������jD<��8{6D��f1��z]Ԇ�t@�lӵ��� ��%&: O��U��n����}��wsO��{�+�CC�Q]�lY6�i����^�u�h��cn��޼#�iW&�&0V�~�D�7��
o����H�N����C�oL0��^��wu� �$��.4te�e2=0�����{�'\���҅�bu�ߕW��Y1����R����Yu��k��ii��Iy-��#���M���I�vg�ߚw2����j"^����.?������/z����&�48ť9#� �����u��W`��;a}�9��9ԅ�'��_�ϭ�YO���!o���}Q����ALF����o�\�T�z2>�ɪ��f5�'��V�t���u�Ù�Y2,��K� uO��O�zt�>ן���	�Pk4��;E��b�*�
�fR^e�����a�j��le�҇��S�Gܳo��Ry"�.��(�4�Ȏ�՚_�8��Rx݁CS\֖���>��y�lH�[��T������1N�(�S�Zue�� K_��:�)ش�����@���A勥�.�|�A �����Q�RYP+�h!�Tmٚ��E�.�����G��I���.�@a��e�8����3T:z�y,(Ĵa��E<��MDI�af����RbS�6��K�cs��?��S住$�f��׏��i|�	x�f���)F5� =RE|��H����^@�������L97[Lw�x�����[�k��4���?��&����|�r
�	K��'���_vsm����=u��¨P�P��&��c���9Z�Ʈ�_(m\m��J��<��"�0���s���BQ${4���c���M�o`�	��Y���Gง��ONx<�тG,�IqAEt�rP/���,$��pZ[�<q�I��X2��8�m�w�������s���#�PKT*��Ԥթ^㕘!ц.���/��Mc��G^Z�Tg���ú`�!�
>�Ӆ��B�V��p�C��V�f2($��x�c�����CoҼs�(��
�-��ݯ���J!�e�_Si ,q�eabo��GpQ�$^�I�m�K����6��DhOI�7�r�Q���FS?��]�k����s�1k�?�xs^4��IG"Y��t�k�nj_�`1�G��Ț�|���-��"��҅S���މ?��>�-����L�B� \}	&>��m�'�����(3W���5�_U����4A�+b�R�C,��7܃k�����Ԏ�n���%�n���*(ʥepLd��w�n�����@��<������w��L�G�E֭�j����u���]����|�u��8NVf�%'�3	q~A�O��c��%/�Eb������n�+���-����$����z�DH-�fi9���іٍ�H�I:�N�D���@�����[�	h;%F��k�LW�:��`v,����M�[�R�V�F�~G��W):��ί�W늮x�k���G���h#�$s��[��C櫵�����n�nEF�`d��B�������q�����/X�,�Ɓ��%��Y-��L��mJBV��c��:0u��2]^��j
�.�"٩��4C��oh(A�����i�e��3+��\,ߟ��r |0���b��?x^�R��<3��n�84F�&��._Y�Ep���ѿdC3���m���F	8��=�!�s��X�X����\ߵNu"�&_b�٭T��P�(P�2g#]q�]�Za/й��n92�������Y��g�g{��G��"��%�͐�U�ou�Nd��psҨ�AdC�J����W9����dE�eۙ+Z���U�x�x0b�4�ސe+�zn��+���XCk��E����
�8{��*N�ˌ>{��#�c���Rj�O3%������\���;F惞(Ė�C�,��J�K��ݲ�G�<|�����(�w��Xj���t /q�ɟ(�����Ц��O�]_�������~�l�/B�bP�9�G#��3�\^�R�Җ�����h��-�3����y�s�_t��^wX�=�R��_��'�؎T(��v 	��#(�da�/ ���M<��Y>�ޑ �#��+��c=�C��*b���G���riyJ���ޝ�H�˽Juq��Z�j�a���PuT4J��ζB����y����	Κ�6�F���		E!��3���2%9�\�a����}Qs�bU��ő��+�m:�f�=�L�������	DO7���U�2�Kr�	�1��r�5}��	���x3Q#�3���GA�N3������	��iC����l�$��.:(�}�@�������c�+C�ԓܲ%��u�UtȄC��� �w����0;�+ơ@�x2�����1vr.�#���5�h[?�r��J�,L+'�d��;�sA`�ɫ�*�g�u�؎���L�Ϣ�.+�F�dȹi{�}R*|��*��4�/�S8�kI��%o�m'�<��{S4�R�<E{vq���Wɰ� Ze�5��(��_%����{�	^���J��&�
���l\t������m�J
�0�?�yRϤɒ�-�G�aI��� �Vz�cK���9����N�}r�1�0���M?8�x���!ָ=*W-�ȸ�^�]-)k����� ��g���p���$�CR�%y��aΪ˪Q�OMb��k:��#�\7�V8I(�xaE'�AMy��a�swrj��H�-l�t�����F�������>e��%M'��+�D�0.w� �[���`p�{�Q4�d86R�.3B�v�`0(%v�yn���$�q�j��V�cj}��'��^��l���S�� �7�K;[�$��9p��x O�ܥ�����ל�Uv"���3�,��In�:vB�`48*�d�7н���u:Q��h�%�GQ�'�L�H�ŋ�;��B�ܔ��IV��Q��mW=2 �+e����M]R&��:�нX��]�B2��[Y���dt���'>}�r�b�)��5��m���A�q=�	�d�#"̖��d^��8�1��Ր��A� ��4�6��|D	�X�|�"�.��e��9R:��XHin�7�Y~R�#3Y�fB)�n�/�sv��w��ۍ �!�?~>/>{�&���z���4TH�v�)�<��OPB��;��vT��W�b���XǬ���ďE�o9l$��Ō���.;X�z_6�OOn{z�|A,Y��s;@�yc�Hh�u�oZ�ӛ�4��r��G�|�O��:W9])0�-L{���B���c��й�kݥ5A�؄q�˞EYɫ>R��~93�e:�Y�S-�n[u���*��NQ�7g	'iOG$QM4�2��7|�˶�\����E6����4�}�������^�Ȏ߫��^N��77��
/����sT4�^Ye���!�Է����2o�K��~oPބ��ˊ�8��q__i�s���+@\m��گ�U�`�����(�dS'�K�@M>Dsp��ՖkYm!E*X|^��ڎ{����3��v���2:�7��������C���;@���>����$�� 6� ����|���g�K�1�Hh�v���(AU�_.��Ⱥ	�˓`���@u({�椅97�az�;��z��dGHp�`��ԯ&T���ڥ����Av��'�A��*�7���I8�O�kC��z؅c�zM��GjJ1y���)�&����M�<�O��w_*�i'^K�h4u49O'?/7�x ��ӃfQ���&	�	�
 Y���?���Jd�^q�>v�*Fb�z�'P/	��A�����o	gs�p�#�+��Bԣ�{�>����M�� �Z��+-��E8Kr���"{䋹��E��a@s�e����g�2NM�B��i��
�6���	-�����0��y>t:ļ�?��j��΅UX��c��p�S��k����)6��o�g�� �DLF�����%���3c\VS�X{>D(�[��F3y�}3cUYx	�_-��mݼw�N�X!��L(K�[s��u&�f.j����0����:��0����oZ�>:U��u��0�o�x�ȧ�Ov1Px<e�Iǐm��9k��\i�o>�"�	+��%mI@M�:]؎]U�ڎ�<!Ex/1ntf�e��s7������[�m��������
�>�ž����]e�,e3��S�J�*�İ9��6�uf+���yf�%���i��U��M|����[(�����}��J-{�~`�4]��)�e'B��T2�*��d�q���`��X'���9��1��D�:���Հ���3�Ij�*�A�؝�*
����`�T��=3��x�Kh�݄g�����&��S���O9�G�醡�$=�V�]���s�ӫ!:�Z����<闙&���l�?��j���~��0��^Wk�w,�bȽJ$O3������ɡ�<�vQ�P����<$�ug0~����:�L,]>�>�L����*p����TF�1̃��s�t��������r�inf�HO| ^�������{*�iu�c���Z)�����C�#���b��/�W�hV��k�o��;o�W� �ͺ�=�o���V�
Kq7je--��pj����/3�;b����
Gci1,�����-jPf�M�q�����ǉ,���6nZ�������#�7XS5�@�����(����U����/?<4��ɉlv�b�T�8_�?��S`�~�4�(m�س�B�߫�k0�R��w���Ȁn�
Aʇn�>��H��O�|n�������[�O����b;�����F�(' ��]������$����Ŕ.~��]��r*&�j��:���F[���d�M��&�E�v�qn윐��21.����ɮ$3���.�_�4�F1(�|:~[9����lU$�sĆ�=,�}�u��g���n��o��MӸ�}��.P�ԓ���-�=]��g;d�* �"&��y梷�~�b!��VYQh��E���M]` ]�b��t�`N&��Hq2�~��adxkj5�MP`Uh@��\RB������
3��B%q��T��	d$���i�mb�(%.쪩�,"Z��J:bv챢��m�bz�Â��6�Ŕ�7E���1X����V��c��r�+8K��75`�g<Eڿ��$Z���{�]h���޼��^��3�H. �������7a ������9���B��[y��K�[�7`��W��?� �i^�ک�z8���\f'��+���1���̡!fA2]����:�_;6b��v�В�k�b�Tqm(�Jw����ڰń	&�a�o$�O�9f<T^*]�O����m���x��e��5��}�*o���(o�Հ��+�<�y���D�_f�ɱYY
��S���^���o�r��-Z	XK|�xǽ�[lɂ\���3i�O<Xe�ז���� ���[`Q�)FR�hn�T�[+>����̐�s�\Sl 5��5{m/��G����x�	�����`�ȎaV�=��V7�6t�ܕl��H�J���LrǦ�+,_"�&8Y��Ժ�X���?T��)�*��X<�ֿ���6���H��|�/m�q�FV=>��/�Ο^E+�"D��i�nk����n�&@�L��Ad�IB�?����,��o3�B��ER.8�?�0��C�b���0��22r�a��4��S����N
���W�jT�X۞�Xu�ɘ�i���c����xv�J�L�Z�|�Ș�����6Is�#�uT	�N	��g�R��O6[(���1�	��]�;��c��C��_S�t�����O�d��������vz(d-��|Ca��8ΝVe}9^E�-�&H�`vٞ�ֲ�rlL�g� ��xK^לA���V���lp�j({U:2g�b30wX��D��/��#�4 �*xJ����N��|����V�;G����Qz��X(��x�P�ˑ��?�B�V���8CQUY�1��%ǻ^F�.�<q&��=�ϛ(q��jYO��xd���d_"�t�3�W�����qL-σkD�.01�7S�y։:��TV������6,@�|4x0�$B�?A���%��L%d[a@�"���!�}��K5m�t�2}J}�E�k~Fk�]�7�p,]���bWb�� G0(��O6��=���Up����/|���\�\�����V���.y�����,�H�i�d�yn6V0� ���8��/��w��%����=EVB��{�m|_�U�����;����i ���P��x	�<���6V\AA���j75o �1F� �a��=a�Ya��\����~�z6Y�4���0�$Ŕ+������Qc�����T����fndT��0V��!�D�5���V�={u�c�$�-;�Q\lF��+����w*E[����P�i,|�a�EtD������n$��N��5{�cC�,R��z�D�āUd���߸$B�
 ɑ4m�c���f�o�0L��Z1fAlnX��Ԓ�@C�xO�n���A��]�D�0	N@p{P������c��$ըF����z����	X~u�E4�M�yOi���dM�w�:N���2o!pP�E$�*y[�u!��D��b���D
�鰞�#����Yٗ^�Zl<��1`�2����*��x��F�I�^s5[vBf�R;`ҟ=���vb��m��?�.�|<R�t�l=�� ?�����YC4�X*��~9�]��Z�Zؼ�� ׸�'�o���x ���/�uBIݴU�y;�Bt�V����C�����mw����WO�Z�U|���0��S�l!��<�T�m�s��d+Y��иzԅ�R�ç�;�&Řk���/�>� 5ku��])�n�|6���@�O�)���U_r�H�ꍟs���N\����Y(*5��$noG��kh{mT�5��^�Ǡ�ঞ��`h%*��ڲ�ύ��.x�E�%��ν�2�6	~�@���g�m���,�4R'X�aj��qM��懲�U������v|�z_K�����r;�r��Y9s��n2~UYv����ާ-�h��bF�x8TaO�U�E�Q{�˟��n%����4cР'�h8�B��:a��Gj ���\v1G�ԫэ��+r|�팪8�~IB��Ps3;�\&e&/��R�~7.�$'�6i�\nt�~6��q>��wu�����8l��(��r�w*U��G}�M��)vj��������;������cT�9��X"�����V�L��C����:�����/)y�!�i���H�鿵6��vN>�Ġ��������1���XA�u@����[�,�)�Jͮwdo?=l<?�Bj�sUC/��ҥxؤ�)'u�mQQ0=�������⠾��a�wo�)�M�i�g��MD,k�Mt^�)�c*u�8�]沉���Ѯ��b�T��Z����c�����(OA%���WZ[��$���/�ˈ/��b#�!���5�R,Y��u�*������ �$��h�-z�[ޚ-�? 2��ek XZ�Zm_fi�ً���K���b5�+�p������S����qx����_�s�����6����|P��;���Oܡ��J
�r��h�:��̋[#�4h؃��� ���g�jɛ��>�rj�	mԹQ��\��¦�<D��@/�=�=��z��M���W�<vQy1�7.��Q�n�,�gR�m�,�מF����C?�>~I���2�[��_�nb�t7�c�Sp���ɿ��1���A��x�X�`U\2l�i���z�4u�C�.;.Qi<�3���K�$���-��7,�6��W�%�	<o��{+� ��R�T@~��C0.p��*L�-�W?�x�L��T���tp:8�x�AVyY,%���F�W����k�F��I�/*C�� �\R�b
�=orn2X�4�//J7�[M	��O*#7b9�{hS��kQ_?����"��T?02�����6���-a2�	}M���=�	+k�ȕ3�Z��`쎈60�"�XE�W.oc
����{ 	�g���sx=J98W�����֩�������+*�Wn�Kϓ'��B��By��we��F��{|V����9/2�@�~�'�����7F���k|"kAhip��b��a�لj#����Ҍ$�b����4��ҡ`8�J�����E��WP�s7=.Ăx)��)��]��P*���4n�q�)�;g���(�go�o�Q���̖��/�lxho���CNӍM��{2ǪP�\�?��$8��8�ܦ���F�����2�34��똠�^��E>&-���}f�F��#ҝ��
�%[l��s���}9��u�r�R�b%!L������c� �$�)�_BJ��M����[�t%7�U����m�WQD���k�㋐��(R9�d}�n��n���R�6hC�_{�a�)��ɺ���^wĚgЍb D�ryÁ��'2�\������(��K�hH��G������;�-�:��
�On��<5W��� ���`r���U0�J�D�=�]V�S٫��(Ws�*���^��w���΋�lC���|uZ7f�U}K�c�>�F�^]�A0�RQ	o�oLH{�J
�����%-��&�׺E1�Q>���K��j����&�<*�=��i1��-O�i1ĳ��s{�m='�E]��E���J���| �@/�t	�,ڞ=���9�a=�͹~>���ژ�����߰~����d��O0%%�!�&q<��Itu&�����TP0��!A&�U�LFpq�����Ƞ��e���B���[We��B'�)��lU1x�� ����6v���-��)�`��O�0aeצͤ�BG�2��?��nо���z<����%˿�ɑ�9�u��#�{͊z
ש�%��`�+�~�������D�:�g"x��٧��xܒ=��7���_�$�L�-��iZxDDS��%��$уq<R�)����n+g��!� 9Ac��l�N9ga*�z3�6�[pq��pZ���bg��d/������y��hM�c�$�<Yڟ#U������.J�ڀ�����>��:�`k�Y�c�E#�V\șz{���x~��i��F�D���K�=�s�>1{_|�Ն\X�C�CZI'�;"���0���Ή��O\<�9j��;ޤ����o���4�"
�o �Q$(���$���|GM�<�8'L�(�z&P��*I�Z0W��MYm>�n��wI��H!-�ż��d�φ���5)T��թ��I�(��L�(�ȺK�3k�cb�38���������Q,[a+.8z���|Xt�s-�B�LK�=U���^��۵F%�Iuø���'�/4n���I}T��=�e�*u�΀����m��T�J�� ��d9���ܢp,)�G�����|*��A��\���K�5|p��v�b��)E,{h%Uf�ח���:��I�;�t ��+��̈߉%d�C����-�y5}��@��4����e�q�R�JJ�G�.�p�������K1��	.	v΃�Se��7/i��l��Wi�pڬQ�=�ʋ3���r��h��2jg6`!1��گ�\��i�a�a�=iTSl��<T}����+"�QT�GI,���Z�.���MYp�y�U�8)�HM
3��DĴ��V�>_��Y�'Ĉ��K��;����XH��'\kp��I�r�=����{ng峭@tQ����:�����Rxg�T���;�d�9���q�����8�zt�é������k=ؤq���ێ���?QjrAMe'��?�k���X{���9��k�/��Ѕ[}V�����XD���W��:���S��G���s� dG�vB��/5"~{�U���ݲ��u-=�LO�-�ڢ�f���+�h#��HF��z�n�>��wcYt�q/�x*[��懆�`h�Q����?K�|c��,�wV�S�K�"��Z�x� ~_�E��u_	�;Xԉn�јT�G�R�m���d^cǗM�9%�2o^�_[�3Q��� Q5~��e����Ԅ��ҧ��s;�8�Ti��9 W�Gζ�r���k��9�����C��RCV�q^��{v9(v�nϬ;Sv�o��S%�6�S	m��p_�[��������Or��`�G�0�]c�-=��j�ӻ�Hۉ�㚉u�m0��<��L�9� D���?	Ɔ��䳡����7�@�%��U<�8����-O�1��f��-��G+�,�[���d�s�w��7�|A�ܥf�}�,�>m��"�u�ٗ$:�Pjm��\l�zރ�] 0u0'�CN�^[s D�s�����0��BM�o1y=�x=m}����8'S�L��4�����u�+�o`�}$����&e�g�2�{l�R�ى f�:���i52!�{>o] �J������:�&ͮQ�l2r�`��K��П�ܱ�� �ʟh�38�U'���L�l��nG��Xt��0����m��`�����O��Gaҋ�,J�]�&x�J�1n���KK|.�6w<`���� �5a��/o�ܻ�b�uɓ��zN݄Ec�
~�p&�E=�I\��ȡ�5��
��b)8~���r�������q�9��"H��f�� |Y�R��ӎ��PS����iR����[á,%�o��"���qD��+�`����[K�,�;D�e�V�$!:S �e��Lw�`N��7?�׶�t�`�����M[)G��hec� ��F�P��d.�>J�i�=+�OT~��ϣ<K�U�5Wl&��0ȃ����e,���sxHϭ�*H����@ zCv�vy˜M"�8��J����R��<�s��+!��w�4�do�]�cP9��m:�Z�i�YI��-�~~��u��&RHN轀O�X��k�Z�����n� �#���@�2FN��"�N�߫w������cem�_]`��qun!(ɝ
'o]�P͞&����5�Yqo$���J�Թ�yq䉞�n��M��a�a �ۛ:����}�������X��E��16����_5�dr�p�Ԭ1h��(
���
��E����������L�jCN��К�&L�m�elV	�	c����M�!�8����/$"+� *{�!��i�����6UW�<�;�ת�� I��X�ᑙe�tU/L��7�Vǒ�[��r;�	������y��8��`�餲��)&�4V䇇~��m/[X$�o�S���Q.H�1���O�H����"��6n��f�s͚z�:]]��m�q�xM�r&?K���a�'l�.�o��=�>�4[8<�5�.DGѰ���i�o�tR�9������~W;�V��V�J&�1�r����.9�H�:�.���޹W����޽��B2���Ą��#u!��U�Y���4�ZQo�7����Xp�~�e��v�D_�9b��!��8�w�Z�rd;��f-��g�	�v�8���G}#Y ���~P֗�����`֭�������yuak�2M^�E��F���X=E;�H	uK��@|fM@P�u
�n-|5����H�a?&CdC���ۛ����V|r*��!�M�v��� ��%K���G��ژ�b�s5�F���d)��W3.s�<P+Hy�e�{¶��{����X��$T�|�����cՇW��>�X�/��;�&[z&sU���_W�߰7AT��`�� /d��5'� ��͔ѻ�����E�'�<ږ�_�s�itKM��q5��WKy�¤hTĜ�VO�+X\�֪ ̡���Y@�.�`h�+ȝstO��� 4�f��=�F7t�?���\��)��[mP�a�����E�dQuI���x^����Y�,�uq��A/í{�����[��ŀD���@�]�S��Z_��	�������
[Z��҇M��K��Tu����jő8��=>=^=�t�q'�}'��Eц�9P�TtAJ�U�)>Q���uwe����įL����R��e�Muo���[)�n�r\�|WN˯��T�,�OR+nQ��IF����K��j�]�/ �����\��&�ju�tjA���档OGp�[%�)ךھN��$��=�b�T������.4>�%[r�*Ux�"�ќ��[�v�/2��!1���<S�)R��L�6��̒���Q�d�@���#F���?��v��Ys�^��� n��+�������1x��%�h��\���C�x��.od��J���BH�ڞ�`/%�&��E<��<��3mu�V[�q�nU�-�����;�����֤$�Wd��y��ۍ���9#�HPGd�U�FTL��(���2���;��媤^�I�ZբL�)��@�k�R��E��5#�2��h��o��Hk|��`	+1����v�B�����T�"�oWK��Y�É!0[���u�N<�!�����O�V��e�i�6�k��3�"���%��#W��PN�b,ć�%�)��.�ru��b]B42x���6��g3���b8U�CL(F���7Шz3�����F(�����F�!A��!�8�R`!j�l)~Jt���?n	fഄmP��Ե��c3��Klls�G6}�I�?(�3[L|�%_ڪ|=���4� ��ǒ����O �K6}�LC1���'�F��/El$�Z@?�$��{�U� -KU�)}���|�J���O�Ԋ�%m���ھ!��xժ0BX\��K�o��T��(�^�"B�c�@����N#�h�	lG�7��&�V�/	�.)'Ä�����[B��Ƹ�j�J?�����C;ғˊ5a�6�if��8��pcO8�Fx��댉���hE�T��j����������W���_BS�T�>%�w�5Jc���^�\x�4$�t�Z2�m��xM'�ȣR�	������Hy�f���l)��?�l�%�.�Z�9<c���m>�r+,z��=�\Cb<����_9��MN���п���PaJ�h�6��W���W��s8�˽��{�yN����
�_e̜�L�~%�u�w��z�Q�Q �n˳�]�{�"��g���
[�s�r��Z+r?搰�\^���Ĝ�o����ğρL��/[�I�H7� n�p�3lP2�S��t5�󄗩=qn��>D�+��<�F#�R��r��[�ܿ���U��]�~�"ƴ�}!�t��OSS�b�3躥��"<�y��>R	o1��S�3��OѸ`o�7�>�ra�T���`sQGH�#W�"��[@�Ba��U�@N��s�4��W4y�w�3��V�s��]b'j�I���Q��`cX3���n�$	O���-��
;N�m;���|/���<IK�֚��$)�pگ�1�Fƶ�O%X��E�sg�JL��~� ������ݓV���-%�˪\U���H���� )d���tˎ�|�]�`k龦�����[�K���,Y��>����[�]�!bcȸR�*�n�f�75�s�.�����no��ۘ���T�*���U3�4�]������
wAM�����8Ĭ�����m;>9��KVQ���A��#n��d��E|��E΋Y��+��A�� X$�p�ݣ�|7��_�6t�� ����5�d�C���P�)�UU^�dK���C��یɾӝG͙�:�{)��&+(���-o���-�B{���m�̵p�{Dm�<��r`L�/��t_`��:�p�)���;+\)�'��Qt��o��&r2�!�4e�|�N��E��ٻW-3CЯl� �ƻAO��,�g'�'O-y�������8ƲÇ�L�:������q� ���'����ϭ@� ��������mV��]����B$:ę.�.Б4��˞a�q�rZF�L��k ��Gy���*�H�U�/�2< �����]d`� 7��ߪ���c�:�GGE��57�����!&�4�^#�T�<�h�A�$5o�.w�O�c�՞,���L�Ik��p�|�wZg��C��V�POEJٲ��:��>�B�؄[u'�����3)y���$Xt�o".ۼȵ�AaV=�\��Jr��M���c��';�w�j��EQ�(�4�����{;C�$5��ʈ�~�n�f�w(�{���rt���<a�E<�d'�u�ј�덝���e+����Ā�<[\N-��|�K�Ꮫ��sC�Ǟ���X����g�?� B%j���D���E 5I&ЊÚ�_��
E���4"��\��̅�@�]C��p���h���lM��MQ<�''��՞��ps뗥̅�	!j�\�ΈI\ܯ�мr��p��K����
XX~c,�N50� MaR��@������b��3����؊����8+�'�_��5��뗏f �-Ҕ#���x��2�v7d�#+՞NX��r
���f|���7�L�1�����
Q����?��g?�(��D��=���{��6����Z��V,}F��!�:�yZ���K��e��>4�jDrjO��%T2��(��9	,�����e�F�"�q�O������E�m��ߵ�g���^���E��������}�br��j�<#�����e�l�m�v�.�(�N�;�=�1�uQ�C��a]9b��p���c]��!h~XkL[��ҭ�X��ۯ�j˟f�3iv0�xRIҠl����Yt=��ș17t|f�'����5}R$*`OZ������+��9�P��������m��P�'����Vm s��L�
Ƒ���ř�aj=v���Ť�ᦱH��M�����5�Z�W��ur���"~}q�U^sU�k��Nt�0Z��F�tN�H���iֈ�!<k�Iu��Pڊd��N��?H��O�IF��q�Bo�ky-`B&	c�b�4�_ٸ`�`�V_�x�ߴ/$�
=�h�0;(q&�/����/&zs=��8%7l���5ѐ�<�P���ۡ����d0�����_c�G���޻�^I6�Taʨ��Vhp���:+�/P���!�E�j�k�$_����su&\�[�o��ԘdJ'@2���q)6&��	z��9y���7t] �_���>�~�nI�T�:Gi� j܏:M9���4�&>�+Z�����":�z���m2�}��쵄��� |�N�(Z/)�c�����E����gs'�Q��[v1ŬG���e�?�5^O֯�����D�a�b�8���y�@9;%����¤����<�d"+��^M�IT.�Q?�pޯ�L��>�Hh�|�Mr�<Vq%�7���aU}����b���7�rg�?��S���JB3���r�vn�T���DB���AOz�5�8��E�댺l����ŗ�a�1�rD��T���r�\@Gð���5��K�ϫ����6�	ƞ5��T'PT��gm\����[�5w���K���4>�M�YX]CPV�X�{͵����z��8�2F�>�T
�M�W�"�b�ɽ҂�ƴ1�ޓ|��L���ܕ��^��m	Vg�� 0�P]N�-�O��y�.�m�vU7;�Ox�J�ok�6�
c�J����\?�]S3PMnP��g���A3���#hv2Q�Yi�wCm������	�9T�����@���2RX�әv��A���^��K��ds�g����X��l�E���?,/�oKY�D�B��6O[�'<���@F0!��d�J���2�
O�K/"���'�����=�u&�H"�\�*���yC����d�C޵���
�� �W<�֬A=YH�1��"�]�zs��^U���N���5m���$��;�C%���k�A\����m����hi%��i�f�>� 	6�����\Ѕ��u��қ��������-1h	���|<u����	K�E��/��d�{�k�轄�m�Td�hg�Yu>�)Uw���Π��A��YE�tG9���@Ԃ(�
�O�8�Y�������hY(�S�	E��
�Q�����R<�I00T:H^�ΗlKѷ��ɀ�>�S&W�J�/m���R�dh�ZkJw�p���1�RH���t�.��>��{
<�.�0��a<y]�_����iV����\� �3遙���a���r�6���H�-:ev���]�9E�+ݮ:;��A��Hiq�|z�V���| �\Mt9���z�qV��h]Č�@�	�;��i��MR%lӛ���c�s����#v�=����[�b���]��f��O(���`+�߃��r8�à4цd�Q#�C�_u�x���,i���τmt��]��H�O��2��d����k�r��^B�A]v�4�����SX�āM�F�]��ʰ�L�����4��;U�=>�UgK-Gź_=��� �`�T�1�2�s'�*�Yt��{��48Ҡ:�x�\�����ޗgS�7��4�f5,{��Q�4t���V�rȓ����i����ޛ���X��q��Hx�)��uE�X0?��95�t��l&���b�F�K�M�z�D�%���Q�;��;�=�����
C%2GDQh��?�9��$��]������;�k�QSyu0�A	�<��;���ԝ��3[B���}q��o��H[�l�B �:���N
���&=N|����bN�$k,�8f� S��V/pNw�QI�9�S�5k��O+�,�.�i���4�i������� Ŕ )'�ũ��ytTT��X�7�
?N��䚛�m�
�������d�e��b�a��,�k�ˠdHoO*��'^�J0��B��3�} ?F�i��>��x	���%W�:����I���3�lT��zUv�oÇ�q�I��N )̋i�Rp�*{ �[�-4ݧ|�C��^�An��6s½���ļH��3lP���1_��@$������Q��c�'�Dև[�pw��m]�w�B�l�
ۤ�/~�A���mQ92�2���쩔�8�% ��&+�Q�J��K��/u�N!��L+�z0�ɺ�<�g�Ko׬���e�UX �ɳF��=.A#��`�eHՍҌ�#���[H6b%󣃣v\��8Si�tթ.a����<���^��2�$��+��#6C�r�����|��B�h�0�g�P�b�廏���Mm���� �

���vj$<D�t����$9N��L(HϷ�߲h��6o� >n�i\T%�_9��$�@?ܪ��-;h��U6�P!_�8&�t�7�V�=6WͰA��b��%i����y�P(��L֕��,ĠW,QP��΀��yۉ�K��w�ެXFD�CtB�W�T��ׯ�b�\6�و�e�k���)�ܚ?Z|�Eՠֹ���Zh�I��obT�HQ�ms��ŠQ���+c˞��~I۱qf�d�\�����Wg���`hl�ra�%3�T3����~�5@;���n	�gN�t��M�{[�*��劘�; �Ћ��:�Sd���9�9�TOZI	�Î�l�x�경�N��@É*�jB�i�Dڂ=dn�V�J�p�F���NlMo��/�� J>g�lMPԕ��y���?N�;���w�Π�+t�=9�`�5'�G�}Q�{[�s��J|�'q	���%Z6?Jc�fߎ�����@B��F�¨�Qv�"D�m�ܕ8��W���a,WH]�xX�啭u�/��;'�M�!4H́������ O,�TT
�Qe	D��s�s�i�j#Р�m����y�G����Jb:�]���1���#���By�3�h���Ÿ���&�ʳ�ݺ�$?�곑���;�������'Dmw��f#3:%�\��_�Y��;�f���b(��8��[�9Ѭv!a9��i���?�1ߒ�TU���bs7a���!β����v汒��l�����O�`��q#T���8�oN-�(�elBQ�2�s�
��n����[u����|yO��� x�Ԩ�3�W�p+Z '^���s)�f�����Ϗ�8u>�f U7K�|h��15�k��� w!!���T�v��T��&�u~Ao��|�ӵxG��$oW��^U	ơb�i7��3Q��dv=(;�F_�
��.*5�[=Q�ZZ+=�,����T�] "d��V�M4�4�hH'��V(_S����?���w�A�����<r�h�&�k�Z��v<H�!1$3*�w�~b\�����Iw?t��okuٿ����ׇV�ɷW-pj���35~�z��
f l���d�%��G�t���6C��ŴB��X-	P��z+"���l�{7'%��W�L����婫���>Cvn�@ҙ����U1��1�V�Ɓ%#�� `�U��9�0[i0��P@��׶��Қ�)�T��ޭ�<d�D��2�b�9�~`��%�Gs
Y\�>��ۄ�����Q�wD�EO���>2i�!�I�e�1�cF��#�ӯi`�[W쟮��ϐ�>+�)�h���N`��/{>CWx��O���FS���Ҫ��2�*Q����{0��ǝ�a�x���й�3h�asU��W;akiz��q}����'�Q�=�	��h�A�V���[�ѝP4Չ,����1�S0�/�1�4�MCV��RL�C�p(�C��������v]�ؿ�P���V�$P@3�%x�L_�ϓ��yˬ�ǣu����P���E��]rmi
ۛ&Do_4��Fp��|^�����Y�(y�����qz�DmK��ZԊ�OΗ_�&3�H^�)�i?���3�]Uð���:<tV��4 9�xF'foZ,4�y��]l��́�hA~�M=Ŀl:��*�wَ/��_���(�K)�RkF��(fáUy�8�*�c�ǸE1�>"����W
�=�4 ����Yq��3G��@f_�י�Lޜ�C�H���z��