-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
l1Yezcvgco0LHB35l8WtxWbmPfdxQefBHWPqyOh9nptBCj9SM7ik3uTKqgfW5W2pNiDWgQ07S+80
SxppLZtN2ds+gzHV5YcOpRBFifVQwZCQzQFs+B6zYzWha19cXyK2ttM1nwpKZGGgfUR6YY4hMGvl
/O5+iYIvSe3PA68z+kkadMqCZzichwpF/I9sXniLUX51ot50ldzsS89za5wg8IJ8v0rMoISWH/lM
3UBp9pggKwR+QwlMUzKcY8ZjBJKMfAegWveTM2i08qfd5o5LyVA+JjK9vf93n3mMajUddCIgHjxD
e7mf+0qgOKVtCubJfTzOWbKFh6O/pa8hJ8Ub8A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10272)
`protect data_block
Y5+OtLJ5UY+WDKNRquT6oMNmITnspeordbMYUb84eEGgIeFdUGQXJtunN7DSHtHbSj/9mi54UPL1
5s3sIB3WUGbzgR4jzSUIrRk0YqsWVwEeWoQtUllj599QCSYBue2FUAfvq9i9I04Ljm2K5E0GbKR1
CljowRLY51+iP6relnydTkFSUsCahOlacKl2Nj5ShH1A9t6Lb2Iv89rAVfM4+ZhLYIUBL1nP6zf1
uunVy87faOg2WIU/hAgIJHZVAAmh5BztAx7GvT1YZKZcFDedf4foiXNGxSBl/m/mRuxW50/ZWiBP
5Brw95G5B4Zk0ufzOkPounkDwWCRZiOOOgA+ahfgtT0NyhnYxrY05l9DhmqsKccO12rSee+ffM2j
PWay+1xxRQ9GtIEKyA7bRwK6SnPrlg4Z9k9UOswlp9FTYsVnhJrQXr+EMEO2wfIia//jusxJbN5n
J2IZZzr9COgqPD6fnXR2xQ/PefvzuuthFUxuwzIvMwYQ7okWm4h52ShrryiCAVjmBbDHR8ZtAINt
3liZT4NFSXh4gCskcI7NW1h9mX1sX3OwrIPJtkAINvlSGp8WOKylHjH+T/nK0nXFyuuEFRr0sSsV
FtswSJYjbGFiBQtiwZyt94x7gNYQdN/BqqKJ0F5jUMH6ldca0FuySYGxHMXFDanKVvqIxfPbe7iq
4driPSEzE1hFJJWPZG3yyM+2cE7eOjXgNvnTYM7g8JokI8xE7fQk3/6ItGAFxCHblTqS98FEed1H
uQOuXKEyD2P88MtqgeL3QPyFT413i+BPJiZx3gS4Py91QJu1KT4biEABGd+W4xQ/0ysO39dt3nd8
PIOT+NeVXbF1U0mxcgVUtRmz2sVsIfE7UnyA8TyxeAyqS2TIAc/NxKHZFcY/iDt6Bf78LDAI52KU
xl8aFxnjMFnzqqVxGo807verCXOR8a6li2C4IehBEXB9zCqYeMlid7thzFVgqXlNghsIr5qDYc8h
lBrvzGr7iHIe5Iau2MhBDFiE35hWXPvcbY1TnvyDUDPq2BWQEvEzn0KYPZppekD4PldjLKQg/A4P
ueMTA6wZMx0NAKJSZLXJBPCljF9eCodPKslGYLYh5hadOIxbCn235Z1nbsW2s/0sE36903jnhv43
2D98FPEAkjBHm6WViM5SKVOL21542uA4h6M4KPUftXq0n07U23EeSPaxnSJO5QCBNpjeoaVHeqjh
02wEqjaxXSo88DCLHXlNU1Xdy60LqH5Emo1yYj8kNJ/S6nXUPmUkpTq2+fR2/RP8O73Pu/BS8Imv
GZ37wTKT6uMVQkEyqRN/yjPFxYqeM4+xqm0CaBrQ6mCAn1tJ3/w/Rb7XRGUP+KudXHpfCpLOueEh
wPZc//buGAaVU+W2JmOUcb/uk/WE1gyBloVfKl1D/oBczKKLAAIVBzb8M7ReZgQi0PouYoWIWtdq
MZMN7ntQZZ+4mYbfAbMyH95gUDoryrP9EpeV1fw5C9HnN5SNAoYd38cZD8RK5tx+0TNSnawS2rw/
a4xhPFzGSIgTdMTL03Ckm+kXYZfrwgiaiP4Gcy/vJHHUDpMBirTPslDHj0eivK/RyIDuaA902TkL
nbcVybvZQLI9bAb/KgjJDySaGsbXCYfrNraVKCWUJcvi5TDu69j7RPCULyhH11S21FVafp1kWBF6
4fcqQzVcbbGQ1wmSkAiO57ZpUWrfJ+7WO+D0bkWzZQHlYfPOt8xgp6tTVZDg2QPk2HfG1CGGFKus
9Arfyt2G7JPJHyJV3p3C45oeuS3aju7OVvEoqsZoZ7MNKdiw+Qxiq0fexv2bb4rDYAUIbChiFNHy
oCbc6hc0oYMG3z92FWYpAFgeTiBKdi4RyO/edzPL7/RwuGsZfbwmkBU1Y+sIT4Gjb3CuI394NQRj
GmpcSGQqEUyDnOuBA7MTmHk5XLlkt0+/vDfkA499Koy5Wv1ajpj0ahtVrxajDAmOvYmsuZQCmqqf
01DVDgPCynljGiIsruUQ6K8IDNY7iXeeGd2Ux2iU8VGoXkNse1t2SE63KOG25xre6zBZSV2hDlmm
3/KDltE5YQjfbZ/zi1NT4e0fHB9LK6LV58FaVesfzDGBK7Dn4xCoOj12KrXWXCBYGR71ajlXzVTM
O44JsCFQgzttcju0Z3VLEdo+82+pWZ2HSWoaVPCNk2gC+stRlKErHdugcq8vZgSpOkP5VsSORJeG
7rsKqX+FnSm4KePm/UgTImFMBBrZ6QCm2taKfRt2WwgndNCrHjdoHaoDZziLWRMmNY7c5xmzSjPW
bKXArGggAqkJO7z14AjQn1yF7I4qtizGK8piFnsbZ8DzzN0AAD8wC3wpRQXE1xZaI+5iDEqAnoNQ
l2Qt2zUCElQ/7itIev3za25MN3d+xXzqUnprBDH2guincyuvY3S7RKYnuaw2hEnxxA7FaSB79HjB
Ow631XmeQa3OkbOTlB1bGZeL1gOhnnB/0toBJy97XDwBELvzpBfT11TtM0SNZI9VEi4Xp/O1WXWQ
3J4gLBv3HfoP5mNjwnApVKELji2r+JsZRqEFrzwXDK7gvfpKSqdLMV6u3lkcnMsXaFq/Y1oCN8Fp
uzq8FlLXBK+XGaJli2QFgIR0OatR1o2CpMOvIRsJ1FOrlmFEcEQaYamhjWWAHMaBgd2sWVqT0SjJ
iKVHGakxlbNuZemxuba+NE7joQ3gq77yoUFnD40yhJPZQuFhxhGlP1KYyICRaZj/eK/swaFuzDjm
dpEMIaUVBoi754DZIxT8DBN1/LdR43FoxmTxqzQ9gAoqpPCAbaeLOT9/zgvrOeuce9HS38/cTfqY
mtEV57S2KevhTn9O4EGg9az+StF3dkJEUeu5YeBlLtgk47yhMzJdxJ5wLzmDGV0/JcNDR2qxGObi
3wYYX0AXxufwtwBCgZVWk2zSLJje2zHs6ClZoA6fBIhjWVm9xC2Gtq3TG17g5D9XjdMX4gNkIK2k
/xYsJ+dZY66nF7l+/WWfX/xJA9RPMx3yBKHVrTnBHnmZhLmqNW86r0dTKh7SzXRuVfpEQMOLg9Nc
kv4lbN0LGOiuvBAAjLka4N3P1bUOqfidS5hvMnCPJnai3Gj0LUAaoe/nbyeMcHTSr3mcF2sGDf5u
b6A9noVkdF3tAS6EzXv+GfdTlUfVI95xLsnR2Q+QmWvgW/hzbP8U5H1Mdqko71xVOE+dzy7vc1C7
lRJLJzCfnvLl4VnjYqh2BnEfwoErx291DusMPf9NvQJ+1g3Ff88ICigZ3jyvjCWHifed+1RgHEGQ
ZUfT/SBV4lvi+8JEtjl/qkLmUGQr/Uo1xbxaeIJCcGcbN4zHpG/E8LT6o1Uzt+Of392ogCEPLMU4
dryB8R+W5ciyB5jX/RdJwRY/QIs/mqAjGmWwn4C7KZgdyP1VyMtnsC5FD5kiIk/PkwGMu3i7VCfB
TIYIuH3hpDAeAqpN4O7qnNG54tq/s7zJ/hl9FL/VkRhABGBNmo4YMtXaKHq8A8jcbiNNX5A+cXsH
oItSedVp/wlEJ2b9zOjlmLzOnS1D9hZ+WQGxdrbUVeGmr492SFdFYmFG4eRRsIyMKivK5J/JMCpY
Jzv1BrpeHK1yaOz3N7uQXPWfTwWcf4kOeAHUPQpPFT4RmLt5pJ3sKl5k90gFae9HLWYjTb/m17rH
gn9XwsYhxr04n+qAVLWn2KJrncsQADp5dH+GpX3LwT3j5fLPnUrTa7ftjDo2kX++EiF4UOc5vWAa
Ob/ZUSBB9kfDiSxFU1Rkli+JUoxn5pU5tUMNGpMO2XwiAyPZGbhAuw1TCpetOeWoeCXU49anf0hS
b1MCtt3xlQiiCrTf/XthxDSGkA6cvmk9fgyS/8GZLlXVMOphvwjhcFr6uuzoGlFf3tEbJd5KIIGj
UBA3bG79fauE1/Xn6WLeBqq4ndjvybnavEQdzR7hB0APFXj6cfxTNKNqihn8cripAXpCTh3belAW
oeJzT/TW4VM9pVxzZG6PsyOfA7qG04SOYgUFwAO3GWWjunEAjdGi4sMPlpUlzXr8KJO8bUYv27M6
1DgsdH/kc56GUxztn1/47ocMHOG+JNefqMZiKtijiXjrviXYbOkvAJSo+VoQekZdGKo31r8AhM8z
2aj1qhvVQdJhdsdh+vTUQN3Ilxsz49MiO5PHwBgxxJBp9c0R/xkojofO8yzT8F1xgOsfRPLhfHnM
hUvXfRuRJN9qd18qPVqDkGDs8DC9UPT09NEOuRt8Ze/A2ru305Y9sGjVw7Az2KbEtngiVNSA3H3Q
pscOYG1wmCJJ5Wr4udGTrm4py3IpzjBM5s8L0BhZMeXovnXgIxx92r91Gyj6lx3ZUVPZP1nS3EXg
HxQwmZA2JEC+3ilQX2cKFnVI5RvjEH+tD9AXLU6wYEiaKhnlRxGgdGuS3ee+exJHScrZexAn6POV
tXa9Z0ZGnYlnPfG9TDssipQCZy6O8OG39F7aN8JeZEsckKoIZAQcTGGYXS3Epu+Ng8QfBn293oae
LDl4p3q8XFkXOuOVe54Hgwi6MokZAcGyPIilkmGKvc34DSCSlrHNlCNyd1YC2NXkp+09gj4mSrVL
jilJb5EwQUBcetTicK7bfacOrgIpzsQM/nM7016LXhCaH8OIRzj8ir5uDvTez5xNe82UMlg2ntRF
jozw4jWqMX1A1kMJDy4H5rg1XuLGajnC4Sc5FASs0/qMr+SCHbNLOhQJcAvdMSNwf/ivfeFUcpEB
RL901ml12TjHmOyHbjM9v5P27KjAiK9HGsPtybGmntoqjXaM/MPKc0codq5hwByhCQWqSo1vLYgd
AY5DakEn8jtpwjDb2Uen+SPZja2RcfL/4Ptv2u9FGxbJceCYsiBbCOJVrzKGWMkPt8yVMSdPMi9Q
Jr21V/QKeqKN5DgXgstT4e/AmpmcnLAwBB/atGQkV5WX+k7m1qex9baeSeWxjFIu3BezgrDypjUj
LlYNkNngTAeHBwPhTdcN/6Z+/EIol7cmDpsvXH9giZAXLQhcRyyr9Fa5Kz20Zd/mv5wQG7OZun6Q
qI1ZpamXH/9qOW1sD/hhcqvU2pia9btlx3Sz3HdBa20qWEJI+dz06rNTL5jR7MRIqzfkjblhRync
2wQrVykcwelYAavzjB1i0fYn5xbBdlGuBMGVYrEq8XhIa3db4kbOPf8YGRCw2at6NrspzSLCW1TA
XOcGX3bUfVkgP99n0Az9vpweEkFY3SkAj40kxKXoQCrN9zRzGOu+mtNVvKCE7OmHeAQQfdWIGy0y
e8nD0Rwc4d4V8IaWNa48eKZlemXNqUUVqzdJfEI3tKrFYuHXcq1lnTNEsfg+qyG0E3Nn6dhYEgFs
sMtht5gaGOfpkjFyCb/C7Xx1I0AdmYyssMgoz1jKfpj48B2DM1/T/4Htx9wnSpeG9hkDsUDHpjfU
JrGSQf+Scrxji6wQb5FROGJx8+fLuTL4JsMAn/fPC3z9YHDxvVBz2nGHoWr3VLM/GnYOvSwxW7jg
hCK+rPxDuxdUkBlAdO1dIcCeP7feSOVH8SejYQKWu6M/+orZFU/RXVihrtsVyT5i/oXYxcGu09nE
p/RBl2mLXTUwZN5zczOQfcMCxZjBkTqRzyUaTTpN8dWedLqdXej+bjdV5cyHs4Dh+mDcdKzbMSEn
Tki0i0navh9HiqwsS4dtSATRy+NGsayBoaspnid+gLU5ZEZctGcDEFjZPmxS7xGaODnigM04YL/j
95qNIZ4icPSslP3jkqyxbBQeSpKdVwTQYRdUnYefy9HW5nchiCq/rrECCgyp+O4aSZgzA7O7v1/5
lvxdXFkTAu11n+wmJzfCglsrUhcYM0KoTWsTTJuQ7LaUa83vhhGNd8OIrIAMcXUR4y2SNjURrQrb
mr32qaGh8n+Aq0vu9Z7wfPCHQSditc8cR7yectHXmyKpdYZYyURV/c5xTOMzkLeU8V8uHeuPy1Wd
BZE58SJiSlNuJcHqorytucsPoQrOz2L7RhK6C2mLDL6ns+W8GtCtKJ+sMSYRzfsmaZK2oJZBjvn5
jhhEd0/phwdmWBaHiQCuMg/IMoxbzlzYEeCsQxSP5kE4uxXecEc0grcl1+KXBVhAcF8JkSJlUUDO
JCgluX58tFc6NRZu11CdvI4TfKPBBG5GmSB1khJBR7/VF/lUz/kCe9MAYFIDgNxjTdEk0eEnLqT/
XNDI4PTO8bKdknyoGJ1nl1/TENfYel9KqaaqZd4p6/TQIQMJJfMw+/Xs2LMGa6qYyCL74NGX0ct/
5VBk26IyASra0iWfatrOXetqmsZSfSv8jovCMGOJk/p6zX14JzrUKA8bu/JnVaKM2H291QQrQ6vH
FJrd2T938zxJxHc9fPzUvLNivN8odXbn9JKBjwjqykXaWpgf2CxPlJP/6Pmh8gap8lkhf8OA8NlL
BPzMaVbNN8SwX4ePb1UBfbqsoa36j0LJCZf0H5zdyDvhJs0Whx0tu2XoT29upHv4DOI1mSLUjWXL
GfggpUyQ1N027tffDOQpCJwBBAs00CZNzt6nCTT7L/xwacqYp+Ae2224JDcKp9BMSYziz/uyJWoo
fu8ClAFVd07Q2Hb2giZ0WqtR1uvaZ7DlO40DzXOFIwVgBoLO5ClX4Wf1DzUp9ZnuLgFzkT0bGYsb
WwGUAp2wesySIaCNvaP3dLyYve5H8EDHG9VsMu934+OcIrw2R1uW063qEjZqT4UI1dlRqucoNmis
udrlb9ET9sCu+wEQi8VTGsSCapt506dxB2NaOy4xGZzqvMcTwgZkNUuHlUDO7NPCvzrYi4eJzQ3l
9T+3+YscMP8jyo7tuGdtQUMU7nGYJkJ3NC+FMc2DeF1wMQAMMxd8Difa8EqrsK/mR0+CNNPv+hL7
zdoAyrT3k/oIjNj7HWv9nm7BWjg1JR0UhCwurCFK4QJ88T/lGX8+cHfGP1iUzevbWANIt0KPaVOy
myXRj9Qh2XFkjz+EyLVKys+1brHYFXHVIp6z2yk9A6IYuy8LTAxoxdjlES+4TnfnnfF1j15ZVVhY
OdW6w3Bxu8auCPjgRh+I0moxBu4k9/izSVEPntlpmLGwxCtvMiivoG+DOQyOZcFrnx5iOm0hoN1v
XxtkQnSPCoKuOEuPGINm0AvvWdVXIKELVV09MTnoJ44GwfW0q0Iuo8/th7PGHgBLiClnXC93VQT8
lTyhmAyk+wZSX466sQ/ruLZ77CWBW2pQq4aUxNU0U+JnVkZZgqlYB6QPw1LaGLPZ7vjSIvCwCmAY
0Y/X/lSi1e3Q+Thk3X7AGGfkQJnJSIWX8AAxlpsYK2ThHuGs+PdxixS4C9Ds0ZdQa/XylgeLN4DP
bdd8/EZnzD3C7mNZswq0zryFt0yMM4Ejo1ZCQRYH/PpcI0LDFCUOcMdZIVlIt8eakwMS3xZD1Ju2
rUtQcf9ZQ/Htg1unAHS/1Xs7MQyVW9EcBNMTJtQu5MX0uGjNS0odOEFh+Vyma3utzfESzurrbPhX
kkRcaI33/tffdwBpNTuLplHmkKxgk5YH6Y10puDqOyxyP/oo8ldPzWdSUTx5hpq8iIXYL5R2pV9v
rVX9UyrBDbkDYjgvm2DaQGHZJnWHwmA6sen1Pzv1CqrkYM6tFoeIy3+ujbQiWMi1PKwoPlRX6s04
cBMfZ6t9Bxct9yiZfn7bFmlx7tyKj67JfE3cyFO/TPi0GtsrP61xdSHkSreacQHHeMVVZX9ACdUj
/pDxZE0yxaO7mKypqwAX+oDoiCE/WgH0UeqB0/6eDU+7RvG1NRaKH/22mo7pb2zn3wGgEeFMyIsM
c75W3agpAeIsLcNxnRYGsyBAyvtJ8CsJGScKkN2p7x/g8tRKPpCmr7hj8k86u6GzyukZzD/FzjDN
Yf5LpZcML/OgaWamdmRhMCwEIB4VWJ3fPMneASpfliuY5nDoaZk+D+8B7tXOdEkD259tAJd26StJ
foQlB6UitmwekEi4pJ94qfOrAT0LJSu2DuQj0tV1Y9fj2Vb8jiOQPHeUo6JKKcxCges5fBkGu+23
5sb6IuB2WIrZcOdRpLdNjta9kyNH9pCprfSZxxraC0Ei6waxovM8ng+AUCI8+7JccyQctRKP8uxF
jIJjPWlKxDwDx+bDP8jJfpRs9xJ0JWD2QC8VsekxvfmVAGWvCHVIG2FuGqNJXaD1lf1SAbZC81vC
JS4Ge3e7eC0BQ7+SnDXFDsJytrZ0svgn/pyvImhav+FWFpuQRHL+yCEuVeuLJD4A9+0hx09nN9Gw
kPBUqcdc7HRQ2LxCFwtvDxQaOeF4GYSmqXHhHx8HdrUMjwN73Vh0MkCQxX0kTTYbQob3NNBbpJ1J
AY+hb0SYpYMOzU2K8qzBkMdHG39/LvRCh1XOOydDur5MRRTcHyG6mvjduJPXrl44/LbeM31H2eS9
qXcB1vfKRTNzkfaG695sD+fP4e6QBM2c4ePq6eRKkxCEq1AdJ7q/qxMX5nHdpAm2QSeFPzoxXuKe
xLPVI0cJiTgzoUonnp9aKn+WaEsRK3osjXjzXnMpS/AkjnU3uBXNuVlPSkG3swl7ZBTXlb067tvk
v1+2QyhzNpUmrjWJHjbrGD+9J3q97rH6wzr2MrHsIOlo/CfGAwvI5OQhtWAngUwRZCmt0eI5obAa
bVa3yqWVOQ/4lW1agKlVqOGPUfPyaFczcPMv2+168sguP9czvGgMSAhC91ptvpkNN8TFuwPEUdz9
Y7JI+orcSM8cVZPY5tmoNG/pRo0nibgy9Udgz4+PEfdEX7wh0XBktWsldewH7rWY2qTE81pqdXqs
rAd6mqC3ztGuV2DLd0U9O7tf8wu9fUnwSHivp04mZYC8zbbdyKUJMYnAaSgDCW5ZqHvmeVzXvBJK
uvO6MOdc+96aLOV95MlJ631PXbcidv596SuNisNZ0gc3BC+5S01mjrIaNVeznx8EMaZNltTgXxxj
vPtf+mKKXNBI7fwrOeUOpZcs/J8anUwNXna6NjDYfwaF9ho9q75rE7Yiq2h7/81SPO4+fbB7fDae
RSReBv1LcwGbYZdyPpDxdja+WVKTKHrwR3dIYbsIGKYWEf8ioDJIF9CsW8t0mqOmF8VbdG9BtNsz
P3cQv2kPA4jiIsdBKvljueFx7BioDopU/A/xk7oX1llIj1jfinAMYaq2t4eHR+w6pzGeD9sDhdMy
/WAw+4tDmWlDR467ddfewRgx45P6k6A50ouD8XSKe++KK/KWeBKSCy3erO3LlNT7TGYl2RqShX4t
oSElJClS5Nvn0qQApVuw++8gnnTZTt4vuXjw+MZjWrJO5Q6tGNpG+1RA+2CZE4PHXCIymOjCKde1
2DUTAVzxEvjIdi8gbGYI8b0MzzrSpiENnFFXAgbYwhLn6YgkIjUB4Bx3VgLSgA49YmAdg5LOrvtd
af3xVfJBVdHt94DEZUpX+znojgdgxzpQX7+lwXHuBI5LZLzysH79RMAVyQvRoZ3dQwnoc+1bnGJH
/lrZJL2RX8SvRTJZOEfsPAeuYJgvwGSoz63OoZKsmf1nz8d6kknxTmlL2oUFLESV5H4x9icFBJb0
WAkPi7d/ostqoTQygAUBgwQXofdJOyN62sRDhcDlXBQ7lMxTKg+4tcpXX8VYlkXvEpK4hFV9gZI/
03XIIAvDmEDg7c507ZVpGvrBvZsVEu0uEhEsm088rrTNuVyba9unmFcVr52cnat81fEJt9RIUrHt
SD4ZQoAIcxLDrbU/96RDVpvADEMRmIBh+w4dDeRUBssimBkLN/VGYplYf7IpUkdMkh+QSra+YHKY
mMTPpWfayb1Bdowx5T2Fyh+UGynYQMe+VmzzxdmMBMDTrVLW+Wvc3vUSIsjK8pVieEWYwigqKLni
TE69KICQgjhqw1O4YK8s7+UKkYw1iFyWzEX/ZkKyL0QUL82XmTstAAGnzIBOLj0zNo54lWnsG8p6
P45QlJLqMD3Ia9D+rzIuLqFEN7dJUBRPz57i6QjogZxXhgX+ZvAzFr7U81WvkS1olRNCiQHNbucZ
HavZVJZ+9VE/1ZNghs9rCN2SivkKvN9ELG6ZSMk8TPG8Zk9cWyfwd2CKogfmvx0PU3058ZjkE1vG
eeUE6cIFjjVC0LE/NDhV7pYjr9uGmhlNehK9I98HIo7dvYqow7KCxXDlD63KwGjffkY5tLRaeMzi
HsGLF5SrGIUHMk33yDbaUi+p8sjbdzbLwKE/aoEiWGpLG9ApaCfSAFqeRol8+xlQhhC0oJyQO8G8
yrCBiXJDK8UvOrXQTHt9wt3BDo6kKep86f3EgLBWVOgwUkO1xrMjLTj0VOErQNM1ac+9ZVrJTsIm
pu/c1ynLfN8EbPzfwIee40VeJIx4cnh5L1YvQrutS/opg+bdYUIncNyK+QRBJG77pf+syryrsrnl
2lYw05Y+NKaBXDwcc0Ykpw193URQNlsG/xMJgqRHwnY1h89MayQKE4H6N8AMTvyYdGbLrVBrIkQH
tBtxxItbdiSVPYJZFBv5RG8MFxDkwcjRzdDRLxEfeVntljne6m/qjto7Z5RcaL+gh9hJZZ3fe8Uv
sm1tt6sSJBudnY0C3fIuPV5Jc5Jlk7LvVI341S0vsjWlcruLFEkL4i7YmMAAkiM+FIZSzLnY1d4t
lerMCWpmP2Kfq1KWgImy7dvoOQ2c82YSepszU+8oCbe8oTDyPsRHWoWZOqDTWAd0SPrPeXweCily
kIkoKb1X+KZjxPIip4KEd684gCRpnW/nWPRmev4tzkfc6FDW2CK978FFZJg0QNUspHzh4xBfVb0u
4c9drOJHBXoRnN2XUtikoU7/7ccXBDYm0Hz/vPKjgF3x+5mHBlKXIBR4PdgKJZM0xq8zsqaDt4Dt
FCeYeumuJmACafIt/DDPX6fZnEhFYAliJW2fQct00jp9Zri5WHRHzDqUPtQjOE1y8L9gygIdPt6U
uTL4nSXyJrVZOaZF6CXTsz54pEBVx2JimOQbcTcLKkxLmh4U1CK4otoov2nIKqsR8ZfB+ZJugXe2
dSZAgkaCkeDR/5u92v3czPCE50lUSEEpOAsCtc8WFE0n+3D+DZmemq7kEoHUW243rFsnzz0vf4Lz
qGHcCFtN3EjtNAQKEk2pciXAGqg9TP+mm7IkJQ8bmAAXhBlOAHN+ZJjymE91wKNs0GdmKZH7tKrc
zyOG9EdKQBulOtFiEd+bXG85xuNLqll0G188QDVi9YLvObBLXy3VCYkTH/hRLTwem/U1MrSl4Mey
0vqXvyOfuf/smBmCyDMCwluhS8OBHej1ab5tPcwKEv5hg7MouGFrLvgQZLymmf2SMEApnph/uwjV
SSpqoYZrXZ4Yl4zVv0YKs+XwVw3T/UezitsxgREDU9Cqpwj312Y/3dxBcPONk9zM+sQpXiFmCEhT
n/y670W4vyEtJe9RJTkK/gmx3z8my9A7bMrtEofEmulJfd54TuPe3K/7EqJemUh9B6KP+CQIfaic
SPiNhr9yuO2KQXFvo7cYuZsSqC6W/6QzwccBDHzwVNkw9v154h7PwD/kllj2I/WKUJD9IoBuTSEz
ro1Nm+rwZfneu6PsKqPY9JRtGYC/9pliwOXazz2AcTnciJVpHu2uOPWsvJAMpmqtUEpaXhfuwOv6
zBGqCyhUZvA3h8jI8+d8GEwVFCRmii3B2tf9v09VbHT8CqjzORkvTX3/lK6qP7uLKC5LCnP+yLZG
u92ye9wx7JEbK7z3MgYpS37JPIksAOm6ilPHYMhaNz72k54DHduhTia0ucWqBtcdB5wmFt9wZrXZ
IP2L8yiweMTa0udV48V8008lxGVsfr+liyj79LVymUlCnaTtNuxxqNgNpySCgPqPSeA6KUFjtAsH
3/aTDQpUN/TCPl6keHPUX42FLJ4UKLxLuqpKmCcqbtAy9kdkxKXjkuTYNUmPIjgLNYeX5caYZ7AS
L5oXVDFs6SsqKteamwUy4lHPKCz8w/Navz9yLyZqOlfTM3jbDo3VAjAQ6wpVBKZPeh2M6CvCRnJZ
OzAgCYIo/V6yCBic6ca8+7DYrEZ87xd6paIWyPPvCq9uRgE2qmxUo/KiiNveeUaxrfgi7Q/TlGGm
Dc1U/MVNPUwm2+XMtYmyuSIKlde2vCY0pH5qik/9I8dbouifJCKRguZE6DfzwdRW/fE7bHnwYImF
ZEtd5pih7amN6/fWRFw3g/IUQ+R2yYCpZCBCH/0ufhbZ+BQw/x8dWUJziDcLTIRaf6abBo4of/LE
CXRw4DbRmpWE4SlKJj3u/wx/mZqqvmqC4ABCkKGeH9fmC/ZcDV9Sm18PDnm8+q6pxa+fgRlkIcyJ
jrv2JR1Chr5pbSQZvwhz1uhXyzEwHL6N3MiDvQnFjUQ78VJW4wTW1xHvO9G2kcYxmrnGl54KX/BQ
rLGBG+JjbqBAY4ZWts278CTiWUI1roOZD8uRo1dTE4PIpdA83bqKyAU8F95ZEDT7firmWOHAnDCX
+wlfs0dofRfqfJt3rOn3G5LMt1w0WipxutBxga2clQ/XpT0Sy//wPToWmF/lnZgcVufJoNX3xdVz
Ryd5WDJzpmvBglQbjxNImtoEVly7zsHXYAqKfkDnhr69finr99IldzDi9Tw26avURHM0YwKfJv6M
dsLRvT6rBG6FRao5uY075sQ/GvKLyHzCQM/Ko7uajd7X5CFrsYox/9eg3IUjr2UVSIW2wRrAF/qa
alR2eyrpvTRvv0OST+pwlIPU1KtEBxGfbNUoVfA6AKFM+iZgAvq1UtXlw0f8JhVVuB0Sw2bYEJcv
/VS46ZkmafJLS9OLBXT7N19IKR9awJaU/jzv86A6lQcp5DBlBTE2YOXzLCPucjkBx9X1eO/3GCaf
0BsDWQH5gS913sGeYoNvUvaEF8YuNRcFds03EpfHQ36pMFguVusbuWP1gQg7jt7qsPFvLeBTO1/l
KUnITPshEf+76DaHK0VBKmV/TLAwuWA+NYEllHpJt2RTSqZ63GaiulouHlpk/3APnAyGHWLFVtlC
det08+zWklCACH3Pu9oQxnR/2cJnUnPJpI13rEyOc9DeZ77H/7sCtKZY5CIP2fcFKjjxUQBbN648
z2f8frnj9dVhdpYunJipKauYPv+RydFNC2h7otx6Xncz0gUFQIplRh9dESeYhIezlA7iSd273zO4
GiFnc6JMn/qw/qXwHIzkhs20JKi6+PmJTGUdQKmpJzuYfSr24kg4tkWBsoOB9AW/Zkpt4C/NPboX
bnbgeZEY4Z6Vk1wpflHFuPBz3xa1olo1R8HZUxF0y6VQtF+CIDaTsStkWIzmQ5iKIerRSB0Q2yUU
SzPAF5QyQ8y4x/JTYpR9ucalvdP2/PQPGd9eelswbNAotRzNKhfVvF5mq47IKd/DHj5t+OIG1s0B
oj2c2wEtkrsPjCtbxR0ImHqV6F+1S7xda2h7J7u3pe7qlC9I3DOCTmP+nJBsMMzU5MMc+wpiMsE6
Bcw0ufYePmdBhd62hMqBBhnbHMK19GAjT53qN8czHyexWdHPvN+e2DLhNHrJkLaDXCrwtEdbjRm4
6VfXAajkXLyLiwxxXe+RCwDmtqMwmirjMelqMFBs9Gn3StyAwwMZrhy5acvrCiCnLT5pX1mwUMyO
Ax6V/VW/fn/BFiKHPvsKNf4muj0BckyXhlQf5kqrbsZzGUTnXwjP2A5+LegfHwbYz5WB7HarZEUu
vlcP2K3uSdjOBvD2sGQr1ujupWRx1nyeKofN3JRk2DeU8kHjTFdfvNnL9MwSlDVQ5YYI6NOJtz0D
C4ljT1R20zOEVPr6
`protect end_protected
