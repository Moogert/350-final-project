-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NZNrYITehipAAoK3u04AprZJXxkLn9l6ckD8CIZUA8m+3znmiege8ViBYs6o6DdJXi2Su08NgMmB
BCmIH5ZcUylRw0hgAFv2Nc1XG9f1jFJ7ixfFtOtjolURgWNW7ZZeyg/bxs+kykj/QxpR6V/WzVW9
SaCG/AQC+LDVwjibIdgcsuWY8hC2cxY6u/hvYJNWQDnJkHbdVF2eyKQ+ouTD/kQsweva8mMBzmLP
w5BVf0dI4h6S66KZer1SGt68L4MK2xWMqfr9tQ75XxRa3G8N1kbd18KgilMNQcq1/FRZsXzm1ZK2
xvQYOYnsLgSJAL1fUYdtIP4qzHNXyxF/owUdlA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
c5XJQkNhEaanUhov12DCc88p41eLL2w5e/aZ7Gunmv/IsxRBB1SpBlPBd0pr2DulLnlHGROVlREJ
o98rfwrvf9c/SLwRcBFPxbnJgPYVy0XTUQZ47QtStS1mxND9lU5oX4xe5ZIl9RhZdQSfswbY78xx
AtK0JJhzHqCN03l2osymmoNsMnQerSy2HeimTOkSCcVG3zzVcvWog3QX0an+3629ouwvFPQKec34
gNhKcA6o5KFsR7Kv89LNlbwBylFcd66j85oaUVgU9xsRVv70j8gLJDBZTPkA60B6EDsecAQ2amhd
SK4jZlYDmS+h+pcQhoPJaFitP9Ye+AizhVTEcFZSRty9MXWStR67eIZkg4CdAVP3fDXZM3DeDGCa
od27fjmX3Pa/CuNXuhA5CuFQEH0xPtuuwOr4byGXECL6l9+T9XX1WEes2iMAcSi1xvt6jhfkJloz
nNYk/8Ngl+Z98Idx63im5MDz7xE9gKvK53AL6BnAk4ShWGEPKhTOreeIKpwFNWuHlqojIeG+LYq0
gkFY1Etd2XgJOnEcUOMCGuRZHKGDgcWZLlf29JP8eGzRPAdksv2wlOoQLhHf3RCzqVAZy9/XtRUg
bENoWq52P41PrFBoNiiFrS6sYlkCkIxipPqyyuC8gFvjiE9IpKNE49yjT8nm9B93bvi90WHv+8ED
Zb455gie3Ibcu3goN/hMudfFBS9YGA8B9CRvz2RYDLZkHBOXKaxkbf//EqoLMfje6CNJnlyQwBpH
4el2jT85QAXbBuMt9ddZTdKg4hgqUBl8MgGkqvwhqw+FznXd2VxB46he03ThHs0npKj+nx3Qf8Wx
/95IAB+5y75BZJR72pXWnXBIXvS7kSiSqv4e+93H0FdVZpvwe65WtX2gh/l9jfMfFRIEuXs2YyBS
32xPg7CI9o2Fm+ghKYnxrKY1ClinccNV6TKcdluCvULuVSYDHye9/In/qb7GbCAxCPmS1c6q+5Nh
mrLHT0XDzHpqPJVEP1Z0YhF9UV53QxeYzpkBA/SN/pqMs0cCZm0oRMJOq/CI12P++oXFmyrdxn/+
/+MEDv3kg67+6omn9BkbOCOBbUhPFVI8pT73JTX66zqMaJ+u395qtqtPwd+C10l1Z6L4v3OnkfD2
JJ/r3Y6olH+GnIPAI5YoxmfzcSPYR5L+pOLqB73M72InDzEx9KwJdS1mLaLY00KRcwuge9jiW/37
3osILu2jwWeVHCs/Zru9ZxS1oPjxrJi12zCdMRCmLJRj0lKsW4SNFNNCAFzM29Plb4e1BfkK+TnB
FP1+SSZSUpP63YMexULcC/39AnfUcvuJw5kAav0aSF9EaoB+kwPL4MNx21iLeZT1GYYuc88mOACS
djDHHgAdGHM63XFaJ7oVRisLXC+M1A2Qfgqlb6llOcRGuQwEpfGqvbBJu49E1J6ueixatTGHYvyn
gP+gHX+HlLx12rjcFnLePQTEBX6Ihszoih6ueyf7lsmNCu6Eewx9wPn9ubr2ovmzzDKGJqQqFD3J
bA7K4bnUKEZC9UIp/ihr+JBQxFUAhUAGAK1nTJBZ8E+3RF7AaPN2Pza7ivCO1RFA5MRPSltAKwwP
V4XzeZd+o77o4nEfWNkforck4VXkOeyMBsjc0EBJfCQIUpJ6G8D6ihv2RcboHRPrcW3thEdWRyZ1
nrNBc8JNr9+5TzN+2447BBkiig5KMcaAa1bNWOSyqLsqEtMgT2BjtSQSxGB2+JLzbJ7MlvB4qHWE
F7Q5Q6nRlr5TjWTQ9BL+TQ2cHmwm0PLzecriMp51rmOQ6uDfgo63fmbNmKAu9sOIxmsCs0OGKiWd
VUTmPUeCP7n0aj5sNb1PpCJJZDbxo8ixvIearwIGt7k5Vqpg0NCoWLtBVRek4Ry1JVt2zkQIyyyi
SODjbFRVdM7vt62flDyJJaA+35CKDmTqpX5limZVJAVZMLqeUTu26t20juOdoK0jcEtNgm0hjyya
j/labazGJ0maapRw0LlkRMuKQcI7OABtfugKgsE7QF8C8nH7lP+e7aIhwYvHcofrg0heednVEEft
piR76z9OO4Kn+BAEIzT3cQKvo+2dhqw1TvZw9metfhhTikaHkGgcW5IhrqMkDaQ92Vx8OO3Xt78D
7LN1km27Ovb3Do+SJQAd5nxp9i1MsKjotfOPPSD1Hv63EnsuqpIvPBEC24lo8UBZ7p4ZmQJyXO5K
fE5xMEULnHJGfc+9JNtO4arf/TgFOoRvmcxztoLS1tZCCxq/9VzCpbn1ORgebL2RMHKXBgd346tn
tyRBKhljdq87ZXBNyN5s88OnCwmrirtnaDtYsKlP9AUz6u2HBf7/BEDQFilERonY9dgnA4s8pCGP
sdl8tWUYRQ1R3hSSuPxHxY9vBUMIXn09WEGet3OHgk/uOB4yNn2CSXZy/ny4EOdYjcHCAENsSq20
GgpDtVF07BqMvMt8E5HhuVFiLTP/ikDLzeSAQPYSghjAj5U6Syt8SFC0U8xA1Y5Zd1tfqz9coaV6
sl0RY71clNKk9DBKVQZK4pzR4k6nfcJa7/7sXViWhWGilDfTrPr3qWK6ctEG7iVKVgmSyWP6DMjR
SzBQOcgbeKIqB7mirLZzYNTi5hWs+NzyGxaZ+TXv6jzBxKQJUe+zkwZGmmW1E3AXIP1XXb8fBZF9
2AkYi7YWqaj7aAgKPIyVFW3OsPglph2l5/pYOR+tAg008vYeRmhzv+eXyEwNh8Vwz2PclAFgWdiZ
lcUGRsRIYjAIUdoHeTd342BaVrkMeMEs34c9nRcPj9XS8eekV7Vjd6RHewPK86D5sS1o81KwsxUa
EYidMPo10NzhD2d6BXInm+hRiwTFDfCjNaricUx1MODOauUMenITzMaBinpH4FcGsvPgRFXq/r+9
CZnmR4DNqD+r+PL2bKuJHV6FTMrHm1bw/GDc+VQCEQMLevvsPj+3z2SUYoSmO/e9dEL8HKASw+96
vTkccioFaao5oCaoZLRdcu8CVC4cFwxHBYbNjrQfo8EsiOSbc3egVwJGe4IRTg5W7CZvytsFx2DV
rvb9erBiwDDfS0FQwk+zLq9puyxQww5zT0VlceOu+NraW4sM3NISosp77e45RsPbd7j945DRpd3j
VKy+g9YfZvn+h0GioLHYkzdHklOI5RDmtywoA/Rnk8DyXyP7PPTA0+0JjGpRofkAM7hoMYAmkFVG
KyIZiXApYUXKP/z4TeAWCx39T27QNeDMjEhX8XjmFsYaeKU6J2QcUc85KQbIXsMCj8EA+03lOibD
C3ctVT7wFC2TYBESfUGHeo9IHpsdtUHaVUASGLTrxA4liY/OERbRtqmWuwiLnqeXk+/9mw8sW6Y/
OlSVUQn9x1mYUqdTad0MucQfcvSQ078U6yxzFpnTxJNWRAQcKYQVdHOrCJG1EC0l/f3sv3wMzimc
1uOaBXZBkH/YSBm+dyeeVMcb+2EiTBDUqT8yWbXQ0QqhPDSnCm0bv2IumAQddbS3Hcn7ivsN4unS
1c6fwXYE5TeAjWGQLlWVYauWG6JtlX6PB1ixUdBI3PC7lzyHlKt9uLDM8Y068BBtYAbZ9swvBR07
mZCLcZve5WytSsecw04buJekSWcWNG2IIM+TIpG5NJd3WdlL8+4Bp8yNNPGj/04KlcjSEPs7xWZZ
eKGz0LCCvTJ5pBO5YNY23EO30Omvwvi5vKiOYWVZQPLgjp5bgljquKWglaAjoTfbnfZSIcG/a9dD
xfCzNUILgFKmZXlGTwyk41bhXhRY7DJ8c2SNqsMc77y5YSdqOsjHG5Is/iM9mPp2aZdg4KU9lwtO
yTQ6dWIBCBmclx5KOIf1gnT1VS6RzGQ+TLq27uBDKAhYY25tp98AcuoKwJ48uP2qjm65EtMc1T+i
pH0Z8ONA06e4J6u8jfwJwG1wziN9h/KULjy8xdE7kfZ57ctWrwZ+7rUJCRcdme1M9mYhA7wZ3Oi5
gkXjHnyyVNAx9oYCeW8wgVwhqdrldxjOE68kDtM8dYDXAvzzwddsQOBs5yW8U1ZoftH6adZn88sw
uWaKaDdxCBDU5a8icsY/WgvJOgFmMnhe3UjxjUbn94R0ZZEWrizFZTEs8Z7UEy4S/x4Echoa05Ey
YtxpzoPB9R03NJ/Q19VAZDPOGWN8i7wxbR6YXdeyQ6HNqH38bcvEWejFBFqRb1Zg37ywYPU0iVfM
gN5zvmcUImrhnysDGOYlXiHDNB8PwosRzS+ON6QMXW1g64f21LNUOP4Eg89hC1ZMZAHrhzcouoDH
qPdmWwHIA7qPqhjROo97g7AgkUce7Xghc4tlxjlss3+DOBiktUMvOaqfS8iFzHrf9aGUlxbFk29I
9ZKrgC4gUn1pKHOSZBsIqN+ldZHcXHkyWtAACiGJiVYJ76FR+nGbmJ3+1RCK96TJstg8kjZsCZSK
XzxeEWkiHVwrOUlC/vc8CUwrMj1MdsYIMzSFY2U/wgCl0IKhfTlMO7n/+xiHZiJJfeabXDmJ8Gyd
d2QpWCjaQkjJLBEcxqh/ns/jdZYTPOpeZqf5imTdNcbeBU/FrkszKB+G/px9rZSKoQTRP4sMFU4l
Olbo81lzn6j0qccgSJH9r1lE2qhsIC0QOecJt9efYy3vMy4S411ng2ueH6yBRvIUQo46Z1OolEtp
e/v2sC5EZB3X5rGipLofvugSUPFoY8KE3GkfnbSxajGzksRJY6EhwJtx7c62wkm0asTi/iBjRCmw
AphqGBDZhICjw3pA1c5uLbNrMTXILmBA6N3auYWWIyyvaZxT4ocQ1HL2Dvm+LFUc2ufy9liNy5Vr
OsIfvQpd6U7CaJ/+y96JQAXQySWOxgv1OOeeW5SBHK0f29+nycCcDiBaDVfO9ZqGf9Y2bGA9TVod
ECoRhEnTlYyWfxWdUGixBHBBlbIKZYom4lwDv92rqKaw+tBJC5+4P/nwvafWE1ekpO/kiGITutt7
MM6M0bQt9/Lymo1NVmc7gXJIw6e0mogQY8hlKSKxL7cA6PjJVbM6xISYqrtrLCwUPK37GrY2Z0j4
WoKt0fCH0E6cBQBAQJfaw66fHQ8W1JbK3X8nkIaHsaFcaK8Ooju5xlGY1XiIKOqGK791wf6NhQcX
uceA9bmQctBZOHC5q6N7/HYTlGAwsNhyF9DZag2j1zDSlrYVgvxKDAj98C+IBMlVSmeqwx/cCGk0
Uap41N5O4EuHZH4BuCl9lnA1DNiMElmif02Cz4Whi5AVzPn34tvSgqTbcQ8mN/n0CujqNfoJkkMp
g9LEv6AipI7G8ViaOk/0shfhgZMcyTxRypsp6AeP8+wCHhRWqIrMF2XuUZ1I41/lW5WkB0Z5x257
gfrTPFcHGEohe+AzU0rbuk6PqRdzc2kRA5yZj050+V4Z1UQyb//2vtFbaKbmjj6nXXuqDV20bReQ
kV/vvx9SB65VQEctUeXF1eNY7MZuAOfgOScCIDcoiXeorei7n5g4eahMJq5cG5LsKe/h5r+ukEOk
akWRVj4TM+LJR33jYv390VkHMyULzYMpU4t1Bvt/OJFPCaAUH0m5b/6vOZjV7pGU1wxh7lt8LvTj
ex7Gdbod7jj3fu2fhgrtY6o2ORVS1BDBtrijhdRABB/P6+iCgqwC/W2fTeeEd+XBApwPlAEovK/I
KU3OUSISPqgly34chWTvjl2FAJXHWjwRrT9bZBPmdUrpYgrfMmsWe5tXLXdIuwDAvukUU1+FHiNa
ggMehGzrl7+zYrpYpL3Mwi/T0J0ElPXlF7BGqY3sz2IYH7OfJGQNjI8k+XogFC6/ta8XeOytdxW5
GgYgg8v+xPiw2WFp7ROp3VJ9DH3WPfD0TEurv2hHQReAQmZ5ekoquH4uvav2vfQHptIt7Pp1fBZN
apcW4Nj2FywifjK4AGckSW2a37uX+koD1AeqB/n2rlyUkCIYDR7+RxMJWQgPJqVxgs5DnoJDrQjF
tTZ7ReYN1RpERaop3jJibevanQLd916mAisrHYcoOwC85kJxTEJtrHy1DCE8rX19khRdWOOHlV11
1kWHxFwPcciY4uRgACVJQMJUAAykaWFdx90o4xhlUmMa7De4mb8/3VpXozOgngqL3ZywKU8EXdGq
hA1u5n8hraZaTmZrHhN4ZHPUbvHxp8nokQAW5gHhCCbdy/dZVanbaQXK44L5ZwSP5QvAbYLnBLXs
omNehSN3jOc8VF38kYG9tc32rLJ6xT0d4tGiggJ61OP2ejCsRAhcpla1Mc5mr1h8mFW9E3GNJK5Y
vc6xmOV6TNAM17XQgZEywtkHV2dDFds2kt3UrD7doWUTkcuPKLS2k1p0W/9PholwF9ZQOX3MixHU
3x7RieMqDBpby7cxuqewQyi9egK5guLoRh/ZQil6RJr1cU+CGOzcM1fm1K/MldG7Rus5up2A+IsE
b27+tOOPuVVNLzw6kXbSaKqkdUD6KxMssPCficxJGRP9WM94aa6+0hoV17J6QzDo5q4nTF7+SsOk
yG1XSNE0UmFHmGvRV+O4pDPD+CHEx/GISHu2KzpAAcXiRIfNs/b9FwhOz3JsjM6e2wxKTUq5gGTY
hUASbLUUcxqS/cqxv+2p9b4YD58PyMSOTx9KpeqIcqLB7miA02qKmWZkF7Fr6QMYIU6MAdLKR2hN
az6NSlGSPrk4M3JW6TKhN3ooRYuGKsGDiLUU0XfCYn56qYWYVUVAz8xLQAFzz+f02IWAeI2m6QgV
J0l2PxARpdo0LmVUUD9EYh34BUdd9KnHWvo92+oArp46mEMKu4OJxc3RrAONXTBMsuzmDadngNm+
9yboBDmztl9HYm45Ad/mDea6ffRgTYeqC0X5A1t2MTCkUhFHR7fQNHyIhhLLOX8J2P2rf4dcl71D
FspU/6yPPYULrIc2rrYg8rEOQc+gPL6xd12fUuaH1Y8y0yJ39q96RdcW/mTXsMw/PQbBEGsOZZ9S
yjH+GzHhi5yZ4JwCvfzFk/eoKYNTlD/ZINrRIDVUi0K1v7joTlZLfDb0NUXPkaBiv/0n3cleArAq
E64PtlqJ9zCp47/0GnqcKTllMoAo35jCpS4edOe5JonWwV/V8b9SQsOhrx88wMs1WvOhHh9ywGRd
6tf4LhtolJj5lqiHRY5wpQUiSfcxRhmhy3yT32xN7yblZwtaFEvmLDLmfXmqO04mTZoTTpsCqYg9
rebwCQsr0JAPl/wSbrxEXVsDBRQuObglU35mbpvH7nrW6tnRjlGByOicA/hg8KgWaUW/YF0cy2Y5
EdlxfFuesQ8vetHicF70P4rqkaShACqgw/Go0/f3NUINVC7vaXou6xXA+jcOJIz5zhNVkrKQU5SA
LKah+UbOD0XEimSYT6mgUtF7+S3hwsro95oDBO6oONT3ItzfvczxpfbMCDazrB1POpY4tsB6RwkY
/awaiLlsunQnAvK6PoovL8mqNkDYq97Xg/zVXP1c80DtMIdSADHbLwc/0sCe5nWKrggh5sHrVMVi
EIDlHh4JH99cxqvlpbKGV1yRU6e6mgpiCYKo5pcPn7OKgXOc6aewKL6CMUZSp9rniJj0N0Aih5og
agRin02+Sb3n8zYQ+XcW9ZBRmRsG46IS0Js2cvY7sE/V9qu5/dl45EUxcHNqzOI5NGirXY4Z39OU
Ht0k8koIEo3qS1qy8Gora2I3tQKxYAuLXey/oyNiTdw7uA3rykcnsAvbliIxqAJtpJWywDZYKrCP
T+cWSmn2N6tDKO5gcpdbMNNqUOX8gSZ1+qN2M1fnTlL5jA3zMPOgENiR3JzFE/XZ/dL3Pwgjcru0
Zar3K6O99Cp8fjKbmqwAOpeUo9fu0lDVzVaqhyuhJpTqJBuS8pynPbGoQ4pHkm6Q1V9VSiydAWec
TXtb8HAinH5hilmnJiNEz9T4Mp1wkHFLVZBtY+4a9ksueYcuyAcy8VJsLnzo5pxsMiL/64yBhzmo
WqGeaICjF9ZddvkNPQhx9ocBXNNcxZAE7PWTKa396nc2xczpCazEUBTvbdknMXKVtckafXuoCDhy
1VX8LIp7OhVozLv8gazjDXnrYSXmGKwKNIclxJHk12RaT2pKbdfvGaBv7rbmubgbf39Alsh6yQJr
rDcweVn4cvFAPK26AQTbUTQBUMYv2dGjurXdmpiq6dqplTXw5EYxWksmpGhMurDYirwq4XSw4GTJ
dn1E3OHTv3JpuO4ej4UXmpS6i44IKLZfLjrMIADy2GCQZl8DvFDZ0R9OwRZ6td3ZALRWpCTcPjxw
OAZeKnc0C58KfV76itPeFnGUAORku9hmLw3h9OuM1OFrVMd/EXVHCXdCnMeQYlPkYwoHiuNBFJow
HiUsJoZyNTsSXRmKp1dUX9c55nDASpV28La5vM4NUJ8IXKOg0EH4hlgVapKeh28YyDZgS8f+49VV
FSCHfVmoQi8RS892jci9m72RkCfcaiVg/DvEgsgww40lImznJTeV51dsYgwNNbzY0Nk7I1lLIgKE
x2pJGbW/ZTLMy1HZPsD143hs5j7N+AJDxbGjk1HclHyazgucKguHqrVDQNMfKrHFTD1roEViVt0D
48EIVaNE5eCJUPui7vfBnfsxh0+oDDZe7dtJniplz5DU4GOeRVEE8Prs7Ok7J3fS4cLnxNZI2d7g
hj6fA2Ifx9cNsymkRtOcUvo57DSRxddS4dCn9JhNukQ5/IsKUYeXjGjMoKNrR3fWT4WjUYx6MMUp
UoVUBTN2usVOLmHrlZhX39+aUh4MF7Tg1fr5eMuUqGh+e8NNSCYo4CdFwNRQCyukau9Z995gy+kt
RT3sL0ZgrUuZdSSaot37g8D+ExcX/o2fIuQO1aPPGkNGux1ALIuLOSoB6KQKVlrXF8Q4jh3luZ6h
O41J9CJQ97HzoCRdOH4vu+0atedBe+xfqZY7UkPfBGeKABMEUxAaZeyVKwFoRA5UGa9hTsMWyguS
Gok8MgwqWZIGKzDJHXIackditptWc0bMbquRk7ljoxcq9/kBmUYgF4wRSx9rmQC5V16E5SR/JBG/
TBrbcZWUwPde6wss80ZRRH6FKkoNMalBPyKtJHGXZNhu/+lPDvVRIffTHSxuTENCPnZHMAoESQ1G
vHjmRKGfHKBdPKBgjGnXGWUnQAzF6/w3Ra4VXM4w70l+ynrhERq0kBdrhA4961K/ZFNCc72Y5JTs
ygdE5c0xyYadFp9mHzV9699Kb/m27rp6gB5iBuhcpMJ3HIL9jHpeawL4XD7YMQhm+KK3x/nhOKDa
kOljryown6QcAb4PZlBYw8jkCWuGyZ+1SAwMWdEWSYpvRjnAPu8YSMHINfEObu71bp8vHPJhtObf
gLEBx8OMHy6tgKXWreunCLN+9xH4FNM8v/DqbZI/jh7V/2+iL7OewD2/yPZ0aZIefIvN/hBuQIXB
bDpAdIoXD2Aaze1eWtQeFf0mEjbf6+BYXWzgeyF2JI8W1svNHvUwLTaa0N8fV58zpeMMMca6Q9fw
3nefP2HeqO4aP2hMkVG8k31tsi5YnRq/TEWgqifPx0Rcc4ygD+XHI1K5jlITj5HjfJgnbTPkjDsD
5tyHYJFWN53Lg39UA5axS7RiSgrHzoIRIvB1GkE1uVT17m6HPlQG7uxj80R2HBwYDhkUKM/+7hw/
/N5qoMVMfhsVQD7XEY6xSIPBU3Z37tHXWl9QcTOCEJqlv7NyUJNdItgvrpig0BTMk3LaqMHPEPgF
jS4TNyeb1ELV7qfVjWzwlOXD1q8gxp5u2+z+bbuVK0I6vefw61GSZ+4f4IPyZz4+Di2pSOyXTt/E
FuBXof86eikK9AHolh39kV0uDV9b2jMixVFNiBOnTk2cPvUdYFxG79HbemGQ5caWO7Rfm5i1fDxm
v8o9cFGoU7ZtOxYsDKCatDGAlwz9YCKXVFMcSnLJqrxEV5Vf+OyCLyDzu+XSriY3f2mrJmvGXwLd
JEjdSRhrm3/7RyIU9FWQNqmcG/ncFtdsXDzMFrWYDD8+JKlu+2o/LHF9Yd88KYe7HsUgljj8XGYq
x6VCLHl8GEV6RFxtpyv9AWvHkgpzKp0A8vzgAV7TSTz+QAR0E0wXnh8t+zfDruEh3MZ9G3UpvnDP
LBxu0eFirwpMoBGHaw3N4dV91OaIqdP9oHugsbowx9B3unD8vW03BiUbdeoIafQ3QHuseH2UWfPH
uA5wyp3s2RzVPBD8kEzEepKHdFQfKM+aXjel700+KOEkGiWKcc5N81Dycq4o9ZH5V/lMBGS0onlY
5nSomBBeiBP7aqbKAg5edRoVwkjqtueUivz0n6qwDzyQg4hZ2VQptnqMxtH71sy2P1kGlA+8umnZ
pnuJdeW+wE+yn4tfJifdITqT17Y0vPFaMCnByVLetf+JaUT6v+Icj5KPs+JGEcwKT0k/0p5DMBBs
f0MAUdzV4lmJo6qMDxhl4KV7Mm6MGVJoZgbVgt7g5Cf6cJ6h2Lt1VR3IzlOKs4o7jQHvKItzaf4m
m2l4qOMyHrGOiD7NEAraAld5KytSTTfoC5RxlXBTHVF20IFdtGj/hgcGnGSL8yNvDY8On5SLC1b8
O8txAdYoEWW+RQ1zjO21GmyLotZBL4SJfOH1oF28ep/wXErkY1R6xUbBT+37FT2M+GUCfq1PLndG
+Cv5P51qGRonxCxLr3XkxyZ0aB7m7Sb7qc/0ZsiWTl60rW6PHCcJS0B8MCT3ldwEGw7j7lONryhF
USkuBJqFpteN1ew3gvVmqZTbDSzgcVUttdqMxYDJACTNXHjAnUex2Nykk29ruYBKioG0c/KCxOzZ
EbhGhhYpowSlbma1x0fbSKo4QzdS7aEstr6Zu8cMbbUyACt+U4x4a9U6Q7cFXR+lFH6TNK/qA30L
gFfxdDzhQpMhdwQU7BJW3KFR7JnVXbNI/ZBHKk/hgmGXWznNoZI2t6PexgZPB58+RC4wIYFKeajO
nAYFLbvUZJtZFxLAQShNSmspoNoURfY3yBYDxiVuuwr7W8dP8IBta1LydIDkwXYXA8LDHIFI3nbk
5cxlLayPKxcOHTLJKqEutiL+dRplu9xpBcpfA/W9cronVl7sMGjwBoSL0HMhlPrcKjo89OynHskJ
FUb7ptSM6gkgqzs6Aky/yrvQUWuO4m+pwEh02Ki5UqKUDDOwdK88IH54DopZwkqc/S250ZYs+buv
OPJFkXPKgS/+DMDd2g2U9+T3qC8K0F853k3vp2NLvWrdWcQh2IQ1rlIMsbjtN6as2Ryxj/Hz7/2e
Sk4XVohCw2akrWy1UN1+Tz45Z32hxPmvm3sF4MLDsqBnLSfdXj2sppzM4BU6mUsDydmEH9rNV0lO
KlX3wocmas+06mvp4r+deYcKAxm3aPP9gYXyWTT7DimNjNnjjaGpn9qC5MiR4g4k1tbXDnlzM5Ku
PigpPRKrcsdoJFPRVNq0Sn4rYATCFT+EKpVuqkUP638/j0Tz61RtmwEGS+b1EtofXePX64LlJIX3
/jICMh3ZU9Cr0TSLYjDHsOUczkDKTOzZAr4RlwS+Dm5WdQzL3Q9sIF77aiiFC1gUuyfLI8mSDf9f
AZ5/738RZWsceozLSKRBrsce8KVIM9NTtliF1dJZv/ZvZYCqNSnCKqddswPxtH6qFoBsNN7M7SW+
oj4ZBC0EdeR2FpUh0aCTAi3C1TRKvO6V9nUtTCN2D48D1h8uzugC6AY7bWcVg9H7daRY0z/XOerK
iS0bghPOUVK2Cl1PCF5YLHVRKhSSl1Je7FLETV/1brCkvwkQzliqq/B5doSQ+9QU9MeUWYROYYde
VQNaoxQu0B/iCY8Tcd8eiwLwEGjTTsCM+AYf8hKypxNIxSJfnels/Lj9TwxYdK7KkavkKYtUM2u7
axrPiBrA1qDq//kv8Pcp2sPJsiBi/+2oLzWG7fnOyijyWq5B+vIkJYD0gbRvPBQVGKi2Ztss6SPY
2j2smpqUBNHMWP+Fa946JW5pg0LemV3BC7NTaKi09XyvY+eHbiCtiqwYsCqTcuqErg+1MPrZRDih
ZdNZBKsCCJWrmrutQIVS9LA+WrwmlQKui5ZVFupm1exUltulgqJKloOXUQVQkIfOyS2vzmw92sBD
JKp5Sj7WdjDDPJJbRarrZd18pl8f1h2NeeA0NJ7byZhilUL262PEHWazTLAhyiUXa9949xt0u6Pf
dJQrzG4GlWy74sO1U7z7Sg1tR+4mTk3gIMtftx0X8qr1swi28mAj3CgjRPLZdREAK9MSed7a5Qdr
4ka3ERjXXrw7Hi2EK8qMmWhaN4ata/qxlzbwLvGVRByag0DhG+1QcLuCPf3v1dfOiqgX0iF6xG18
WkEEmmFbkb1YT3tn1KYTh3k/RnsJe6t11rI1UTxpM3CEqWpeeEmyjXzlZB+MNfkurj/4FnA+iKYZ
t49nqhpN3nmFJMFen1qUMDfrDx2haM5Cnpbc8/BkOMqN3VVqQ+nbXzMac6bUjPaorUep7/v8Mj3M
XoPz/RLmV9Q82qKHYLjo1w2vzhyzLPmFYy2xVzds4wNUsJHsHfyce0HcgdBLH7wWUeMZ4scOaiC9
/o1RlJ4DkBlSe7OTzdBXhMacE6CFVfylhSPMbVl0v3QiX6uYPlnsBmxmgWgrFGmmZzK8ddius6/W
Y+R1mfLVdjiH6SgO78mOkU45jLISgpvBYpbuwV455IE+Kx/c4NGUD0zssVoX5R/JSCdjQHAkL8f9
gx0if54xkEEbeTMxhOy1n8RPMGwfjTbP4uN2i1kTRUCjU4DSbB40NvTQZS1g5rwIGwcJSXB8Srtr
OFZLfi71wCA2DWQ9+YgbGFJ3kAO9AX96euRge/X9NTNlug7m+XdAW8ENUjup6Xosp0yduv8x5i9n
6uG5eTvA/1SRlThFaypbed+uVPOP6A3bjkk0bKyYcYTnPbBNke47Ndx25iVAhvb/wf7Q3EJYSWJC
yYk3yaYXRNJDWH+shvFgCMgWsICDVMBuRmIJgg5AxwVcLm1Qe1J9ER6hil+aNEHCil9OVFkgwJNC
Lq7+3Qj2jH0qvdIm3wxpYPBc1G68MTJT0O4DFpkb+wtf4urKYXCqJQ8lQTr5VMa5TDSPn3rY9T+6
Ea6nyErbmbXgXtmy3JaMgAsEVvV7IeCS46UY8HVHUwWN49Fb97Alo7xPM9EUc/bfxhkY5P9Tcm26
5ihoeapLMPPC6+ueUmKi1yzbKKWOmumfhsUPjN6jvlC6umqlh5UHe9eer0NpaKgsHPXBo5UEfdTe
0Elcn3+BXFUjR/tSEqzwGw2NhyE+WxpZotEiAb6nRtN12muMZS9kACUsfb6Bs2Ewsz13XUlJQ6tV
dw2mP9ojehJKvpeIx9tHrNXoxH96vRTu7MaL70ZRRSf9MYea6Ajm6N9UM+nt0O27l+Tvv1g9Gum8
If6H/zlL0Zs31H1pQrm8idUo5GBz3izyqKYQ0M4w1N6uIeHcWV9R52slFDIiPlMNtc1B087G2zaj
zFen3mAf4O997RfOW7wy2nKQWlYwWJcxObDkZUJx66uuMwr5zApgvvt7lQPOC8tq8sOffe55pf8c
Bk7sV4pQEh5omaVp9Mt8KM1dJ1EHUvg0SvQZ9aWAcFmbo1oGOomuCvkHc2wgIAzenHJqoouTeFPz
6fHqzuXVW54yc1zYbRA7peADIfeKYUWmjHvigMBYWOZJo9cqvnNLQtgzBC8A+MDmjtYvTnbHyK1V
wr6sU9KnZVIqnJkYE+wIei1hRO6YhSNYMLyPvJFWgJ3sGVmnt79z5yzbYEMjakSMw9UCeLt5Uytb
rmsdsZl7goBkzpXRVsXXcfIefwImKm+lPqNT3cgKwCd4cKi3lUmOL1sl/V8s9cRm7VHDvG3AiX7R
6u1G8O1g8PvCxVDzKLCl3lVxOPx57wE3XO98jMnuUY+S3OM7vmljG8VybwHq3ELXTixAW+HEqo4Y
ki3pYhV9utLgkrm/l3tygzJ53w1O1uFtTvJOX7eZOAPfoD0zSYX0L3aeHVTLYjcIUGiO086MvwKZ
GFUCI5KsxFaLug3kFkeqfvEh6He4Ouh2RvqYHACdxgM+3Livgf/QHzfvk6wJDVQl9nUpLoj9rekI
mVCWDKD8RR777UOrDqlV6wB95JzJR7cSeJs9nxLncm3gLAFFcqG0XObYpQZ8XSsg/5+HOKHyM71H
ePFsoIljNNPkgG+SdBh+Z9t0fh9VtaBqLbAWGQHNX/0BlIWkvHnyyQ52fUqaw8uY4kyrUaTVX2cU
NuuURFQClEa1SssrM1RjM3lf7XP7Yq/GNw5OTW0CiFD6Y7cuL83bn0bj3Be3fHQcCiSf5gsLyJVC
e0J0aYPGe70HrnJEtbKbxkStyqzPoTEMxXFziki7AyJT8jF8dr2hvPSoXQL0J/lWxDUVTdjmsNBB
kV6EVLQ2B5yiJ/8SabQR2mHBt7WNrq4t7Lac+7qhuIxFT4ADKzf8Q6YHq/LRMWSKHjgxEd4dMZ9O
Y/U9PbJPBEQgL4fuuNWH6tXS+p/zt0BnyyVYnBFxsOuPS9zvuKNqTMzo0zZtAkIQP/klOjtoYw0t
l4j8j/kcNIsQM++KOt7sFnuGuBuO1yapL+xLZR5WfvlOQdrEH6aepqb0lpQ712j8xbe8ZgtNKQNA
8V2IA6rQCQGaZXFAtVOAbIh/Gvkkr9kTaLdL0mALwi2sXk9XYMIAPrnXVloV1YUFC+5TX5HWX/+r
sIgUi4nBcHpEAD+ln+sPOgud7yX6QXf4j2qpG8jcrc4CAA5tWfv27q3NtbOjvSqaDGqJYHWhWnhA
66S2JwpFD74xeHKDfFD07CVKH8DhWYxqAfP+wJdchx1dKTIkh/WGk9d0tZq3A+nrJLveh5WHQymi
t+wF22chyP0llj6VCxn5U40/5SFZCGWnaqGEFZ9zv8X8LPYMOzguhbRRPf+PEe6yBnxCQl6RtlBs
/jBmdUADtZfUWUNIq8CjiYHblK4z+kzdWfuG96aBL6JIcTojN9kmUtdBAFYYyWFhR9ziZNP/zd/S
ln3BSQPiffCoVQaKx/QHxTOybAcZtKLlg0Sos+sgXSRiLknJD8F/hnlrgVTmVxts7UQGnK3siuMI
mAtfUmQ9YayG1zKfa8Y+LpRfZmEUXdH+RBv3Zv05mQ8g7qc0FYoBksFPwkOoZM80RYX2MWT+VjuG
dLRDQ6ftANS0brDwsT/JWr50A+nJ6EtgHcQsDDNi+Hy6THxb0KwdoQ4tyj2mdjZD0upV431bwjsg
WyTTMLsdzYFsTVaEaTsXrnGNZheQ7GaCPA0UgW3n9ta/v4X5eMQqOU33JZBB/xq8fwNRcKCQpnkE
TD9C2RU7wlNPQfum7Fj4/XrsDjEzOUc743X75L3S2J6PoOkS+hDe7sh+GX9Rl4CWVJUHYaUxv9JA
IOEEgpEtg0m0z6OCgDmb2tfOMUti+pi4zrqmM7t424qvbpHEe6xg/du2mLT69YQjGi9mEoqmvmk8
kMWwHFDnMvo8qVJYTNBPrrvVt+6ZQ/glXea3KKwyL+KcOspcjZEasPWDRPOxdmUVh3FW2N4eB4kg
ugGSLqAJPVyJeiCWdeYpMa1UtZfCeNbfYsDH/h71+zgmw4x6v2oOZzIjsCkKcvuY9cdEriT4hEZg
e9wIPeAmhbcxcdgEo3lN9qqsHNXPwryhimp/rIWmwISAIx9MSG3/HPIa7MnGGMRLPctgOyx13m4h
yHcdlrKtFOEtmbxENON2wP5eHZnCnsl8brKjilEQfHZ5EI2/L2J+QT/8bGF3GAKJqy9cURcp+19Q
3rxwNMC1IPXuSL+CuDAIwfNptHxqQWICSzcYRZ7/sUOizaexFhZfyvxLmk879UbOIHyJTM2f41Hh
oAkynDBRzc8T11IUjeSdROJ76Xx64pi/go0JelY2NUBy3S2+WkVqh4foSdpLPfxbxh8KckVDFEut
k4nXJzbmy02yYlinaJUStz64UiVi+9ex/03CZoJoAM0vCb68mUsir/d3l5pAnlYAUPl9c3xR0OdD
0+/7vRHCVQcqDoXzjLfceQRW7gOsanrlw0og7ICOEsg4Xrg1NNpTaatl1S07Olfh4PVj0q7bBp4K
Z7YKMtwOK47np6B58MECV3c4Rn2l4/QqcT6UvldB/vm/qLY9eENMiTHvdmAW5qdigSgt8v9pO+C8
wPrSqhLQnsi3fT1uRH2Bz4XtP+RZo7xQPva83mQiGKxHddTnJqfiC2qphRNq63JsEvsR5ap7LVq6
J/kK8eGKBUoMbcqYVegRglrizuGgpgnMGYHMKduGrsXcKHPda0Xxyokbiug638IzxQzd6NvbLnM9
ZmbxDw1lXFd+fpK60Hpwi+jzDXbNsjUYPAbObAmfYqN86eWly7ZVsu+Px85yAEB7n4szNPMyxM4N
Fb4aADOIHJhiOXoB5gGM8kIyXGTjaCbT1Aamt61Ys4rVyPODtL9ztRUzXhcFyWwQ9lLl1Y0Xci8t
T+ymnp5XLPC62bP6JXzhFMO/Fsht7cydc+CvftXaw1p/oGVxBg1Y6rF/oib/ruRLo6y+WPbs/8qQ
zBqEIhMfZ0U1dAmHKOEEjhR6f/KwJgWDJPT8M3oYVxHypR4LI0ih8nX3ApiXyNFo0XE+7C+6dagw
GOG+RUk5hmHMY/SN1QN0jq3VlSkVbIPQOItrxIHyKwx8ojUSp8kMK8OtRu1qNx7CqVlhsJ6JAR8I
1ES6ED3dNSgUJ2cPgBCZeOd+PkBmE51tQ+dQlVu6ne+aG04MLsdc3jndwfwlVzUOlV3HMkd3GehN
+aDsIenZMNU3OdaXMzf11LoZiza1ThQq+wNqE5bTTx0VFiZ3pLRAsoqn9hdWDEJrafzb+Y9AJhZJ
NRV8/LtlILzduDBM5IKIWtEFvWN/DEhMrSd7FrbTDC8LM+LxTPws+BZljQRZjqhnbZNHKAgwoDJq
vpMBG2kPrA8H5RhB9zOCrCzbUslLr1bIJbubqBDumj5CDxWby9SkkkHxv3tB/07oKx2d6gJ30NHk
suqcu+51pk2Q7yh3CTe+bxUtzKZeEybNWW4x9DqBR6k0cwe+kdGqDR3tEfDwrknKUW4XdjSh+AqF
2xVNH0RTzpgNeO8uGY9yQU+39/WLZaL8jOPxzYSJT/90Bc/0PWtWANljXOd6OnAx7Xspy+M9GWCy
HFhG/ZF21pkrhkUiaoFYXtAbejFn/lBN39arKsHsB0WUo1grmW5uKI4DagDZJsgZbR8E1wxE7xPz
jNYEGcl/xbZCVAKH3XsJfIEDkf50si0APq8Jd9W22FMIuuZhtCE2ldNAv7mHBPIVvwMBN4G2XN5R
U4pdgNOmo+lbg+PHDn8DywyOmzYp8/ep1PwRDsr7lvAMiIFEK1SK99TZ3i7FHpz6rEHMv8wFHkiM
+rXxWAgFQhsiJf1A2dkqEfm57iiYBv+fPxoTwDaoHCPDlcAk7EHiRErkEJP2T5/i3Q+ftHGgkiMI
m4QQ83wsXdD8KsEPTvuZ/DyIfrWc/OamdXsdhuQztsPMLgu6ROu+jYDEqQC926JDEwnULsH12fdb
q83269UUxEBSAUeR2kNcJkV0VcHMj9FOZOUtLhXr/tyJSlLKQojT6i2EUjFDfMZ3slyvREBI1ukX
dsN/+lE9PaGbboUiJVcrfHUGLJ1XesMZpRVpDEKKkL6wMFumN2If89PH5rxGbcFsgH7PPM1ssh/S
+VqizV9R8K67PFzKYX/7xlVNO5GyqyQKB1KpUzQ0I0YAZ8JD4iaIMOODwt2bGPbeiH8IsGT5zDvT
lQzm1dBv2xpNzrqckM3kw2qjUd4HWdNVBnikoUjp9KjxHNu3/mA0XQ0jA3wzyTYWiGTVS87/y9Lc
d5tSVHiM+7VtTxxoBIuZctktar+lyHem43CRD3BTdG/adebTDfqfTdNE+tM0CPsx/PffWbbIyR8Q
K1yWbgLC4uDgJJo4GVu34/ycbZYnMu31qmO7QGXl1457VcxGgppGgjd843J0QjomBmk1xtchcCXP
noEweILRmKGJlC5GhyZcUshzIz+CbGA6yIYcYgyiPNNcRE9eDCk/dyIYgx+jc50MeYEla3NGjJ9Z
d10136m3LQx8v29glIUY+wjzreNVwHoOHjEjcEw+uE8hFoGt25a58+E+NuDwowOiBhg9kR7HK+dA
G6SLi/EK71ZhqinjqatkraNKtA1L2qP6AdEwzlnABcP+oJV97Qa2pmpm0H3gapoKyOXYBXtB6aza
enPAfZLlL8005j3L6nSU4XXInWGa8wZv5pAQPg0HqKC7/K7pC5EIBUXKlUwI56o/FKPJxTx8hKHo
LaHudjPcjas/4G/P/Cgw4+09Y/MW32klhCbohPommvFHL+lkmo4QHjGih0oxQbRwY2wbFGH9abiq
9igr9BRnmom8BlhSr4L2QnKWypXsWN9t3vc6E76lGpa3+Q0SVXs7bKwKDhK5637OFyyWoL0QiHFh
wLg5HgQWSbcM32ADraVWj2C4+HMISx3fZGYOGnpUWj5YKjGF2n9dTx2z35+q51Hf6ewUkCfSju+Q
i7BXUFngdbQXJsxzEJPnUbjeC1h3zcHETj/xnYIEWuL/XxZh7Vd8AywEmZ8LTY6UYdSBuqX6rgRS
5HbuoLKg9zAoA5GAGxom3tny8bTb/vpz/U6CxxfcxGQsqC9z6nSMlDHmeQJB0pr0lrquJi2nx/Q8
QFw83gKXwf+/OLBkh9qwHbeptGErPm2Htck7v+tgKQcvvfdGp+1XALEvwd/zBYUrPPo4PNczX4Qu
e/I6nOVS7yexyyEFzMoyeICvhQFEyDcMi0YN7A+VXiUkjfg3izDCLgh6AbVuBwHwsbqrSCFoQFBr
WX5fJz9RvL8Yim1dE/425zxz7hioheE19AK7i/fnfMjf6TRx318v7Sf0qasody3kDabcRMKnPSRl
Cc67Zcinb/jU1cgKubjI7mv0RhTYf1YPY9b5oG+YYbOMzvEuURk7ycnKcBp/+dhdrU9dWKtK+bm1
DJ7y2CQhvf/xIVYzhaEKBiBiV6Z2GRlHQERUDywq827qWlzg8v3ddbV1eHCoKLtHCksWGOC3J240
L2qhCKpnBVaqj2ktvzxOwx7vfAywl6oyl5ns2+H9NYnQb9/QeSpietyRz70SH5C5Hi4H5g/a+3xb
BDTO+xGkSFcaRWIhs+R3dbqG0ectQOnucNYyNkaylTmi4gKmnAxCXPm0GlJ1RgvrGvaU6c8SjfbO
bvqhjq185EmvkpZNFD2A4+SSSnVhOn9h5WqnWGdWOmmMQIxq01ekw2AV6yh+LHvPnMpjp0ExjKui
HlvZ/FLDwI/baHuOO631rz954J9bLfTo7y/qby5+FAGRpfZxQ+FcmlGiQJfTu5ZA5rNwaeWho5qV
3TmxjxCknjOrutHggFzuWFyL6gebnhEBhSeIbK991Hk+wPE5+Xs19kup0NCK6Cr/fqZrV0bAdVxx
Gf9aTzVB8VuPjaHNyPEE/Jquyx+Ba7LiSQ7rHXHWRVligHhAMnFmEWnTX9qINoVB8skUk2WiTkqi
JYF/hPk23TaSBNKEeOysrJdd6w2lN/kGWg1weaXsBJANnC5sDn0IJh78G2KKLlvk4ik8XUhf/FZI
yJ5LkqJrWCx+cpOvl87/HCGyMHN20QcsbP45e7QIPR1UFSemgh6JqZmkfMkvYStM8Z5oyVaVQLWG
abPokERaMyzz2Gs4aQ6W7RFq1lNovUOZwSr0Z81az90WHUz/y3GX1eutrFzC5FWZwU6h9tBUnKS4
5D97nRC1bD6SSpVgoOmAkfXViGCU1Rw2t9ohB+FAWqKS/RI9WWCyfSXT+n2j0O15j/OyyI6KhnZx
npCtM//D5DPx20FRkWjmp0zQ6CEifRmCTWOSpkqjSbodsxgKeN3pRDrlvF/2pzPLGfHu+psVnTcm
7oDvrSdZEYQxHbqVaINCS9r7R5/6cY8gd1c0Btglgbszn7HhyyxwZdRkA80BuiaZTkxabEscVskY
jq2se3G9gFFd9h00xMmgPbUhJnRQ193Dly0QTOsLU2HBdVozg6G9axndyTSeJBmByS7bNdBJfvQF
5gdtO8uH2vs0f5ee4miP9y/JfTMdcbih+rgMjuvWnudXwTTXLLCbC4m9CVLH2F7sOtRItMNvHBIa
8GGX66uzS8fu3PluKE9wS/l6rMSKoI1t/tIPO79C5AVpopsOzeQ5nmp54y6kqMf02+tCY6G6gZmV
cCfK488IMGfl2Lbiv2T6patVR60C5V+SnzjPJGz9Pm7bbxpzM+gZ7ApjEKFWk6mFtT+SLvHH1WHX
KQCR2w5aoV2q+TLnxfIdUKDKK7Ov1XRigrclENbmulkPR7+QOQ87Ds9L+BYRcQWwm1jar94wKGGi
M4n4i/KALg4FTUH56juCxUPu8G4NpeYPeXB3wfS3OuQX9/Sg1NtPGZ/qxcbySTleAOzbqvlQhDu7
yZH/2aIEQ0RU7wyoJzJNnFZyYfayUGSqw+iSJf4/+U4oXbu1UeheSInjUJqOUSXAZOmu/6OXuYmt
bqvnGttELtKzuQwgmt2gOODuP9Bs0lSAch8VM/Vgaf1X6FAok6XKGog+sBZy5ml7zh9qTWWJDlyc
1mqxh1LthM5st0WJfCAlS4qpTmBOB7fwSPx1tlSCNBNC+be/z0Bae9WhbI993BvzbJeO7N7YMSJl
JudjoBhmMfbEwVTmCMIal5P2wxkh1S/v0eaob5uECnaSjhHMVd5qR0n9mDh+sxvbVk+cKZ8l+5Eu
Gr2FPhUuNOI8676BkYlQOLOg8kG97YORvtkmwL1ohJrW8+1OLW5HBgudVPscInUm5puTo1Y+05Rl
uO9XjiE1FA2WUJ/h5y1+ipQOh3T66uxP64azKH7JV5E+tjphwqMSsRe2UCMLmZf4Z/7dhfScO+iz
ieR1+dyPmoUV06VycaNbmJIlRK5OFfwy/0BkFBwwVJ0C7s74VUkBe5SpJqWAnfqZQYtPV/itIY1E
dQYa18npliNEKlNzF74nQDs0g7QECGFwQsmSrzgMW48Kx1KdWxmocnB8dF5gClTsjSGT6HzKHTd8
e/2yUkzQUDp4rLgBj0KNeao6UC4xZJ9USH++Nj/ISxCj2SxN24iXQ0LGGnLzEoOgNF6VFkPECFgF
TRNL5Ax4Kf5qesiPjE0oFCEbVzPuAhPkT+yUQoNv729Dgtdz9qMt9KEYZ6AAgBBTMJlU4FeDwlGz
nwQQOUD29pHNj+E0Wzx9cIMeRs6Tuhf8p6ryFI+uvOlWbOsU/HcRVt90mCH+40alHJskAJ9MUYYB
3dQax+STIQFRrRccmU0IZuNXUL5NWHZVKLLNuQLbZK3ApdQ/CCWNK5Vyj65bviq4OaCbeLwDyuM/
cmv5z0WOuPxpm0ENV64hX6EDwZ/xgdRvt3dXMnqyM5syKKAEX+NnqiEECeSv5P5j6yqUcxNI/uQF
djmaMDaXvB0VOyCM1y4AiWzLbL0q7YulDF+s66A3MS12SnAfB5JPFmznNXJttJ5k+vQog6rz5bNv
R0RyxeGitguRMfb+w8xnb3vMnQttQ7fS/NWuGF2aDtL3ApviZRzQNBPT9x3us1wRa0C1HrRXvQWm
GDiFk/ajn98rW5lm6gG9C8XmKwv13nKpKBuruldLrRh/cQH+12oFv/MOT8hpn6VJ8WpFtwMmqP2Y
igyZT0Zm4iNZ0iO/Zu/lK0Px1K1UoAuvlSmi6gJsebTxQnaaPP52RRETN9/XefTGEQuK74Dt3z54
8/WvDQcqbVzf4JIuzIkInesDCV3dyK9mzhygDhwqLbv1mCmgXfof0vkCXwdnjrBdhkPHQz9fXLS+
d/F4PIy5dCgxDzkSlS+Wmid8WcrAtkAmecNo5tyJMsBXmG3b4vCF5FJLdj/QVJI6LZG0ztCEi7o3
Z8OE4EW2PmilMCu9f+bg7tGQxl0PJOxR25b/z+vd2FcvGN9T4FFAOQmkuPgFAtLK5Ryjvsu7xv5P
8kemmshgYcDSwS+jm0chwpq2d96brjvQbKNLoiJy4vI69OLUe5eL2HX6VLdvAezy1Om9UzmzJD/+
St/uHOobUmfI7JSwaOoWnqkKIgSEAlVkkXZWsxLt/+xJy9cEAqFHS89HeUWe39xjfsbJq3XsxxrY
ge2Elq9ANFaadpVG8IrKRQOWfR5DM394pSeD3ijwD2T/xoZFZSGxKhNuCydJxfOKvErhOtg1kK2W
T0yPmLe05x9HuMPbyEPQoNZEls1cW32dF0f3m35cJTtOzSIWWHI86NOJVGc/DbN1dZUV3X/h1cxh
SHxTdWQ+0NKxEcNXDDO4oUjx26Z317f3lLwzGDMC4LOsSZNk3M1k5sDQiNnZoY9DWI7kzK6JUY4W
EtRZZK4n21Xj7gTvJ/SdgOn6ISHi02RcCnXybLxnnm1TlBpDjdhC5wkty780PgdY9vpt0P6522hz
3A0SEZYsAm5dJHJwkxXa7TBpXFmH3eK4xA5xvPr+w8dEO1BIO02TEW5Iojw5Ev3gYGg2ko/813zz
ON7KoL1NUOwgQ7YHJFBPsyujf31kS3/p3y4mM9DkN/IdzJWVUmo4XspBDQtlvf7yf5k+AIXJ+pum
UDlvn/jPkI+xVvYFZRUZAS5CjysndSmt3pS0rfLMiHNLGyNrewlp1geamZoeuCObt19sJwZyPXoT
BGlWVHJHbpXi75PnDQkZ92R0urJKUdQt3DCKnwHkye4iZ3wCTtGj9JFDaVlfHAwXOaPeg0292yLL
Fizt7bsb9uGRYUzyVWSVMr5c035w67c5jsuDaxMEmHyhrY1Zod/tezJMjMtzpoibOD4gT3hGaDyl
FUo7V+uvQ2CexfFNVBWj2ha+3uCI7sN/3WEZEJIZmAHemPdU7XjcWvbefnZnxNlEB0a9lryP6etf
G30XwnRnm6CPv9qj/Ue7PubjI0Rpt0KKdt5F5abWrgCMtyn9cT7TThmGZkd9YolHhdqCET/qLrzc
mrADcs0CtjKnZ989vdOh11dMXM0N80aDtX6mUmeHc65aJf2S1xy2bU9KHw2cZTVuEOcY22PLHjGF
c+BxePC3GKlvCKpF1Pa/nDx9z8RXGWzeur50hl1VRTjxDeTSfuF1WTQYzf3pbex2ano8Tem6qbJx
+hTgDLn3wtDJI7Jb9/3maYaR+8a3kCvpcCeVRbF/Uj7JxedDCxTeaCFBaaAQpwH2jeeiwVbrNeLk
GYBQE0l/zpfzcye44t3diUhr2GLQZgidSiIwrFNwaiz40PoE28iNKnSKbat+BkhXhYTK5avoo4Vo
aljVdVq0lwU/8kZdd1No893K1novOH5Ky6H6lt6kzky5zlPS/pGQbjz/mSlVRpZwG9bfr+P60XHx
rGW/dfFXzbgJsWwrMi/wBTVUD000fiEaWzPuo4CQjpGX7pwsLk1t9Ad1J0flZ0yBXVulw4VjBPg2
gk9Kf77Ou7RnX5JuOIbuJ9zHemzIpHn/bKlfLI1Fgfti0R9Hpmgvhs7oSaLvLqtNelDPiYnzxlbY
mp9QVkdcriS7BePG+PqFjNz/+pl2Rai0TZhE4MK7f4p+TDn37zckMQMt5RlsErZQ4hCKf+ZVtMoh
VM5oU81cXYfqcxBGR2xFhEKGFc924Edr5DbrvjI834OiMHNO95M5TjXwXzFrz60KmgBbiFGa24My
si6AkHY1F6oG6+OcNgMegzf1O9QPdYQ44Hsx+S+zCDQW5dmlrpIvGIGBiMAHPPZAiYV8zkTtqlbe
v+/4ADknlv2wWMqpuNigqH1AAsChpRCxwsYNFI7QMo6Wk+jC1BQxLQZ4C0N9YB6lqFt75dJpnG2Q
UGuu7fBN+5tfvszARmb1LrGyw2GJy9GkPPaMpcpcTE+/4PggFk8CPTHeJm9NHgxWdMtGZUwX4WnT
WDVaD+2AANUt/qar1+pdn/PhztEd8RFDREpVdclxhTrhgkJwwLOzypPAi9lyYuySy6q+YVzHfWNk
jeAXugQFAMrBdI5S3I09T85/JjPdWNpPLYdNIA1I9/5YjDaKqdgj9FBmyxPj0Saoz2JoKxoqQFig
pNBUEYTU2CC1cGNPZT8QL/xvmg2XnapG+aHWya6dheP5qZvy/fzQZdFidAZ8J1ACyYwFrDbzXH0z
7FmFGLPhNISc6WjphigETXF4NrvKKR3OholVzRkA3d2oxYZwRhkpx92b6sHKsH9ccWCuTtn7veLt
IH9ik1k1LT/Bye+lY2fWAWwkSYFwvoUhN2f6k0obYKhLc3Sh3fqlrGctxREQshEpjis6Kj6AY0Zd
frKxQrQTQM1uPcfdDa4ixMemiJyH+6rQyfMU9VvH3//BIsGYO1E9utuXIkM5aU2YBMJK3VegelBM
Mrcz+j4sBlgIWl3/S/tfvuDtRAY3CjiqnkcPBg564EapMBPrJRc/NbZSl2qUMuL4zxQzc6aQ9t25
gYgedEB5KUV9TmdbGXphYnVt9PDCuPlxjxoH/Ws8T2onc5NMuf7CJQZd2LKuMnMOsw7YM9iCfG1S
jmgNYA7GLf0tML48HtGmzTOnCdBOciNcCoW+BKfxo3PWtco+lZx9nUAiROwKxmNTnf7zAmcy7vim
ymFZAGBws2ZLfqS8XStajOR7bmhAxjLgD4K/rd6wnn5Xkqv4GYmCnYG3oOqnopqxncTyrChs3r1c
qhl6dVRXHvFmQSf69mzYd85Adz2l0USJB79odtM5o7TFvcFzIfIfRKJCherfOyw+u3lxBUOnB+VC
B0hsm3N8qGYSAY7lIzJl479hvuSEovMwUXc/eQsnM2aL7p3zXYKjXLl61xQRzfuq2uB2rTEmlfUm
uihr7A6G8ZWYZ2T3QHfVKlQ0SpjZxBAJl0Zzk8kS0XH6/TAAHqe/T+83iXEw5H2+t+jcsughgRRk
rxSdW8fhCSJ2kqvTnakBe1fQqhLeWozqPcjDGr7euNXQWhck1aZIC9c+C26nMPZm31x+tnD7AlzA
/I5SLKo/N5WeAut4+Jn31XrV0+3nLIlHK5R9+yEKq69y78c3P95A4ZuiMdUkJCk6sBTT6OIIUiJV
hfunr0Vu7Dmn6EeeWQogZp6wzFMDKKWpfQK7yVlepqnBWR/BGHPiDscVwD2rpLoJNGGch2lUT8Th
CoTye+CrtK4mq4Dgy5A+vtas2XWMDEebI8LO5ZoUWr1Rc4Q6dYHRipBUeP83jLKsgi6wCvSOkkD+
tBtNzxtJ1dnSnUZZOn/xK7HGDjLTrpNqr7xSImBkMAUavv4dskHNlrDdCXxvX7X3mvr5VoU9h4RW
r2b6mALnuzIsgFNJEZ174gKex1gA/IavMabiYx2ymdfqlAkMA+a3legUBUbB4jOElFxNT+EmOwwo
Y92MLkpn5lSlPbvORhISGWJXF/otSK5cO3GfIWBwPwTHD9qV0dQfv27BrzyrokAimYU/bLppOoTc
iYbYvG3NPntlhnOzzv0Y5+qxsGyRPIaPu2DQuqcY4k+AzAlFsONUqM3YkQ+92nom2wiDHBp6M9Yo
FsW/OLwUuwDfOfDPYGiVe4qWGwNDymStn79p2dRezep7LodHID+T0TRt/YjJVXOlCBFcLNWNYkTZ
ETAcQBj8TeBSshAny45nkjHI9uJefCfj4sw27RhcyHCMz69+FjCI5b3uD/bmj/NZAicyxUxSWYX+
gxvlVg/vR7HBCKpDetZ78MIN7l9yHuKR4H4QYRMcG023SRTMDEvZx/KAybGGzffIxjaf/7bWgEa4
i4UmDmz9/B8dpEOB/k9Zpv/c5K1WeVv6rWYXW6LohiM5yXSvetFQSmV/jGx+Vy+71oxvEEPFnGMZ
1O8KNC0v8oWVzCG4xnzX3cmiAwUjitsA+uM2drKPDuhk2ednCSMU4NHpzfezBBuwkjHvnRJ2hirD
cF97Y/xmPvHMqXHW4EUueDIG2N9wajWyKkCw/FLBN8Bn9qaLzxfPL4QW9OKGga1wY4xUUuBGO5+s
7HsSxeUjIfKqsV7VX+3PiwZxc8f+eyWPsYUZBLHZDst9+LM7z8z3J7hHiHFvW2LjAmlIJQP5zUUZ
IfIs5AYG9qlolGOfSQYAhdMU/9bEYNO+o++Tg/7uVB3q1x7UJg92yE9NTobZqk+gX0P4E3omcsG2
YOnIBMEYYjwah0QEHgra+OLFeIgBbiX1n8HSs64V08R7LnfP26yCpk8viqXTSuhUy+AIBB3qisat
nc4UZ9xUFZBPd9jRht3bAqeH8Ihi0Fn7SvB70VSwh/VvuKL1zs37X7ikGSMBD/EQOK6mPUoxXBCM
GTWd0rCu3KlHoqMHApHDg3q1XOzi4UwiwWqa60NPG9AGVMvZ0r+hezMJ55uZ0oHvUOk2R7rP2QAZ
ymDrq6Ie7KhTJ+93txpeN4zXApRexMu0wkV02uykf3bX7k5ito6KYRkmI9ly0cZ3E0aLppDcZllX
+OVj9MJIcsYuuC4bit3w2Ie/SOkVzfKQNjFBWdVu/xbGPHJqNuhmnAb3noR++uUZNb8CSVlHgx5c
Qwvs6P1ai8JadEP3QqAbcupozEZwHL650iXBuTBnxHHcs+mkzTRtoxpsKAroAxNaEkQzjV/yPj4y
UjQ2QPTmhWWcLYejxx2N0/BmJB1ODbw6soMXRda3MIYYtGY5LGAXR+7m368tcBG5SzGOBY/VBZuz
mN4j3LBJ6OUaFquPcLPWazbcPKJgM3NJOUi9A+hIi+9MUpK7P2lfY4toSAOPgOMexkeJQXlWTjt1
TUdMWJaxtlff7zaMcTCo3AGrxz7HuhTihoTgT8cJ4mrN+seqDTaneTgaLrjkjV11qd43gQVU8mJH
wODzCKRYEi9/h9689t67+uUGhoa5uHulF2fd3mE9MRfzyFBpoQ+ngMFRyjac+36S9qeUL4nyEH/o
DrheAcama5tpFoQAizyuEYbvEn8jepFBgBJT3ofXL+CyF4iKrHBmFvLFprPUOr6Z0xYISW/XzTSL
ll7p2fBk3CNhLGdgKlQyETahQwWMr7Gkfgl9v8OG49TyzKslpCwMXbigQ0DeB+wZ4ruIvyFQTupv
HwwTpguqtrn8PY7ZmtLPJbAkWI7qWkswLcdz83m5X+ebkYTFGoerGt3Xbq0Cixn4v/VPbG/AtKrK
L31ZzYmKSt5Ra5b6qnZnb2mnYyBRGG/3x/ffA05nCbU9Mg68zL/VvJJHgytE1CffLfhtzU5nog08
gt5FV59M/ydX8mxZyqT9WU3QPcRq5yWfchZfikwlbTDfoNnuFkIGdDX/T14qzahDQB2zu+8FycJM
3IuGl1eHEqTU6+cSEBg1QXCL5s75Pd5GgX0c77YYTytfAjZHahiKzLXrgxAkXRSqeFSlgYIxGFNp
yE3LKuISB3Z8tfSJ9G/OEZTJCSub96q+Afp3zBGi2hNJgw01qW8ulCMNsaWNZvFSGpwP1zm+wSyl
bU7YR9KvBjFxCiy8sJjhj1dP+3H6r6Q1nybk2ia3rOeRKKRUPMw/zfv11lTUkzhhFfMW1snli1ok
so+IDZ0h7hTgVva3e0lcljRr/9RlQW8+/rhDdPRAURWTbxsotRlBeG07zb994Yx1fwNDQyKbXPvd
adZ7cwWEhc3MvgI3nkhp3GrbtN3/tUqbmntf2zI5osoG719IoWZ0LW2UbhooclEdAcQDMPjUUaH6
gJN8/RYutoXpbO5S6blq5Ue4aMqsGrJzbzXbYblWekXhjmdSK+c2he5xg4jB84dyncamx+vwPQnS
ybJalaVeU/1w4BMN/WzAc8nv35eyFTipgua560S3Z6DVq+pxuKGfScY/ICjRxh4Th4whejCda+32
/PbF9zAselowTqNXQ95+E4rPiMnztHbFV0U2NeUaWzwm0/IxlCwREJft0L5LNERIe+nYJqNuu8GE
GyJTQVXas6nv3VLd5s/GnlkSlTEM6jhtvhg/YzF6lR6xYA56tEZvya5Fy++hekc1uGi9gEZQitv5
5Kpr3Rkb8SRVao3P0LWf7gShwG6Bz9v+ETREjl9N6qMBJR8dbeLZuOl4qDk9b2g2BHrlfIi7fmWS
2JPovzIQgHuFsrtFvMA1dDcRrXy3ixQw8LYIQbr71BK34ZQyPYg49aMsmEr8HzwcwblOISAf25Mi
U6F7jwSkRDrVvZ3cbv3tRMxmAj58O621vFAa0OPqfuF+pKjJC0awtrld6yZZVM6NFWnrrBduiIcC
crV8LvU4Q5tgYTnERLHY0zGvyqSdvNL/1PYkHZeW0wdI7kXQDBdQPqgTbeOe1OhYFm6VoKiBZ3w5
tQI2vXCcNAYoacJU6ucdf/v5gaBk8XGLHaN8r9nNltUnG+E60bTHmLHhWWkTo1eiTMZzGbcM6kWn
v+hn0N6AP5DzMRvV6jWOsvnwntkM/sPCjPlkHjsF52H3f2PFmo3e0UfVN73HMiocKWwR+J5MEemr
U3E9AcU5zWmtOBfPPQu+RER5Wou7D2mqo3N1RiDlsbNeSMQ0zX0LAxNnrsWIetD8PheaLT/OeLuY
Chp19zvV+6zR15Zs2xbeUpk9ga6JZLIrMNmLOjfC78ldXV8603xO30w5CkDcvQ1uMk6qK/ccFhsk
uEAkniAwQZDw85wL8hT8z/bq4Hln/5pnXmxPwWNlQGUu/CukYMYVRcDyda0QxKdV54zUrXxmWgYh
QSnRzHecZYQedLA47C3kOh/LuGtzWrt8KBrfclyLLXqMAXigYe3cnNqkrT/rN1fFCMVc4M5Brh4u
vyd4bBOCxg/X/R4Iqg5lRnzUGJNi6coB7Wi7YdWPIaYdb0ZuNL5e05Sh5AqcFAPQdTgFATl92KKQ
sY4Xik61HHqacDr3Z5FvzHg9WKOUu6d3HVvMIQuToYRlqriYcFAkn8ZKsd2NvVXF+t/7tgUZ3GTG
l8qFWaWyv1nEvAFAy9g2P66J09fNBGh+OohvoligXtfBb5AHvDHWQMthc0ePYXZQXK6S1l/ko+5U
qVbkoxL7pi4j48dF6cpgh278Bx359S7PR6ZM6XE7rgxru/vBhkguAi/68f2mPKttg7xdRxg1Z6zq
kH4o3CqqGAKmhpx09q//iIgX9A/30CT2e73g39op9yBPQ3ewLf3Q8WiubZzVs7ls+/bgrADzfUmh
UM5Sl03Kvbt/olSQCF6LLAENAQr62CF2wiRTA+nIjFQb5ktpjGtAWOtDN67P4rFfw30AiOHzP3wn
6WGpEkHOZwwQB4iKt55Wx7zY2w+233weNkRij9OpdtrOZsWaK7kYw2mx2Iokjq+y3JZlC6whyqFz
/tBrtBvCJoQxilOSepyq8467/Tp6qrZVKGhG4bM/fwnTknETB4lGXIDiZAjakt7mzkSKagGSNSeh
b9+Te7R7KHB+K33sJ5CMvlS/0X4nLXMSyLnI9gMHTB2CRKSJK//bFyp/2yKf6alSYNTX+iK0Q47e
PQJTo8e3DLHfzmLHw6/hD1DScoGfqoUULwavp0zSkMBRWlGTqg559rcawwku4pE4M3ItfvP1RE+u
6ciLfDDvt6+PLdiQwvcv/OoupApCaOdf3GDvWhBYe3Uz2a5B+28Or1kUIjPx+LhVSwWfAiiTmwWD
Wi63JT85l3U72gnK2UNZycSV0JBHSN7ZKXOkHMwpafFw9+PP7h9j7MRq+MPpL6Gq0OTvlhfFY3RJ
xcCWcFqQ3TUlBLJeefU6El0aVF/EbPTaUT9bSHh8AuVRasn1slAGsZItXeEsb/mTStIOQsw+5Vs6
q7BMoFwoTGZdQlkoqj7Rhgb/OnwsEYFrBwh5M+v2R4tFjqdb91/i5oKIMeLMjJJrx0PWA35bx03e
PSPFtcN0NJrtTskirWmvMOYWx8wKau18tNeCjNlZfIVYH0Xyd4wNlIwUP3NbJEotSFdl5rH3TUVW
YEgIELm1DP7tCsPpgvrW8VPvOlGCanZ9nS9G9ThDf0SkCyUreXVP0eIVIH9HnZxFh0nx6HVcAMH3
dSllTFKELSEkirsMND9iOSleneJOLPwxkMGgGR+8ljfiyaUrhJ9WFetieYfyS3ci1IjtOzVH8FT4
FaRIVfCQ0In7cV4Zz0D2Er944Ukg7ReT0qto8Tr6kp7MXOA37ZOmN5JSAkwybQCJkg0lceAdu5/d
aJJ24we1uT4h3eNG6MhBwjy+XxjTblVNCh5fQ3QjfineCZC3fo/KgK37wTEa6ildJvh/k6Vz6Fkt
Vw8leRyZud7Uf3sif50jTlNmZfMSynz9kHgoIaljJ0x0aScDOg82qFp9e5mm+K6GBtttZRb6Auan
/ENXEG1dg/adRC/EDchMiY6dA14PQPOGwzO7SUY2qql/WwYaC4SfGaOgsrILkmx2bVleFlC0hMTT
qLzML53+Dgufr38r/6s/lfZvckZAoccDnVm/QUiZFmH3DP9s3uJI9IjWAd1qvgsPbOg2CC2fjBwj
7Lny+YcJxn0WrXw2l613TSWEPgh6gaWCsE6cJOJxDDtJ6nJc/2RAckUt9bA/ttYZZfKrjO1U1o3v
+AQshBU+lI39XqYZ8zdfvvIHcS30zB6zdwJE6Xk4HfYMxaGZRCCxewYiYyQdcc+/ltwSdzI/vtiD
7hTtAY3MAtdROVR7yxPpTH9LkJ1l8Uc4JbarCdNRvtOx2ThCPOLDSDzYfllayoscKOwza/ysdCjw
mIgkLZ1lfXgKBWSdiwzwOilzok+QsyhMcSkq8vgnRm/+3cKKtNPKGq4N/IpmI/l8yLQppCugYngK
mgPW5mKIG6d8bzpiGGWtbWqhU39g//TaUwh7GxbTePK8iI2i4D8saUsU4OYtfR+WX88o/94tfxEO
+BB+gqvlm06j+DMaITgTDx7Z4iUHEFb+OTJqyFfz4aVM7EtEgI8/ItdA80hN6UsoFhWV978uY/MO
iakkEnU70/Nd4MCn4e/AVi9Ub6fqrDr1ycJ2HDA2+R/JYtjNEh0LLqJAgmwc2CcwPSDMs3Hgvq/g
ls4ED1aCHSSPIIi674zgH+xPPM9xZ7IEyGhh/vYQcdqDS8hl/XuI9ASHWCxr9bGTZgB0ltdywrFy
NKCatkY/jlogY//eg4Ek6tGG524A/O2Nb7r67DFZENeaLnHkLz8GMbYknXTbk4DFWps8zJnFuuvN
1oZxm0QM1P90245lEqPMOIOTnNf7VJ5NUn3Q3f76y+A0ySE26lW+3HB7oRYTYZvK9Cml4dLA4hQF
INa4Z+gBU7b/3S0Yd/Fk2SADidYLZcH6/1rcga0nuh4rM3ydeT13S22qARUSWNdeMwFFisqQE71o
zpvZGMl08IlUCKQ5j4i0gGoHunSkovIl8E1lC8ABeUS/CC1cveC1y2Aae/bfYtLvtFfBtvMi4b5s
fT65Jp+TzX9LHAfGPRdnIRfRwax1wm4YvzyDQLMQ6e0JdQFkackviLr0AX2nuZYWhWmckER2XFLD
JJLeZBslRS+uQ64CJJEZET5FoPVJ+HjoxT+unaNLNBGMeiW/9XwVK1u67OHWcKdLPNQO4IRjk5yw
ICdEckVDVpwMdGRAp2BIUvUS5cgjv1mrVVLJOubX+v9SKVZxpngk6SKsFcdHM8sAhT9wvxJ5ni59
F9fcxjArLviG54K2QvC/pjctOyS8UNxLbXBLvY9bIRmC2LXBb/pm5aDVSnORK1NRmNtGwgjxjpji
Xf8vKilUybPOTlONfMeNGSNCTCSA5VIafngUzESKNzlX6jXs4o/EQodnMD+dPfMhs54rNChBIL2r
MSxz9c521Il81s/DxLQKZAVXEpQb/AYBS1P6gjGlzwlFsvfqfUPiA5V/KZp4TFRb1q4Vzc3mbvY6
6ZHAup2CRpRxLjOq7Ix3yggUn+bo47yoqYImLVKesqIUFhgNhygbs1l+y8aYkFHwSAYr/40pYoJ/
kMT0cFbeK4mmpoFlwFw3rYYkgC4oQMqtVyjZZTRzcllkhCK+yDjmISOBNb+DkEgtgEj4lDKyo/io
T9XRkPVe6fb1MMxV6atJXnTgilV6zl17BqGi+urPsivXxSh2QcnjgGdIVTS7p8z32nw6KmyI5Tp5
AFj35nDXsseVI6oa5VYNE/ZaJEf776/wO6xPrODadJrlkHuYKcEnTf3WSVfyEMxt2QKc7XOpJWiG
jFhP7cbRsE38SsOO9HZ/B4HFZMduZS3fukBPubiYfJplNdsSzzTX7YsWBEPdg3gALXVM+eKz4NrY
uKZgrbqAdqpSkm7o2eCQeV80WR/gFttBEjx6LpZ9/Tm1FOmrf5WThasZbLrqC6ATeHGik6KnChql
U9OGEzDIrhEaFNSJyc9VNUEBfjm+e78iCScpZU95zBFi7nUJdfNZitOvfDSyEmBPiLw0QSQkMC3L
lZhl1CdFm3VgUYhaN60WRKpErRJDFZxAGbni9uXTqJgdaqVKb0vqqqtXRnxvJJOgoADYEiChYlbx
jxMhQ1xDbO72TP+Qt2PRxvL98IxbHzdQxYc8A30o77jolisK0Zj9K7BmOCFrwJg9op8fg/KatgOV
jxm5SxGJbEGp2u6pyIm80A3CYA+5M12XcSstlqpHYKgzwV+EY310vRS+RAWnlnHRUcSGDBBDmC5j
0ZbibcDOWU1AtAWZ80obu9aMtLhWtwX2HzCN8p8lhB0SxRabo/x+B/mysWoon9ymJyBb8pKYreIR
459asSVGQo9UMaJaDegiez8sO72drUDu+PaSlDzvS6iWOT8RZ7+vF1RPM1L+xQfefu3oxdKo+jiD
8t2CxQUlffYJJZrcd+B7IlG34TiYfxja4ATag9Q+nPpdkWQBSkVkc5UqTLhhlBMgsK3JU+rvYjCJ
6QaiuAggJB0eStBIPPXza0tN9xzN8YVfI0LlQSBeKq1B4Z76h6G55jsLPC9YqghEWAtMM/Y4K2PQ
K5coFqfN9ExQ/YLNzM/ZijjIaWfjaOFXvTn+LqYZ/XcZWsq49ytVSK7aA7DzLAYxXoclKd6H9eU7
Fh1RaqutKx3zC+y2PHqdUJHm1KuWsc6qBL0J85WwWUFKVie9V+X2yE8nEG8ovHD0GcwoLQDAG0rz
CHnPztaqTiu2cWCcUbClHGfXRL0M4W4G/EQHn5CqREbMPhJbsKYVt+1vyO8EDNqEv62DB5r8D14z
wB8awA8WLvX7ieimaaGAejrarHHpbtNCxn26tuotsbIUeu9oN6L5psQu21kdxG46HdbQW7Phd5r+
tuoHJ/Gx+7o5KB0jfTR11hJMOILwjI3uf0I8h0oqgGVhsK2o4id8ryUohrK89RXpd1yU5kgA9Xg4
wpyGlPTP0P7SEBzZkiQ1U2DHQPVU01ST3mRKEzQiTwJ8NyNCmxwFXhztYE7ydNGn7XRlkL9Zb7rL
26uQ//oei5sMv0dXMRKCHy3l0AM+nCayagna9nrwwbaEU6XAsB05boYRlaxTzLyAA9VYyNzKAm4e
jjxgDwBp5db2rUMRZobGMLqkb1JjZR6CBbWGavRYBcBbBeBc+5phqLr8ZsVH/MUYxDrJd7r0GHN+
DOxvG0eehjyXYEvgEf1K9IK5lYY5JSxyw8IYUtLc17Urn481V9d57NnmXgPk4k3eLkG2cdonDVxu
bMkz7PPWY7cqwqUR/dnvPkLy47onGqO77VOjFMfzuu/XrHSdxnH+emaPmGKhWvIHoSv0QlBqsjvr
NUquFVgS/g6SISqhWkWvI8tE4kcWfj1/3LpaWEjMyO6LLPEA5FpsLhg+BNUEw4krjZ9EDG3parX9
GrwVFDMhoWQm7+0/160e6mtXCTWo15B4wPfNgFrkSjjc5qVkQxEomk/aavEZ6lm7V+fusTqrewQy
kqUSsgixtTTJ4JHScCnGNBXC9UH9oV7WfRyEYOM/P0Z6dpvNZs4TBKjf88kI7OgpP7NuELTN1l9+
x8BXJqNRdRdC/OSz3PwVE+6UqUl0dRnLk45QfEj9A7js1CcuA6VIin9GlJ+JpaCd16aT4aM99e3G
rGuMbXcxMQ5Zi3nj+Jfra2SlpuX8vQp+NS631DyR7yAvXWHMWReblNZd7NnVNbFVfDlaVLL6nfaY
ZW97A/e/aDTRH59rFCopf3uI90R4DCnfdXn9vbT0dNyS7PGeiZ4HnVbrmje7x2sa9wiWREPyOuRY
OEJrMWmmsnQODwSx6sdC9i0LDsvG8CNcVsV18Uo0/q9k86wv/TakApIN1tvjayOxAScad/Em2M95
mu7F+P5SLUpCoqhXgUDbpHbnrIawE1kIa1GkkrrMPSIEzbr2mkHpAsrJEgketsXCD0Sq01RbGM/6
W/3JMn83RSyTJjEdTWCHBe1h2FRkJdlAVVNxvwVzBQQsnfg0t7CSLmLbSg1GmX7V3h7yD1hME6Qn
VrHHKFkncWlUMEJTs7iYk38DD7J5jUoWiQ8m32YN2hs5/XdzxWl7Ps42zHy91rStdXIXaiYJN+PF
rZpjZEoVNKxCa5GUyJMO7+aNntxHz6+uglDkDJY1TSTKONpIjWzzDrueMYlUmPr+LAPImkg4w5O8
r1YNG7xEIuKdSPXBIa3emwmUHM4C0ulHSq4QiYY3kf/UFLWLZ9UR6PtLTVehbz2XPo81xd40/NYr
J1kx03yHmKaLI9tyAKS/A9M7vZXMMqD0QulDucvQPmH8bTe5BEF/R5HPcC9Qmi1ZL7aSllc4v3Np
OMDFZaWUgzwBZnYXoT39XBPGW65yueZ8kWNRUGXDVzGCsoYeUu7F9B5aShqiXxIxikPITfnogsi2
8bxbC0pBJ8PMuf0q8r4c1sDcVM1/SLBCxb9T58q7khlRNgbRJP/2WQ0o10PgzScmEuVzxnjazRoL
VnrWnasZuVRMMCWfDliCQKWBy7Ep13f4I5YeylxVxwEEon1EuQ7VZl0pucThxmH3eRbPzZBgpJ7d
NOxeIDfQzNJxo1Vppzh2T6YrBFyVcSsKkAh9hgvG5xHM6yD56xevfrDx2xtPeEYRJ2ChoHjm5kJP
ol8kUwzxaybM+7g2EcnQP1pG5kTJX2yoK9yMhGYXc/CfGTJlcJwHCTnz0X1v7K2LGhNMiyso5De4
LUEnNJuzV4pOOikwP8XZNLNF3I4zov7HSqL3e0sJ8xsg9fdT0HH2x0sYIBFQIAuH1eOPmAkj6FhH
l4wMtvnQycK06PQZgBEFmFJlx+k7OgaYwG27DHrkZsN86/fTqTBUe1OoNXoWcnbbQaaat3O+RX5k
VMfLpE3DtJctmQFJqBUpWKRc42Srs7j8Tr/dBPMN9PumJCSZh8NxnqFmqxLkUUuLQhu+gcR5Kxm8
tCup18qExjzXQ30J/UQStti9dl1ZywE6QAqFxpXyWguv2SfhxIQBu63Z9YXtoM5/+XVMsWSHOmB9
Cx9yW1Q/JjAx/5akVzQsbyqkzHh0h/PvOVTACd+zL1D6V5ydEaboXdOugmP23QLS0BRdDmwgfXRy
HL6K6rZfunPeBp+1ran1SFLTgA/ICTztR6bOX0eviWmfFyA5nh5vZ9swlQVq+dwAMXJ8yAK+GX4m
EP78j4CpD9GhV9D/Tbhy9GidATHFzVcpb5KBL5mrtV0Gpa+GzOK6VXr/bNMycdbwmEcSC4I2x1RT
qvHwpRQSYroVxW+bT/2WTHSH84S4haRv1iwop/Q56mUFvoQmEWM5wJtX3g1D0ojPOmNuMjU9qTAq
V4FZl3XJ98O7S6TXm27tKj0eymGVwZvLiY6Spa4e66QIP/CbUsH0Jfro77h5Bzm/LfLFlFkNpzFp
CE3iEs4JlObaf0X8zZzThRPZ9SilEhqViFssQWF7qVM17PqtnF7yHueNu5bi2bx0L/6eu6yKjcNl
7DXyhP3wAfIwZbLOGy3BdM4Q0pp1+hOd+n4t8vE3zBUgc7PfMVqAS8KI2JdldK0NtkREAiotGL8p
nvTmeI32LQDFYVkeo1NMqqsBrolz5/KtpHISQwneyFw/4THzInu6b5DdBpF4zYI9QDiLwhkvN7h8
exVb6JpqBUzuizX0kC9kKMgGUWyvXJ44VBo0PenllhNRKqjwKfF5izkYyW/iO/2R/zI+aJCgGiyJ
42L//x8ozHlfTZUAqNHjo7QMtxhUdYKc6zdYXFX9mcP2BMxu7XAXd941Sk4raJKMuwA7OaT6KBP1
iXUJq3nye+Q0qn1icuXMf9jMwLoD0iZllyZsWuemVhta
`protect end_protected
