-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zeN2jLd22XiC7RZfqQjzjj6t8ERQksVi0KGwMTOCDR+hi05cfaWvbQUXSHHFADw5tR1iRrc/uVmD
3AH+f92M3TQtApFdGRnh8wfWbYb+CV8MW7jdGchTW2vMUh9Bu4HB0e44wSTiAguWZ++c2I/hIVfj
4BXp4CFk98Lpam5ivy77BOL706wtNGUYKzRWmXqydgsJdCQ5TmpyZK8Q5/BRyN1AjBISb6+vnde4
hszP4+nc2QEKVx/50s1UJqw2km+Q/U/MpWinPGHIUntZXQZbNDQGWqn74AleUX/FjogPi7r4E+uf
DmqIfydUezFZ359lsAkW07E3e9GXoDlQgZU/kQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14672)
`protect data_block
Yc9azbU/+JL/lykcpJ1hrWQjyjXgveovtQsdR4zW2GHOjvaGpOriuv0L6bBU0lkrpMeYYrKpgd1p
3+KulJM0PaRGTxGNT6AUd0QWr85D2FY5yci+pyUlZo/yR1ikw3MMpCAsWFApbfyNvc84l2KJ9V1f
5XLys2Y5KhN+DXEpplJwu6vELcwksS1XNcFDRK4Ak7FmC/g6VLgw9yv8aDzfJdwlURUhntLfKd9O
8ZyqnNK3Nw8rJG8pM+y/ewp5Mw0gnkixZVidKh9dOTWqSZOv6SjPSrVNKwQIi5eP9VllMctonQPW
o20k0jQUukucK3B7rYzqyKfRQqcu7iJ+hsfFyHUo9G3BwROKuc8pSrkixWm4OZ4kPf9O0RPLo7g0
swufrVM7QPdmsiD6T26aw2GgGOqQQ+LglPfN1TAxmg5wNsuEAbNCYvqGWaNEyckrz2XKxWi85rLG
MIV0IFxsM7dRLgvs4ihsKvxSPwJ44ZV8V34TWXzBUAF09W1Xk4J82caIOHIqw+n/FRSeda5aBhAI
zw2nBUqisHRAj4r8AeGYJHo+i3AiYY7/Jfss+47sYI/XPjPSj6OrHbHZtWvqzlmFZlI99dfXHzXz
0WAeKH7TYgNGiuB0xfIR3Yn/KhZZeLVuajDJAgkDoSpdIEiALNOCI8EduWefGmh7rabpTh+CcYC9
MQCs0eo2m0Z7abJWQlpPD82HvNECRpQniJ2HQJexaM1OyQhWnS6gZsrgfe1zB5amR8FE/2ylozNX
WtgDxs4Zh7Fv9BsyxC/u/9P9lDrsQ0A3hg3RkvdtIv3uz2piyM22iN9T7Lx6JmP5pSfdCmfO7pPx
pIHZtbW22vd9S14ahKyZ/ZKt1/UMls5aK0K6XyNLhxVXOQXkuDxTgr0RMHEV110LH8QYMJ+NoUmZ
1JKd8SiDfcdJ8th9VJ9c511bPX/o06R9KBbD0uBYaLBcIcFS7LWVlVFQlqYpGATjVtguL70QGLLu
zhYFdIhl2c0hBCMIxFSaF/iSReX6xbk4Ms0by06UvDAiN6aJvosE2UnOLN1uFOJJJRQqYb9mFB2e
q2Ajti88rP9Hec9NMaEYZPRJyQ7TcFiF2IzyNgvdTVd9PzEY4jqki1y+Hbuerqzk+hS74+iVzoZu
L2XY3/HpdKqjTxUoyEeXB2DULzyOiozKhvlYDMSRyHpgcKI0adkPrdSx4xwBKjZjG11NUPDMosc+
XzDGzvsjIhOPCxp3BdFUCW9kbVeiDAfg1ZCLjigTU5cUOOUthqPAtA8XARZLDqKlHElgpb6QrOyJ
ofFypwQ+/z4T/JPmR8qrJXoKq/v1KNWWeR4VZ0W0v7frsrbKRMgFFzm+v6vVhlbYKEgkW1zsCRT4
YJcCyd0wVT3FhM1jDo/7pjK6SSZbcuaSOFpqv+qbAl7YvrgXTTjbJLM1+i2TMHBoQU5FUySnymi6
/Ic8qFOr9prjC/TNMBmeOLpgsxfTWnHof/S2OezlEgW6yex0fiV0ch07fsbWljRHjTJwlwatgbUP
U1NNGKtio+0RtResM+szYV9FAICpAz6jV8/jZYOyXDj37AUJFBdVrWVsheNMHwmSX+qAJG9/sWfQ
QW5+/AGKw4Ug3jWQUkQEpl5BNL/eU6LtfXpwZuUlYi5SZwCK/RhRLSdXKlWhF58GXjm6TW/bQ0rk
MQorCIZQH5Dbaf1zUhQFt528ghuwbti3YCJLbyx2rqGevpJaWI7uXgjIKMWRleNsxyd3e6x2pyDm
hhvkc6pC7fc5Ex5UaRbLT+4TEu16LiWJLAIR4VHavbFOKrAueeLD2ec1BZLby9mzT6arXzjggN2h
5tVxTWcvWDT8HKFgUGqvfevXKTN/0xgJaNfTY86yD29jrIuNNqsCAg6gT8o4mnDBzB5txHZAY7Cd
s1NuXeXDzALd5g1MtLrbzSBLz3Pg0NmmCzDQRV1M1uzAcM2aVy1FEde/MKI9NZfhl65PjwqqrHpi
Ef2SuxiIBzorPOm7ISCtNZB2uWmdchJW8NWDoLb650YyaoDbkedpq5rfUumHfmFb8eObWYObjMqK
wIwN2ovYijq+z8Vm2JXAkSzsefmf6uZEiTS/9AsvHm/ebL/nFeYMqub2/9gqOBBL9HL4pNX1ibFp
TaM6SyqF3S1lFF2U9HGmQs6+hg8Z8+GBAGEaenE3ZArgqJZoyqy1hh6FCx+r6QgsexIESGowS3AA
q6BfrjAfJnITvlqRqvspbTy7zfKyhwdsFIrTN63aWa04aYwPoYGkP6vmp6UYpSPhqNEPbZE/6PoW
VfGc9hxf/Qk0qQt4tCLSw9IY5ceJQGqyQTKKrIilEx/lN8oPWsIDWCztu97rH6tBXhOydtg3uLvX
5Dagoniw80rhRfvKgHJ1XMQIFuCXp5LgWCG1yEPkEBsugTLjkWekiYddhxxORSvTkWryAp6TfNCV
RfckXF/W/0ovsjONiqaxH3eCStFQtis7zjnzu3EzxGB3OsWRbuxYBlHgybcaxAt/oqUJcAIQdRtc
vmkkVkxLf5+AdnB8FLP6PGASn3I3HfoCfbHQTUXYG7lJaievlQEulZnNWZnrQO2LrqhIANAUD+NU
ksRtDULgZ2u6DG5tQW4GdJ2YsNHnNy9FYxdwYZ/rs1Aed65Q61ytPxTwGXFRlfdkEJyTMP+yNy74
P/Av3PCELD67zz5XWCsMgijLO0hS3oa9QQFFDu5Uxg13iM/Q9ue+ZPHywQWH3zv7xZiBGgZfyasz
YRlE+mIcGNVKnoJ32EKepVoRC90V3doh/YD6DNJqf+z8xFH56vn8ccGChCIVGeJY2Ps+MtJjPqIA
YtNWlNY7vcLrq9II+PnUuhmD8KfwW4ZXG7QBk2mf6Ga2vPdThUISe6d9vJ4eKhiFwsMqDniuLhWp
7ReJn9hckkQxrKXF3TA7u6G/epegfVivx9n/Wx2qgjLsa+Hf4rYC41fKEIZT9VRSyo9RVMVIhVgY
jaZOmro2ANPgHTSCLnuCIbZC7Mug7NkBFR1yCe4zNGJXCXTyRVCpLAFIpr12VLZy72b5aMsxqtA7
G6viWHWwJyq2sc/paFOz5SAwHc9FiAA9NlGIlY3dRckaNjQYj55DiatnSzWI3DH4NyGRqXGXUEwP
AeEyNYHY0x7a1G2CFkpFiFbq6YIHMT6hdyRTLUcvJn0x6T8jnV7V+2gP1m0+EEzOBtIygUClghcK
p/S9dONBFPKP3LHtYPtW+3qpSW6vkdYdegc8w4GpH0z2eAsWwCJoux9ypCFRv5b2C3vhLJOBbOzP
O8lDDFAgt+uf4GvTAQGrJ0orlALK7x51vJcve+2C/cawRnIQuIuLIm1lymPpmFDhyJl7xp7bl3ix
0gVyTNcrsldiVMk1DqRgmcsA9gRTmZYR+NbWt9Z4Jge0zpHdggIpvJumb+lttd3087tqhZYAWxbM
neMZ50vsT4dDqV2dhdDB54awq4uh82+ct+GlsHF496s/EkwNtg2x44TvrMx3+PLJerlSSE9Z6ACL
hkH57btY+5nc9lwDNfp+biB0SIUZvFHz9x+d6SQ34ToDQM9pMvt+qINTEzymzKIq2XxY4Ry0cn8h
35+tO2OjzRRaLOktE97PmRbHTgA1h1vYF46ZJ5oTcDvSI+OkxSCRDOsqLMfrBThYXtMkusOQ9uW0
xSYjMUhCsfU2jrkBWT7LsGuq4xhRWUCxYvgC/QdI5GP804tK6IlPAaSxAmfPTjz/IKsbl5E/h9wE
zrVv40ovxG9SZcuGIAux6SYzK/IZ/8OvrDKYVoX4sbGbRT1IASn8fQKUzIqTIq1VBTi9wViRrAR2
wThEh3lp3frFm1QckeevppQio0p3TzRzqyg03shm9SzkthaYXv812fdhz0nTwlK8dZr8A1kdq7cp
/Aljz445vRf1RVTJje4+e5UBUzYBPCbDIkYvo+ItzJM/nrYa3G34uVAVG8/dMRabEdBA29jcxO4K
tNBOfiPpczd3bXVvI/TOlAVoFv3J46tzS7WhKEovcWeeNuSHaDb86t7Iu9+Zg+jyRPK1hSUjkvPY
YrJ7oP6fo721ZTk6IVjxbK8kqnZjvjRS3aFvqCJYGAJsUNgBL9cvcwFPFlO4WIhH+exgL2q7+/tv
sy185Y3K9wYqffpyX2px60PMG7xfOtZPynuFGl5O0JX6o/S5gEGHCCwBeGeVn/O9ce5cvGa4NQol
2SNvAEOaaWACD8VvzYHmxgKvcsP41/zmXMqM8O597wrA6Hz4zNOcN+OnptuehsMTpld2VJVtloq+
I6D5s9tMT9uYKjnriGXUTgygW1NUT0xOnr8KXX7DK1zxItsWMmSBTipeepV56M3rL4WxYTeztxBV
y16MpPeKGRmgbkJSAzbLMpip2dtYy45MKlmFhzEaKv53ICu8bMZj5K2bfaIHO7PL/B9w09gx6xRc
e912cB/Zcwb3+M2oFA7ANvdhbjRJYn/FdYkC9+vy2U7OJ9Eneg9t5faT6+90andRWvQM0Dk0NZuW
uOu/sXpV0dw7xQGtYoKT0yKb6Aewhpx6rG6NsR3HgqwVloAU67OvAld9yopl/2oZUUqSfvr2I9v5
mGbXukk3lntG/Wbgy26JbGrYXHUBF0FaDtKqMtozVg4uni3kQO2NAyefpgXQEesYWdOT7WCxhNzf
CAqa3V8ad4g4cFA//qOP4Q6OzOQfqZweT3Ex3ps0ia/Fa6qo61EV+CMcNU49+jqS/aZjuq12hrUh
htlBO08i7XDO4n4eIuGf0X2rJFPmWyMc5Wl3tOY+8P7hcD4fWDvq3DilNNuUgtk4LKixDeaRL81Q
S23FV3LTSPswOMOIGr4wjv2HfQfcgeA4gzVMM/PQdBQlEqlluVwgn2z0dQYkdiGxHEpcH1YesaeE
6xEYqnBNhHxooelvze8avaA3xaxyghpG2Vp2uPvhVAfmH3WpPCVpgV/8QNY9mN3jRIPzI2dkHzYK
EyMgdt5hYSlNornO6IIizxZrQ3H/3To5QRq00MD23JoTUYNnQBxLa5GO/ivNH5Lu9oThs8K/705p
rAKVRjWq2WLq5eX0FXVXrJ1PayPMmPIgoy3p94ktT8vuDnhDDl/eNazYqdQveySuJgLAa3RCA4o3
CMeUNWm/haumCQoSyqzE7mdNrN1dgTnkgdqpC+S6PNU8NnQkhVU0h1xwUCO2+l8ia6w2nfFi3QaA
fOHi7StXpY/Nh2JplFef06onnTSX3V+iaSExOz77LRsgnvKUDhcJyzwgw9uSJhfr6g/DQYuNcTX/
VxO2Zh4rkLy4lS5btmUPuX5S335jT4e1FBIEjaEeNshSsR+ngC6frmlnK131zx6twe5kpCyQxtyB
OVmLI1Yolmj1mQ+9yxMOs3Q9y8Nvd4uB1rkK5KSG8wZuqfVdUdl0cFr+IIPlgA2pRvf61l/8hS0m
lv7YgGlTSlSrGY9HVNCu+Mt16tNTjrI8qH8TOvZUdYAheWSUIHABnCpSpE713wBn7DzUZWWbI618
QWiuZBG+yB+iLey+OVjzwl908oWBeRJ+Zy1mYFSffppYIDCM6LRmr3c3SBUYU/vyWjYwSE8j/+Xp
cGDdOtRc3/D48I/8H+CCxMfMCcHDdYxdUN90v2aJFI+N81hbbtt0N7UxI3KwZTnBy0QOx4eKaGg6
ROzUPPPSjhD82RFL5Epi55rJa8rjsDorsZOBh4v5D3pEi31BbS3a/iD+yqNJfVRwhw3eQUSHEcEz
P8pMHQzJxfetLwZ9ECUn9if407bixz9Img6UCFlVX9vPAPGlPTUoFuMQiMYGrhy5J9obQTFl9Y8K
31znlolLWnisc4e+z5/0AmsMTSRN1GwviDFlGW8e+GVgDrNYmwvdrvEOOoHEupgb9B4SEJhyIPdN
02+UmQmSEchjbdlQEezxAH7SoxJ0QxHvXK8Z4W5BKE4p/Pfjt4nwzqyQ2NThqtMRUVnHCS3FEgbW
2yqIjn5WqFvt2PqVC9O6zXaBPt1vmoIN3hNrtQWNSqgVEgR/gbqRYoJbu0rNOaKCr11fy9uJCn5i
f+o15Ufso2zd9nEPJFjna8E7wPFw7ey/0JUdYgzIDsGMDQTkfryfujqSDNP6lbXeKWoPJMLFMGhl
1YrQsdcbOllbdbT3SmRsTDjl/f8yorbhVFwbSeXIT3hqkAqsnhCzc6co+jz3Y5nyeVAybR8+/uxx
yo6mBscMVexKeE0bwPw6zMX+qy6Em6eyuJ+iJoB6+fTwY/46mi1pZl9JGKU3A1JAPUvEbcifOXed
kMu55o8iV+AISzcq5EWQeENsvDj4fS83S3hTbYSJy1iiDvVhAS2Hox+X2aQme7J+p5y1Z0MQTNQp
UsHkSLqhz7aBsG/LuOMaERymeiSUl5EtXfSSGda1Q12AwusWL3R3686h/xX7U994SNc0vffeqbJs
uSfIabeD8APDfLpIJbg80lr7V2C31hbw9bAZ2LG8j+6ZjNRiA/137/9mLsDMFOEAVFEW4seankcy
SqAauMnmoIX2f7KfWKgYjjbXOzAuhQp6RQBMs2uPrZtv3bi2+cvf8WYV1TcqmZgs6o++cRjqNpMz
ry6BqcgShGAoH+gnpgGjm5wZzOS/cuGjHbVwko5FNhFcXgryUi34G3xEHsAJ2GAuA6n3cu9GANGJ
GSGmzC5VOnXCxbWeibm+SRcMl/DeSPfd/lD9TaS+AeQDbuET5kRqxjhAhEFOIV4hET6RVutRGjaL
KNy4yNgeDp0wMahX/SatJTrA3YDDWB2AVEDdowu45CM3cgN/gHhyE//aaqhksDxpKR4cxFdbcCmr
ffpL6E/Lqf/mheV3szGqV8HeGIeRlSKn0mtRUuEeHdG6aAAAxqO5MdnNhhgYURnk2X8WVdP2TJDn
uai+E67Ols0UT24vIiaJ2VnAEsoarGqagbpbTv8BiUW/1ZHA+ug+fJ5bangWfuZv2pCTL6NMdk9q
ekCebOCbQE8DYyAHyiXgY6eK7/H+dk1WuSL4bVxmWW/zSeNYNDS01mrXmukLVzGHmXZjdezjVV2v
ZxLjk7XcdboK3xW+3YHfftYHFToMkqgeRxU0K8Lu09tSXJqa3LZzn45U7k4GeDuoVDUY8ij2xkRV
oLvtTWTgKAFUx/ESxIf2hHZlE5fEdLLrYuFUiDzse/URLtxppvkU7htkP1afR/MQcJdvCd98Ii9J
4ZTYBTRdPNTdPCjab31F5Ielzfo1dOVUMGRGik3K3JExHxQ/j0TG0rYniWvcN5Acv1BlIvlH9K9L
MrqOpn9wbc73pHJeYJHIPo3Ra2RlygVevELQpoD/F34WxJdobRqKLR0mRhbZ4VBmBsVX6hhpklEt
d5e9FnuCe4uGFwIDJwKfhRFjSnUsSOBmWEoj0E4/gPEmDqAXgKbQNlClg6wpuu8f9k0Ze56jBAeO
l1Qp57oxu0PW4xM6OJ1P/kv+C2v/8nLbi25wdJ6Yxn1O6MuFFA/FlSDn4VuI8x/rjUs4Cyj3PEx0
gdnooYcE2AhyWuyETEijVQPb+5sBOSRJpKT5ZxOR4yq5fWpThBdT2M6T8oKzDhMSy8GRVV0HGL2v
yjHV2zvvQVdZszPghcrOCzRF1Fp2CgUhh4oaRC/lJFyXGisSPIb2QZCg7bY8xqke5fJuv3OeCO7K
OkWJk5kfjMZrlt0GO9naigxoQRt3u7TJZrVnFiw305tWh2KkLYT61fh4qpbcA4BNyLRvBuwbGIGe
YQBDe8fugIz6UP308P1V0QVrCRI5mnHijDQ53u5Vo8VkJ+vcZBuTL/w2CSHRIiGfC/Dyu2ms9nFt
NCND5iZgn5Pp1ZI8hlk4tu6kyyBQFlePzwFOjdAJeW0FhPyJCqZcPOIh5EVoRZ3eIyuuIUC9fvmw
r4MTc+b+rWVump5aVa/Nmwu+ZOjHYJDUSWWARkcKdIGUPZYt1b3iBxLnTJQ3j82WwMSyJh2plUHl
u24n6S/zLdnxIuHoQIEpu4N5Z/9qNhqzv3TOSfC1IAdsIDrZMsPc5/w0FZUCIanbi5estdb1e6u3
EL8fx1jsM8AbsdFwI8L81eF2PveMsCbmarYuRtqQAgG7whvkXxsFmgmQRfPwlWoEGS8IiFtzQaEE
2wWnKoeh4CRx+WqLPbs5i9eU3xVEll/vUAVUVjrE3AX2VOcV88ULR+3Kp7XYJRy+b7BKtrykIXu1
Rulvm5MIpSxvYoRdlxIS2mUCiCfJl7C+aQRm+zn40OQvGpVdfpq3GzJ4DCUi53OX0EmMd5bTSbjw
7XeIjHbpvRXAy3eEIDcAyxlMSRj6uFrQZXQaUMRJb74k/pY593ghHf+8pIIZy5JXl6vCyOCwqEiX
6ADxB61OvK0aZqMBz7yxlWJhPp3p75NEdUAH9lv2+NaNEsJ+4lMeA0t5azm0/xb0e6XEPH238H5c
KeW0uuiOs1FmIo4OkeHPl8IrZk5ug+YF0tSB27gKInHUxDW20F+qUbTg04xj2g9r/IL0ajBvoBI8
15vPQG12ckfktjMrG5MYnQXe+TuX/byUBF804hsGRxWqJQsLgReZojrr8EhIgds2Zjk5brpsUDLi
doWJo/uPbUeJWxMq4v3WMMjXcimQG7rLjRaUZFxwoYj+icZ2Vio7Xi7zUWuuVyP010uJrBZ37pND
3CuEVJYlGN7t+m56mdLku0IohL/ZRpxifZmtgrw1pLg0ku0DYKHy43Xg4+k58+yx41qMD2C9L6Y9
5hqkatZXnY9KqPWI1id7NxPc4pbr3d2m4Ko5cTm7ow5CF9YwC0PObULiIC7Ed0n4a1XxUhd3qBHS
TFprSV5rt5ZQXXcOl27E3UdMTJsH4hmyeLb7XYY16Y0XTPnLxBsRjtB4VIMAJqIGDNVYZ4xUZRn4
YxYw+EDD5uzMiJ21Wb4GKbYd5uIsP4O2GPdry9wTcGR6FagPv6vXC97Jq8tfb/M/fbNLPuX0lkwz
VKg10WqlsggB3KV8m1/yrL+t69uc7QnG/inQyeRb8D5cQ9x5bpBgQrUxdnEyNo/7MDszmtPwa37X
QClC+UO4ymzYsmvDSMxHgWGQzxBUWhFLOYN3Pea3TfERfjFmr3GLs+5lFRH7yBfh3lNOKR/BCOQp
fsieVEcVIswjbZnipjUNgHYLNub1XJ74jJtPGNsLQHmPNdaITGlKj+23EJ4dLpLRSPlQclK8NzP0
1rtgg9wiHK3teY8u0+h9huRzXQZ7KcBTRhr2Q0n1Lt5wECH18/Cju0H2yM8dCqituuN1hTPh3c42
SFk2AhcpIvaUKQKkufVieFswQ8v5AVbsYnZ4sznFbN0d9S6tob3C1eL+L2tsll7z+N6tGP8ye+Nr
h4qLMhuNy6PV+7MHSLZ3Iqs2xeA2fhqHCU7FC0X2xLib5+friN9jqraelf8OSyeBIgkDP2V2ZONz
GAnG27nKMgZertyQJ8QojG42XJ6oUj+RvoBJmvfPzct1Gx9p6elHPPAGieZw9NFZLLDRbNaKZYwo
HzI/q/DHfvaI0qUbIo3tFjZ4MF4PI2Tt7B9u7dIrq0YY6hItg/D2G8dA2t+54yu+ciVPjF3zr2WQ
1S3ZfL/LNdzFI3YCP571xYpDnhcZU3/GRg/x94Lm/ZK/DvCTn3FDmcZu4imnp2vGzt53CtpyxZx9
PiidYLJgZFfRV5xcpjXhKe9AsB9TE9Lf2jgY28OZe7M0R9x4WANcDybKmQVpsAqCOPRKlxcEpo1b
aUjlZax9/rsGCh4mtgab56z564EknpWKsV9EyvHSlwEgnXyDdWvBC/qVDGj8lmcnoLprcZjDqpvK
8ljlwoZ68JXYyhwWx8W0ZvEf73iI2qlkJztWwaeu7dn78118ai1eXKszr7EDBnoNP+CGiv5gcO18
wXF3GY8EBodbBFrqBINyRB90lPB+HxRgNNBxwhRpYe+iDDWZuDdJlUSc8YD/O0tTOUwXX+q6oI1R
RStdUFWnMmgHxB5BDqg+SfUkkrC/OJgyAvTyWA+OwK4Op9FlXDuKcWv/KE/Veyoj30uFD16Ea+HZ
2vqAM6DWjVaXsKGqFBRN/P3OF7uYtU4o8+yPKbArzCo5rz0jV82zp6OHodblZUZrzpdrgQ0uaMmL
/vbvQOvpFU/7V8FdwT20Q8CtbL6z3WqWSgz11CaFU2f3PugdpgK+hhV5ugGpn8GKTiDqXmCsgAdT
cuDmHT1OD4Myy3qU7md7iN8rfo3AMEfY5CqsExPbMNa5kvpkk6+OUcqMKunJbymz0x4wZWp24z09
2fiEczo5zRWNMcwIYeRf427hU2vgtuQS8Xpf+OjgReBF5wbwgoYaxX4tgX3938L7/+1J8id4aW0H
v2hNQYN2oxJzzXfCyU9fNNQUuI5KMwIUc4HimcLWJ2uugQXPsJ0qILqwiPFs7Z4ZdV5cAW8QOwlv
X1O9y/jtY/sy6wLtOUVTszhtJ+LHcMfAx2ykbrVkTFPrCa0j8gsJF5MzT4xAnx2FWZUDZDMIjBR4
sFOgUx9YMsdSm/1HMTVqwm/sqxRrLg48S1Rck8krLHFtsnHnhjaJbB6etLKXtA1Txk8VA1yLF4b4
k6pQ0WLrrNipIyssnqHBloXgU+GHi2yCrVcbKKr5c2TG4jYdB+z2b24SHHA4y5CXRPl/dZH3iJol
kgqz8ZXKxmE4jTEPIIj9Tay0dL4+l+RDuFTqQvHLigdColuhUlkwZdRlb/17yhmPk6Vr3jgkP3AJ
1JCdwkJTP5X8GxdFHvwAednwJPcwN3OYcWzpjpDq44z1iSeYQvCppcYBFtXp1zscDhGpi7uddSN0
VWh2ORkpe9X1DxliprHzSNrz16OK5mLYd0aaH+boST5Z+3siwexwCfARLpQFEXr370+WNC+1YTow
I1Vr7KtSvbxmtl6Au1y0OkKUXjEpCKd8XKvE66ynovb1lR7SUMAVfIQ8arK1B6oMtPUQCHmIgC3B
K9RrKn7VYci/EYbahsS29RlnOOZhEszEgl/qTQu30+m3VJL5ph9jNDRg9LTGz4XZcZoFqflh4Es6
WgTgGkn1GKkjxn375POPdf367IDK3jurxjedpfxwSkKJD+uaPu54oQC770g0FeQiJC1B7AEqf5V5
dVcgnkIPKYMth62BS9lMgFQu+LxYuOsroYMZniXaJeTa/DpC4rQgPw9opPHYW+gdzYt/n00AZ4Xf
PuXris4J2WSXKUEWsmgjTlx4UX18qJyRGzGX8FRJp6SD+ObI4KtmvFV/OZg0VTaxY0wzON2mg5Me
3FUkf0CamMeBlzoPoCwpDksa6Fqi9kmZaOXzxcFLktLPNtnsyzGLQbvz69CPpekzzDrKrjK5fSN9
e/f6mX5lsPzMxOvm+uBCuKdTCpXtedhT3IpNQXlwqXXByT8iM+0/W+HYwrtvZdx39UQ+97uuyC+L
14XpSPk1uA6ZRgLBAlgLUCq4tXWqE1Mwt76qL1dFvlqRBBHbMR5CCYPZhJSJm7VWR7JlOjAs94rt
Od5QdAJFSK350wBsQu2jsqgi2O5f/nBKI0S9tCf2DTxrdrLfnEiTyTe3/xyhNHdjNVoTAhvHfoSU
/eulkbLi3LkJb6j9IT6UqibZz2xaLNTpCfjSM7bhMOuPaysz17AnYnhKMxGPUKQKdT1/sy3IPFv7
Ri2oO+wIe43bNgYjlHS7mAysbexQuQSHiXbg7b1ILqbalMskbWlcBrIhL7/ofrEXZEcuD2K7C2oG
iaZq3wbu7d97gzI90grWNYNwYN/N6lrzEkdPm4inFpgh6BojmUp+I4kqx5WaSJfdlVB2QIVJeJWi
9NNiEWKdfq68HIN8CkWE7etOW8bBkKzJTDe3DXZSafVy1gv6Q1oeBo+5hnNyoR6YyZaVRBr1nJXd
epZa1WmvcM4AW7YxcU70AaEmQvgVFHjzNL+QpiGWmriR56bcz+Oqs5iS1gZseO4Dwpa2gFEja8oC
g0P7/Lzqoaxv2syQSrs85ehu0UTxUiuihWEUXRhhbuH62Nl8/Cf+2ISg2Hygd8KQUhgLHn1pQ0P5
c2B0LNUr0WfQ5EdEjh6pkz62SWEWX9nuwUpNbzXIRX09/mGJQ7sXtNt4TLQHEi1R8xCaBq5Ha7di
n0tTSryN2C5YUu9XtBj2OLTHroatIqkviG+EczTjLTa458L5+hG0Aui1orCfPJZiotHMX4VcC3X7
PfWiJH8InxePaHlhQ6ZmCoqXmAQlL4a4e1FwGFtLTWCklwHFgRS6N7JO+TQeaIAWmkgAePMp16EY
kdylx2ta2DSCWnk1ANvHqS3JGChHjQigW6mHLgHUQTnPu4NuG/vqFdPB5e8ZwxrWpIXU8wrASxJy
hWxqzXzalClVpHwvl4bkfi345tglxeCZXmMEzatM85spP7n20HhR/Id9FA1X01YZQ+D6RtsU+qIl
8UaH5gp36jHniIB8RGTC63OmAryDLu5yHAQSNhHnMmphF2vH2zdH+V1u1/NhUfZ89ADvw+i/tQ1N
1dyXqebdMTmNhi3+yiMP3rI1cPzZvhuawL6ufbK4Yl2S+h1w1bhnVXXDaAP3DbQdht3CtbxWrgE2
TryubTegRH+GewsE5BUDiMvg6AEpU5m2nk420xUObHcNkDSDgkfWwk0fVEVLD/GkGRK9ihA4Y44N
/0uICannTKjGdM0t97UKEGcwUnvojCz7nuqCN1/sl69rqScjLSIPl0i3dJa+BsWQHfj+lKSzAatr
T5xbzpRL8LXE0QdCYRppoD3WSUdGQ9Xiuys3CNlfH9iw3N3jYGXe0oFZxmBNaZAFha8m0ut4V1z+
bvFUSFH5Xzu10uACuQVj/uv4WTWeOEPLA7cg9Sisizwwzapp0394AGLVOocnvGt+P5rJbbz7CNvf
25d4Uss8AcbF5ZEEBPEiC8+nUdO85tcA6q2VZmzewzE5sIg8YhV+10D+GBwjAYLt21PoNeUOl0Tm
2CVMhn/wyjJmYws+jgHI3AkelSPPNXlXRf7r/WeuvL1buzeTcd71Rmje0OLoIPWkewCWORKUuMAU
djVS/e1JOL68AN62bX8GFoFZjhgwKnzDXCm4wKW2wUuahU+acwW8eQnxt5o26trCNXCSnc4VtN9F
oLBd6YL4If5QoONV5l1R4MO3FCXDn9IXRy9ljN5SbUMjelA0c0X7KkYNuyOgoLZ+Fvv5wl3ui3om
XzhdeDLH8/vNIUWMBPkOufzOM78c2u8k4/rMkWzeM+2UMyfWLcOzklOJuWTzXsqMvy0rHRy2RwJk
G5qw/p2L8Hn/MeBS/Gl8ZJaCqle+rZlMUkJ5ht+XXFMuoq7BhLiOLrwwkYEUJGTj4/Ly9VicWqfX
kGUmQ8HQD2Ze9VF8/dpf3D8ao5ov4ADF75Y+ROFj20Y6/9RbIK1CXrWcJSjLSQ2VtPwWQZy+G9JU
fxZDUfuaL6C7J+acLIJWojtvk7bPVMvABdff2gz+9BN3kh4fsVR4gXBAipzJ+2ik4UGGA48RfEKT
XlnqW/MyO9MrN3mwbO2VdWnLovDNZXJX/yx9heLWMnk1zLgb6KtXF7m4031bEwCzRRvXdMmu+ShA
0x6I+1Bu67KZi2QRpzUajrUJXOI1lTQFpVdgqslkuoyN5LmAfALhLpTBOUf8WPaEpKYJoHSeSJ2y
v82YhvdgAcUtQIh+shkU7n507ytpyCDtHs4ttkSSQdBgx3zro19hLGeEUveDN9VvqQqlTAqXqqZd
BfcyHDIfSsAMD5dYgNU/SSWD1qbKnB0YmBVb6LRVqVpcG8DoDIe5te60IR9jJUQL6Qtj3BHggD9z
Vqe8Vihsv9GoJnKlutzOmVeU2cYyOWqWFzbcvz5McGbncR3VB/OMUz4mCgO3XEDHj++BB0Zts6O5
FpjRqlwnrcIF/yYWr0RgLmOOFxT0IlwnVLdY5wYCU5CPN38EUNEanUbipiwIFcRmOAQYlhFsHrS+
22ZxKk9+04g34F2zglWvB3qnN0Y7D4hQJGsYfqxOXWjN8kvKdk2znax6EJ6zQXcA+yKqT7yiOIhk
GdESOQuqszU/wQpWZ/7wPRgxs6KRph3dTUM5ChCsEoz6IPqYaDGWYh4Kq5LitFhFXKgISn9GzJFM
6N70KmbVtIaVKYvu+8rZPhnZ0n07xMEFimk64Xar1C9zXvPo4344TH9wBVgNLZmvvtt3AeXtr4Bl
uG+WS+18GsbcB+RrWhuZB+yqk5xhW7k2FhZzFolUsd/qJMzxOInrR0dhtrEKpHYPfZizG3F9Q30L
WJy7nzTvIfpB09UrbtpxPPZKo2CSoKCRPGw6OagXP7GHW6U7PVab7eDiNzv68LWiAPioSzfyjD/t
onfoJowSjSNy2HYyTSHrOe6XoV55Y0Exiqcl44cOAj46Fjs4nYtnjNQAyrgjSlp7I0uJO9Xod2fw
Be4Jua+X8mBbeEO3hYDk6+6chKcv+TnuwrPZL9loqLXveN5A4w4fXmnp9CB2PdeI/Cof3Lbmq7i7
HhF0I/89yW18UpQR6Qh5/lrWQ8q72Nix0MQsKD1x5W2pqalKXYcyLML6Jaomob7M4e4bcL65daO7
Otd5Bu7YETwkZtBcdBvtG4kehWE4W+Muid0a7sW+fm9liXMKltfl9N7gg8IVO1LGG/6y0/RiqMaG
aHIlJ6B9gdu/GwK6AXeiOVB5SLtPjJKwbrjjs5ChS94G0qoT1rOUrhs0Esy46gGa62ufAMCh3xpV
WTPI8MNCdU65d9PyAZcR7jDtVHkVWtRpuvgPnzNwLuGKoDPz8VDJOKhojWheJaRW5lptUr4M3R4e
4FunUbmJE+aiRH+eCRBnbKu90103bqPLztf1Vq9oWLGedoyLuob8O7L2Oz1osq8w0xjrsGZ6pOmq
l6RM9bHCqoE0NwCMxEbrkU6eJfem9ktyfUNSvrDY0cmm/bfPTqPmiIjRetHStbR5GXoWQhBbM2wy
X8pf3A587SCsJnP8lD1ooc2+R81mMSTLxlWd81hhQ59dFGDBulJshBBkVOT+StLncG+bnD2bzO4c
xC/lnex6zCE3t5dhWXcIUeS9SgBBh+WgLfAE+JwEN9zfW53om1w/fL8QxREtkx+PS0CXeFa/9Six
WeoJViRIqausgttu3sTLW+qebyjs//ejPuyssU0w8CwwKj+qZcQuTqJ4Ao9xiH6ixqIxZCRjGI+O
Ug7XjfJbYw0n2TUwjSo6E8ceTmMhrUl6WbfkQtaqLJBD2SiSkxBZ9zTnFpCM2ZY2K8LH8RcD7zub
J29QKeotgYQIndsDSF4DDOo1tyRS5YBZFKQP91BETowv5mOhwLcBZEYRFliJhoUhQCpuZiFInY9i
1yWZRcpURpdurUyKGGqSlHABoPXdC0WOxK++3Q8DJw9x3vl/d1ujPNqN4ryfSdFtErSOPXgmReVL
9yDtsp3s/wI8hXiD2uio3HeJVZ1HvYSI0c3y4OVsTZmDc1PphiPaBaPhm0kw9QeG2rmCOsSe6om0
Qg6BMMroHEok/l+ZULqvPV0pqDoAcBm4/nZ1wHlqXXxedm7Tv32d0SQVSbyR94rjqy2/ee9lmZ3w
+9jm48ih4qJrGI85eFWmlB0u0u4zidPPZruJQEyRIQgt0bQ3SS9kpFeoppLTrDfB5APHCsLIsN67
71S2vhjQRxFhmwRyg3tlCaXQxyX6V7RUGMDEZqLWNr10p8yG5HA7TbNcDKMXzL0jKTbNEEtmTMvS
jh+L3e5PCQxhXHQHDzzrESj46AVhXVKY3yd8tbfZDd2pgRXeMWlGO7/uLeliLl8oKSE8NZrM5RN6
s4/Qb1ynxM5yKzgF/zPiJxbyvcvBUTLv3cnlq9uO++WRJ/hjJTnJu8+rIvXXYFWXdky2zqFKUWsp
CyxwEk4tUcRDUNk8CkC+0/mT+3T4O2AhiEA6lgV4FgZ1ZbTA0thMikm32GlfSQOMwX49SvUlfHqL
3U4YXJSym5C8pQb9Y97rDBMGQAN8Qi2q6opYHV1myp47itVMwngHwSEv1c4/iB1H49Q8wjY770VS
IF5IBFZDrzkO40ki90yku7iEbQzISTyjFP0c5A/Fc5VHENK3KBlVmbnHVD7FEffLghlGvEkFEN6F
KlF2hdr2TRvT3qbD6P2MO7kwGs2SXfe+MtTcC/lpv70twqKk6UKfqalis3SPC4aROMB0mRtzuGpV
qDVrdzzJvjLdDG5FBFxJw2UBd18u4eNJfZoSBNxOfVg9yOi0rRHtuutXxHpsA+xWP1iOjkzwnagb
UtvkQtSXUu6NFvae9lwhpH3zx+1n1vLmuPuRKIkaAGbUd6vjIpJsScSt61WOVM/n74ll/out83sH
3ko82U4nZ1hkwa9hnTVZIVAuzVi1TgFLCUS2+1U5Gu9G6tbHo9iRv+NuNGyUiFXdZtWwfU5GY6E5
7ksvPLXuFX3wLQ598izFByjTnkksZqI4JlxJJsTuxmaLWIwk2Gw06/kvk1aV9x7+SaQO83lqfVli
asnFAZkSMSlVZjuTjo1BRR/6SjkPtnzCewlJOev62ha2k+RSEVMyV5WAxPo+v8ttBVNu60BgnMZQ
UDPxSFplgzwqOnwkut7IjmiNCQzw6SxJ/xMR74QM479+Bg2fdM5QUrD+8XJ2HTv2h1OF0iEbiOcG
iljLXEnDA5ph4b4vAC+brC2euWJCWEsp90K1BwNCEsa4uvnWgG4YyMN0Ih+OZBRFjzzkQIsa2Q4g
qMDssiugdBgmFI31LkHhHgqJyLTAFJ0Zqb1mhuHP6Wy+USpgypsdAF4szhsQ1uF1wut85ZiTZsTh
26GlP149wftneM1FTg+HtMkbme7YuNKTzwDueD1efGC8Y0Cyq3t+UT7kVdBVv57n+2Wz4KnwEurQ
L8L8b1l2Wg2n+udKmxf4fE1yidwl8meN+mJkZrhnLuZb4Q4LOZITG+0KREZMFapZ9uAO1ZApxEZt
KBgCBIDRP3GPXAUbbx/iKj4FY3rmhSg8SKBzmPVQSNdhgroxQxhO802S5TY7RbO1y0CQhnobNs5b
/VVQhVWvT7R5NKYiGQkGDwGnv5RWV+vwqC5DH+O4lS09tBdaEBawtGrSEbI11D7uM1VD1B34Ivzk
bsqN9nwkcUXVFPsiz0wbC1CSyyHH8F6/QU8NobxTQT9ARbjPjK8f1GC6B7nJmVPkE7ar4uGqbTAu
poG9kNvJPRg/qdY6JHTSWon0U29tyb+nZ4WDXX+y+mSPc0Piia/8MsruIkE6saCYZa1Ofd3lgDta
rAKLpFgBmi7XRUVNiRPPQC4iVtXntpvQ3ULpcZcfFs2fdI9ryBmJstmwi2gHiiz20XR7VMwCVEtq
0IProbdwDmaCNrAvj73OsszY+c5wc6wx1j8o0YHxGkEw6Wu23+LgJTENp5GruRqFWFJ9Stz6yVVF
oHvnGlBmoDrwlLXCd5dSjB2J7DnpgYMiL0Sp+xgGPraFdJe6axuQKgnTvcVJaYzPONYd1/aO0AvQ
+YLB7PBkKAAGUnPxFbEa3MOkkdoWOfd+ZYmU5QI6nQLZX5r2yaELeXGcGmzv3c4poSAF3sV/LXnx
/mw2q08Octwou1g045Uwfc4xKC40a625GRGk1dWstpsturluuR52vqpOgPH/2J/Yc6tJbvwBmK4u
xMRNsWbfHtKMG4+HdY99DB1JPMiiIrdwTk/5loUW/NUQCuiMrJWCXvQXyJ7c8/QFJ3KH38EdOi5D
LVyxBFmxy8PZGV6PnHvlHYUkG+vmjbLd3bpnFLDnNxxybl/RlQI0svC1RYRhGwilUWrw1tIhqQll
EbP1E9iZnx3etXrLIwEuT295uatPjxItJ8PeH2JJHhbiIMNlWrKv8Fk1bs0Oj57ZnfsHP6EGyjNw
PKFzF88QsU7etf9Gj6FXmumIAmuRpYib7qXDf0WrerMF/ta72bzlyj3d9OWa+noWpwZUtH8FcwlL
qRuvgK3pIwy0mpA9COW6TUiKvvkMEy/KFtBncS8NVJR/7zQFWU8FUUZl44rDLMmJ5WHYY6a9+Eje
lmQPvxebUykbjkpeLjs9q4jmdTSFrySNUqbuN00+nbWUd4mgM+lZeSU7QEzqswdh5GL/IDBtzhmc
+ZjshhK5Ar0aZ3ygCKjLASq+oIITs+tWJq/jve5w7cMZhyQsL5PVezK+/PqsB4S2PDSW8hCCreiB
r3kU90G8x8nKhWksC7znnaEBqLcBNR/zS+e9EDVxoKI720coTc1ZT7oKP6KrR2waZ+mx6l2y64m4
/u81KBh/t5v21AtbVo89I6bcbEPt/xQOSPIbasbUXe7Vn41a+n+Ls9Eusqy38Yy6nUDrCFNy/ueC
GIt0zIxoomhJO6vp/dG6Ch9DXWoM6eA+VqaqKB0ykvMovCyrkSBgfwI7kAjWOra2mG2OIfZYyvz+
YzzOEXvHIRNb7aIwpwOiZr2k96J9mGAZvaI2PeOG6AEwK9XWznU2HXnczGB12lBuLIo9d43dwzUo
S1cKTvFd2o1fYWPoYdFjZcmgXi4Ks/jT2rVrzUrZDbwTAAg2xrC+mBhEVrOsXny3UxtqmGxnw5ON
60Enij2+UYlklCedioQhmrQQIG4h3+IA0xDslw6PeJJZ1yQG2/c2hgpR1a6MFZMF1UdheByIOPsb
lyQblejU0S6iG3UE6L9NZS4en/c/KLFl88lITN62Z5xpwICNTH8oHCaVeZKYC1MUsAPcpKM7NBo8
54rWdR3Cjbj28K9l9wHnHL6FkNLaNMnfMD3yghXf3Ty3iOcE+pUOFNRzk7l7Pco/T3Xfm0Bd30Pu
W2Z7RWQ/KByNBbEKprLMl46MBn+LpBKBAry8mCjPIiblp0mvTHyIaEwMwhcsxXGTGLFDu99LJfmB
57hn73ISUtZF191lunKwR8ug+K9mb+2nrkgyeFBQRzmd8we25a/ph/V5mEe5mKUHGY+eDgF4gdLb
zurTIWaAHS2oGh4AuBUs85SC/4k3ELXib3LCveCzn9+hCcS+TDHtD11xfxvjj5gL5WJIkeaWQzXL
iYU5LcTT01wIU3neRkuXYkFEg9uQChncYRURvDHQP6d72Vziz2/1SD6yQQKI+TDLqkq1VVL5iMg0
+YLj2I8cDaq5WJaX/Zpy1Oe7tgJnFWvHkCZ7inV8Zq274YkTb6B9owxXFD08NpsHH7PGDKm+eyNd
1HwkqsRdZBLqW8/TBJCizng9ZJP1AdBzhIvc8gZIUPINsr0NEVY7xvBrfaxtSBPtkUot2u7J8LeR
BZQPGSMom6P5FLB2SYv+bsj7X1+LF+s7Q4iF8ILrPVsuUcHe6tMg8BhUTAbrS6hXUiqFpykDd1+D
hXbq4toeACOCeciXW5Smu1klsmiRfzLuIpNDofIsgUEkQ0k8FayJgyHzTnL+11ulhKnHjIVY76SO
dJdT7yO0QEojtH7jxD9Dv14drGOtzn9PzL3RvLF6SwqqCj4f3jsV8vUR9XU7uzc60KC/jB8Mwk/u
Y9KUW887UViW8vf9o7EhayTVDgqw3stBWY3v9iauUcL2RciM1mIZLuFxf89/1rucAzanS2VLvQ1R
0hzlUm6au65uBV6Vd84FjJ0BIkBySxmYAgShf2qDiNcOccgVOX/HqulSsr27wxK+jZkThFyvV1hm
HMjrmhCeu6UFCMA20yiGYTxktQcOIhuaVIFwNwXvIgBnRDlZNSqqxheYbb0/59fl5HKzhMEUyQDn
QM18vc8S+Wa1gSrXb5rOiLYts9zVyCE=
`protect end_protected
