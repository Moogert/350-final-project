-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Vvj5q9Rm1SPHQeynCErgvbQ2YlP0tJWrQAjzpwBP2Usii2qkDUoZqai8llsQ+oPaIqd6rBldYL8x
b25SgNL54EXdia6Eqk3KLZd1m0TxUaN3nTXWRdOJRCmUCvrlmri5+jPn280wWzdg4l/EDiZWXFqK
rPinzl7MycRk6xI65GqnjManTQKJT6Tev0QlVa9NgHTU7/xRaxxwZLTORBf1iqrsFE8CDLh+f8a/
XpInWWEDb20/n+gYrWAYXonHauTxQD9JHNcjh4tmACtjiG0bCcCr8QakIkwTr6luUhUknG+403Hv
pIsEtGpRFQEKk0CobT8Bqc4fgw8tEGEgeaKTzw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
ktYwvkmQoNRss92vjIgcL/gIyAQ1z5PVY3TIbKM7Y6vkkmMBiGI0+u2KTtYBNpSaClwEy/OSmWtq
/oewKFqGIyCX6qzJQu/g4bMPMf46SbdiJ60jjkgHzLeQAnGv1hnCpvijMTwC5+WQSKt2kr9ubZIb
PD+y4Kz4rDvsplA/g5tFos3+p3aypXTJ/h7uZ+Kip7HG1UrCBG7WBVMZvUoz/5L04aPhQbH3qlA7
bC4eRrf7QCIb4KLlY+NypP0njlNK8664g6CDW9P5WyUNt7+OF4sU6+OtmIB35AbQWTtlPxjZ+Wzf
QpxKUtn80i2LncatXSrUdf2b0FwiJoOn9NTIBs9II6NAkx5iYWwF+ld1XPdQJERbQRrLQHyr+KvA
AXx14Z+unrthlszO5NxwQErcalCa4eaVd3pKaXmjbTlTjc4IxURvEksNwWlnE8JkC3vSFWxHymZJ
UuxN3gvVCHkovAJhlzwUKUSba/o+Y5t7cBYmRg66W6FK0vr/0yslxjWbamRG4lLwVKp/5SBzVkOj
/VrX1/lNCyfGRwEBc2VomCkMARBI/pAQT4/2f3mGK5KR8gq7sFGLTuWkWRG6PCnSsPd63LGlXx7U
U1TBOLtwUFmoUdmXRyS9TMxBZiVViz2ITq4supF11InWwzqk8OugFAixXFkXq0JShdAoJCaJ6X2K
rWhFZAMJPwz/6cZ9Upn3rSi7Z6r5ZcwW8ZW71yI4OC5mR9lcU8Cvno9CE3OZM5ftmfWihBffXJ2s
tf9iBzmX6F6GIJ57EWzrHGCovjsTgzFWIzsAEoYMMhvBYZrVEhreNjtfdd1RJn3r61p3vczpOxlm
C8lRfve86MbYJzd/VoTS2eRU4i8Hc6itktT0AGgxneSMv9DFa7bvO+Z0nED1qr1JhafZTuMOGgtL
Arhb3vxGR06IH4wj4yxsDNCLXv/aQcJNuGS1Z5g81h09dlnBFAg4G/47/9Mfkru8ETkwiggGDL9t
7kyihn1K0kW2aPFWC6K687sdGq9iBMj9PqZ/fCo9H7kTxeHgE4BwB/lYaogevlhHAWpA92SDWcb+
wZfZDxxJkLOd8atZjUjbVvLOMR4s6SjfRvfrKqQhbzrE2CUCDAIljlL2PhdDFdrpi2qv/YRp47yU
c63w9tpIBuRrvse2We4/d4771xVWKaqXFYQy7W06gNz2c3sPKgO1lbUe7wW/Md+Uer2VeoJwxet8
eaMYaAeD6DWzfqaHh+I+qTbVWhACX974fM2SKpHZblka7YF0YUb+6Pp11cAiTfbrN5OWKDdIrC7j
G/Hu4zrH9bcBh/YI8RqI63X9DzoIXA9HZhZWc7Bnz0CHGzxAiwp8x0ZCXvtCNZ3Fnhc1wC0ZuKaD
t/Dsqz6LVa8krm//IgkuHZbz8MouX0uIPpmktqxyngI2/fBQ/lnL71o3R5GNU+cML+rJrsHlfyBn
HpioYNQQHD+S57/uEHHMcDU9c5hl5ELXgA3c+NEQZH5TMIBoQ1fgRcjs2CG3YhMEMzKGjCj2hVQ2
/Rt/plxmoWKvKWISC+b3dSSus+zmKSvmk0AKe9wc/TmpyDGsgQcXJzs/X+EtGHRuTfw1YZLv4u3O
kC0o7CUKCSGJ8RBaW5jzMPxVdpxQbOg8Hnu02bfojPDBzzapNMmAtKnfmwojBRk/YsZfJAS3v2Uq
enUh0veGJaiv3wkAg01qNt/VDn1bic56/7u6/aE7/l70yyMh2elPEB5OtwMf+1uwK3aFFOYAmxHd
H3RJ6a/75QFbAs5jBEwIWYVadgtw8nu/4kuimbO9QEyJG+xmXqzsM2bPj4cuFmjQ23dUqJroF06T
YLXFxm6qDRGv0TnITWZFY30MQKUgIl2JbMfGlxt07uRZWgeOaFL8TkODtDkwy7m8y/t2COKj7LY7
8jTSKglDAmhRP6sASTxPG/IaFWz3pkes37BcsDGuTnloMKY8Yq8OE1IjOet3fb/OHzlfK3DAqIZT
q1rGsRRjTO32zAZINSQohfuVid2PaslicOdyxL9Y9fsWv6/VCMp3XDFlSQDjU/rXpcHdfmT5xpEu
taNeirGScNk7UOm2p5yWB7XDn4ogazYECN6S2pPSOKSIau4xvVTqx6MAawJQTPCmo8p0OMu8uG0g
y2EDCvJrakk+AKlDhyAsPkeRj0HcvXmfSQ7CLW7BYG51QZkAdX7W5aL9J0pWP05nRzO/iiZtnaOD
9xKzY8uWLKcqh6ur2bHGEaXQD+oenarO9tPzTdEryUVLRddO3ImvwiDt0LlEV3XOBw+RjHpgDtJv
OwbTpTIr7/vTKUEKjKNnymNW9u77NVXpfhqMBSQ2AfI/E6FZt9Z6+QGg4tJE8kvQrVlHrVS8/Hht
9SGrCvseQZufIOiedqwyoxFVQivAv9t26xZkc4/ltVLEH77cOgo5d9ihAAp+gC5KG2XeMYnodktP
z5CEi/Yy4gTt+XlAswGsKT9l/8rXiCpn4Jxjs8oXnGyQEQkkLM5J4ofs1Acpkpg3FegUqaYFK4V5
LwehYHgLL5zcgUPxo8/OHWElL5sq7ZnQyE8qOCu1MKXncYpMKVsLDqUlJpEqcqdeqVPqqo/edRbM
Hkr5V4bIBj2yM1MlRUNnsWZAu4EcZZ2ifQ6Ok2HdT6LlKNEMQn06UnViJE3UuD+cbaWyGX6JS4Wo
DMRwcOFzgbFkafRaCEf4dL0BF630nzWH5XCdpeh+o2TYfwFp7wmlVVFkSByEGdFGyIjIZ8n1q/kS
gTtzC4F1hiPL9cBI53jFr98E86dJgTj7os9dXH9UFSEETqKUz35hiM/pnY20Ma2fUU9SLvLRMwXb
etI+S4btzqi4P1s7p8vi7XdfsoESmvHx3ivNct5GALlrcedLf2v/x4oI6HmabKc7rO34u39b4ljo
ON4WztF963Cnk3XpPEWtnFMaqqzHNnDfPqQSsdBFoW8TqcyK+YzIHHUCv+F8kVJRTtCpCng8KRuO
SPHNQboxnF7uNX8lkZzMRzr34uXmYVmaZ/E5krpXrxb9O3qOOi4HITrM1NogMjVZ8c1buV4myhBx
nz0VX/+QobxZblN1eFQkMUH3kghVIvMS7SkNeay/GBQxIzk4rbR3ymew+37JSTjkpV7bnPui7NOB
2FnBKtyG1ZpzwZmF3gm2qG6HH2pMNvxqM4vZhiNpjoJ1pa/pxlmXVnir/09ZltfSJ7Sxiek3CEoJ
4ZOrhadqmHTtLKdyozQCUNOWlmpZJW+hJ7cjL2PqXyZSkq2L7gb2awa8AYoZYAGwKf4zfAelAAzP
07wVK08pVHW5I1vsf8mWMbVbz7g9sl4PLjVuGUNO+Lp9axlLhHCTGV59KM9/ywFAEQtGsP5HM3t5
C0UC875lWx/upauilv5pas1YJ4wSp9jtukCuMsb0Ktgeb3GcLvNzEjqdW8XfWdCRiPhqoMWinNdl
Y7AwFDVlLbhfU2vJrvqwMQCdWYn+xgrCI40/G39GlwQCkWasSmlY3zqS3hcRmlKuVqn/Fq2oGmMM
B5fEgBPDNeUnk+2U8fI2qC0MI8FRIMNhr/YeLVxEGLp1B7F77zC9Zcnr9nFmCPCbK8r1OHUZPUnL
NlVCi2fwzUngQmmIAnTlfQhcnQ4Fldd22MH4YLuJ0ojkaGoPFK0IXK2RKOf7Jgpu0T1PBYbo8/tQ
3jGqEcGEK7f+B2vJj1TdOhHxMwwYglBN5JDhEjCwukA4sKEuP/wVKH7UQGSucSBrpeE2qX6uMqt6
yhi2K3aRLAZHOXXQ1af0a/RhC8JBrIgN2/Y8XmG6zT4qmNV7MqX4qxv3CThsw5ydUoAY6TnntuF2
Zvv0B2KShBrIv91Cby/rOb4q2+XE+OVfHFk7lbvpJmYCMYfcM3qUP5BM0ZK5J5DLTQsPDGt0nwtc
jIy/tSQ4u/jUkZmSd4jwyyGeXiewp5gfjlTDNmoVy8JEdaVstG6Efn8vMuUTyEYcdOD8OC9P1bqz
X5U4z+tdTA/8Jb32XwJoJ8fTty2C4jW4GDLvg9WsG4UQ4wQcHFkTG0gKVPRxzteT9wBYXdvcXFrY
BQJrJcyyF3UKBpgVI64FuI5/Pa06xPO/7iUhrCfLy6dKs4//37R6q63nZkQ6COs7Weqj1t2H/C9b
B9m5PQgt0xOqHv625LFqZbBZ4r/V4E57V5Vz2Gq4OV60of+xKNv7SWsyg7cenQ7vpV67NYWue4u8
n0Q0AiplpcEbhar21nLwysADrTSbR9Ouqr0S1HGI8Bs/paixhbmidmRtm111MWOhU0Ehw37aoMDl
ZtGFNAAiZ5lFTfX4ubOsY02Zc4H+Z2cgKPxby1gHHnYcOBeGJZIsjoQvzTYLEYnIvNy8Hiy2xi6m
EfVEPHyuAcAFFoPpcFBRRw6rZhh3IB3gkYSQtL/sHVC8tgCBFjF96B/bPKu6BrnpwLoGnyzQqfn5
zjMdPnvG7SQcZGS+SnMhUIKejyLSOPvaAOGmw4lYMJPiv6sUwH1ep8U/jjkNiSL6AyCf33sdhr/S
9ReiqxVHb3e2pC31B6cmEODG1VordR+S2q9dbgJ51PiYwhua+u1EB8U4nIlQm4k0502zGK0mUMCL
YhP7IbCsoWYp4D80JY9BAuUBStPkDrdOwvEtWdMbt40W1NUC3O7fa8WqMlj+Zu1D5CSul5782h2s
Mq0o+ocaImbazQUJNMHxz1MN/F+kFxi+TwgC61gK5JM5m/IWM8G7n6eLSAEM+XYABBBnBDVlwZ/9
8jkoSCey9NeL7EUVD/G5tRpPBakfoNEcXZI0eev/W7Qr/o8wZ6bKRSTF1Mg2Ma3UtTlO6jsfJYf3
Clqv1aZQvYJmpug/R9jvAMWyZ8z+p/aBEi1oPTCizshDR8SLty6zMzqjQGNchBfhmZC+fLJ5NdpX
79LP3veOQh8w//fBgqDm2241TOdn+gSvjcKM3akpKADm3ZhnafAtKW05d1vda9nuwjtq9JJgq6ft
/tD8xFRRvNDo7Nqyu2PRDnXCqYTDri7luCi3B9t42mYWjeEAVhSqv9OEZw4W2o8bGSEbUTeqmdQV
4bZGFraYU6+QpOrLwtQVVk5Mu46DWnFTYk6/i18NMROGLQcFTn4co+XxZ4fPaKgbVXmu/7Bn6s2X
YWfOgxengJbm5YAIRNmdFa0RPw7X098C65rU4J1jQDHhUJ/t9xoLxfW7yxECgypLXNBs6JkqoZ5x
yqfO6XONyB7rv8g3iUW5Hq0Qzm2KgFkiVrSFlHkfrZrYem4+iEflhJFYDZefYLhdLN9sBJoSqm4X
wn4kyT3CTKLhyx6V3l7oXNE5q3pZuQBKcadDBC2fsYg04++ZL0Z8i9JxcXIBGQubwshISFIe5vVt
S+mbOrIAzLYMbuXaqjiYRMF8qzLGsemSg2kp0PgMVSn7gXSLQG7PFr1aB0BZGouV/DXJkjMXCK8e
dVGngHZfannRexqXS2D8NhucJ7M3tsnA+rhTA/hVBkS6+ZU4yVJUKYLdizyGN4AIRxkQitDVHKjJ
OjGeZX911uz82Lju/EtgHNMx3IwFADhThdqh390i575L4OBqkb6flMyOqc3c0QnzhScqK9W47pEk
V0FxV780HjSG3QuRgnZy5UFmJy7ZbCAYA/qdD4BYQi+vZIutUj5uepDf9FcJ3bHBRGh2oGLc+mka
8iEXLN1bxEWEjPhxNJfx3FbZAKhNKjT5DyiNhOgewiiXn0y8MlOr5pqdwSrQ+UrhpJ2LF7mErFv9
Yh43/xz+JJrRW8qWNaLU2YyKcJhZEbcN+B70R3YUgEx1YH7fkULhRC4Hhmcj4LQsgrhpdF+2a+IH
0wwW7Wlkee5myDGCqKZ1m5SM9saMhFItAeWm2dSpNVvNevR5V6+AAx3ecEDqpqysZqwVWz9PuS97
rEA+fFTbi2HQx6kwC2PHDvimxtfzqrjDvsQuy1mXE8LUpsgXrCg1zx2ao/qgLelJO/pSEgNV8S2K
N8rZYvnah1LivOMQV82Oq5IKdijxyD8fp6J9SiUPG6EQyWzfuPEIp5U+t7JjKmpODWazlKxkZDgJ
d2sIo+lwaS0dvPMv5Ax0/cJtbSVk9Vu8CArWmYZ3nINggbAOYtHBgdHYb/Zs+7Lf+9iZkGcckcY1
Zvps7TvehH+2eE9GnrHTD10AAZx+9gpD0wtulktFEjFfWlUNedXRRoYvcRTeo5j7SNlq28wr/lef
bCTH0aOdfy+3eb0Gu/iw0x08sagXtEMJBaRkuvKjukURkk9M8pKEguWyfMtx3gJ8DW5MbE8kIFkc
CFIHEofehnXr0qUUFzYaP27CF9O6QuHNIgybLFynOkFuR7VVvmeMJ3HMzMS2KCF3eJCnapEo5eE1
sIFSFDB47+/kqycmxl/We8r4YohiIc+XorgtLwaM4CdV4AOU4zLJ2iWExQFcpboJ2OgGwIqAkST+
pTPKElmGOXZQHravljWxTK8qCgSzwf/SmzgH6NI2slymtXvk6d6wFVq3qOVJU0uLImeQ7wLja7bX
NySu7I2Wb2w4+P/VyID9n8QdM1ezhUOEDfeNgfjUqyjN+agOrIo/iZ1r0yNmiFBSBLdVLoxFwPcX
RBqxqcGwHEQ5hh8Rz3xBRHApbFJNBduVsXXTsh9dOEWwhuOkPnTjnODMqj2DJ6ULvBlOTveob+U0
u27xHUDdpat0IhmPM/ttZBOhEFOERDuaFZ4eCE3H1CcDQPLW4ZNg94SYClLR4p4c7gcv1YIp/zYk
wlPADtOTe9geZeOSYvL8QJQwXSeI7KEHcbMQjNtvcBi31MpagQbWXBHB1gpAm5bWrdSEgm4CUKLa
xpl9qszI6cJEsV3XpXSwrTk+pRsgbHaWGTfGs7XUEVpWupKJW6kvO28WtJ2sCkCUbajXhwTRwICG
IZzzdN+ZdUBJBJ6Q1Uot2bfwzIJMGvFP1X01GOl81THbPzIpHBc3ro9/T/TEHmA1CVIULexg5S7X
bfn5Ws9Xen5b0QJKChf+nmQvjEGz+rkeFkqGxxclcLbl58CnoqRtc9SB5EPPugvl7v+o1yl0yOT+
/8Y5iTD9etDwicsHp5SmkZQPeJO4ygK5WKeDi2k4IbOu4zD3wJG/JL4I0RpgQCnYPR5sNkVI0C3b
NB9hplhhLXeJeI+ePTVzpIbtz7SeD9/VkJClFE2mGllFaKIhF7u5QuGgfFUTCP7dDx3vmQDAICTN
3GE3f0sf365pZRmr24nl0vNOLZ4WVcByqRn1cLQZEA9MAi8VRIg+2Rvkp8DfUnzNF4rXQxrTNxfh
Acllz573RNOTUj+kNoGt16i7nvojUobJTIi61ok4big6v812AMou52m3/dmHSWD3hdWR2wJuFcOU
Ng7wTlV6yBoqy3bgp++tfe5f8fbFvkCpaFrwdFfg/Zx3m2DwrIFBeltqsKX7gOSDvFr/Ey6hWmoE
wVN99Rwh9bhLZqGYQwRJxa8X2qxmDgv/o+pQsbnB9LjkR6QIUOmHuq7Fld6SuvyqII8Tooo0HKUP
TaGDrKfurelgR34OMMDi4TpqQrjbY5r+gPExYdb7W//PhI0jBXO7CQ5fGzET3eG0szSVgAf2C5uf
2EHryZ/3ViAVdIQcWwRFGUuWnZMkmiUx98Pf0ionBgjxOVDG88QnWy59Vu/wF9w4Zrty1mwzLWMb
9G0OSNkMPv5dzhSeGjab88GxWxATWH/BicEXjt4Ffy48jA790+6nN3ENuftzKEuoO/EQsjYGA5wz
riQses3YNZa5hMOK9YrAK/L2wJutDQICaJ96dju4sdo2r+cXdSolkhcPZ9feiYY4WATmkSxt9/bz
dwrGnloS5NyP32QP6gIdPpTkS5fNYWVTAgmFomZ85FTLuwoNKwolq/9TfX1+PICajTTQp1F7snua
qCM+H3JLywOe4L/cVikRJOmhI7MqR98vU8PMD5mD/j0OAI1Gi59jxVzCyB7fP/bQLMeYr/XKPrsI
UPz6F9apiavn6S2jcSj1x8cBMbDrq84imk+a6M+GF2PxbtyJDWx4Vb6AmLd4132ziTVuRZbQhRvk
nvoZOs7ry+l2OIUQ0wd730QS2T4Gxa3DzgW20Ztc8rPVGudh5R/KLSuR7GypmL40Lfb+AU4ow58l
St6R+H/UjKRUL7dulMErE26sqCvxl8lCb1U5cs5oPcCOiAtFNM070sehxx7VXTTMCUicwpY+5dnz
eaxTVD9mqNOsaFNPBZ0WUttjzD3q5I+d3LXccGjxAOSUw6jZDT6oXwbNUNwrs7lea8FEW6ju7LRO
kdsHmUxjl82Kx3yeuqhfCEBCAqu0Zhj2gTdP9oolzFYuGhSC06RhyPJvM7hMavHVxRtoSgN55sgz
CxOEsBbi3//pzxRuj7IWaRMJEHA7oRhjaSSH8rq2SGkybWAAg+RbVQHuAovhnoBYFypVUm/m/yMt
Nt2wiF+jqGCck7iFzHdWNslyPo5sTAfSA5GVglSg3nDrfrP+wSgbEHBHWs7i9WmeoHUiewSyM3U3
j1dlgrZN7KGKymxCcVzHqZtIiMbEG5jQxcCJuhjcrk6YuZGZCrsNAbAvsVjEky1gUVyEcVZk7t6N
tW+PP53JTDDQMSP8Rl9poNOLbWJRt0iNoEnJDxavd8m5D/mnyi9suDamT9ejOe86pZag6NnqNOPu
SQ7hVxutVSzqaDm6Pn3uUxIXBXQCIPzzOppKdcAwYLmwsk21IpeiesI5PZZLKuuVPnShvpjmkzKu
Udqj76DSdc6HmqLmbKlERD3yn1OazTper8KkodRFH7SlV/ddvytZZKQWR/H7SLUlf+KeL8fvqrQ8
tZmp2eg7UjvK5Qv3TRt9vWAVgrqJaJzSsu3QRDyujsG9ZXS7JaSidaye4HmEhIXT02FjHbOqOpwU
1u3IDE5OOC3+MWZVrwN0lKcy60OohyXgxr7E5w1w5FtFpCjS3G67S3kmoas8aPlYM8R4BVKpR9Xd
lujMw9KxigUTw8Vcq0pdnq9srxVZbW/9rW22FBGmXcu5jaQhVqaS/AL0543aPtJMZSYMJ7ZBBsbP
oc9fhwhDj8+iT99GwUiBO69VkdVle+XChqsu5/a48kmdfpdVC1SEhvFokHNsNAtPp2fG586RWwSj
7oXJCV7Mehti/4EclU64YgbCDZGr+uJE66xD6E2EHoPzWxcbOir8xxWI1SJbYbzIiKBAUS2e0OLi
1MM/nC+hL9ek6Ro/2erqOgtzSz7cYTATm5/ahcgpKS37rOOwd22yA48GR7UPbSZDuc2bWEY7lz5I
fYuKohhJdxWUDka2QmYjRCF7K7EcAugl5YzALZQBunAW9L/ASHfWE0iMlbLBDcXMvYrfah5jKM6B
mDtYZquQGEJLTXv3Rw0BfIIkS92lQGVz0Jnk9NXj8Gn0G/UBiZClUOBZbW1dVevSjWGxWRJLcjw8
cpjkwCaOmilxSJJLfffMj8I6mWAh5wNSFhJwyA9URM7SddNZQ4kKZea8SVNzNjO4U+hZMwFcBJc4
/28aXxPVn/WgrqnN+j3Ttjo1rZRRNDxClbZ9hw8M6Kq7ZWs9b9pPXRNTS6GMrS1PhrWkr+zSpvhd
Kd+Gc/vpMuWDDzB4l7L+Ra7V6D4b71zQntrF0Zn29zXRuLPM4RJ3jImTWCVifhuawTrTBJQqc/80
+2hiLu4b6PnPD7s9u/EUpKWOSSrjRCFGOBfxJSYRrh9KfXLyKZxOnNgtEP141d9HdlFYHuvWlChM
6Wr/f1ZeogWTHRA0DldyNnypRipc8VyBfxTqajcvek8Cv7paHBKLT31SZErEUlAoVhziO0WcCkAq
x53sYSJmHXBoxRBYY+aBCEhMu/UHj4HtDkAT8OZhIRQS1XICyCIIPkbXO1OcJGgFNo7uuUXJ2RDd
slB6R4l0QlDd0ijSqAijmDGwTBcUQSnFMHW5e0NT8mA6ldzc4QGCy5b9rqUUEjzSjkEHprIC0lUK
rlvBvbMKN7SzpltpDpfefNK/MUn9eYnjigDizvTx8bkUiMzJUufSBpmbETsnYDTzJmSwEzzpO8xH
asenkk4qs+Ju/gUg/EIviUcNa5OCgJF6jjCoWUl1LK5iIhHrVZO95e7nbekPiz7JlWnc/Jny3cZX
emMEhIqs+IAWbGvYkxm0Ga2Yt8YhlbDOnx/Q+PvLgWdKidMXGgoVKXWaHd0lcpytNUJEuSa7Wxwc
OqYQVUZJcLPTvkQs5Ps7EMsq4uO65OIwk3/RdyNPYdyw8yfi38yJu85I+sYgjO7hLkf2PiZq1vhL
MDWUwtSmY8aPAreF7TXEAmQGw3lsHx0v5yKGShLDGl2y20JyiRswjPOWXKQLvQmm3u2ooXuRcABf
srX5NLOoK5GMYSoIUlzFMtTmGHbCPLcs1YrAec8NF/UsObuW48SCD4YRxz4XfbO5MbPkWHtiPJ5U
7nhGb3+hR6JxbLhtbLLB3A5yzpWFlDIAwNRP6bSZid+k0/psi1s3O/93HzrVZjwmj4g5NQgidhGV
Xgu1a38Em90shnPuklph6GWHjKMLNuKJCZ9F70CaIbY8znmBqp4HCIUBT+I/AOcOqENsH358XEor
TeClO/KnXyJ3iGUOYVxNWJVvJJosIU7GQQ1UU0N+6yXabft7CbSfOMyeQ6UELie8sHagvpV1piq/
h/u5IaoUcYPBfh/5kpRzCYeeQuUzB2WPGTKzkI1xHKQK4c6QgVok4txgvmXBgYh10BLutApEVrNb
yYyCSFVGL6l2ITSdYUzmIG4nhdeQ8cRcFY5lCnK7axAho15HWuzUPk4Ez1qQzf8nFgXgmJDhpWjM
GW4oxdOoCs/nx+SVPvsvTf1roZadma4jDbnKIFiRiVYK7cBupaEaqYAXkEpvAk9/bRUJEgaYXCq6
sGAF0ynY+gKIE7MJneHZgjucDaNIaE+OjZOGOFX0as5IUPtRQS9jnADrAT77PuiFPkaOlyHtRwBo
HiTsIzwZ6Oq89VIFsIIhxkDrnm96oCHEki/BobvXvEa55XWF72VDgtc5JD0wxdPgiMvUBFLEuHRJ
AsGji41wxdKrJSE5cx7lbgG9xVjHx7KSunrSnqs6oCzY96qPvwjYE/OnWZJs8fYDp45ZX64nn3JA
g4V1kfb8ucNNXZx/VeJzznX774UvbVBfxdJPXDLPFcUn83bJ/Bd6IBKG2VK2ZS2f9tFBGiLwWLGr
YEckuBH1qUzSo+auLvhWwAn9fhJV+HRnYDZCmZY1jopRpxFJQtOYWx8+7hnsEugMKdSm7icFwDTL
iv+PQKY5d0FOb73F5BBk2/z6pO5lpdHGQL1v7T8kbOALNzsaeOoVD7TgDIe5pN+riYrx6Ceb4T0K
x1QO0NN4qDIl+FoUQieFROrz7Do+y/2Gf0tLvJTtELFn56XpxJyQBrXn+TGEquLvSbczXRiYBgLP
qI4GSH7aDvzYXTRo4YdRbkzB5ESpiqTS5OK8asArcBaQPeYuKF7+BPnZUuQo16EHeKDfWtWZGLkl
9zEI/0IUBapE6hNG1ZpzS4WAH7I4SVEzyKqqiH4R02IYE5cCs3JswvU9VIhi1HL3kqL80OG8bZOd
JOkLgxzorxOcCSvIhSuXr8NTOUsln13WQpGXtOXskwU7PlKkVuRjxiyG0qaXfMIW41M6IsawwEHY
5SPmC2YxM+k6yIQfOM5K/DI3c9mdUUzaF/ly2nRs7kv0pbhvWYA9RzYq+9pfRd30F+vIkm0BDZCp
7F4El5q41V7tWc0XoqRoErYcIdZMM/Yh0j7K0PhAM2jNUw5QGpWte8BTbDNHDM5orNJw1rfYwVJH
LfM2A5U8NiS52Xn2QhHpQsjpj/SjHRuH0LNkm+Q+ZrfLnjl1tkgzs72gzLKCyOMGvhErgCmSALyF
/131tDr6lHX8TOhb0HVUiQ8MNw57DxYJXvvSVROJU0omQtbTlPrMWVfT2MpGGZLxGq5z/TxlwOEe
nUkAKr4Iot5Yxr6ReKUf/4WCVKxZDxyLHIwsOtUXa7ZMLzdrrWDvwf/EUiibHj5pZONDIxL2JAPz
9VAdMA5ABiw4aaUKKSZTCP8lqcsJ3ODFUiXiGhfnilsjkEtn91WmEYDLCvr2zPZqvujQSsBB5U23
4+4S7cqvw/2SUSMHwrv+R57kJfGA0NsE2waQ4IpuecFsHJEa/vKbmmQNM6ehpuN186JJ+8EYFfFA
T/WH8dVUNKtMGENcbdhDXYh93YZfV8Dl2JjkILpzMBgu53E6Zo8GznuCIll1rwe2y/EpCGIKLHNC
Wvz6cHGymnUYx4FrKolMqtUgAECDRvtshO4YFjwE4euOyLPlnQT87NzBtEG9E/hrBBgs7xphgNro
UTIk0OlkbDpqrWDxTTip6zdkbZ4zPZupPtTWSZ8MM0t5xTkpk0/2fSeDml0M1Gps8RkJphhAiA9X
28tnFLHpmCo51E2ppEnfv8hpX/mrW/z9C24xV08ITgDZvloV7h9GD3lPTHFpFJqzfnVkOWGdbC7z
M0MvRsH5gHYi61RbCRwMck6lxoKsM09XhMXYgRIAKNZ7Ez25Y9qO61E3R/qFsqUeGRCjFB8OqcqD
Af1JOx7Jq98ZKWZjkuN9RIKxPMKb5c3Bqy8HqoE/nIHdVMiEB4dF9VNy+1rDo7OG1M5W9QYCjRFw
3zzSeGchzK0dT7CmmU5/x/7bAJZ/21sw/S3DQ1DYuhelEhqno4BwtQHeOiAe5tTLOG8+iYqNTdl0
AkR5ysC6GE4QDLrmJUT7UiQOKW6zoSnSSQqvpcn60r3mI7ZRNJRilIJR8Wmq396AV2pT+6vNozPt
bx1NEzCodkdRY1OZUubJqOpx+Vq4Z5jfS52yClSAJ0YTSvQA7ofV7vbSnO0DvP/f7ISPBtXeIhPk
wuYvzkcVKyKRPsHNIYe0KDXrwvAh/xTMxfk7/Qdk5cJFSIYaDYf02PTBmIArMg2o48T/b2runRzQ
9q2+71ZxMm48//dIYjCLlRoLS3dUJhywVouxFD10CgCseOcpV0vQe8QAYF5Ne2y5FHn5oNQqCu9h
TE1DdG6mMSlsrj0y7oOokUPW69HUHPhMZ60TWr8pdfyRp7xg3OdZ8SIezhovd4j7zjIqp6JFJQJt
zwG3dXKyRs7vwMupq+I/mkd77YhE7Rdhh5pRk/WrUOdD022gIDT8OwVarG9SrL97Fm6GD5mSzCbA
33vTLwP1tALpIvsTLVZTfV4IR9O+wZ/jcu+F3V7jlTXtWmu2jkkE+cdK4d0THVIM1YptFNzEGBvc
MIx8XdYqCcvuwf9UewvZn5kexWySuYI7zMue2YHDKYmvHeP0F9ayhV+juTytyD4Yw0Cmk/OMTRe3
fds=
`protect end_protected
