-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M/QtpehdzK3g/X13kk6YM3q27GCOEXOzm0CrnGj4QAanz2Ej2Tu1EB1qcLInnpQvtMWUDdame0+g
Ow4SB0BdI338maeszXmXyHCElaZcO9u4xOebAXzZNT+ozvT7j/u2+xrD4lnGpS0ljdBbmJ7DowKZ
8ioNl0H9Uk+hp5CgXq0Pk129MjmlItQZ6xL/v7qctCYvzTKY80fvqKqy/YMjW2yY1pYeIJr3w32p
7dSRiPkR6dDclBh3kJpj4ACXP7BhMcSMtURzyWMLLGwM4gW0ckBVG/nFI+0DkJQoI8bjAqKLMf5F
MIbUHV4yL/3gaygvwQP2b7+ZGImSlSSCLdN/BA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
06C3x+t6N1BjEDBkFBXVV2OXOhOGbmja3oCul0nwInJcDdguDC0I2s9AfKfXZWEQTmm/reoFWwm6
i0EztTJBiH1H706eo8lpt/tz2dhYoGAsMOK9NpQ6W/yyZVuNpn9A6fcgVJCqWiWLAbw0ZAgycGlG
Pk4E7kvllmgz7JvrFU7gtUnGYI0oDBzn2CZUwPUfPVTHSPH/Zu86HavA2Vcpps8I+vlcmP16E7lI
RjbxONbsBh6fxUg0drWSfVjQvwsgnVefOL1T4MwLPwQ5QYqFOB/5WEpCSTr9H8EJU06aBezPNmus
sWJ7FJjRsTqT4/miwn7wyEW0DLkDTjCfPzr2Cmv9AE99BqTODzYQYY+7QKQQqE7kZ+B8EA2oNRrM
3ltEhWzY1/1OVSA/qyt44KWlUUfpB+ggfrRMgng9Ezmd9H3/IZ0iVJy9jiumbZYUf98bI/L92vWi
nx/UDkCPbZ1rDUvHZ4fQtDjMMICwPMJflSOFhMsRhN4chdHE4e8mPhyIigW26+CVQuQhlOjgs3kc
sMFTBz6WN1XMwX6la+NmcKCwe+KDQfymg5Uwrkol01CWHBqWdsfqWpG+871qGByPnwi4iqG4M90A
j3oK7megk6B6P9v5WUopF3lt05JTQbigEGIl/5CuIrvwjfv4gOTTwctaUrxm/+e/b1qCMyABoSyz
07V7kJVl5jAJHngOXkJA0ctuFUept8H1ocV8TksnBk0inJtyjEjDS4JCpZRzpFJJNd2n4kVcosqp
zRFOgI14xkVQPbGmfzbex8KLeQIcuaCqMt4qKXWi9pdIcGqS5Vc3H+yYrkjpyjJH2aREVsGU7EqF
psgmi1jnhd5ezXPd8xRpDkQsMYsERAJyK9aeX0YKxsuHT1LAp7Gl5qFSJ3x+twTIioiGno4+WlPC
akfK2WRoEpON9RnhnHvtzwAeNw4DWbn+wTaQmZvwx2P833WDDQBw9M8SKLNd6HF++9rPQglK/k7x
qTNUvEjCxuTZrKMJs4ONSd3tTeOEtG8TYJDbowDuf955f4IairGZ7qx5/mVQfl72rsox7giUu/cg
X5eEBe/WCfJMw53shtP/eCHysi/xQzbwVcPVfa3Lk/tbChkUSWinvCjfHes4bHOyVKiWGA5imgJ3
VQ1mB8/epQTXfwMwLKicqEspdMsomnTz+z0ySGFzEVQ7skShSsbPEhQpREQfo1g6K0MGEGb/QaVg
8OdZM79cP40GrRj2NxyA8Xzv1ItDT/N8v9uj6vmaQF+xVQxhjevNQZn5FCfPsPPtgpWWRFpi1dNW
s3Q1GtNT2DtXqQb86C86LC5/cQZqj37Nv3GzL82OROy9SqgXmCF7mVTrJPf4J6dCKmmsHW6FjehY
Yid2RkVAU0qk4PyjSYEOGoc9o6LEfWl1g2vYBHFD2l7ZNGfIUX5wzK9PCtmqUoX8/PaDKDOf9IU2
10cOWKOtsFDUbD/05uxJcIC7ZG5tNLxyOPKRKoqtY4LU9ZgYxoNL48YMPzbdkZ1PDrM4UM/XW9bh
IkGw4GpMqlCyacnSb47LgXkQwmF1JAu7m8nS1Qx3deofUR+bjdCiTXD4YrCfUHkT5JFcGDi1S1/o
kz6wrCxJstsNpxNhbPo2FxuYJqSQQR6+lGLrXgRc7aEK15FfvOufBIKLLDITos9+N1lEDpVAY1YM
w/zB5hJFVj2ZHjExudkbsvdW2PPb+OSDHe6moRyudBs+EYfXGgRsEbPrZz5zgv0SDTt8ng9MloGg
89rJHa4E5SmYfeEZZHxy34qCerGHgg9ghfbGjsHFpYvgWfikhIlKFwHnhLeJ6UHGb5L/jySZvNfo
gYYT907xEqO6+BkObbNxu42RG0pNxQP2jm5ZktVOYeLKpXakAjWMvL9dNNo2M2lyEXma2gsMR5FS
U/RSZGV6AI0SjbYBsl6/YXD4+jt5w0HMznZd8O1mNiHb7B6xlA46CQfVhQbtKMhVcgoFP0M33kA1
CE5ImRU93dKRzSBVnqQ9PBLy2k2GhI6si5V9BX2scF2sODKp8UugtPAs7+OKMUKv5QlYp/71FukN
47JiG4LQ/KiqRWPGkRb9QWr2j6Q08cumMukQlGbqy/2EPWZ12jhknxZ3jdXc1mcA5Zb1Yvua5Lbr
C4YNspMRdH/ngrZxIXHPnb6TujAIcQDiLgERzRUjzXvzEbU0UNOBu+EUsEibkjpsyjoKE1n+2BNH
rc5ZA+kUwH8tbIUUu8huDk4sgLZtCEXkKd0fWZ8imtgW0mYeG/uYYXg5Ji8fldBBJVHn5ukGjh1y
kPFmmsufaYOE4Ul2/Ok3LIY+sDf+eF8PK6hQMLxzR61cA6NhY9q8f7pFpA4wmbBl31z2F9A/CeuO
VupoBKG/PbIFVc/P7115kDu8FQe0CDLYOUdKnjt6BVwtTAqtZFEUcpHSwL9MKBFnUW3wvTOOGSWV
0WjhidACkNHWM9XMHsPUVFcZ//Qr3iNsAhpudW38MACrmx5/7g+tBSHkTXhJIw13+/Ovl7t9GDtU
jnmtt28Q+GFNDYLNLIiZq0epM/M6y35TXbOc//xAEkpjP4vZKS62bJCnMqPbUQrhpTVDERj/ovmJ
PDgyJM+WVAnO5tnEepg5ZI41CMAmXlbVo3xXy8iqpg6CMzN1jx0L0xPgd6MZLQyn5Db6REZX3S0b
4NAMOxLOTnT0jS7gY9FvP7hv+mTgHBNcIc9P2SroF+rNTt+h5/muwxFR4qAicgK/48bzNN8/4zxK
4lySFEbt2he21RwQ8zPdhPyx9lv/tS4Ium3in7lt0A508NKUKMAF1IrK9civ0jtr5ZInYDWIqF7c
qThPfA4cI+QSyTxwkb6AcwDdtty0B57MJAZ0FRL+7OhkD7HFyNC22ytK+ET4BjqG7IqVOTa9pBhb
7UY/tgJXd2qj60hHu2lpkGwwDEaPdZUzeTHQXLHoOZjh6d+Iq9vtpmLK2VJC6HSwHyZnmXolijoa
+n+S7mTXoAXHCgrh22a+tnBbi9b5A5PH53Ux9ta9Awg2Ae4r51m4Qv7QKl5yiSnwxMRR8VzJ3Oc3
8QnbXeoId0j4aJLuOyrr8Sb0B8sk44uIuUtTisN4+gba1GLOQvuZDbB+isrvvIoUyyGNf66CK5ao
9X0eBdiFjbodZCoLGE9qdUIkC+TkxpvIb4aBm+DLkgLm1wyaHlG9/pCTqWIUt/Eutf2MXdnpKiqt
wUM/jOOGcQV8NxOBHJmnNA6+4csNmSF+4i3Gn/7nvkGrOX7pqi9d+UKgi5BtL9UTk0Wh88FjAnww
zPdVIXfLxCsvrEC4Axkxqsr/b/O8TKsqtRPQISTnnNlDOtPmIzbU3ZJroIRMhK+0cjyAa+saVF4t
TeRMqYCIHURaRGKvGuxoYdw+6kmMZTxghs5NbjJ9+NUpt3X1j044Tpty87MjGY0iRJRlHMj8DlFT
QV1jBcJXbnZb67Yp340MV3KM1USnaVrsqKx0teK6P97T5ZXHm7OC73DNDOApnRXzC3iqb+DlRneG
BOs3IMGvSD8cYXlGsgIaaWLp9MEQD+v4NS31ZzM2i59jeCjjJksajfJdA0rhMXlkP+0cYSl/HRx9
RNMmlAVD27ToISIloWYKISTKyEonAbuaxkuN0vWCJPf6EAzga4c5tot444QDQbPqWfJS0ttLxRMo
K7elsNraaqEsjG+OYcddISxO0mKA1ztZqOZQiF4n42m2bk4inda3oPeKdgsyWXpzFSb/6nqUzLai
OvHlXOVHkAlACJgVml6bbEWxr+gc2qzk9RpBn7PjCL6FQI5L+jGThQgdMr2M5l//de1OP2m1PirH
ACGGD2AuZAxxfpFmpn3sg2mW0jD+B9FJ2xjSz7d53S2qLZJHaSKg5SCx6CX8pC1EbhoaRze/LEh1
M0cjuXwNxFMYyFa4Z8LMNiSejN9nnoDZ9+kVZj844EqJevXTzfpgooJBuTDqwmM95Z3hzlxGM3gW
9Mfu+N5lBv4d66TcnW61cGtewrnP/Y+9b9Q79nFhP81OHmPIJMSab9C/0mqvL6QYITAwfiZvpKzf
stDMpoOnHzBywiWIf+PAHt9qy8fQyYDyVIl/cl+rwsNkOIgFwgbPqqUNjRJCzAFQuequcpDPpF0Y
pmhzLFutNHh9omvB2HcXWF3+Dg/7xqp/4KAhIO9HjlJ+CN6eoHCvFxzKrUgpyUQ1yTqpOs/HBWId
RWN/xFC6/wIq5eKvdMShgaXued1dIpzaPv8A4QL/nofu7eEaYISRf+pa8Oo4ofDxjcMYorWjac9K
Oisjk8XOLHCYCtE7gqvTvBM6xu0U2IBPnk3JAUL1Leds2iRAN9dmrm0JzDGUiEf0A0TiQmIHaMyJ
lzJ8NIM9O0jxfCJe7xCJ9896j+ZPjzYIr+3iVsBdzjD3W/aIx6nbaxOQVXNF36YGvD2fGdOZO9Id
n0U2P/0ODmpWGRLTlxVPOzhFkj6eHuYCV8vL0Sz4F7WEwnDIuma5MZd81z2r8XDh/Fez7VtVakQS
pDA1UJh3q8IIXzTeuo5B2mOvj8qfpF0jfTgRTOfIHfSoSS3eqjtUi7PWBHwl07vgwJDVtyId5ODf
VioHHzWvNA78w0NRz62egYQgomW++OfpM1YmYvMG/X3err3fyE9XFDYHqj8yY1dODcxcoXeVe/lu
EDODBOcahnYxP216LucdONluoEmXZL0xB8GTiQJZmTDd4h/mPhXuMRda9ZJJeVIeanqR2oG9ldJW
kZf4uzNGk90KNeYBVq4P1nHlpnSomXyN8pKeMSBYsrCgUm+9bYK3+h1X6nJ/iTcYyuUpIJIiuqjA
iGKwBAHLuFvnsbZGV3WvS/7W5mkdmM99tNf/3ugJWUjMDuxZbRsmJLoaAyWzjjw59GitErWBtlKF
XTtLjAfcZTrufQmpPJEPZri+1Vf+x/RMOML7jh4berZ/jdwXmyprqcFOMIIqtP8hK29Z6cRL+SJ/
kiv3m1kam8Xr9dkA6lvCQwhYZKeNcurWqowfxATwuPRg5TOyD9sFKiJfG6zLbXS0SegEEArYu6cF
Jj9UExawbcxNmk5f6ImwF0Rm7bncTHDjufGU6y/pwLf6RsnBcuTr9FIlA/Rq/H3TAEa7RlS/siu0
Ib+fp0ojisBWCWYEhBkI2gFVq+lsr1z6U4uddtz95c2q+h71LIumvDn4cWUJ062piUa2Gh4ZNGaU
yzpMKdkd9CX8I66Y8ySURRTDHLtBCAEjjD1IqD6TLHKKXOWcYMKUliaM5jpDVqqQS/vcUQeYRlli
C35RMe/3+G/cw9WBXj1p8LiqjpK54mO05vnzbNM7zVo1kIc9zup2MqoxDN8DiQ8LbYMicOxgm4eg
xDHOtZCzbldyP/xNtppImPDsWyxfxKWaJoFyEKIHOfTDy5/Rr1GNTE3tpdzMcKE1xRsVmvVJv8JL
uDHGE2xC/moh7SG6U6zvBk9EZjJBC0t8sj7/Zoc+c31A4uPYfFBrhS2jNf9Gy68xFr9whpprkqtY
so4Q8aM7ImU9HMYYXTWW9FduA1LKaNJucZ5MuP+jovkoW3lvb99LbGWyezM3iZsg1nR2LwymJAxS
hIwf1Id3j4xLYaACwBozqZY+24XfrWVmJCqxh7qIVTl5vkfOJEf8Bin3qAFOuaxvnVb2r6hGg8PS
OaLOe9dcma0lHRRR8hwKBQ3Kk3bOoCW9iqoQ3LZFf0frq7ln8E6zrwFiXTeICbG6oRhIksGhG7Pn
6ZZqIE7KE490jhUc1ITSm3yAPNTRwo4lqxfGWOKP8lnzMx9LqsRsWDvxQgXtA+2eOftiRlh7kF4/
zv7qh4FHhfIz/IxzEj+TlQIdsxh/BroKrUlNYtCB1DPJAHwKfMTLEM6+tU5/jyUAGD2xL0tETZOT
fwD8QAeYIPwBAjaYNCSzshLX1YbyiqILfMk0FahQbwt64aRkUaW/AgMXL7hIm2OxLwLOMOvwUCiC
OdOzJyUNZvynKNzQ7wI2ly0d1k16xVrqOQHSt0+OtPFk8rL88+gvZ/xNqhf6wXPX+sP0bczleypT
xSQ1OTmWHQi5CGC7NLR7+wWwkqD9r/x5lYiLEH0RU50pxaeHr71nBuvU67sJ7aMrn+7fGr8dFMWS
z9LZkS2jfnJSmOCYBabKLEN+2JXwC+Moex1DePE3IdQv8HJ1iBTV2oMoRw6u5nHySkiBcHFETfS/
nGRyljSRlRjiWZlN4NipRIL0DTiLTMTMWmZQ+YWVaQLness2iOxAqAq0iHMx/q4vDgRnkLzdcFVQ
q7xod2YwOFpJlUoVaZHxrixrsdXIQlPNjhY3p56yRISULf/ZNRDpkcSxnmBDs/rKZUAg0++lAxHm
JCTV9PbFrUDZaJ36EsNuqoqpSJAruaehfDLudXz8HJwCDCDr7yRy9LKBPLsToIVZIncfHlK3yFTy
5SvsEiFLR7MDX+7Emvf3DqCaEVdVQluLXtwzQKtVAH+91rEtpuI8syfLfD1rKenaPN0zY2d2HtLi
O7esj1slb6ktVeGM18y4s7jTIRLPOIYujNUSOQ6GpNYlNb690sc4FEWbJ58Y31cUUs2c1Xx16lA5
jz9hb4Ckekt/D0fUf36VT/frLL88BpjqJkzvFrf0PV+lDMkT+yvTky1ED8OHT0KMOF258qVdaX27
qlRMfzx49DnHHXozv++t6umkcKTMLKGWHghaopJCfdYpDGYNxEN1vNw+kX7JddYt1BH9Z5NyfZ0R
Ci9HYwm9Dx03z0tf87Q0jpLPQ/amw24Z9999P5Z7+/9emsusLFLVxoNCWUar4n4EScAMf0ZXwIV3
YXRjip8+zNEfFn0YMs5IClpwWZFqGEd7HaVzXvDq8jCFSjwvgZQgiSH2RpKC+LuJEuFJTcQawq5V
2W/y6sFAYs7st9IsEtlDCgW4Q32df5FdbACdZwNLG4jYXfY+Vwe2npyRJ6EfqRdSQDkSAxHeB877
E+eU2vEq/u15I55MRyZAIaw/j22ehqhtCX5bJdSdGl2cfDLwLXb6uLdraM+r1FPSKGYDv3pz+0eo
qMGLhZrL9ruFjzbLod6iHhHJ+UD3Ea0NNSZjlI81qMW9Dp+LE1/VaMekSD+OPpAWgFgVkB5DDjK9
bKpW108+rdu9uKhCmhETdCCO46tiMqavFQFrGc1U2kV3AhqyqIhe+B10bQJUuP+uvu14SOYo995J
i91omMUqfb8TkrrpfmAxYl8bVuKYn5PGEDRUhduNOl03Dijp86EdpkuA5NbW2mNqqmv/GDwicunU
iVeQN/EUsxpWcrSxiI1hblOK6vWEl0NH3P6Y0V07WO6KzZ0RR3yet5dWQ7HdgRliZxsBTOTquLOy
AjCM68NL2WHXoPBiD0eI6tNqqGMOHPU7YG/5Xh5ikfVWwKeoYCCFDNybVkjTlb9X9NIFik5y0cif
Nn6GHj9ZN5de/OZjnwC0weRNCT/NGXaz8QmQDSeBFTvy0RJ0plyqc8eoTSLoM+hAq5cRJ/7EtHz2
9DXn3EUi+iWL0E7f2VJMullhKUUDt7wR/GI4YgpVKCk0lABPd5q1EvyS8u+EdpLb+MsT3wVahhgX
nTKcHi9vHHfgO3WTsZVDmvmeDAT35Hcj0cs6CQIfRRdX778MYWVJ4Vfwn6TSB4cHCk76D02XTGlG
h2QahapPNtjDh34DvHxWzwlzvdOJ9lSkYRksNhn7EU3jFcoXq3pHYP3x5NJ2jQhpjC0Xza+WS7z8
Ecze54WisC121DS96l/CMOro49BoPdK06idh3jKkkEVtCXeUfAK9XjEIVtXX790pbpuk795c56g+
snLrTvBmVGfNSfNFeeM/+py6i4LrsVwYtqwLP+8vEDUDadZvjBiOo3XL7k4T9JQFK6l5TYa4xQrL
oBXgbvzRWLSDnj8YFQFyGtszIZ8qBt+zfHJKe/+m4ErmCsYh07wjNGYQJr5AGoBda/mQXMvju4VM
gRMPg4yzq7t9oTbWv0HY41Mqk1D4Kn6fzA0U4WpBSzkKc2nJmoAwDw1SE6D38u9HnZMTxJCrptI1
dtIbwTbvV/8qx0v7a5GEoFVGjDKLKFALK7IEW+Vr6SAM3UPGRD3QbF1yMSAzRBT3RgGZb1qsZGdq
qFHCmADnt2U361A+1eStRRHmQddszBgeXkk1f+psw0erGKqiHeK0IQKRyeLbTPgVK+4VLgotuDo9
DsiViRPIj6t5D4Fr1ejk1RBLOcaQJR13ZqgfG/Wlz32DF3fKy/cima8Jbd8DeZmDFVNXgyZ+ooZt
JMgcI6Ku/+kujAlClV/JDcDQscDVGt4Up6yRZDJzBCxgIvNnkT78ol7ivxs7Il6Gj6MsLBJVhI1c
OpnZZ30noXbgGxPTouAMREwInSPrpwc+I2LGFFBAq6uUI3QhED/SJuZhZQZC/kjE6WYDqay6LxCM
G/+bnCteCGEdOwJCapKn1GDt8wQa+LmItC6zctbbMfhQGGXbsZgiVPq4xpSBYcC714Y4EFbp7ezw
gOuUMkYK/bBAz4aJnT2/MA5wcsYirK4dEoMxW5CyPqJQEShB6teNR63Ubm3pZ1FPE6TqfXC005mh
zsHUH8oYKu0pRyyt6O5KTAnxE2BkqAWVJr/Mh4W0l7uneNS1GZxoCJMppg8nEaCVLV5n9HjwCqvO
smvBDAEsmeRiVB8WRuuv1/HbeXxXHzF21iNI28fVBT0BMObvs6OlF5EsqJY346OeaAepzqz5u+xl
WkVZkil5FG790aagbrFZEjA426u8CEFy/wqD1CdaSQwJ//s+niUjtsFlRM4ksq5uRwCq4F58K6tA
5PU0sHsXlhEwubW9pX8zvoYEeeTZtnOo6z/5HqcG1nDB04KWoKThd5m2OgLrnj2SNhh+8wjXxrdB
Ko3pKy6+Qzp+tFjpV9RZGwB7HQ2LsHnlnp4NYhYwsRSBLeh84OOJXRryoplHlq9ShfSpmxWvITGS
z06MaFR2IvVSCSfRdY0kfcJuAW/FF4KQUcS2rYzpkJgqdJ52b9PET1Wj52blNWEVZkA0ygdZj9YV
IvjgHDVrdQ4FhIt9uSoqfSpjHFivdunloaLDIMlkjSgquibnUJ+kX5Pv2lslotNq5X1tZZUWmXnr
NbEGByXYPVWKkxkzRdiXEBUfvwzE3tNaTBwCsxq2zH+LS04azZ+an3Ss8GyDlqpetrnHwmFWFOs1
FSEMZi+xPLFm+SMyroARn4MYRh4j7VdANqKXpBVFBXLCcD8Tg5TMy7gONiGH1YohWhkC6KPXS+3F
sIIESI63y72zLNTwmKDGlbqexCxqoFin27eohPXblYZF2LjSDw3i90SF0S1hkhuogVYH7VZ4i8hO
U5x7AMgoAwUDrk6uYwqhAgDDsMsAybcQtlwStaUcksWIg2lSFOLHn/0vYPlKWBnYKAgPBnh99uD6
DJNB8+I/ZYB8QM8TdMfRrDbxLVHU8Zx3rYS6jaXJQQfyZPdyJQKqElpKdtUEAAyObMNA53rexkyT
AUFpzVGMjDVylnJIQsXv7dteTSdjn3aI+g28BRl2mJS0cn/JbJbrWY/6zOGbxl0zsObMqd4I3V2y
dZFbTJVvTHjD1Qlm/azO6XxCwuwtlYEhmgzPt/AxuQvraP2pKgINpDriNf+DcjVSDiEOVD8gFEwf
ZVdxPIN3SM3dui+1R+5+f/saYRc+mA/olLZY0DXVXI6Uw5onYjZ0JsiZT8E0vA5+zUePKHKMwZyL
bmW+gtoK/Q/aIwgUjSpmkCLg/wL8UX8I4+8GWxa91DQtSwWkKX0239rZ6AoNTyAhnzLyh0TgxiDm
q9SfHgnpGo2G1sAD7/rNtbTT7YItYsJnnH92kiQ4LaBwjW5mUbnf6tUyGAQGEFzp4cRS9iUkjyXf
2OMAs+eSLN887+fHax9GYtDlimI/hOt6zhaNj346T8SuGo7Qz0cgvOUEF8aXlQDQ/9irthzsPF7z
ronGQAC08x4zsBHemX7ovcCOEQEEGw6FH88+ko9/zXAH9FGN4338E5WEbbkq5m9CdASjnVHNXfAC
0YYfm/OPRVeSEnqsYLjBYgvGvStHr3GzeOx+/PS1tgq0KpFO1tHdiNZaFeuCYe/aTlxN2SNDcGrY
UZlCUb/qqGa3wmuKv1FZOF4aVBI2Di6c0SigTzWsYIEsRtnHkm9moOe3+w7eWp9yWhWcFl/+1FrU
CLbi7p2Vk4G30qSqwD/fkXbiwlERvCVnkglczo7nsXXopLzT+pPqeY6t7incFr2Lhz1JQMbTPKaV
+TKlV97RjZ2rX8RD+XoPhB5XdhL17Xuy9FVdzXMjTPTcaGvb1tvUOqJXKU04hhzhP1WeF2vdhPsu
cseL0aym7PSJN1X57beJNE4abVEeai4hQXqp/Eu7mNBPjGSDPQnau6J1W2HOcPv1S2ZP8s6lRCTY
o9f0HjIpnQ+cOD5MPzZVsqpqwdgk/DTNiHbCXHrSOV87pMDr7BBFNbj56zrTi6l9kPGZoqNMlkcs
+x1l8ueBf1Z53GjeBX14r9GizLo6qXrJnkJWUn2cKEtBwprLDE5Pdgi1cDs/ZSu/VJUA4/MrXrdl
5FK+4W29fIqFcE2SqW4fs263GWJoThc8vYJC+GeWwBfPGWom67oFojlEm4ub/dqokNS7uxl3YJn4
Ax/1HGlc8qaHtEffsegb3n+Zb1LMMTFvGPB38q++lxp1ZrKqwVUPkDpU2NZ5OJinWHNGtvga6EKY
XGfZi05+5kpH/NPpSDrZxDvf5CTxmvBAPQqAVlokCAEGqJ3esi9WJkGkTyQF3y6ZeqXaMamU4zOR
gDGrDRLqI4Nu47CKEHwuqf8GWbU8aamb+3helAWx2C0D2mzcCiu7G60SoWqMJ9AFd20z+3yQXCIT
Mgcs98SfeOzawri11hwSPZ2MafHt2bVDiHc+FHAQ2ZplfbRIt6xA0kPdTDu41uxRb8c9L90R0Mh+
pl2ss+GQ98yr8wmzCv5iu5K/rK67A742Bk9EU51mxG9mIaDw4cnAshut9RAHFKnKOCMUH0lVYsxb
ZVUWbPhWekhX/mcQ4BXNTD1FXLl6uj5lhGu5ialVqonLUKmNWKGx7kczdIU5lO30HgxQDlW7sZm1
AcPZFNQhV8MGru//5FUhgTFh/Dwl0cX3+3l6P6aX8OU0Cw8JB0HqKhfEf038LAGm6BqqKVLGx5AP
1v3ZVlVDD8MEtCzjvnLUOuh7T/3fmN74ODg9CG9xhl4Z+RuuWLAFiB0CEMQ+ghiiKTeDp275MwTL
QTA2TGEpWC7rSDivPqRX/oYXdrwCdXPgjgJl9Fnk9eaHKSl8Y8+23LQWzzy4yptn6csRZ2BzUfw4
kh2Se6UCDwKl3QIOlAQ9rnJd/TzYjRaC/onuliOfn1cjNLG1TY5YhN801aDpor+R8bkDguJhnuA7
Se590CxTrOhV1CliQru5Ezw61S9Fbx+hos6nNLbQNVPLxMlmGaJEjt055mqjRvw1nOSUl5/TtP0m
5x2M14zgCeSQRoOIHphgPJs9dJXlMFLSstKmBJxyFoFRXKZBRb0EqEIhv0bYIrcskTyl0T0WW83z
VxTUUn1g2OJyGzwxyDyUlosKrM+Ovg4So6/T4j3uCrS33NUYxdpTX7HUfX+5g/2jDQcHR+Vn5TSO
Vbut11VyviF/8P9uRbeLoUsejZvsRPNLH4JS28OdTObqyxLF5kg5eG1HjP/yFzs2Blq6U0E3tKHX
yJpog1YF9I1dNPhgGopBZ0AeI9rf0Er32B23nAiODigAqlJSM3pvI0QhJXoecRsBMCRSM3cfNJRE
pePHWYMaZrhb7REDTwcaPin3TQIYWyjfYzvLDKXBWAPbs5Khk70ivL6RvUexQzVfehIXS9hq++/m
Z9zq3nXSwjObufCO3GzlKdLvt8ZRZVXrFaVebrpgn3+0/PTxQ4rNoW0Kh0Pn4e6jWYgRm4mZnbYe
dyUEn8dEfsg2JAPAO5U6+k/vMHWz7m/uvjW8iZOpVLsERebRp60/v7iVHM1eLLH3pSFYt6cmpzws
/mjE+vfBlZ+U2CsXuTaRuYXDlEBtmy3sMC08eS09h4G+3WLcMERxgWferfSu/zOtG1XjlEPnljeB
e3s3LYWNXHc8Rhde6lblaP/C9uRmLmYP0mzjcwzP+G4xyQ9VGHVpO/hUBAUULlanDJapbiQPDlRH
lxervySoJ/O8OIgvin0KEtqILTOudOJLHnrTMd6A7K8VN2oME39YVqzvOdPjtwNJGmfXZ3EVYIhv
+iLEL6Ll1tmDK6l5EyMPOJRKZLoembUgKl4uL5XG4SeCoxugFzETsKfzKDc9bgFiuqyZJUsWLOjw
PgPYcnUVRdapTFUTanvz9KLyDK+OIPx8OCRICGHmX332Ox92p+I5JQm8CEMswXXCs0VEYl9CDaLm
C62Vt0FVoajVr+8XsFPFOeEXvl+k6RTYJJVxv6hjd1+1fOzPe1O3bdysamLASUy4EpvwLrSE9tKb
xioaBZpHRZriaUvCQcIdbbbJwVTkqSHYG0MOghpmFY3mrImJyg6nZrwxo1voyDbhR2cqV7M49cLE
kdKOgnT2+yRvkRDoVJh2jJrxZSOf+L5XHH9sH+AjgjH6jhumVkdbhWVM35BLAtRU75YiiWg9QNM5
GtiiqNw6grsJB42LC4nbnZpvJvZr77vqSE+ceg0Jwjx7c1hyNUUkmU3QbzR1DD9pve1ueJ2AK3zQ
tDK/Zc+4a2ui2VoNKJogWlI0OG3j12TFhmusC4dCLIKxT4EVe3BPnN5Xf8XOqvUa8pP4VBljeQRd
2DGN/xieYYd6BuCxCt/6YGfdph9U8dGDFEJB/YZCV6HWweCaGlybe1LvJjYnNc0FvAIvbXZUM03F
cNRQy4nk4l3dym3WubcpNX0oDAQhY2NpXcVgxT7tvPyEvo1PGdqUTniR+kfpEqSYwkUNDl7qcWG+
1abkauf3MST3SuQCjuL1v4MyvHMpaomvJ3UJotDwRuwB7WQTSbLulGkApVdEW1X1TiHF47piTOfm
B7HOOwzdI2EDpMmd/WZlX4+TGJWkE9rOBIGru4mSHwV7v5O+06DXKAhkarCrYvBuzGTHMMugkjnK
2wESGsTc4qeOpyegN/vzq2cJBGHE1h562pBJJD1Mu57doGZabpriKC/CRka1tlBpLP2rPDKqkOZq
Ky/q/aZOEkGROU5ywztVa7y8ogy5+1+5vo22CXPuwhe6Dv6XjHKqC3GGcGxPx4EL4/Bh13dVUFvP
x8toIjnQyPAwawl28djFFNhRe0bQA1raAuevhJKPWhAJ/rPESiyhoak4j5IVfzYhMbItJRTRE9eh
5YYrOK0yySRh0LlM6wFvuV3JELyAjC9NrJnxuifFb9UJogrr6jhqX9zIuCJ13OQYNz5b4WnezQbb
fRSk0D/mxeCF8qtUupJbner7QBaDP/8T2oXZTgcBHAI+OkzzKcI3LxFuxFjL7Fcm+OqGfp65R4X5
725E1WMxrTBs3iU9PbMqsstcscSR/TNclWSwVgHpBOBa4hHKCWXhekvkM6TOwT58Rud95OTObvV1
DacNv9LynUjmJLIZ75A1eD3NZPGOg6DDCJ6vip80vH+FZyleZOEs4uReSFdd3o0vXiulz7e34baJ
lHDhUirpTXSCh/bsiseANUr5DWB05mtarhK4jM3qAGmsThKcxEOw/wqz7v16ge8wQVoR5aYjoGgZ
q5IRdsLpIsZac/OMxtE2n9J6M9y40aaOGtFwqfe8HR8FwdUYBBma2pt1vgfd/9bb5d74vCTAsBjk
+h+7mNR7mk+Gr8sCqKgBsBmKqcNDyGjqBZNP3RIIZmFxMS3QcCmX1aUqH0ugfmgc+uo4JaWnwEXH
OrAQPGatViQZg8w8wjX/rSusTIeHoL8WgOIrzTAil1bjkH5Oh9YOVUA13aVwKOF2u+uCon7A/wqS
zmWPqhade4/2R0dAxY2XnRA72i8tFghQKIwl1nwRLFR+VbOBbBnjQ3xuCMHyuhratMw3WuvDexId
pvnagS2qgmmdXbe1tZaM/gss8VtCaC5ho3+FZ8X3krw2ZNwa0QN1OlE/C5lfsWSItfYW2bXqasUc
fGQVQSzM41WiH+tg1tQVPTbKljoKjWSozXX9U0OKP5yz2q9+6ud/LLAMFTHG23pdMg3EhrtVucH9
mtSxZBqN4e6GuAwrPaDhKEFJd5s84PXMrkMUcIPJf30ddSl2A7YAl5BwnLjmni1cmP5RiyGnhBSd
kF5yDaFgt2jUBbT+rgvbSRU6KFFthoIWex1TnqxBn98SMF9vPhHLfx8xR//sgN6KXWaxxifBfnSb
f7tE/AOzL0OaamGmIPuAk3FxpeSDgPsvBvWas2LYEoz6FZOe7YPi3DxLjdVpjpQXxsJ032eTYCNX
pd678yOwvNdLZv6T6rNrWqycI5mcm51w7lZRgFAIkEzyBUJDLkAyUl2Y8gHrGJfLAmS68/h/9UVZ
+CS2joDeJovWJD9YScwokyMh8h4QAx/rUfx8NhHir28zzuuZJNVml3nPMJbLUWalpqif3DVhrun3
T43zBJz2+N5bJ4T0S50/Jfuu2z93hcx7vqW4Q2N/BGiTrKbrHT1iqCgcBI+YHkcmG6zJ0U100Cyt
20A6SOtxsWKZ8dmITvWPKcnkL2rjDzNHFvddul7Vu0cH3pP/z+0pQl8iCw91z29XuurFpWgCLZVi
nGu8yVAT3hkDfYx82C7e4QveOWpo1fGbufcYL+If8HTQILD4ESzp6YtzQpU2+0c+lwv+zM3xQsqk
HeYuYxLcVCN00RlYkbUn7QCOH2LEUAU5q88dLBzHYsjcomuzBF5i8+D7K1AfHpWwO0IlgQ/nANPS
Flk8p4aXCbEPCa/PUOXviiLFo2Hcb6e4jOTb+bRUp40OunYW51PXR8mFwrsuQWEzZ6g9LSMd/cZf
M3J1bU+npMbr2hrmj5Oar5TYbErr3VjGN8ew+/P6Vh2lR1VtCzOhXVxNMlFil7ZEQLcLHw8QzP86
zS0vq3F7+QOUh4pJuNUEKZQHeIGhl3O6u1P5Oyiq32XYXfMK+1Fhb274iDG3TmZhD91F1c6PwPam
b87CMJg1UK4JpSFCEb8qVKKOroAnE9h4cG9ZZrDE5GKjzeBjkw9qieIKIekdwsBPmZUqzKrwoVC4
n6P4eJ3O+xwb5AnxbAi37biZZjdccvrq2878j0dsR3yXvZ2W/+j9YAOnvG1LG5Vyq3oP4mVktVV9
hTRjyc9OKyhSNljiyEsqjqDieV2sctvmcUhUaWiHBKXLqy+y9haH37HWYaVbvT/dQHjL7Bb4beNr
zmZJ49KPYI6BA19e9ecdHMLtDaY+Fz1lGuUseB6dwE/NlWqMS9jOkpCYNbAeo6j8o2ruJYwlhTqb
mE9T99Wj+wob/6xpdNbyghNh8qLKlfQUZj8Bzzo+SYtk8d9MB+ki/XQODt8N4lAUeauN1BTqGFAF
CnSeeSmFBLnKhBqBzS87JuPztBjc32iGb2IBj63ei6rVKBJvC/H7LSeKXBsxR5CeMnACeXK9WoWk
9yy2XUd+nGvC9pHZYPseVv+41QhlOVGyVOzlwM336AxFtgmhagUT/MQqgRmXz4/1YuiwmwXd8bb0
1iBeUTlVW4D3rfRumCgroW4MY5OPfBKyvm6wuLGuMICnmBK9/KQAZSD8oh9B4jZdKODDsPoZMfMN
jXQDkacmoWDRSeHkqoAUxcjQpLECobz/lzkD4SAgXXIO0pyHUft8F6wBe7xBB1lZLqsnFARLulW0
mJqbHeA+j19veHRR8Io5g44cEX52FRpus96Bs0KMHabPU6IJMypVCaYkmDP/8Mw0axAcvK8JYftI
Ew/lT6TdovGylQwRKtURUAY0CrTL2QakbJzxPVHOdtl0XUUfsI1VFWcvi95huc3QM3DSpJNeKznY
j5IUyb0r/M3BPHAp1pW3gqsq9g45bMFYu0Yfr3BXtbws271BaXIhlgzeVFj6wUn/RjXT7qX3Q9iw
RWRYmcobuMfqag6s7hEAy4sLeecuuaByy4wzH8SosGV0fbd/RybtU2rCsbvuJ2pd058l6Ugk5Drt
NKy83Tg4udbA6r8hpuJBx1w/L58JcBQ/eozEb3nIya0mhrEGA881TpWdnXXezlXfmP7qqUEedFe1
c9d0aUJrGkjCnd2HKFhfYI54uV0vDnEAxG5UndelzBFS6U94HC4vaK4m4+Pezuo8oS9h7kYB+0S/
uvPowwaYJjZtJs7+8Sh+A+5ihq5Tti9cmZZftoR411IrRWnhrdWjp8ap3wJPB59Me08krzFpdZyW
MSZVLB5fzwOtrTjRLlEFZDNMa9yiX9WW+zHlC0QouiJS6Qzvqv+hepEo/1zIYGDE7LH5n679rpg/
kfJ7smlROkJS9pnSzvgZd3qGYQg9V/O64PEI9lZnZHiUh6ZKNwmjTY1Ju0G3eNI6hjFTusYKrQLx
k0SbUNr4CiyY4CaZw3L6lgStNqWXPdb9Ciwc9zFg3394TS3NkUlASUXQu3PEKfDgXvPNtRTbl9hJ
ndu9abecoIkf7CHRANzyyIuYRnt1RqreFEUP1KMAcB9znK9xPPvz+kOZtuOpBefz1MBihmZ2FrG5
ZZyONgs6YpTF1VV59d8YHOrDqlwV8E7ipNl7INtc8exePSkZ6PSbZ6EoxwmNfGrmXMpHPMpN8a3s
EXJ1MWU/ymOvcV0R3CaknD61zyLIGGpv9yRtTw8pewTMsX6Lp1cLEPS97J58kCZaNgasroJjZVeY
b6z8PTgmtD0trLvCtWnle9nAT1PMb7Xh3ZCNUhOBamDk0EmRHZo7TJf7fVkD6RCql2PafFMMONIH
oONm0eRvnWl19AUyauvlbQEzhyrJzF5B2OL5dQHehXHG5NsVcdJoTcII8D9g9S9C5smB8+RFD2xC
210CHC86R6Iz+N5Is88QDmFgVLAXu1tb+PE2KvQwbq1MhCWAGXG8a82Lk6fiTGY+nZi5rVs+Nqnn
geuaRSDHX4YuDb+tNBKyBDWajzE5UOuH6AKirMSxZPgKTxI8kDnY0EWJX0L3AuOLjTWWlWvsbJtI
kkXfXpbU77tDgI4+cQ8gvBgwRFFQmla9mXBRU0ZZZfTerEbjnPUxRaUUDiri8t1iE+zZsbNdUyzP
s7jylSTHh0oVhjTHYjgYz9tWaHH6+QqH/bwez4MxQafKTqPtgEj3jmzskEU97N5Zh8i66n4DLQiw
Q/MhMuSZmZT9aqbUrGoCAU+vSxyAdTfYPe8kY6BDxPcsKNtC7lRwO5xb5l9isvhuOX2GiJ0P7HdJ
2pDc7vmwrmV7YR9taoZ0ZWo+cJatJP3skO34TWManNkmhuLH9KXWk9GdR76n3hfVLG7TehtmSS1c
F9lHoT014+sZzlI5SsT4EXDwC2G/v5sbrNq2ilTQLtKQ0kBNJGpFp2rVpYOMRdHMmq81jtMLVa/I
qgPNVc6biFJEpzsGX7LMCHkxmHDwy/rf740KUTQ3Jbi0WIZKIKkb/QPeGXmLyQsJ+bqahzK3/lWn
pBOZHYkzQGavzq4y60OtTFreeoydPO7vcmqL9Xru4QLDyKwI4v9ui/QJvS71Pj6xqEqeppipfqXG
9MUdrZMfs/lW1g9j34fc+ISAnQ+hN7mbf3dzwWdVurybL9NkjwlN/Q2F0X0C4CsnS5izhKSaU97x
l8RjXBOcR6X9JtSsPuQhKWv7K4QOa57sR1YqlH+HRu24E3MwKoC8tPwTF90iTrAk2gsqq5riTFP8
6GmjfQzCq7reu2+UM4Z6qm4jqWcm9rUPoIF0zECRXL3gw6j2MEIesUpJY0C4j9IZWCSh7L7Fcjw2
FYy2WlywQHkajQoUxpZcq0kdvMQ4HIPRkCmK4jL8qDUul9312lKNjc/AiVhdhu1jWfzcYcZnl+yG
usRroPXu58SSZjj09PtqSLSsn9T48wKwctTcK3kr6SWdlvlLZ3MLDu6a8ewkwTeXa92Ax7uvU4DC
lDT/iRpYQRJDf6t+Ue+S4NxM+7ReyO3wrxmh2stozps2myhM26MvMwdVtVHbUyvIXpLxetbTu2oT
t1pkb1QY4WKvsByr4ggNkLIV8HDTPe0s9sfOp3rHWAPfm2AXAatwzQzVYsXed/my87RlfLursavn
tBiXXZcxjIDzPWQyWvnAbUDmbz6XUrdz/ZVAr/k17j0T+4uvMkXWBKDN9RMlQrGkQmrSTqsO7YMA
vKXCoMvbCB1w0NYwKGa6eE+T1gT7yWK1wzRfPhGOatLx4uKQecMr62h7Opse6wAyJ272XX/1mqKK
PhEbzVqQ+c1iH/SSl1xT5WI1lv9Hwi4lJcmprScAXn9WkWiQEhFn86I4D7RQLJdtg8zmT91Rvt0T
lTSp9GGTzZDku9ZVr3nlcZ0l2wlct1mej5/bazky6tYFVyLQyLRTswxyqtKyoFI5iffVa1h1X76i
oSP0YFVSXMPnfoj6iMXA+5ec5T48+bkQ2nzbbERzk9JhZMw59z2RT0M7h+bB12/9PUTrkoIK9VxE
7dNko0ZNYlzvguM7wfjvDHkxXTVPfP73ozED4XBfJkX46Rq3oscMU90IbclnzU/mfRcSDUiMwp+s
5PiIbpL8Ko7lS0vBk13eU4AKuDJd44aNbVG81h0hZWm752Z1rf6I6+SgMrpGH9MBpkUyPqdZGeWA
bje9QlbMXigH0Q/Nyj+X6Lt6CYKL9Iq+8FRjLHnYp1sC0GWJJS53O462v8pbFot/OQMewCpand0j
LI0hflR0jOpSchaiIAeunYj2KtqabhkGwU7sGltPq2BA0Nk56MrNa4UrAGQzEZTNhu1noJrcEPDt
SLNqIBfkMS0MuzxMHP/ZLf9K5NVCtuwXyN7Us/KPs9DBzKu/TIudcvTGh5BXNjrqio4ty6E31sT4
eq4Ul82tQSMHfl2rZzDknepzcZIDf6LmTgoJ7SHYVX31EODaGrumU4ED00qsEA1sQ6vpVxQeOUOa
K0ohEBDXeumjwDABjJsJg+s+bGNlw5k/mFx5VmIQZgiX4RlOuYkaUmZpWHuD+NcZnFjQGfyFNIhb
kk5RX/fVnSVVC/UM/fOUlbXBUhXv4Nv8HWLgLOxNxmUOaPcF0s9A5CZCEZJg3i9nEZbns5sumjww
lJFS1GHtn6BGgPr883j/gS0MkaTkoYDkvacobULT45dj/8m4pksb6qPFvztQgJ+0terkNwlKq87Y
fQoDKYsZNkfSx6WK2j/8Lb8UkclUnngpZ0t+SpoP0bfT3dGFUSKukbNir4H/jjVyBnPPvhuP1ZCd
fruAQmuLOTOsUz8fsVLWIlHT+P1/QsC0rDn0Ke2k5HLvhV6dPEKPNhngG4gZBx7h60EjgeNPN54t
A3ho4UCz/ywcd3dvKHsE28V3NjuJfympC8iHdxYZuPTh2Nb+Ggg5LqKMbwasKSUTEZ9tJa4CwkPg
fx23seWHYxm1/ChoPlVLYSgl6Uqziku7lEbEfzsXEiThXCAIHjjT3h5UNu+v9/HByn9gMYTrhsHi
Rt5bxRNbpgOFqyDJuz/tbgicIFlgPSR5j+368wZiDAmMs/wvc+DkOfT8tJMcLpr1mvR/EzXnHwty
Qwi0p6kIbGjDQcqgRZFijqwM77lPPCMGhSWHx0cyg5R367vlRWGmn3uREo5nOqAw8lFMOYoCbnYn
YXJOrPzFVGFQgVM1+GaCEs5FjQEMzGADukAijpIYCIOzPkIErQaK3jdEzE7dLdcFnKX2dFNFz5hh
H2PcICO7ZFxFdMzAsmxxjytqHHD5ZbZ2cRr6W5qqhzPUUVJakMMXbFZ7crFfnllBra8FXROwirus
WXtiC2dgVWgmpXFohh21l8npSHS0HuyATni85Z9sNIvaLndfc+YgVhcN2s80FVB2xft9u/JUw/9f
YfV1udyp4JH1NO2oBLrCyV6Stk9vwyCQRklZQWLfs4NnKtLPRRNCLIZyOTxp77lG9CMD9vVid3/B
d3IWGD1IVWO/gbuXRMJkQSdESjm812Cn8ymrE+DT5mqWLmXDCmB6qnp1YQ+bz21JFtghq1gLND2V
SYRHJz8dJBEVBwLJzxMmFwsHclSHvCeC1+f0IbYcYzuqWmL9hcVha9e92hqLUbbGxlAMUCAODBjG
1Bk40HWyda2vL3sDxxs855t1UpxUSO84NYGweO44B2D+snSsOa9ClJ7VE+r8T8XTgrUYEc1DKuY6
aDP18OT/26meqJ2uIGC7+6+nwe/alJ67KHRilS4mPpGIpgXujSt7ZY0FlGmPQBY5J4YdlAJERX5q
LbGgHQ4HTdhS6kQji531sEsDoM/pwdBws9ks7/KGHVrfq7uNr7KJLqLcXRtde4SKw6Jj1EDBhI0U
uyYGkjxRf/TYpZdNFwvnjCFVmcmKGBYnlDlj9hUUltmo1/ZBr97G6fF5jObH6J7G6M63Nac7bQzj
iwQ74D6PbwKVid0/bc4lyT9tjb6woASHz9yEb+yglF//F6ab0EijDfECpTnu4obtN7n7ZmdOyst7
zMwFnED5NCSWogCvTsZYygSAtG2z22/5VJBoHBCrxGLFi5HglU24mN9Zlost7OGGAnF/JJMt0myK
+wjL+XUl09kBTMAtwOUqKByqhjU/cvLTS1h9r1aCgVCFOpGRb/tiJy8MY9MZhY9+UUiC7+oJanXt
vjTagFv73SRroqpe/TQq8NaRe37MGB+KEQXzRWc1wLw+byhXeUDMifQd6L7+dWKStVhZj8U3BN35
cGE/bCIpSSJnHG+PYlfK7CNG6d+iGyYGRqZtNvN3ezxivTRg3N7+Nf4A0qx3xreZT/rgKpudHLB7
9gL8YCURqKL7BxhiTESx0Cx9nJewpuDJRA6muqFSDDDMH8dv0CaV6n21VhzNO3PI9D9Gd5KlUbOw
+jM2r5artpnCkZOfu1Txwq27im3hcs0VNDajzzSA2d+X+HKcku3Mb4lMpfUZoyMfSYLWH9isX57P
W2CVFPlcS2q+Aiuqgge301VOZWFDBZnrMRV7zb1z26kFMUwkPd/JUzELmap8CHvWPUV1QOjAtn1T
j9wMxiipvoXQLktURZQSdJO9v4cATck7jgV4TDokVhYCfEuM/clfocJhnZFzMBD08eGgbDX9OMG8
E5A7sJBVPbc2RNRKSpZC9ZV7x551JsmTaZrFahh40UCm0ptcVceZlzVZFKonCluBkn5FFnCARdYZ
ShcVj6UeolssC7vz5hPk6SEArEvKIPSzcz7oyh5tq6oX9c0etW3od0DIkQxTY/wbYVsY1GSFjTlu
ICFC9i1UxI7URNTDN06sEoO4qgYDIS9JYZl9NSX1h5mmCKttdHTbmbLuGBFjD/XeUNKepgyapJFO
9Lxu2DNo75NQyeSrao/VOiIJZpVkGV8l1wWPHLBh9ywG/jzbyYO+LE9OaTwgHA704UcxoJALCVNJ
o0NE+0H+F7TPe4atobTYXJCNnTnDjQBdVlbvKOCT+Scue1UFpR7PZOL12mJGvbPFp/QrzfXdczI6
PeLtyz8E64WddJiruCZlkwCnUlr2/cY9JEKPgSs+f0HB3azPV/NahKTXnCkUWdUjHWOvfgHy2fb7
P8n8j4tBizzkUiUMslU2z9Ul4ri6l4BCl9CRv5pqZUpzgWhfLTmvSMjy/GHfSqAt6RCev5Xmwm1E
jxEh0v/UjRnzHV8/vet1V1rsoSFcyTdcNTvdiwOZJ4M9b1Htt8VpEb124WD5LW19w33/oZRKFnda
Czl2aUgvGS8hZLS7vaLmvuekAOf3sS62MQE5sKKgm/QBhRFDrR5GoBGbcue2Ri3QgiY+Ach1+tHj
m1BokheftGBvApWQZx1yzb3IfDeww1fsgkQqtpshGnYh9KiHGG+wIki2/4M483cBGTEIFqoSZI43
H0lCbXLR2CDX2wsGhct3DL5YieLGkC2igYsNHKbISuV/X0r5aJmxDlTOOrov/D1xBs+6CqJv9Xsm
m0KiaSqjEplNS0VZtrE3FtznHB5tUFGAEwfGCH1lTriwNwb1+M6rGK2+b8z+nTRK6KBLlhovaEDP
4Fo3ry6gguJwY40K/fxWret/YKdpmuBAsEPzRaWmkHPYcjGxNCjh6II1iXWhhkthaAE4WwGBC+vS
Bc5UDTE/yCVJCgfnmu0SnyTz4KnD6g4MW5PdooD1XOPD5VbDDGLvBoULydzSrbDlwFE7gjHfNfaz
w1P+NDTBkrG7BRXGhHNR4ih8Lq+dV0+yY0s2JmNnjTZMmQd7ZOIzZKphOF5rQ3Ql6EwbFSJfJQmL
QJe4Yc8nWVD9MOJkpKcTkYQu+dEI/zXQAzyselS5SvBPWtIb0Kc9IiWniy5fXUXsuyjjYcLOepGU
Q/m6tjUkaBs6SlqhoYEmXSFZnyHfmHesC1EhaEdVy3xx9zhzxFf6GsMH1aHDybS0vomFENW4CPhf
QpQY6KavhwT4gIjRnpjlz7fAgWkHPPbgPwE92Q3flyNoBJ936zpyE9CJUfh+/sPz5bfxE6c38cHt
5psd84koMKMyMiM6C1uClmBLBHxJUjHXDmvkzKYISXT/Zjp5vF2rXiJiqtfnz7KTfImwrwJfHWnh
tPdoz2XVG9Myf07jUHBp51Jme0BVv8JG7izdT9zM0x9Y1jHjK717/OClY7+2LywAfSJrFzeVptmw
J16TJk1Hx8qEqFbr9j+jWStM/ykKa+nXfU9gfx++PkLyEIlsEjV9QkQ0EvhdFW8Lm1JpbjDqxFlx
c/v0iYl03nSEkT1jaItQ3MA5WE0I9dhV2DmYTgBLATQ3T5AgVSHIxkJ39QMrIF8TmVoZ3V46DU7+
EV3aW5pqnQ06Bpv1IXVrKMBgW3hMPSmVoB+CRBjWpZtSiuzPKn+6qunOHeo3/f13fnhJnaHFt/h/
XZDXxqlb8Nd4BekbFxtdYblZg+KOHXA/WuWpc4Ln7Zo2TEc5nisIYSeDtthmwC6BDhzM09/eGGDD
/2ZaDs4IXqFVqnHwqKBrux5Hy/FR25Dh86yn78mtAYvtVbSEoMZCLu6tglo5+ARmnNbAbwWIqkqe
EpUHjDoQ6NTPaVTMP0AwFYlFWXGYWzvf0HHJhLhjgCsRP1aKojwx3E84SI8iGzgRfzfdJeVxkmko
AlM2UORB2SiKUKQ/3hOumsZguTxHUIXVzVtAewDfhin6FgpbjPG1NTX93sO7IB9dFS9MyleIp4j8
r4M1y9Gh1ZbCj1tBDO3pM1LRh0FIhISQP3to/aU+x8SIivH/iOkiXOZB7755D0mv7DexrnpPG+9o
5iSiFJCV0p4YW3TwOzDSjVYDDM0NJc1AxJ0qEh33AEmusqhk3J/eCRYTYKUys3ittxBbjGPdu9Ah
NKdY246XykNOOhxcWX0MQIQZ4fNS8jRZ54sbHi8q1Kmg7VnVYw42uds/4WLH7dy1DuL8QVgaTZU7
5MpIOV2I7nykcJFlCnpulCCVMr9bs93uxJu01bSjwDimo1ZNymxp1QjLMCujBBTp5eCA7wewr1Qv
1kPRqShNFJHSz+4nDtSCVwiKPmAsrv9rPE2aN+yQgZk71N7/nJ55wkbJJXMplWANcAdf4aMpZmG5
oUDEHqclSdP4u8rSiGmSm9TXre2p1LTqR9SFwko4zdPXWjE5GIqu5uGgxi/yuJNvRQ71gLIdYzxC
f4NdA5X3ADC1RU0rrFcJq+rAciMJWiX2zlGWD9jmAwC8BuJIQKypnICMSUsy9jC0cfEHlR+Hv2e4
dHWnJEugWlpPe+Y7o565yHOsrWwGqbld7H4s4U7MDfQvQjikZFaS7oSGg3sy/McEY5qoX0TbrTLT
eUTz/QN+JxSGcElD3wpCzXCwXkFEtPYAxF7q7e7e5BnWV+kzIpWQQjW5rXTi/ggd9MNXg95gMz5O
RHS7PQVv2unpTN5VLSsnOhLJKPAkC45W4pcG0kX58BAIjWuX2VWI+2OaECknyw5IjdSIhy1UQMDB
a96NGB6pdWwWihMSarWS+zJO+f/C46oKhI6iqzdohxcwOris1polENR3DU0NmDTABwki0WfB/C5m
D8KSkWRZBFas66+PR+qEkAR1m3XJo3OCgXJ1nE3tlg1lcpkkipRPogvir4raQ70HiYr4spI0QA/6
gTY030nrU0Yqx0tby4cPH/bzoiBVUnd2T2VHlCml/Oi2BZ1deIoKJLqSiZMov8HlBVCS7k0ITOzV
oGCxRLzGgnhQ+10nZUBHr2bUCQJwR2Sow5GYR6w4uBC7/nMoWDXstGOt824bjMX9zi/1Z+Ammhpy
4jVnC53Uf33TDJpIH2clJWthyexVA8geCQccw4kVy8ycCU4lbFeuB0X5y9KAa/CTP+oagf+8Z4qO
DwrVZBJHOABcyniIPhi+/fNGmAXqxaGzJWppuweEpTNTTe4YReT3OsvKFQrPxgFjFD5C/xr92lfQ
X8m/dsJXlg96hip4ArI/MdTkeWJbjd2fZLIzOaFJVfgXhKLqvyfWiIeTMLlbOMD/nNjYXnLHbKeE
Py87TLCg4wA1bu+QHTD2nEgUyyCkHWJnq6WuGVlD9+jh2fctHFeS/voxHfcmj7IkIHtZXrdq9rrE
LSz83VuSFpqfFekeJv2eKEbPdrKmq2SZRb3n5f1gM+tujRFuUZIbGObWf7qHnp/YBY/X7wc6nfOD
mvXMgHyDETRBQ9HH1fejC+89E1YEx+Llj1p3bZj+JES1IqBPqV97xUtSpACiRz0s/oknmIle5PqM
lOB1tFqb1uiNTa0egIT87rO4vfO4VGuaYqL8BQAb8iCjmm827S8sU26SFYTCiS32CHnt1l2UcY+l
0alqbdvCJ3F2pFJZ2LuU0bOKRlfxjAqejs7GzG6hMJf7ZpneZge0WStAVJKUCh0Gwul55Mvb+SEE
xdBEypGXjpJc4qjylTI02DzhsKNAEppo+Z7UIS7jV/HHXjqML1nl7xE80oNZe56Wwjie2uJmGkp9
ZKfSqDyGHEKroT0c5gTLZgRObgCbMpYn7Rho9l+xc3e/l6zJrL9Fu1JYKujYzaxBgcISU9KVOmUh
Rd+4Wdc++HiVetOuiuMs31IfgUZlYdtmZKi4oWG44EN2398G7d5wAO0mpBB6Hxs8O0UUL7VBmWCW
9fYq3bBCDuTQwhPbl4/JUEazN86SyYjsCfyGvXkwig2THPf3EtK7qK5J50TBC5Gyx5cdKORYKm0T
Rrz8jCIuqb09PbryK6XLvHY7bktwYxwxsvq53p5Rz4evRAlQAZGGv9CnkiiV8KR+YMMZcWHlWpsJ
a7b8ZQJYfrGyLtioW47UqPUjozG2OUclPSAOoL39WGh97IxDFV7kKmfcqN1VfHkxzW0SOSuuHq8O
oUx1eYdVxv9XzRC2nIzSpxqyg1wjG8gZiktDYnlA3xpxbj0pXPeEi9luAZ/1M9DsUcm8OIWm/Z5m
KuqGtKqOI9yz09EjzwIaaqV7YW2GgM0JEcDhZ43K8HL4QSQworbx2AQxJiKseRee18iBjhmQT20w
KDrAbnTqWI7GBCrIW10uJbAbykUNSwMZUdxGZ4tyWkoRVRu+rPTtp7h1TbyNIGpCOMKWgiqFRRVP
txaCXIDiWoVGdL8TzxcrrKToozrgQCNDj5TiCT44KC7UuXm92fgn+bEN1vV5mdbC+nwRlYB4D+zb
46Md89Eg9eSRjTkScE3W+aSt1+jMVki3PsIbhfuipWjKUqc+ARRrBk53xEcp02uonrJ5Mjij3cGv
O3yqIaRj4RUZ8IAOEol33MY6jo766s4kjnxVfn5P+yUICxiVFELggbxTNAFLYFM6/klZW6hUqwCo
0bLDxwRSZySPgTjmK6zSQQSeXhk1gt9RJYBJxrzSTUQyud1yBqZkFDz7CzFelHOOdTFjuzyFLKja
EJhD9ynoJCjqbvqKJvZqxssyAJlwvZy7277XuJcfJ0vRBzbPraC/zO7zSrA920quz0yr7hGCT9mr
qBtU8GUrhAGMmdDan7DGyFckhzzJ7/25OtkMUjKnW3gZx5y8lhZGCQCXllKJF3fYH3Y9XqHaI/5a
IdoloGt6ZWJLXRyxUo6y55pFvVKD/fYDvnb85y6fp0Z4ltjh/s1Qf3IrvZyRVoAOuk4qqIkPocc2
lnQoqdUM+bFkpX6bX6nZW1BfZzOa7glBwnKCzlUfKTXnR4K25jXPvi0yXKIoicTs7zoqR0Hm9eWN
oxONzvYSyOHTk2fODbxceGDr5Fom750wtBuEJWoZdsaBdW10vvlKqNJD7t93KNWiHOpmY4GUmPGH
jOesiLhv1euUtT4fLTW/jV6u13XZn+p4cZupS2KPJ9pPPZUkHHYsnpNHkbnsIbrsjnSYMTDdBAx5
9AgwYfzVCewvI/bfy84zc5XDmAqEOEkkVPR2r85sk4FvkIgGfARTrdtxwUdDK44oRG5zg6K3gy1E
eMi+gKadxwK5W27zNVKLtrQVwziM0D9kEbNn0krSI9LcF53FOdwDrLZUhgyTUO3vjFbTEopomUqZ
5u0HDT4Cr1GTYx0g2Z4g0LLDypor4heYGFJ+GDtHaQqbu0z9o7iib2aO+g5rRXdX022LvvLGara/
jyW0EZYOwCw9aFm9Zb2NMalRhe3NKRJ9YyZszbR0OqZ9eUbyJf1IVRerqTJe0itjYcSkg8hV89fw
U9WlC3x3MmnG3qoqdhArfhYuAPVpOERFwBD+3bFwAeyqycZ8e6MJIivSdT8yqmrIxCBiYx8SQJYN
urmudFzkoO6C1Zk5UsbBKEgX03Dzj213rFiHyiKaEfGRbHvs9IsxRGsVmXXoC2PJvEx0aeUom+2m
rTgzJMZgGJvyfTKC4V0o0FTns5cbEg7azomhV4afo6LkQkEpTsyb/hMQ1eAqqCCX5MXD10334ols
3VYWbDnzPp9h1urkx9Rz3uSADoz/Rqo0vdP1QbdBqFERaW7bJ0YBjSjdXaW4BtpvMG3QuUtSBXN0
1EBb8a2Do3LWEDb0Q9BVWI+MXUzszbEAIkw2U8Bx2dqtqJOVMlhRFACJvld1OFy2q/5cy7yK1GP+
feYWyMkV2AzOUmJIOfmngVqrgehkColRTGX1MLkSBIZGCKQ4xoknexeEYPvlT6Fm6OnF4hksZSNC
crpzCyY3Xt4kmB3vkN3gUAl66H5L2j6jQXnMp5LLUvm62Kze+B4PN1W1BTjGSgyJcyLNRbouvZJK
q5i+/HgnIagZX2UzKaGuq24uy76Mg8VYcjql0hyOT8GAk4PQ2Ex/XwOsWd4nhZH1Qt+/T8SuQuVt
/Ge7Fm/K5Umc0vIebz0cZsIefncjqM/wrHDOC0NRLuatWV64pFo91CjPB7xtYDNh8sJ1UWAjTAeO
Vp5c2CicRKGWHq6Ft2X2jaBxGFkqTOnOPNYgnDxmpdX3n5XMi3ldSWUd/rwk9GfdU+aFGPVg+RQw
P8At4L8IPV1i+RYWLeSCB5/g7z8v1lllsNwa76PrxEjBOZR/CjKE/Kl2Q/NK8wWS8rx3D38ktqzS
TYkhfuVHxe0pwSEoU/R09HGZjY2zIj6vMB5w5ZrH66riDHjNVEun472yvVjFEMmSTvr4fyVF117l
9MU8/KnruGuF7xVhoqg5aBQaToeyy+OfC2RvTAnuQCfskfSfSC8h841g+Q4sQPvtcoc8BFSVc7i+
5WINlZCYHpYgPzni38+ChWrFemJ81oxiTKDMGDxiSWvYzGZPkyOrOoQR9xxewFJFwqDeLNjgUGST
BVwys3k5rjeQo7vLJ9Uce+T+qPGW9fKIC68UwLZEQk8D6Fz225XFvJ/5/I/7y1J8wdwz0dWOxlkg
CK1uy9WytrygSPDumnNzk+3CrAf5P1REuaBfT5s1enJI8aNyQbY5VRcxZWN9l6g9PJKs8o4PYcUM
J5RwJ1wlpPG7/1fAdezXNCR/s6e2/SUNzyuZ/1ajaFIEkDwQId2kacE7rsr2Erj3RKLnV3rrBWTw
y3GrSEJgVa6o+tL39N6CKcRljwU2UuLzKdBRTzV1Hd0R7zrBu1A7drMCYCSwZ/b2YlAxSkHnk7uo
1ej/alYPL/ig1WLSn8stpaXHmpphV6VQXyMVO7UJGV+gfV6ummjK9P1AElFh2q1PSMLfE82988ml
sT0K8zhWN7VtlduCkR7coY/j4hW7yEOY6SxRIvzntUYIJIqMh11O/LoZ4CVKYdt5w7tTDz1QLvTj
3nWUEsXpLBHAP4lUl9X/bf7yj4H+FXXyZhJ9+jKo4At+fFCLlilnGafXmjHShcid2+7sdYnJ6iNV
yW0PFXSeRSoum6IFI3LFHHfo2Hcv9Yh8vnTYLwj8I4O0wzoOOAcLZvxUuvU945I+0K9Wvr/405rS
WfSaOghfkJhWBLeED5vR+p053AYeRFxsjkeHiR2NamMJOoXGtdQPLpzIEnNvS0GJCAs/ih6DhDvd
Q89RPaGC380GetYMFJdQiHzjFoD/SrpJCONZcuSPG0px0csZq3l0B1wS9XU30vS+Py99pZnL+SDp
pNO6u0U92e6hpkL45PJdETPTO9ZFskTd3dgM83c6PyeR+sU7NH8HsjJtLZKbWRhBsm5y5nnFjVzH
uZwRdKzkUC8K1z3CKYoFUr2R8q/GFru+UYupUULa3cYhsL3MPL1ue1DSAhhm6cXnmIToaO5ZFfDj
NGlucQKQg0EMqqar3dq4kaxwTBNjSsKph/a5q3KbmKOdMHH/L2VHvyWoJiYxqlA2Bi5tqWyS8Fi2
boSBt3f11C3lp7FjgPgiPZk1qInIq09u6CAHZrhYOQu5mXRhQGLjlg5o163Da1aclecSuRF6Xjy1
vISZQ2gAi89WKrRFMtRwkB7dg+yojKJXyyf0VPjnZ5H/TeZDU1zsbAb8wf9P87fg6M7K1gAXsmLs
46rzu3FUe1KaJC0A03jxjPBc2FIvXHFpmP52+/q6tTflmGZCbIrgrp92I5yg02brRYsllBD0dxR6
nh5iN3dK3HlElBc5Vm0UwPYkWmI76VihTODiP9FHroa41u+wsK66KoChDa7SmBsC/koG3XFtzfcU
7LPIeClFHF7G7BEebamY4TZnKd/pvuojo0NW9AS5qTcSWzAnVip3Xit785nXDbyVb1p+oIm54pqg
xeDmwW8sK2zR3J6LLOXRteY+FSmrJPKdDABSFHvV94Q8b2zrLJc/ydQi2isnH0GUh06jOT6Gw1Oz
e5Hfm24NZErkazLdCID9fJl2aYDd1KY3KMNSz0l4aymi8yQiEEuJo16Yo7mut7iIa2n6v/Adihen
pbEinEetgVFIvAmDDECB0FcJwf93/TrssMVkJRJslnbagFKSTcFH81LgTracefa9/I5VGJolThqc
Xzzi8DPw+IvF8Z0hQ+6LKu3hvBONwfybxo7IF9lmY9bgJ8vtjjrI+Q69r9LRBy6LatZBpYO8v46P
SSHDADRXg6uKYgryPq0eB3xZjDPXEkIL+aEU6wa2lW4mvayIt5W2UNYU9hZWmH+J33THH6YBo9oq
W0WzywhUdnQDR8C3MprlUAM4L5NoTZA5wBHPIW5McY8PWBw5njWVTHSK/tRcyk643wZ61S2zAmte
GsAOWcVGP9AgDx185NYU14xh6V3Ih0vFh0kkF9jM6nAkzQmxydmXvlguA8SMa7m7CE4P6sUtLapJ
OzDZiazI44/3e9rKQGHvutacqfe/FGwRLjQTWrJLnvVRJazbifkQzy5DA9klmxBNVHdGyXxyAqur
XEI3FLuJNutEvYb+J73nhejjfJSP/1slfBrhiHNd5P2bZvnj9cNWLxu5TYfvLBuaus9eVlvg1wyf
d3KZjEPLjHaXOhoqsxZIaczC0YOLWrjLDwwH6VBFKg9AIk1/b24z8puaIHh3dMmI5T70vRpP+iq5
3hJJaGMoEPO8+9VmG54GVzBAeU/+m29PFHNaVzWaThD5/oeu50hOBWxOLUYAGwMkdv+8/kda7h+C
ek1AtkqBMIC2dKizy1s4TRl9fy754I3qe8VkxPJY9H4yLFeXdKn39wVztcMmtQ0DIS+adH9oCrhB
lwAnhwIonQe7ksrnRoQtFj0xlVLcgxsIHelPt/wDVDLDpsWMu/TLwaP0Va5IEDUcMLEDIlK2nSV2
J9uTmYuQo81hm/o+5UUizB88V+lWmYG5CFUbWfXoxB/UnsHeqEvw+QEceg8bSeNG7EcJoVt98oWI
Xq4gFOOTsNKpioLsE38W3aEfZfHtEdYmtcCMiTqT5yePH2eDeo5toLClkeEdFDU2vvoi7ovJw6zV
neGUc11cjtX/KMnsF3UHUtmAOW2NYLCZ2ZgesQxuN6oN1bqVmONCu5Qe9ZO12hxQn2FVQzstfAfT
0Gl0eA3g90XO4uBzJBmjqRRz8GTFxYay/fxU7j3cptu+WRdG19AyIXXJOw3B6xp5BUOiJneI2sYl
YEmqcF0kHXyP5qUADGz1/QVmHERsu/1EvIdGXINr/E4b3PKuvqhQVvpn0PMuusVXQUbhrSpwI87P
izGK5lafHYW6OQEBtHv+A1vRyoFwygRqIVnZHx17icU7h5vLTqWlrdzzPKAc9HQW7IcOqWS5IrMU
+qeF73aLGd021DYvBjk3lqThgOBDcKzIOJo1vToIOtJzctYB+L63dy+6vG2oL4NkzA42PwPEiPiR
vJFqnPAhoYBPgdnGhLwmG4b49idCaHtimDcHOmJGEo4O9iaLjuXDC4FSoqSYbVWUFO1IfAnoIpiT
eLycOl3BEDVEFl5dhq39+Lyf+A6B/n5JioAW4Pd0ia+Esucg7P9qA+pBrIDHi7x68vj+34me0VjC
A4gh5jPhPJevxoDRLVn1YGC1JV3tUkfJmynvl4/L127UUawKo71m3si9DiMT0a6C3DiqVmGXOBpC
Wwn1uPqZlNnoN1Cvn3zebbf5rsuxKDaQQacvHA9reVwhaE4GxRm/P18EYG+U1oCMmN5tdCo9szNF
ZWVcvXRvBhb5TDn5sD4rYVt6LNlF5/HTJC/pDdkSOhBuOLx7X9Pyxp7NH5nKrMtXC/VsaTA2UeiQ
LJTAwCfqLGJ4u+wG7rnd9E8vxMsy3APFxWHMevulEAZ24QvRc/kWTXNnmvgvj40PpPY2VYPIk5Om
mix015D5hk0qCp8LDT/b+XPSRiZO9QSInZQVoCHRMjNu5moaFja4E0l0EfhrnE7k9I7CXZM/YtjF
/bfW5v3tLz3gHeL/oJP13F0qqnJMJHM14aawSYzDXlVxgVBcuyt5QKPgWpacrnzUSzOzgzAxD+4l
auCQjiXvIcgvtDfXdlddQrbbLym/22if+04fhuntfBjQephFxPTi/wwX7gk4+rB085OJ1DVtsUXA
jbow/VfVuYGWavOPotkCJUgFkCMkBA7ybsmAhpXsVZRh+87VvbK7TebrOD/dpuwqt/3gAEWsRdgV
K/2oex7mWBiwCH/VxJdsL7CpoNzxXTzIdFSYGemzY0PGbNl+OEnhhCUKdhwXCpWJix/UrIMl5Yxm
Eh7JB32OI+LHj42Q9iPGZVkA6LhVyUUGx1tYrKxVcY1y0PODZX6ctTwdh1xVM/OUOyFTzLECRD5V
xXvE1rO4vyr4wILDVu7YDlCHo3erXKIOaNtPtbJYT8D9O1de1Ti5BhSEtnjKG+FZbyaqC2wEtdfF
P3a7P/yxZbP1z6EJOzgivmj6UUFuNO9qR2u5JugzOupH3tD0W11AzBeOCcD9eIUrG7RURsP85uAQ
nJG7aSsYdCOsgpRoB/bBPa/KmJG6mAf83eDOMGmZJgOzNP1bkbEUDCLJmzMtdpA+GbEoKt9BrbJz
5o0TTMnP3D7HzN1FI1BEtjm38kCYEhYMyrJY97CX5PeMsrS0kDoI4H1VjlyDCglBFIz5Y8zn5FdH
veVnCW3Hpq5CnTjc9PaXAp4Xy9O2q4tk26A+C9jUSUnicZcjkDnkvGavJnJrdqjqrLv4PFYFrjEO
WT/dbL37vNmLasEJbgBMKB0oBV8g0cNlhI0S7OsPlIK07OFBmbzpXdIXQvHFY5y/tMqcdTSG5ljw
pqNzfVSMYFCGqSaydbp4QF/8Mb6IUn8uQr1lbhdKoG+f17xPWRmMi9pWCH6lUxuvGFmVpW6q6qoC
w0dRcEm/9e+YrNy7FT6bPlgKgUFiHeiBoFVRHbdYWb0g/XD8PgwaxBc5s53fvfhkfvAya025CqC9
a41RNku89ZSkaaXSXhknf7bHhJMf6Hte6JjZXD1rjUWkP0Osar2zw2xVlCc0Hzk2qTXatG9EFfum
PgBsQY7q/CfQgdlhx6SDwG6/OgCkobcNcIBXf0nrTFe0W4VY/xSs7AGtwe0UJMwyvVS9Yc23CjUY
lu7dhHdLSNKSHYAdgrjaElWjZGXXJq/jSXPKy2CYOFtwwfNt/MPM0qsLYEU0fZzMop/iE8jDPism
jILupf/D9u/lSBWLCaWQRUsnogPNl9JD9Yb0sU+qWBvmZhkiv6Or3ltnbFN3KMLJwfvEibJwK28f
SZL/ELIfGjC8Eb/2XN2bNl+Pgh2pMTvbXRdms20oqxqLniKsxtr5KpWklNK+99Qc0pE/5SoMeu8V
kPBCBG/gq4bcp95AtuQ0l7qI8sGXnWebEyCpxZUv7FAAlhfto32dPG6OS1w95BdMimJ+CyJAJSu0
ZXYkmiAQowTpCTsFHh4ZlSdJN7D3g7r5vWI6frnLg02fk6c5fgrempu4K7mHuVFgJDrpuReDdMGv
0Sbeifv19YO/f1hsAumOKrQSR8MUk2R2FlyorxzJ/OAwd3RXCw4pOy9R0BB7DZPke8e4gmNOx4sl
DMG7P1GcWCEq+K2VpOm/X5dKP7Y/aT4spGrIegzv/A+49yFbE1+cd97dEArp4TZ40lrVaqZpuLco
ZhrEkdDmbO9XmSFK0Pe6z6qpKr5njBUoHvnkoGHJXVtVL7wa4ZXPii1u7UDJMIPPqtms3RGCb3jZ
GpbZ9pCPgXNMhaVCd3yWTliR16yIZdlOLpXOn8y05Z9O8IDXjUxIRKj8tHcvA42ezWF31ooJet4m
4HMkUDuutk2+RysS2UMVfrK3Q3HBzL/p7qxEaZMnUz0CJbno+TBNrInGeTKshBPZLDAQ/ssDwTDW
DQLyKMtdPpRCYetDAgJfcxROpeQUBPdH94goMIBJ6K0WTbgY7NYTCvd899DqCl4Quo3R+o9QXpvU
eiZo/763FLTQQqrhE1tLQxROYabNnqct5L101qkNDsea/us4j5La4mZkM2DJBta3strbMwovwyJ3
f/PvdZDDHHo+riBC5IygZ8roc8wVFUE6sc3GzlkDSKNH7L7TCQ9/KaPMAZX1blByI38XmPYQOkHG
nwwXm0luZDFIcnqtyl70zrEsZWIq9qdP+4MGhhf5zOj3dUFbGkgBHU2aRxi6wSRdm08KzlBSDZw+
jdFTuJpKpDVtSo6mPG3CkzKHqgV0OiU8uyCfGrHs0TTYYRkvPBBeK3euYTZbFUoIIyl7CLtjmlqg
r2PcYQcl+p7qvBr9TPFo2JIBSSeUuegvHtAy3WzTZqmY9o8rAtG8nwTAl/FZlaMxGOIjiKk4wv/c
tkN3BS4o/wsuEvPc5zYUNKuOQA63BvmUNUAUWF3nxFwOXapbXZPjvGENjl13ywT0MznWHtPYp6fM
7SpFeKbwHObnNoLu0/mBm3wxod/FIy60p5MIckqoYjzrspNVukHjQtrElgrDXeXD9eEbendKiU7m
0fYNPFJ7SvBbBoizVYQpBalHZQJ0emf/AaDVuAuA64hYyi80m0j2N+rwSvub7iZtES+GCpC1H/wN
FmPqFgaUs4anV73Eqqe5GiuQ77oKi/e0ozqcJmKMCo+PeTwG7bPue8Ou7N3DO+R8033LX5l6Liq8
trjTSZwsY96gKAsmjgTglTKQtRU5Mdct7JM77VH3IjiceDT9UOTZNnuXJ6Xq6d1D48SOpdIwTvLl
eXCx/2KNYiaSawYz1sluwNzUcuzi1+AafbYSgjr6qdFKtH7zkk6L5ajXHmfU3Pjdk98yU31BMCvX
yr3ZM9U6eqEPM1lhGr4P9kgU0b1brQBDje7o42S4jK1e/sto98/3i9pmbuT/EoLrdkDWO8fpctiK
XsyKjdn1jw3p0aMbnDh95eu48Ts7xSKqlvI8oQdHP+gAvTYdoA4sdn8hX9pHdhwKzt5/irKfBbFE
2EQWAgZ1wJn1KKwpFCwiwTd2HCG/3++SrvH30jjSxE+YbgGwHxEEsdrXl0K8syF7C5jVm++iFUfO
YzhMMuFwFtLiu1DidvKy+hpVLIj0JIkCWbiBl4mIfHH2uY8QqLPHeY7u6fgNKGH041ica4ne+uMX
XDyNIv2ZufzgVGBrvFqNhHbQh82EthvshnorOSCIUbPL/Zum7Sd/W3X5FY7KRFED4DgAmBO6p/Rv
KPRCmfc4wbuDHHb2NVCgRbxWzpOU/JeMfoQffLRO5+ANHQ/35BoCh8UOau1MWTsSubQMPDIwfXsl
A+CPj6raT65XJRZPnMeybtzuM55EPI5Qgq91ADzFWg4YshSICMqQINAhxpaU1whgGS+awLd0IfV0
xuhHLjgHrQrrqOr/EIBAB267KGGwCzxgUKVVJBUC7XzvpRNvpiyHju56ouNujYR73vpEjlFKUmv7
TaaAJIl7svhasi8thl6nb1KDe3/tF6MMa51cupbA4NcJaP8t0kNpoAmhRLDOCZK6BR0NJR3KbFN6
W58UqxiZOc3KdVr8AuUsk/+rIyEcUn2Jq0OOytrtKtIKj021Rd3y4PtftXTSm8QAOEEr1oyCqFc8
9HG3hhVuLGYzoQhj2iopYbLVvgeQAUFXWdklyJcNhqcm7xNrJYwbs4UsGZKXhkdbFYOfuxPk+hqy
iURk7HYymsfzzFhj48y6gUqM96COEEA9Pcwtkv/orWARbL5F5JJIAN3DA4+iInglZuDVgeHFW3gY
BflH01W9D5vTRzxUR6Qc2otiSh3QhlYRP5UK9zWYD9q0glfJcxcA2rg6+g7M+9v8x8DvZP+Cy6ph
7zVTroNiaoM5jEHUEMLxGlCVTMcU2/34dwGKex/ky4JBW5/e9oKkt82I44TyL+isAX7qaOIsTMB2
6L43404qKqiO5lsQh0rKfkl9/GoRWbbrjI+BpaDOBM6O+4zOqmeRTvJ41wu3inV/5F6LXqNTX7t7
s2aXEkzuV4qhzr8Vgz3qYaOanDmtcpISPyBSB2v+waWVU49ku8VY2QBUPZoCFAZdmt4H2aO94Ji+
1KQuYLxnVWpIdjPvXtXuJFF5yXE10Q8H38kfDfcxAv3D5OQ1HbTPHD0LnchywUZLuq6lFW/Ask06
OOJiX4Dz++oRHFvQuh7OF2D09J+owvcLMWIU/drTBJN/m22j7ySHjeJ+eZnSUprQ3JCvq+ZXqaRu
+lMdu120D9Wxxmwi8dyglQiJlXX0jjDEMJcmWRXE6Ryl2Copfwb4eC3IuqtDTB+V9n/FoA+KeGBG
1oI/OpR9fsjkynB/BjrZiyTV5i2k0yT8DDochFa+pfxm5j1imfG0WU0gGXvY2R/zh/hWqguaMHHp
8dJeegDLpCPAv3keVpTPyZM+ENeFh8fWDaNq5RGgrfsKdIcxHKW33+GP57Cx/sDK6Hr/hkUOGAUy
fd5HuA56Z4x5htnUKAL1oL+qdNlyfhrBtvwIMTuaDpazKqNO7crnevwNZYtuws4LFo0PpoANRjvv
3fO2wQGtCeVFP8y+cV7PbsgIOl95J7BaNXF335v34kswy2J6pmD6VjdlacIKz7F7iE9siFfddyLi
Oo2dTJEpH7uEs0qXgKsp1W8LaTTvcNdOaaa9WOvCgMksc31qWo7idSZjDtjKuNJjJe4qApIEjpB3
fg8rzcY9O6hLBSWukFwSkBe+SWJmGj50cBbRzByF/I5DF/eulqrKVX/BiJDv1I97yPtRlXNC834X
P5HsXcaJyq0GH8vhnzLRYC5YnYLazFMVtqAHlk3pXuyoHMWBWjO+GStdo+VFiSxSmsGlpm5r9UsO
DOPMnACMs8atqZz1sO2LoPBhWrVMiM15QgEEUSxcfdP6YbTNgFJwGiXAAAjIjeqVEILhrQ7pYWcG
NVI3ECQI2ktuKfMzK19vHPHoX1EwGnL0GrNSAyLazsFTxIdxY+xcX32xpZgznzErWXRp44OJvKVx
8iFOrcSn0RH/sXGCG5+hXeE8fSTkiIQy/EFFhDwCIz1xQUARisge6OOkcBUfWoHrZtNQELRfl1Ht
lSPSWOOGe8EGLgbGf29Ok6Aj0ARbXRNprtTViOPkPZiX3niRJ/lPq5mzDrMHx0nOeGTpcmZPHCcj
HreggvZRLIu0HGlPrFA1t6RJUO9Pb8kNflrm1iEznsRJMGYXxFHzZk0U6Miy7ETWFXYXTSU0GwF4
cJq0YJDuhyhowj3M9DBILJY83oRKmcieb3hSW5UQRa8qm99zt8ZqX7y7QjAd63C8adLGDWORAgv4
t+C4pSALNx0r6mQNt3S7NxVxyXbUpMLIoAUbj2QAbgMf22o8y0NNigUfEC0CyeHYNkhwxYWUvvqL
8TkwP7vupnUzYLtAf1Xcw6oupryviUXVLFmW53oLJw+WeB+APP+GfYrWMwCRCTfe0A6j1nI617CG
ahqEIPGm907q5XoR+seFaIqs7lBM+Zg2fYyEz+7N17lJCAQLqiMsz8Ukdv/7sBXj++SJjETotA1w
9qQoPncQdArQOzCZDp3uCcZ2NCkHP4kYBrWX2cipnfVXzic/iynEy5B9G+JL+Ma1MMAih08RPyW1
au+BFZXig7mJr/xWZQyKt7HIXGEivemJ13Ki6tiBJPKOSBzpsIcp6iOV5EsDQavBmVzpMUpEfMuR
2bgQoytwT+W9ZKJ2+V5tcdHgITPKJJIgRW/nuxVlCZ3RPi+GSOaXKPK73v1p9pF9ih/wW2AOnAPT
5KJXEFRJJTNFAhiKIHEkoTf06JP5UwXl60PuMOrmfGeW8C4pz/cjmHynvlbQcDWKVV5TN01g3AMG
47Vu02W1pVB1MoYLAP4+E+WOu5n86izDu8TByzdVVCmhjrZ2pf4kq+b4/A17qd3uIYgdbegXLtX8
IEppkUTf6ZnSZSjOVfwwt9z9mcwIfe0pLybUee7YO8SW1hRlYYti6vN5RMc9KhO2SSsMXm5+xIQf
3p02ZtxYlX+h2fEUoVybzNwEq9uAq4gztQT9xoZvaep2CcCU/cKu80Zlr66QTxDJlXRsXFwa6DxW
PjhqUk14u4gG5Gw7sP79ud6+mbSWyZz5tVnDjI4XodH/oK9QuKGPRShiY6/uPnRS6hUc4172NvGY
NHavDtSQXURUc4EF/MoPxA7VBr4XItyoaM4aMtZUEJGMUwctbPfioE1Qqi4V7Q2G5d+WUKCiMt2z
hgzuyIHNoDdyD4gNx6RtW4spkyW/V1rwsDjLZVQd/PEwuw8OvkFaue7E9kzoiDdkdlb/++9X+PfI
BEcmE7g00SGQETGR5al7TSEkDjuAhH8IHXC8F9TfHOcAERL0TcbwYJ/STNFJhCkpNPkbxZJBxnAD
wuYvI06KF+3fpQu424JPcvDG/j1ahmHVJfkoUSxYQfsX8yPpu16waBe/x9zWf2jXBuO+lVl+VBvn
KFMuM0Iw1SE4e+lrGf6VV5rZNAFGoa0UwTbz9Wv5Ve887kx4Rgng8ho56MpjKzWD4h0gEApiQCy7
cDAmy88KyDAqoJbk54SinklmaPIeMCLt9o6SdTy6GCLr0p4zanXy46ILG5c+sU6BuCAPc6gqvC4r
jVmXcQHLCeIH2FN1ErE/SHy0/8u4u36moMsrnSKNaL6+unXK0ix9aJFrChBqKqm/opYgTiK5iOlm
+XmRU3bLdKIs35vm8EJSrdwf5yFH8QoMs9gS/bExLFTHBvJvaI9w+Z+7X/E33clpbQV/y0T1Y1oP
x1vgHZeuX8LAoEIrrEN4P7xrTQMeBa38R8GbfrLyIzXb6lAYTWcq7NJ0lmFc/HN7de1k5bIxonNm
T/xIi/yLIxjEQr2Pn5yVx7s1+owoZ4IDVAxT8wNQsfJmIiMUhwIbuBnKnFABSZHwlmiUVnvrl9Xg
uGwGdmS53ipxNtuXNYfT9zj4SAYnunDxsswReC/47PzeIoThTvFoYJA5QtdaHHX+dFl3s9+upcRB
/aYcwVdRGhV89/eeOG+NCs5HKe1sUnkU8LQulp5F3tiS0KNXtjG6Ei7NzYKI+5Yl1r9RyUUw5/lr
dK5qOMkpkrFu10WWKFlAMZOrcPxxQOZRpiuewm/yyIbtU7Ct7iwb7AVmS+CTlpi+qmRmRz552j/S
Z1C20dlWOxSf9PcxKnCL3PTgfpEOmPsN+F5HU/USyB2ZVO4ielGmIiY0Z481LQdhV92im1OqLS6L
8EQz69ix2BNW/6WHyghcJVAJE78uJEKygnw7eCL2HUCcQ0uSV21ACiZrgeKJ5Iu+9ODA7dKzbuRJ
kWnwqEYG1nyADWJeUViKIHPXfsaico5bRzlqi/hZAsa4G9AxGSZA6SMNbCIhGX+ZXWeEVyjvVA6s
0ToARvqSUrXVaQWTXj9X2IIBPig+5usMA7nnvctA4ycbUwXsp56etyaiYyrMoMaH9cKFf62uHb+a
pdYBRtZUATkhreCH6fG1oGajrOetIt2CW9IXwto3XvuIEAJbgolQnRdqDW5Efv7/DM2lAQqyFRPd
39AACKa1Mxqj4GLWGBe/tDO5620UBczO7LJUsbAPLSA9fyrwYvPkcw9oUCrmLm7FArE+18By5Z/H
/lOfUkT8YtMe7qVu8jvIL9xEUz6pJDA4JcaseUKjFtVHdcGsM0hg0wm/R2//F5vlBO/h8os8Qikn
OIW6Sv8+zMzNQZMmzdK6iab59ZY57Nx35hv2rtce5y0ofLUrb3jCdpslsmuAZ/qsF9xpPFZndZQL
i9/Z0yXu2oEV5V+wYoNtb8AdyTyl/BypduJU7Oyw17sQjlzjXFTV13kO1ta6EoN6CuZUSAfLb6fg
GLzRlZASfSPSsLBoXvhrD/CY2Ph0F4s7akdXiFo8ka7VrSBoGfo1Pc4yJK28UAtEC0eYfvnh+47n
HAe9kxE93jI0V6vDT3y8UDqMk+cM2muqDzXgmZQjEF3Z0agTJ260EtepVd8jd4hQlHuZ2BDdWA8J
18Yl8JzWsqMwrS1ZpsWTRiLdrpx3apZjpyaKx6X9o9z5YrlCjAXnWpov/2PcDQzofAPUgT6sKf++
OBQIvXk1VNPVbCBwFDzJ434NLmOWuvTdstb98dwpeApBJ8vf1lprSNMuwT8n8e9Kh2wN4Bvz82Mk
2n4OoDl0eiw/YovJLuY8tWfiT6fg4iduaCBM2rH2YBurL5N2qbzil82lK0KstSuhNj1G0nshl9Ai
Y8WqSmaFdhBZx+OK5hv8A6aDpdcUjzIO5ZpZPVk8vQOHK0ojJ+4ntAjF2Zj2hEcYTMlamysuMMrq
53pTLHfyt0z9eHIeuzetvuiwEDfX4iaDlWTaZ1mA+uLO1/6Qs0tAunsWMyE9fQGPNv5bue6pxkqH
/TrKjfUSL/ORqZmK0vhYprNZDXgUeMvqNyoutoRgKHmQ2lTvcEZtdkAw+C3aL99uLAqNgUCEwX7n
MViHIRw/Knk9Xv8AJSF458kzGgdJ5z3MHp6T76n+eWVLiIdlq+Qf+kuKy/zC3mwbBHAs+vU4mPSq
/GD4CjLzqe3xqM1S64sOECFqVhTTKKuQ9SXcYViYxP7TND7OP2miHJTiFyj8zhd5qh6ir8irJ5p7
pdujF3I918Piqp2w2LZXKmor5wH/uxuhasWx5YIJqfAAAovC1cBbNuch+jJFWfR4hCMp7KUhu53U
1JnpHDW7gsmOnLtMGlnkgYarcCIOocdqvCLGe2PHkonOi3c8xRcqpBPBxqCcmS++Rh34NHLYgQO4
CeZQ2YjdVTVMyS0KVhuM/fHKxVBtwAa+fC4TQ9Lqn3Jxah4Jadyv5rk/GyAs+sb6L+DNfhiWUQeY
mexphRC2CjHLYU7T6x9zW7OuvN3Plq/TtrhzkrkHQdeyC1IS4NWelX60gBBc/zXhXc0Gzbwk4VMn
Ijbcvwsmbet0UdKdLUOUvv4vjjTZjD+fnjHM+9N5RFwo9m4TgITDbv1EVNV5mwOt/XJNMrZSPo6c
cTDEn9TxhIroaAbTW4rw9UVFw40ZOF/QzX1fHc8MzdpKjahMfp8qTIsi5XrhMFwDKSChoMWFRXUB
E/Ax7hMTsdXL0yVDafaGI7D0qB0HtyROcZjonm5WobNeStXdgHdFkavhmhgAasj2/qtzQvzgSCDu
6F4UYahH5la8Jie5ki6ZfiWMmSg8+d6eFpz7oG9xDRjdWxrvd3+YD/c6dQMOV4Z97ojSOkF97vLh
4zRHUcA1DG7j0vykGqSWK8PI2DWikd+s1uhWFScNnVcV3uHRT61Ely2t8MV10zc4tZMy/2CbYoK7
rH/olG/o0mKBwQQTIv8bMed5RHTSyHkjzcCp6wLxfCXzNQQn4LYJ/y7TpSKCRENL87VoQ+K7uKHH
LL5y1grlEHsQh62ITSA3zA+7W+S0oYL54cvwTE9FczSxEYpGpxCWN8dH1EYQTR1pRtKhTTsOigyV
/fMQ8+B8iQ6a8CLH5qAe3v7IGEeD83DOjWJ2SDaodARcR3mruYpYDdK0bwU1iSsDAIXjLp/n1/n0
xPhUenkxfUMz262L0BQCZwBzaWmlb6Wed+KboARoozfHc+npppvn8g4WmFrUlr19hEV4I/omqyjt
LHaNehA5P6fXw83uzk0xGualYggbSz1KIa5d1gUobb6o+p6zTcTbWt+lqvhzAron6w81nd9IVnv4
gm0N0SfpOozU2zShOFBU96UY2/fBEDv1m1ca1hUd7pReve7y0JfTHqMnlqwPkMmCGE7UdxptSAQ5
8GQtP1Nk/lavtto6v8s+RnkMBGfouMx3dZwlwf1tMAKrQcUWAlUEA2BuqA7LMv6dNcL9HEZjCoM9
dm8Bc5deo399WouE76g92ISuRXbf4THiPaSycHGHXtoP7jRlgGd/KDfptJRxxClS7ZwZe+DhXfR4
LjTtySeFUBC8ON7czhCqfP/kOW8/iqgopP/xndonvVMLJEGxZ9hJ2PvWw5owkDX7pOeLNWzBpHvt
SLmypxV7AB+f0dJSttlVdmuzBwn12INLBMSIv571q1Gj2biYc34Vp+uv8xMWO15ijdC2iFzxPCfU
TjS0UaB9QuYcFZMcQxsyIieUS+ai8XIpqOTYn2kZ1ZNCDoor2V7/neTfKUbcPHa0eTCwRI3hPRWq
wSSsbGpTWgAXO2rtP7iIVjl3gGcdIxWVux+GMLxZqzAc/alqcxAXk2XaeLJ5tyTVxEnYZFqbD78C
qjgK70+qbreHE2H3Z9YpErQqlUV7aW6YdCAps5TOn0qT+OymjQb1wGh5y6xF4hJcOw/5ihPapI1M
eP+UowyFHUe1OfCZeP/IayXRPPOU/tgKXLfpb/Lq2EHukl8JZFBq6/u6p6jFfVy20eYA84I2UVnZ
0JDzo3QJoxsRDHm+Fo8ednrg5b7oZZHLMM/YezbHuaIuqMEUhZ6iznz0exfYllZ9S1EvIzF+gU04
vxueZjZQyXqTdcVCZBta26/AhW6LuM9ivyBhDBo0rb4zOpS+DLl+Pkh1/htTUS0qg9ww0eygPvZZ
ymMIQ0gGrUkMhhG+DahvjcY0qGmSElRPVwteSYv4lGWc2mG4EISbV/UxPWRQhMM2SON4FnUaXwjN
19p572riplE53dFnV4nvgtCN/HsnYjddJY24h59LV0gDLnPG2r2rtBFlXs5A31SIsfsTXkEZELfY
92rpj7oaxhZmeb61aAGk/23x2blXjC9NEweZD9ZWmA5STjduQ6fCxOrVeR+KBRb0J1tsAyCHVdN6
ItwF/Id3ZG8McWIAVl9JYjeIZbs1wjuPXDu8qkZpd30YpH2ekXaMeGeiED8p3lZPUsRteB4xzj9d
WubXLH7Ezqtj0zpefU71lkvrv/9U8Mx5ZNILDPhV1thMVxgmO+TK+tYnwGKZrkARkkPEmeVJtPYS
Z+dMIztF/OXWFRm5+QKBAV8ZVgo47hwqn7xsJlpQpx3U6Ws3iqSujLFS7V1RanHD/hIPOluPM2vk
NBnv4/ZEX89YXjsN/bs5QuMPkR97Vxam9WGMsUtpHHw3Jq7RWOM2u4qQwyCeA/rlKP9wEi0hQmSK
c1r0jDWAyjPJ06NQ6Xp9UlCejdTGIqny1YywOuS634/GyHOY8x3VyxZcof7cvVBYrBkP26+65v5w
cCCOGYyqn7bH7XUOH9VJ00AdQYhTzOruSBJt5BOxJOQ8RTphTKkntwvcyuIs03EjBxeJpJZ7eEwa
v/9JdBJnFDqzAzbl7ChGorWZiSp+FmKAywMXKiUwJUAFZNQlIeHIFb3jDgHeYB8UEdmLkpMaJaGR
GxPBzJznKo7arZMRdbYx0Blr6exLUBh4SfSaepF2ouZ4FTwag168TqRZXmi8/WTczCopRtsJ+2bb
sAQWLTrtOt+n+GH6umN4v0EnvGO0TCr4/vEEK+58fwLPV2nF1vfF2U2klsUA8AIZH3K8uPdtIvQr
uM2CAEw1FXuZ1XWl8JxYXwq7rHp+D+OLpUb3IwYRkd6OmnnZSC4XaUyyqJNZgs4XynmQwTHBJG7q
+6O/U+jpKJAniYdEZfyxYljT46IQsKMzd3ZHhjxNJC2Nm1zrGiRmkMXcfRhrlfDvTKm5yUZ6xPbj
Wx6IYgVTgOn2gYNbTQpUHTCxO54W+dOhZpp2muDr1GTvxRoxksAmjtRBx5DZ+gN8SIbUBBY8friL
7c7Il138zbbPT4vcpqugXfHffFePiiNUusvj7KiBBLipZ7a6EEftK0s8a42tlsCF+czgSoXMFOVp
YIPnQcl8eWlxDmJMzG8YQ9i5C6OH3Jhlda8/b32qU5GyvHMObkg5aT+gS6Y/u29wXTrpSkL5TbCN
DxT/1SZ8PbGnsF3iTJgDBYJIF/ZKtSnY7OSSwRgm/aEZz9fNhVocgQJtSaPsw4TNcULX5o2LV1mE
1Ymx9VJRjBO/4KHT5jeYYVbj7RGKu1rIIx2oOrQ5rz22U47Qd3GlvLjwZOiuRROEu+YoDvLMyCt1
XS+WPjzZKLJx5a3RiZHFOSaq8AwBSh8dYvv9NGrxMAhIePm8+4JyFlxYWSE3iRzKFdHJytm/aF9a
MFe6SSZJmo3nSlhdmQAQTXVB/7U9qWcFwrpLvnjWNIdMNOfUQF+eWRpkD+iXzLQTT+KUPfyBrnU4
Ty82IR3o3Ce/3oxUr/50LkakLyVkEYeEgwS77FlV8qSSeF+urbr1/j7LokL4A18Oa9dqYWOxSJ2D
TPDD6Ys2hXTXQHtnBcxum9voGh/VbjtqZm9iSkuZPCB0IuwwJAwpx16hs5xt+04lLjWpzjTmcxTG
i7tmqWSX8JvEqPsQAz2/152VnnekAUOh5DAQnfro96wlPUTg2Oeuplc6aZdmoV5x7f+fmLGdaOxj
5D23xnB4Frsme7QWcuQIeW8Rjtt49HCtdNlbopg6k29wewMn5NwcIkpYKcMIBhyOQvonHH5JTHBZ
RevMJ30s6qTGFnUPC+9o3Te2vdGSg7EDxteUrAviLNaU6/W+LrPQHjIOW6G3a7Qe9BsmZXIWiyjq
gvoDb+DyVXeyA0N0qM7/3MdzQpYu0dT7op23Gh58iPHOfjLfqWepN05QSEapN5RT2v2a6kxsrsmO
tx7cRKSorCUOqdzY3JmaecQ79ZQCHzSSexOKuOWq88vGiVBWhUdkqHhi5QOArRVbSBuHeGPyFPDX
5+mDyA4P3YMDAJXIFHx4Sbk7/bCThuK/buCWG5dJL/pINcG3qqzc0TF0SEXABE4yfk1MyR4wo45z
nbq3m83+Xj6vIJHJDaWlVrfAvzNyVN13W86pqpalPKBpyL91tvbggBoOScgQm9Sw1T1HfiQFrirm
lBo35VdAhqi1QrxSX+z1cgzi1euoOPHteC5G9IO1jsjUkzQbcE3zu9UfnPahJGR/nJLt4s4nDezt
cGMuodUXi/C1Fea4EzSRbOO2CnhF/NsSv91yB7mgofPqtQlLmNO8lMSVqydHO4uNSlWbOxXMEuoY
RcnxCwY9oUPN8BKpOrZkXJuY2DgTcSZZyUT4FqnO82FG2i1Ri6BQvITzzLQcd0yYxJFQvWpuwg4E
j++9tWUGcPIdIgCQPnnl7NJLuy2V93sIhoHBLJ46b4gIDjrslZeV3LL4uyR+Bh3Xun9oE6UolTyo
v3H8wRZZ8U1nDaiUIizVi4XIe3f/3xDuuucgL11W8I/VO41yall3ysvTKyVj2ST5ZLVWeyBft4jp
ZU1DLF5WuwPjtzdITTzh/mO4x9YZpRR2JEV363LAk6fGp5QRtlLgyGORtZRNOwwITicUYmNzfguk
V7SQCdMV0Zm/FpJGZe/m7BAeEYRV2uEP5QWH5ucAWiBRhsGTrHAFOygMvSY3wTJ5QWwojTHe1Vgf
j97AIyU6IXimfgivu6dF3/Yq78AGIG3QqoyTyOLlkGJTUr19Ws0VPyyo6am+ip+h2NUj9x9I87uP
s1oR7esmVPQle0G1BcjP1cO3ox57NhjIrpkEc+sSH3HoLwRJV5pUPIQ/DgtdzcSoPAJOsy+KNRvh
r5tEf2Mj2ZmMjaMP4VghTqKtkz6YxThKflAcM7ANy0/60PnSLpuPM27x+2zF/IfzwPUAGHH35QfX
2TbdJsQxdeuuLolnQZpwC9v4o/9eTaihq1LncznJXEUlEPJiZ2wewC61u0NCQxu9sgmuIld8YBL9
1LxrTR4F544wUhKkL1x+2g1DyqbgoygG7BtMK8rv49cYJybL46eI9X199oPu7GrnNWZ3+4DE5Vgx
KT3gNHIoSH0pkpc/MnjzjsbR9A9P2IQlVpFvL3y5OTuTqZwXy/31qF5Az+r4iug0rP71Yj/H+IWT
7zMZreIAhveyeC6ZgrbAaV0YKTbNFgV7ZQ3DG0eaq15SYbxX2duYpXajR7siSaW1zNQODCaq1DLj
U0oNs/ls/Ci/54YfAApZ20Q+/uwKScEec48cEYS7pDFBJ3kLDwFYhlhvTI2UciLbMGBoSnMNUjTP
wlh4eY+30X7X/fq/8IdEhB1SEgn3xkyQUvyxtkEfQSEFxomQaW+9+vf9If3IHTMuunypbjNftHpE
7+EYzOkIyJjaQzoilL2fJH1XwAG0WZYCyMCfdFjvLIsKuq6RE0AAAn0jvBHEa/ZUucJcstkHqGmd
a3rCnZSFZhTnCEUfZJq4zUhSDcbr+qKnIAT2oHdEA+tdXUb3xqHjJyPAf9zb6OBcFoc9XYotrIVW
B4kYTgFB9/6rhpZFNydTcwQYdcebIpr0kYacS7JbNW/Im6oCX6XTAvZoPzVmlms41oihyO2KcJiT
a/TyqwbEsJH0fY0kz0XhuTfrWsd1JDBhAJLwBYoKMZe+aC48EFdUCgvjchmKFz4HpHeXd/bVNXhf
unFQxZ8ofM5XrHo47sOrvJso5Tqlr9PXZQEHzuEzVl/njBZx2LaWA61pNoKMmjOzUNvfxsmJz5uc
Vg/i5Gwo8OW4PtfpZ8k8ZynGFAxmypc5GHRut0HoB1AP2SRjG1aSZY+tSHf4/emEAdjBhNQ08kk8
D/WnOfe65TltbfkDZfUs73UZNHtXEHIlkbso0d27sOSJ2+kuqWXdYVINmJXfvirl8vkD2Ac+jRYS
Zai+fT8qjUq8RIna95WxYRNC0DPQInMT1B7drkXhlmX6cpg7avfmxQkA1LqXMX+IarmW38QOdL4J
5VnWNPU09wypidsKs9RKOGhQ386MTUOtQZyL7jPmxS1OSWbqdoyjgEuStLTgDNK+nfesemPXJ01U
R+dNIXGOKnYaTRFjO+6ntJrBIsYelMdVylvUII3DfAanSsOoHNpNVNArUKZsyVUZVoC12Pa9XKQQ
qeWp5D/Ev+PjXPuRFMHYirZAlUJtn12GPfJ84pnFPRl5tAEeEPnhSTZjcnkZ4yLZMowDv9Bf2i2R
asyp9h8W2wOZmdQVoBxPk35EkFB7KsOPmPMFrPk86fJMhHF81E1MsEcsEM+vC5Yxxtnz0SzhY2BG
Z4YHIdMg9v/p4/LbkoGg1QFfh78dsJFYpDYfiN81pmlASFV27tijZo2tcHxsC4OXfwt9RIi0vEuG
qyGoBcFWdYNDrvh0ax4X03+s3LCBl6uu2L0TfsU2WmPQ4LrQg7XKzqlwdTxYJWzQZn2oh4vP2vA1
gUOheuPXJdG2/8Fpx1pMdX3QKn1/466+kHDLN9jKlYPpC9GXM/P/Nt2roEtAkleB56+VwOnl9z2s
1Ra7w2E4xuRu1feZjpcWanYlFz7WhS3tjnWOgLFMcrvfn/yW3a/751ewLXS97kINCmKqjGRLTHm/
meV2rMtnc0ysztuNx4dw+ESpftTMfAxfk9efYEZxV8+ZcdgOJC3CqXrSaNKXZVZ4ccET8iEeQysY
10ICBXH0J002hGedvlYctuupiCRNiKtPH+u9XKAslxMMphGrI11SSteTxIvyp2nVKOoOqQFM5xtb
MjwGVAY9Yxjl4XugXE6EMO2WLtsunBlI8Il8F8ejmcvQm5W4PoRatLanbfQsLn8ARxZLHKaz84Gw
J493MRQEP9+jNzTjem1QuTi+42FR4yofNu4lKLsH+bL7JkVbIUPJ1BAE4zQysZoO3skKQepnznvu
Om5RNji6e9l5RDIcKL9/eyP556NIlbzJYjS4fiXJ+2F55+ZJ0+h9Miczqj+j3tw8G62Cjnrm6X2b
EJwdDtxVbRxyv86Kv6YJfBktOVt5JzAQCP3wrHDHb48OZ0wJu//fF1T+riPZDhl+DwjWzdRNPAAm
WsJ562cxEdA7ZGq02jeIkfHrfZqgNtw7Giv1wjjj24WCdZjCAbb/OjNowFUAxLZbhIaAbrFFJqvF
U1zcwD9UX4TRQXhaYEAONyT75D2TXG7FsNKpUOppyBoa7tO5RsOq8koAdQ1uJ0/UWinUUpz8ofGp
k5coxGlXwG5SUUd0aBNE7BSs+j8HsICz2sxIRtoSV4MDk4zja3J3IRb4Ss17muZDfUQq/IDmI8xM
9qKtmJItD9doFgs9R7uakyYMOcKxI2WPIkScC2j0LEJVW1EYXtsm0WAX5SvQIIxR0wFJwRYh6BWh
gYglyTpWvqc3OCpkDFi/DHNxbANN16KAm4vhnCws1yy8B8tCG1CZmWJLYxaxksEmxZNMsU66SVkr
j+kkUj7AuvJYyJ5MZ9CLRVnXFL0EUxAXj0sqBvE8iUzznMPjZJ4UCNN+fK8cItKwEEC585eq4bUF
gcVWGk8PWUXLGBZfHRacz57JeWCQ5SXJEHGLz0uicBrdVctAA9Yt97qYZ+mAKbh2yREHa/v5VRu9
lgR2JGRNvb8V/v+amm7b8E0yL6eugMvVoKjcMi7v+y54pmEegvPn95ComIOsmk8cptXLDKiy1Hz7
2XJKBxvQMXDvtJb0x5dgdOCyPSUG8Rq38UcNuQaD7f5dFPgAiAHKHl/QipzZZ5Gkp2cvSd5aueHD
ui8ozd/LHkNROrlIsleaiOo1onMpxzvhnmhz+7u/A0oPIWKngFOIt6xMQddKTT96T5MICTSHmHvU
Go97AI3xSX8tXQhXD6vqPRwiwS/C6InRDZX3ZcLuPPMgKulWSKRW+k+msQes/Hy6nZ4vQ/Xsh0Uf
zzL+iWjseXwh6pKXxHatCrg2a71tPhSUIamkfwX1+z5i4OVQHNC4t9ckVFzqHEav3nmcUZzbEQKt
ylR0fN50nLqcZMLN0HkK8zgI4zuGhV2fOqzWutGmyTPPAzWOeAhIXl8QQTP6AHjxU5eHq7nm/GFk
dJ2h/IomHcA16KGW+ljxBsaEelPYIggC8oF1b7hjKObSLuNzIiE5fmPmhIDv3GiNYNVq6ZNohtRc
4/4ErZtBmfW1mRUoi7/rCD6M7iHLMJsXBVS+1UQtTbPjSq/j06W0mf1snTNCoZpTE09VG54HjQ9m
oWNwGjBUa01N0/pBZfBPhT5mN81v+difjgjWIEVA65v6oLNxP4Gtlf3Lsiqn0KoFcHEXYUAbLnhJ
6HgCzPUeq8ZVldlJgCrsLeM/Gg24ck8hA3W9McBhPbo7EfCeYlvxVMR8NvECZu1XHsfXsUj7vkMD
6fXAJYj2sbfdDH3WWWl6ARxCTC5kHQ7qzqW46MrFJTNmrz7ed1dvvA1+9XNetO68P2jx2rIePAx8
qar+lt3P82M5e6W/P91hPGreJbiUq9pEtxjauwKrfAszVFd6rqyh74xJEDnAlnLjJ7yY8UzELHHz
zIw7CY7n6m/ivCi3+TVAPGJH53aZPW481oWXBX0TgzbUV2MJ/TODNy24QViP3p7sI7a/L2Ppaasp
MO1HsPRnZ6Ql8/DQmKoGqwwy8i13Q9HbQK7r0UZR3JSrTlTr1HWbZ8J0G4rEgY2btXRl1RqTy+Ca
dStLaCEoXhtTgK9uUdWEN1/Z5zfiYkGwgjk9DoEyfKkeDS27S004fnT03iHzskhiKmK+eDSNl0/S
NyRJEhWuIliKcM2O/9HLQvDr0lfCdgjeofFa3Trz8pW9hNuyFB6VO3XPGJhVj3ybD4Jvp6a8/GCk
h9QisqW2yLwYs/r0kAy5LfOXHzYmBYkta0qzjVjhHPLseARdfv47hSYaxsSRs27g5bZ6kJ4CYVre
AK+QBP7guDsfd/Z4x4hFYnf+bZ5VygyfYOS88p3AJRbJ7/Rbno8jdBtOxR62ROA1J04DPZq7pwMg
4REyfq3/5FBt8U9fQXBI/OQxp/LljL6AdpLT6XLQrFaElnvZYeOKE0vrhS1PrM/8EAmnU78QaPKI
vCqXQAy+34/TP4uNsPAo6exPu4oNTRbU9PHXiLvBC5qjr0FWan+ilaw1thSHOxLy6f9uyuBNGYyf
AIvYCY3Pp1F/UCQPyPuoWzWshxS1CHOlDmwl22P8UIdhfnwuTH6eayrrs+kTRgQO34XhN4Z0Gblh
AU/tzce0OpRsW5alcZC6XvWii0fEp3ID6hIq/kiL8qXJepmkQyXdIy6ybLK54QxhuxZUuPZC9E3T
KTIWK3gs8jyqlpxoNifhuP90Yss4AYG9NhlinrmtD4nGeFvJUG9udL5BAnhSE0dzSeBckFfzb919
pD000BoFWRaOGmyEG/7Gx1MrDr4UY8mEzmJ6OTnZoDSHvFZrpKlRbd7c88+pmjcDnOK2S5Ayjr5C
lZ/j1/1uaxAS3frY8NITsZMG7V+9LQKjO69IEPaE8g1qCLnQy0W6OXqPNqaEZsOOgAzQ9Z7c32is
HIZWEqzkL9uDP2/7nD4/CH+pZYRRcUf+CK30NMTJo4hpxXdEmGU0czF23oIhqliRft1j/+lEizCL
MIMufx5XdYS6zZhYio4fMu1BQqPgJzLfxvv9+u+aS8BiPONM94DHQJYoS5jrBKdm9BCq+G5kwT+Y
3msyQcXNMzA+6mj4w7fxdGV8o4X0nsHLpRHHvfnJu8nCUOFq+K6WoUbGvmCIDB+U9mJgKJjUCr9X
ZgNTGCiiIrTFrivKH8k5GNClEbVFynprjiKwoJ2vQAdfJDGtZ3DiMeaEaEEb+IRBZOp6CQQuQNxw
8eYG0I/flT+WF24TnE5s+eeFyYRYqNKQviJtJ1RrgldqSOdFLPM0lkpb8KzV7FLqVUAFmsOc2Zi/
5jqF/8Hc0sTC1EjRmkBKxXf5VLisHPozBvEj1ojtp29vw7cTJVN5OUtFtnyoye9pP1qnL/+FyMmq
3XIUig+Svm2ZnKbrSymEfp5Yg65QCbJR+qbxpIfBgfWKX+3SfwEKOAy8Rf+XyPmNSLB0J2Zj8Diq
62I980DL5w410m1Syg7omEFQZNpe8+E48GCYSgNYVmkmO4XXjBk9mQIkVI0Uo76u/COEbuwIA3CI
c+5nNuUA5gccpIlFb0efwOoWG19FZU9whIhDb8PdYRAI3DbeAmq9dgP539GLq+X4R3x+kZsL6/nH
CkJIx/pSaw0Ri4c12AHxp/qckhRaNBAfQ3ui/4gv5wAEjFXibexyFGJIlsqe18fsXSfCGE82SOg4
xY9GcqajYqjJSvLtvEYL6pUL/a1fx4yyFOnprk0G1+MqajeZcHrDvdj6dZwe8QaC5IhE7GXXGnNE
PjSmEukwEHoGfUnrUXP9ocytlFBsEwKdRsQTK/KC5TRVXqAmsUeayNnP2L4NNgLeoO2vXVyRTuTD
xfBDV82z2klBCOmihoBDlOWlUhRXWM0VAZcqPSs1mmNurkUnJ5IL3dJvwdzXrC0aqHUHJN5UOVSH
g/kEWfurdyxVPi2+VY2mFNGtHdTh2Vdu45Hw2PpdwiUjLl8J+q7G54aIQOCegAfpTRMVax5ZtRsD
DD3MHf0mJTBzEDWie3JQQIoMYy/27rLusjTfLNC1I66f4K8D7zIhWNgYqCjHlNF9Dnix8uYThxQ6
H4VQSeOqSB2T+tyGpH7sD9niICRmS6XoRFi6xYQXWE1s4+jgSOE3hYSJwf8lfUy3nUuHINmXKoVe
5XACu7aOZXbmGY2BAe+W2R9Fyzfqp3zH6yT5d9ekZCTJVwQHSePsO+iIHjxmBLpj8QvM3ChuWKWw
0G/7WDlOHH3m4Jtsw51T8tcIsnAiWIMi91gSVZvsGl1bJU/G4jcxlGYIaGmNRVl9Y+iwbPuFOZKq
sFFQvb91Q0SKUBCSI2C3woQPLWXhYme86j86PKGAowg9/UmcMyuifWqulSfjnqhrAU42uA/ccBWm
x4pcXqRbd/rKw63v55AkEmUopervk7uHXaIoSjYq90Rv74nrxd2mvRuuQ1TauYti082Aan9WSJkz
097pl2cQbXZupv099stFOJIyzW67hxkeKTZ0RD5+TXuMAYOOLcq3+D56ME2qegH9OOy/NYfsQ0Hq
n6duRjd03m3FGWj+riU9JQ1eoLGTO0pnccndm4JXsLjVNBK8JMqJKmk5WQLaxZyMjS2jn8uPDmEx
QsXSp/XNhEmTd1C/cONjdBM4i5ejVagsVHuUu5iza+AoWiUqH3gidzYFU5rZsU41FE+FvuSjzxLX
30nI71cqZ+HC4H46iCGqGI+fKyiaPssfIa/ffHsnbYvB9j/nf4NqBs0Ib6Kix1EOFKxKDrFfpvEw
MVXYyAdJi/tSvsjK+bEzKumCmWnXi26B5xfvfM/OFiXMdN6yrUTLys2rfYCL/auJp+dS/ztLZyU8
DkeTHNUbhUSGnghDSx9wOGtrNxit6aq3WbZ7GulqQ1yUMZGAPW5+5a4YW1lEWME7mqZ+xGJAlm/n
uB1dowkVu3bYdzlK1T7Bjxc73extKoVBp0QgWfoV1f12yvYI0UO8X3FIa0lZesuvOaEA78EbAV7J
sD8WymCta+7vu9u1QflVewPuoGR++4rc2G92ip2sGSn0TyAUrld8fsu/LVb1+3vz7BPUJfpgdzN8
PBAa7Dpm2j+zTXfQNa17IG7chCkoUd9fJ5Gi2Q/y/K+7IzWWlUqpjIfxmJo2lRUVQ5ivuBUGki7S
dAkNOXt43atiwx4sGHtyLaqM74dyTX8RSFulyyIUKyq21ugRRdeG8IuIkJfcYF0TjN1sHOYTgLJe
GJzoM9qBjC220fm08qSvhaRWaOUJeq0jlf7AVvER83MKF4RZGJunVHrcVRmwYzJgrt37AwEIRk7Y
3z0KqW7cV+oVkvvJmTNmjyavd3qjHBMoWRQarjeX51sLJGWuIewHRpycDyxgIMIDWbxsQlb9SB3s
3BtCWNMmYsq2EXNYOVhkFMLsTB777mOTQyH3HAZshXz7Ive+t83Ru9aU/zDE8rHxhHELQsNfmjUg
GUkQULXh6CW1icGNs5RgolygaYaWsNo4RmXuPQ6VoXXfKZVuDFzmgsQIrk6I06AtnfpjUF8dSksw
Ow1Xn94cRwJhAyBrFhq+hPH+csAiFg9eE2dorzv9hoo2fZZK0mJLW967LMflnP2WUmewoKPa9FIM
qiSbqC32rMRDdlk142lGHXjLaZ7nwaOp1OAN2ieUOxAZc3JLSwaOG0+VyS8we7ktkTUUVciYMSyX
npUcdI268D2KxyJ9UEZT3g49CaXKTNVh5PirBgR9VcRwcWDVb8SB9VNW39JViFbohK+ANP57kZTK
4DW7M/qqa+CDRpsdXxKNqyAByoJGkegeG93WMJ+fAtwUafRfRVHtHq/QaE5p8CEpR3j12GETi6LH
bO9ZroUIe+sohgGlUR8dhW8QRC4vigJniI1F5lky0s4+73krO1QBVkgYP3YD6w4owkTJWUfO+Lci
YJ2zoVcMpSABX4FgnobBNKKCXORnAeNLUJKHBVFNmLmUi0ar3VwxrGmfHyA3TP8sjSZzLa+zpLFH
6i/IXjExu5nftQquGt6AnE+vavUKwlHyfCA1ZwMl+ZcbIz61cSqej+TNPlVQRHbpdPEEFi4CVnlh
CJJoc8QGrwfTo3lumIrIaCBdZOA4t068labx0blguKGLhaCqVbi8C9BHI1gj05Zl3oOCBdk2HRxR
7IwrLUfIkGPMlFU8zAmt+ddSQnmnbZ3Bjj84qvKzmjYREQvr8OlAkSiryF+czmwkOFQnobRp4mUi
pBcjTmHIkS5GVgh4ZZq/Y6JW8o09ruta233H68SmyqmOuobDF+y/esZGwi1sTrz6Xm433CRyA9dk
EL+TlOiF+0/JLgjrYF3kxdMUC1sXvRsZlcw3LPRCXgx71PkM90nDoMBjC1kQLOPn+HrDfCdNNmvc
tF+p5TzDniiyP5AMXOmUx72zZ+hfHvVjvVOx06Y/2ZpHvnQ1EbP0xIZW9ddCnQxP/FfpJRb/bj8e
14Ij98tyPyqjoa8WYfZ87rXZNKD+rkjQjCXyhKkg6FKfiI5zDo10Ww0oh6FEUtix69avxFi+oLmQ
lMD87Ank54dbS5Vj0/AyHMyya3hkeoHL06ntugiVSn7FQR3p8gdzfydCnz+DNaeihhn8drV5Ns4U
u3GcTzRON08RJpA9pyMKTa8s1AxfIn8Tp93j2uteyd1T8649lj/zsFqn9Dv57OM5w9N1trKiwey3
D4XOmZPJNxtaFWsC6qlcKQW4ULOFA55/y9lq9Wu6GL5CDBWaSq9cUWNRvw+vRwQm8vAZfXzylwUq
7qOvtyzIPsJe3CABW0dAzZHJt6oFZrms4RgpRrv/V1IPAQg4OYVHDKy8RTygqUJG98TDQTyMO9/k
8yFgk5L/KJYcxl7tnr+Tje3PnJcrtbIPndR1KdXy9nDqnuLG0I21096J9w4msTCBgf+Cb3/TAAVd
BZTzU4nCvA+IM17UUCiFBx8in/aSmkya+XAtJ0dgh+iPsw4Eaef4XwwLbW+vUR+0DS5FRVElSLNx
hrsw+jahk/D9+TwMwfHfO7jB4cRjJ3v8j9isrW0lpPAsmPStdxHpa1W5YLUuVm8OD2mjwk5jc95L
H5N5lz2JRgygvh0t3myGVToUHRjEBpUVWLSkn+or2HMeSuqSaZ5GD0gTDyyo8TKgo3hqoTnfReLJ
xkPX2/OdelTPf/r71QyMH9EQpQkNs208pBuoh/GxWKe4eVj6/g4zhukmu/CrA15+yu4+X2Je95oc
42SxqqBoopb2JW3lmWs1gysZoi9ZB/BLnEpTKwaZALhMEeQxUne8GQJbap515Ja59eKOVZM5RdBy
QQALM74zC0+bCJ4QyHyEF3U576tQ4lakK66x8QUq9YbXwOrEUqlqHxNZWo3kQZj32+Ur+ZuLH3UL
WZlWlt+lfreFXWX093Ri418FkK1nSxTTeuhMlH24ITV2uyo21/Gi09JMRpX3w2KwXreLwDTi/sMU
xbfHRcdQ+gi1KWQlVzHqHuS4ac8WbvgJVuRIbR2qhEc1pBTWpx3dcrOdhoEVs+3krspRxUIaDP15
Oqtl8/oCe2CzwnrQZXuwx2540GZ9hX4NTysyxF9qc5KGWmNXDwDAlHnaVaN/AIZ7fY7A9nQ31NQN
ibuV4jB5/eMflNYt8qBMfA7A2LNZxy8iri/KiWepHC5NLPAPD/Nc
`protect end_protected
