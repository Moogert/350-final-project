��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅRۥ����A��I��jٯ�S�s�,<BD�2oZ�)����Ȭ"����[�n2P3v8i؊bv�:�4���p��^p^W�Ga�8?OH;S�v���������Ǚ�5XE�$�'<�y��Epb��z�^���d*�`�6������r�D� |�.@��%]�9<�W��v5�yP<6ZHa�
��� ��e�K}��q��h9(J�G}6���O�<B�����W��F/��N`v<#wに�gNq5!9� ?��+�ĸcP���O�OA���u��~��B}^W���w5�,��Qx_����GBV�q��g�:�c��ع��p1T{)X!;��V2Yڤ�Q�`r���/b���W�B��ӵ��r�0Eʄ"CS��#RY��ӽ8��4�QS*��6�L5>�s��R[�WT2�]��,��uY����M�h�
e�q�Wpt j@�~���*�g������4O�	�Ŕ���$�+�V�|�7�N�S����N���ct����BҎ�O:�kIV��4Lk$�4��q� ���X�8SE�4?���`��R����. ,`䥏���Lc�J	W c�x!�߸��s�7w7M��[?�N^�ư�K�k�o�����*H��au���C.s��'�?7r,���4�w��/H�u�i��fޝ
A���ʦU��bý����r��I�Bl�_5*��.=�$頯&[̹<_�\��)G
7���������h�AmB�y:|�ߤt�@�:4!9� �޵�Z\"��Vf#�9�s�e���ܸ>�Ġ��k�jGX0��&��ɺ|?M[�<�=�b����T��
�_���#"������~�&���g�:ei-8���;*�F�U i/�Qi�n�#�ݍ�̓�L��@>[��,���@m���"Bx��P)�9�~�˔��t=q�$����+�8�:�),���^�?��B�WL~�(�,�;AB��~��Euᄬ#�.�:Rv:=-z��ÇO`�Т��OTI��yy��hđ��阫�?�^�<Ά^nyd�M��K�R�SK�� ˰�g�U��2�y�	Ԇ����ѽ��D�`���ۭ��D�fz�ztZ�J�j���3U�_y?��ah*̊�NC�����o�T�%�y���7[Ŭrn*�@LѻZuZ�@�>�I����{��U�F�\( ��C�p`G&���U�N��׿�XA\N�F�T:b'RԢ����q�h����M����|L�щ�QqW�@R�e��*�F'b�a�20>^,I|��I~�_D�n��c��0�W�\�d`�#jS�}�m�����L�G�.��n�!��.z�'DHJ��ǭ������/�6��B!�)�*�3���,��q7�a��)K�6O*J,�*P);���Ytp��r�W���#��h�9��˄�l��f���U4�,�h��-�[��u@�� �%��]/�"�<�)������ŷ�N�s)���3)KFQ�9��m��E9u�0P��qd�{��OFh�����n��u���a:xJN��;�U�����q���>,$���u+�Wgt )%�#�:���e�{)��;�S��x��I���R�n��'$_4.ILn��C׏�.A&���!H�e!���CE�#+_C+�|ϛ��݅���?i����&i�sk0�ɲt�����h���Xz�N�A􃸸R�p�)���oy���ir5/������J��/t���`�����1W�M����'�ާH8�.��Y�z�M	���Q�U�q�r�1�28�g�<K�8�i����Bs��֫h� �5���{)1�_Y���6�3�&k���z�H��b+N� ^�NJ���jR�����)�ya1hd<�d�*V�ts˖��c\�l!_���ے�9L��s��p�'���ؤ(����KQذ5��3"�3�c�ST=C���	1D��Ve(��p�����mo�����`�E�F�3U��C5~ԡ�k�3���Q����U�x�g�)�P4˅) ����ǂ�����'7�}a�z%�!��Q��F[��ȁ}�=�h����x�	U�Iᵆ�tL�s�B=L�c�����iVq���u�(��<�=*������P��H��N/�ps=�j�ўO�i��s.lG�j�*�����0E(=H��7�=ُ���0k�D|I����k���˥�ǥ��]4M��=��$[+�s��)6ů܏�h�&/�q��%(�c�4s���@Ir��@��EV��|�,���T��f�L�K��D�'9��D-f�(X�\{*�Ȃ�9E��t�:�	%��o5�9/Swl��?[����I���2#D:��mY�8cAI�+c�O�Y�uL(��y��~���	ºk������/]�^/Ri�'j���N�����X8A$���y��.�H�^��a�S�צ�>�N`p\F&z����|hѝ]
�B`�x����A��JSrnZ<�J��>��$H�؄���nԶB�ч�氫�I�f{E'T���64(�-,l��d�V�v�Ay�l�p�����-�\M��#ƴ7����㦚
��9l���!-D1�����y�f���4^P]�.�q�_�k:��D'��L�\7a��D�	&�#��|���<�����5��Z�4hԥ���q�EP`S�)4KB�9#~!7[
�H��'{�p˴�@�u��Buw���8�~�������29�����|�'�����Qm��uO�t�,%�+�6��D6�iB���^~�����KzY��A�M�R�>���|� j&�E:��!��kv��|IcAՆ��o�z�x���q�S�?��`)=n��e@�X�y���P������ޛ.��j��%��)ϑ��?��)��8�_<e���)�EU�p^�[G<�I9߸�p(ݓ�����?+���t>Y���-Z��ǰ˳|M��X�"^a��/�������o+DN��%�Cr�ʻc&�i���譌�b��A�� G�imΚIZ��R�Otr<�.�D���O�~]ol�򃯣Fp~�6;�OY�t�%�N��G�A{�4}�j��27.�:� 'i]^T��X�F�]�o���<K_'�bO�M�X�ZP��T�#%<�d[2 ��9�.Gq,�yOʷiș�"S��W�1�4_b=eC�����QLd�����
��L�WZ����]�B��b�V� �)�r���X�#0���0��p�Qt)�R%�D��"S,���&;{H�jtY���<3mu�ރvuoi��m�3#hY#(-�tx�3�9<�Ç</s�X����O�������c9O��<@���D>�Y99R�p��p.|Y�1��@DxB2wG{�������#�3��&OdR$�ga�T˔���Ft�w����ck^���p��7	3Y<��D�/���컀���t�d�/k_�Q9�}ew�Z���k8��(���8�eC.�����k{#!q~���&�n>�i��X��x%��\�sӰ��醬�t~MP�H��1��Q���w�Ȯ�$uI�J����@�D��?���õh�/�o����C�t8�*��š���䰃̯Q+T�ϙx��!:�ֶ�2Sb������5�5g�깏����f"��i�����l�rcj�������9�줌v��:YK�v|��mF�	V&��H�8����9�S��a�d��%�����mъ��VK�j�8Dr5N0ӊ���VI_��MD�N�V�<��3�4V�Q.��)�ƍ!l���cF$5!*��V����
"���ә���
�����Y�R�����1��o���;r#e�*�L��v̀��$��nX\O���Lj�ھO�Ȥ ���?��Ƶ�&�*��5�����y��5�h���/����ռ��2���>�;X,Z�*W���҆��P�qAv%}\8l� ͳv��"��@�gF�70tZ�mC-_Zp�����ˑ���zC�e��d�	B�7|��h '�7�~�Y�Q��2�i{!\��������X+X
�υ&��d���a�b_0��ym��cù���DJ�&i� �>�I �c�{�<��d{�ɡ��2�W�3��U,Pu��8N��q��E�T���<��CO&���5x�Kw`~����>9:Z�8k�;;p�T�K�6�0W�f�F�T�ONѳ� ��E�@I�hSk��o�5�~!%S