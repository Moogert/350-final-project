��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}}�jG>�q���*>Lq�(r�&w����d�]��`��PT/+L��S|L�ڐ�S5�7���������!�Ӆ���5V���K�>�6c;�B/�Yi(ȱբ�K��Z</ Wk�3�La�´������ԣE�$�U�a+D��g�~j��<F-NJ�ǭ����M�t�A�H@�?/BSx���5&R�Fڮj��V����o�.E��|e֪'�Q�u��jz-������������Yp��H��E��8�3VX�����4�efi�B��z���j���/GP}����v�?H`ɒbٯs�$��1�L�� ���+�Q�u;j)��L2O������ꏷ�g{���#�aT��*0θ��Qbޔ����O���V�r�#�(^Nz!ȥL��["��^Θ|�T0�5⛝=�8��V'#A������|��k�W�R�Z�:T-.��f{� � ��8��|ï�H�`��0�}L�����l����T��@f����Ʀ�O��N�0w�w[�����{���D�ȋ��
��7�r��*��'qE�.�r�X �l�r#�_�F�&�f�]�� c��M�h���ٜ��He��d��8w�����G��^���3�O\���i1%�	������R����Q�?=���xG
��t�1j��J[BK�8��i�+�բb��UWX��'e8��"����?g$�}羉�����*}.	�V�_7 ܗ~6=ԥz��a���&��؏�,��\�=E��{ŃTU/e�H78D�d!u����$\L����RRY82c?q�xJX7%����*���`䮛��8�V3U5kke�YQjؓ�lk�)���9l~�%��C��N9�w��������{�7���]�5)��F�����o#/�Tz�Pq�g�����<-U�*K�����ڣ�����h0��,���X���E}"��vh73��_A.{gT�]��֑�˴K_��`ʒ'�O�+�MJR�cYb��%N|�! b/�)+hZ���ۤl=�?sڙ*��z�
�����Jt�c�.xF�*C4��S�&J23��m̘�_�/IyqU�}����[�c���HIv���:�ҥ¢�tɺ�A�ڑ�~ H�%O��i��E0�No}4Bc�˒sHH�go>�r�ԁk*gv�C�����ZhP�sR,ʺN�0_���<�9�d;�x3���>z���5�1��P���w�DY��Y�R�"�>X�ҕ`����J���A��6�z0Z����h����c�crD���;��V7�>�3ҋ�x�7���-�.�72F|G�)�c��۝�_1|V�`Oa���;q�(D������8�����XX8��/K����1o��^^6�VI����V���C�Z�f+?�G���3i����`Ё���j���ƝI��A��E���9n�\�	k�������f�c�r����h|��<�}�)8`r8uB���P�Y?���F,�v�%>{wr*ȩ���f�fJb��~�;L�wm�q�S��9�ַ���S���[Ր�9�����L�� }dY�:��!��ݱ+X
rA3|V���y{=N6�ׇ�86��U^��%n��F��x��S|�����R+U穪���[Ɋ�bΝ��?6�WU���.��B�xI��WV�����WLla�&��Y�8��+R�8��D�jQ��e7��9����H4k���(� �ŋPT��z�a+{ګ�y �x���~�K�����aۣ�v��f��T������`�$�B���jy�3�PN�Эc��w�C����1>hr��<GF�#[o�xxف��eI��P4�d�8���ڇ��QH��ʞ{���g�S:F�_�_� /m_S>�,X�eM��sm)�>�?��"���g�/	 �b�MP���a_\r�l�E���f�'�f�1;\����f0Tl�c���E���_�J��d����I��j����A�Kf&UN� �2�B�����P�!&���ΘJ<�\2i���S���/�a���#'9�S>fD�VBd�8X�g���ޠՆR�o+ 
ߋ8b��~!��i���)��F_�J�.$nkX5��gp��Tݯ��FXKX��h�eŎ�6m��U��Wl���&���Ӧy�[�c �\�� N��{jz�D7�p��.�2H���l3t���Iϛ��J�
~*���[�`�\H�?�Q���9�^�����
�ȣ�F����w��L��1/Ì�ddJ>}/���C��`!i�D����X�	wټ����HG�":#��XI��fCoO�PtZ�
plk*ou�.��I�=YȅB-s{Î��6-Q?b'Q�֡�
cO$&�B�e4��o�*ąb.p���f�/��ֿ�6ʬ�'H�!�F�3�䃨�;5Ѥe���~�/���2��5I��HZ�`�Nc����-A�)��
���7�pE�E�[��G��Qܐ#K��ƈx��P[��g���nZ�X�Q7C-��0�-��w#�c�Bi�@��j_�K2�Ɋp>�w��{��2$�Q%$Q!�b�H$.S��;���#̻��0�!�$��Mt�E\���ȥ��A�Z���"���HO��*��^j���Y~瓒z�'Э�*0wv�1rU�l�ߊ��+\���lO�f^7�����6��y�qonzg=�h�DZy��@V�/"pq&.��M�t������Ah�r[[��-�Z�_�<D��8�%�s�W٥��%N�k�uG������r�|+b6֡����Ʋ{J�b���4:,�F��g�Ψ	m�5�����)�ڢ �*���N!X�R����OC~�ڱq�o�Z[��!�"x-uD��:;5iU:i���'�5T��P��H0��r*�0l4����\q�w���� Nf�s$D���r����hU蚔s|�x�ӻ�ź�������Z��T�v����6l���h�z���S�QiN������o�A��-b���b�v�q���3��pQO�����l�yتW� A�_� }�8�U����C��cIIpь��ꮔOE���-t9�;��I���1���Z�.w:2��Rں�����*U��{ܽss�Fߤ�B#��K��.q���=t������V/
�� ɑr��E�� 3�Fo5I�!C��q�In�d�LE*ɯ�ֹ�t~.qƶ��V����;s�s�-�.j��{��P�� �&�P��tdpSD��jG(�xp
��^��Z��3��u;��)���hV&�0��)u���FhhY"�{,T,B"Oɶ�� p؆J�[sI�S.)���f��j��g3�j.r����Hm;;����D3��7���ʜ��,�b>�:������kx�����,�p#&}�k hf.Q���UB$?ѢC�uDs��GS&�3�B)�m�~��Z�,��㸢��\��#J̛V6 w{�s|3s�1� J:H���T9�`�E��s��%:C��k��̌�I�����-����Q1�,OyK1
��P7��)��$�X�f~��q`��Þ}�|�P�λ��4pBySf�^�%u)j�.|���6I�f_�	�:ٕ��u�D{Y�F���������K�����V�-ǁZy5�ei��X�GM'Z�`n�{�s9����d���	��:
��!4�~:jȒ���;TE��1�B�)���A�9$�5Pd�7��4�����h�C4��J��藾^��2��= ��R?�G�.�������λn�0M���1(cg���	M��S	�܃w�(1ښ�����2Hc�e{������*:�� �#N�Z��'��SK��3�mא˞S�#��k��-�;����ὃ��tWn���$>��F���I՗��,���,1�2�lz� ��������{�w(��CY��"��S�������GM�\�]���e��>>V�^S^J*{Lo�q�w�>	�2� @����,�n��
�1�[np��}Xg��)�\>�6K���.dWkq7�f�+���+�ؓ�7��A	 �xd���@/���*���L����tEƶ�MWk��;_'��o�G��g���5 (�Lo�)���+f���q��O�c�:dPuw%�.pR6����wk �!���@)����eR,u�> ��6C��/�^Jg$f��Ex?r�>��Q�e˧���Mqt{�^n���eՐs��O1�)�ɸݧ����v��"P�c��f��� SSc���4����Q��?�v�����x|�f&k-zV˖���00�S�T}`*�����/n,Td��С���p���a����g�՚�ɘDq��g�B{�	�?5>��{�~$��1f�xn�m7�dm�@-��7�g#5��Z�l�A}��r����T`8Y���d1SX`3hC�~U��$�_a�l:���-a�o�a�{-�N?��>$�����z��g
���b]��@��0���甂�M�ձ茉��D7&BÚ���Ǭ�-Ԅ�<w�:�������(��]m�]ՒU�1*�6����!`��x{�]�b����BL��	���Q��ᡝ���ϣ��!�=o<n��`ϴ�v!x�_z��ݞo��"vn&�qX{�"�T��E�:�l�?g�iD�������)�r��w=��v�R����@[ˑ�BeE]��S�a�����_�LE�����&<V�X�l[/����a�MaX�b� �$`h�mk^/X"�q���3�����y���JͶx�`{U;,E���e��CK��B��=��
����[j�I��e���|ER�P6g�S�xm7�0��v��l;��+��nûK�늓�"Zۑb�����08ۢY���MD��T. H��'�K��V{�+}@���F^�ϴ���ם�A`��"�E� ���7�AA�� �c���s�N��	�zY;���7�hq���$�T&�����{P����Jx�Ɯ�
�� �"�8��̓=R�:3*�p������?.gL����2%�Xl��
�	`�"��S
�&��=o-�����\kgr0X�h)�X�����\��j��E ���=2Ý�|�n?]ҏ����q����/�pwV���b�"Ο�0������A)>a���e��>�i�Fl�%0`�bH�{���U�Z ��}�0_����xO�a���Wx��)�4N_%�u��A ���b��y@�CK�|Ȝ����Z��^�j08�������c���������\�wLWfal|�}���/���M���@���S*b�Q:e5�?� �^��B^�		� �_�j=ճHxRZ��T��%��`]cӥ��i���<���[<n{B]UMaJ�J�YF��H���>����m�GeV�y)��Et�;�<AE:�F��~s}6Ma	����X����h�����LQ\�sE:+�A�:�JGݖ�VW�Q锟��f�d�~�F��!0����`[*cps3ˬ��A��\�3+�z��Rzے�-�W$����k!���_�ЗG�b�X�_�;��~�g),j���h��>:��^>^�	��L铬���p@��FD��2�>jA$�fV�'�"<�Q���f�s`��76�������%�I}S��pyZ��H��Y��%<������a5�y�h�u�*��U/	��}��m��Q�O�����vH�6IWJ�]�������2_Ŭ�S$&��Z)S-��S�{��Zc����U�����"$FW)Ml��=ܕC�3��@����!|#��jl1I\b}��x��]�-�*bޙ����{gh?ޢ;�asT�����x�l��Ӛ��Ma�����q�� ��ߘ�*�k�!��������}C(ۍ%p��J�
�e+����|�"�Nxo@@y%Y�����f����j(���l�=4^#�pR����0�����&Õ<gZ��\F���E
����ةu���IO��]�m���g)$[A!��B�U��6�	�y��ŭ{y8֗�'�P�j|h��-m:A����Y�i��񡷞튆%�P-3�B:*~�9o�S��\���)	�y�]#�2�+4�Ѫ߼�%���Lq'7,�))����C.=E�HN��F�ik�P�\g@�a�� ˂�o��bd�{�!`�����������0�Qx����co
O��
�Toc+o%��+ ˝�<���	�P��^*��0��y�9 �:�����|j���9�/�^�
�9믥����I�Q`0#��G�����2��Z_���	p����_�Bg��_)�e�G�W���{`Ñ�Ҳ�흓ȼD�f�K�Y+��?{>h�����_��C��ݚrqqb^�O/��f�d}F�ws���KZpG�$�e����ȃ��a;��_��Ns(,�z֣.!��Ŭ��!T[�em����J}8q�\zӘ� �q��^z{
��]�S�l��tYF�����.�u
n����KU�Q�\˟�Yc�+�!��_؎Fƫ������I2��ժN��y�Gq��
-bĻ4}�1`���j��DҾ�^��c�+���꓈���h�*������`ä�A@*� ��)��,.��Af�W|�$��S�a�a�ubB�#��d��_<�ցŉt廫
�@=!�*�v�<Ο(��~^�%�.���^tMT���iޛ�j��%"�C��>�vQ=���^���OcU�'�� ��8����-<mikW!>�X���D8��P �'�uE��'�8�]p�ʢ��6Ξ���F&�.D�bv����z�����u��y��; �mv@!~��i��o��1�iL��]�?YP���_����/�6:���|aѫ��{U ��a���:y�zS�"��F�vi7a��Q�\M����z����>�v��J����`@y[ɇԠS��D��,�3w���Y�WG����aB�ܪ\��3J���R��WZ�S�z!m�T�Y8ESP��4���F��@I�1��S/�.V�M���&}%a~܆8��VS(��n���̮�C�;QE��=���:g����.=�,�d���AeX���بp3���
z�C���Ͳ���z����޻�F��}i��=3+ڇv��˯nG/����w�:{ض����Mz�I �;Pm��k-�K�����UA�B������qi�6+��.��������n����\�����lD3ɯ�s( ��/)n�.������A$��"������܇<��K���B$��8bJP�u�'����m���a�KUL+T�[��1[�veR�o��|K4��/>Q�G����IN�nm��	������;96�ϰ�\t(��C����wY��e�]j�P%�������NyEԵ�ڭw��P6m��dr��u?`��aP(M�U������*�dS�`|uM�EV\�^ ��u�ކ~|�#�U��p)�"�Y���?���\~|�
�{�{��8�'���Ecſ�Οf�6x��{�_;���By�'Zk�*��)�̶�m���F�L��i�����1LJ�j��9f=$�|@syt�J ��Q�ҹ���x/�eR<�>�%���έ��Gy[�q§5�l�Lo{/d.(sj�؅��2�����)N{���vZ!���Խ�쮎V3 	��O�Vm^�OE^r^��@ż"�*:J�p��J�(�5�