-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
defvIG7FMPiTfICQxJYXr0azNftwsF/Bq/W3CiZZxIOnI53lBeo1YdhtXc7v6ltuOIWhOOeKweHu
ktFm+NtEBWwkezHMwC9ms85AIyIMzhVBZ8wWRt1tndepU3iwYYPXs0bw3VD3TFZKW1Pat99Gmvkt
+ZBjwWFobM2vvB+MnBYKrNyJLi+5WnYxJmWqiJKISFD1fW1IfwpoAKbKlaEs3tiZ/h5/XDyJmk3D
ztwL5GA1wf/OcMpRU49ju5v0LGX+XuphEcVEj4E7+KIXQnfmn1/Uohbddw1k1ecXPLyoIOcgKPDL
Qzdv3ClMaj8zzVdRQ3pvWZG5NY84DpK5mgDShA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7680)
`protect data_block
3usKJjzqiYr6o4GQY9SDM3ekmQp4I8ouNqLGCB9x4085GnAaanr9yY7uCP8517DqNxks0JhecLhu
cCfoEgUn8XAPdiMHczxumRxWh3elKGk+SsJVcBqNoI2Ea9N6sLKVIERXqbRRN3Mam2HNAp97ftAY
ZGHhLQR0T05S28db2mjfYPlkOxFuKlW6oKs9GnD2TCVCS8fEOpv+MZ8bBFPT48i++wSWMWGsm4bd
Odj+za/sFJfoB4cf+ESxDtpCP5aUHGVJ6QM1tEp+GRNO3HN4BQ9+BI+da6uZPPhgfTUSKgf4L89/
BExCcVe4FTvAN6DSxA+wGJLhiphzqJ2CD7E2XuEeedq6UeFOmzYakBo0LOh9C6vxXccKLXZkds6r
gqv0ZCK9ehCEMr42wJF6vg08mH+JBbNacQXwZJ4FUk2tEnDjpwoHBjoHUgboiOOubjdhpjCiWQ5i
g2UQ2ErnfE/Pat/fLveISzf+hbv96eOlS0dHo8iiixMFtciKDy982KEjgUCJxn5d4eFTeNTb6fNn
yICsczNJ8pUDpOO6BOXoQE/eVAXq56WDaQNl5gUawjSa4UGW/TzxeOXfMIDx+Lo9aJEoyA6g2iFD
uRmDEtn6QC8pXCLZrbQRvSWI2enmELgv3npHoGwhbJgXrU0I//jccjzotWsHXoVgUGUbxCIfVV/7
Is08nA2twF6ImxGlo7xEtpiDHkn6mya+6m7keZdBT976ngXkZdu2+SvoFuncZELx2AEC3MFMtSzu
RSAX9QS0KAYrRYeznyyWNFR/An+xR3u2wpWLNxCalUNvgW8go44+hGp9p7WJ+5f50tcB0oX6jydJ
AiyVkIe+7cncJ4EOlW3snGbF3AmzK6wAaeyYe583Z/Ye7N769/sKlgN96ikwQPSZ2n5s05sILkhF
Tm0H9GY/A0UGjvuVdiEw9LUbmVP+joVL+jqKLijYTPx7QPJpdN6nw61e6XmQz3ujcz8JIs9AHzyi
E86lifCsR31m80AntE7WlXOpnl1aAmykkWSS3EE5zuyCueHN16JHwlEx0vDZ6D5ngvONTtRQIbNJ
2jBt6TbG9aATiIYbuycSB9VilDWJICk4d2PWGbjZrT/RoHfr3ul/ozcQu+N841U7eX/PGPlcYhSS
t3lzGoL9Mx79PR5PMq/eRZoEmS/55aCbFhm94zFcfLmn1FqMRzRuE4I4yVZ8huN4qvLO57eI82Ld
FlQun7m2S9CC4F7qZfM+Qya+3kp80aj7luchUsebRaBG/MJ5b2buHSdWA+yGlAn20DEUurxMMZYS
NoRB0V8BghfvqCr73tTiGkwwq6pwO+6S4Z5fsxLDHhhl8wseb3i52LM62zkquxJu/EwZ6hKPLYdm
mSo1Gmgg0AlntAeGhFXsE+98ebwPnGTknAOuOrV1RwHr2XvPHZaL/o/O8C7diz9x/QeHAoonWUFr
gD5wCuJxdOK3uv0c0yiusHp+LHwM7+rnomwV7JBZ2NUggUkfzXRevvzOYQICQyQHF78lEk/wKvT0
VwO4GwiHFeU32ka8Xn7Z4qhD/2mZWeoulflVGgyYRh1YOeIEYwT1fBhhxFilhenV1cEBakzfF7vV
ADkvJKWfTRqbSjwBWZcT1Q2cqzlAuk8VZWKqsqnbmIC2a4d2K8ZMWC0U86YSGplmuw2E3zjUgD1Y
W26AfrfdfIC1zLgDrktmXnloznp3tnzMfzqZ+FWwZ47r/UA148WxblagrK0YYFNDhjI0w2faNX1O
BS2dIliCwXhuHnu6VeJ/41U33SoFtxrOtd3D2CYe/7HltkPACSql1Xki7AbyTzU2Q4J115MQEbtn
5kbBQphc9v18mE3kf3RFWxi+rMTKZ1yS1z6mfU0vHV84oJmC55tv7LtfxB42IULdZFmbh6YikIrh
zOKvz7Y4meUu0ebg9zcr5f97h5L4TSKbC0xu3cnL8z1A7AwWgJ6q4ixNlPpc1bZQCM8kQt+r4R5M
flMxnes5ICc09xv8HxMiWoM4cHLEbnrC0hqHYt+EuXkEHZKsr+IgnkH0ROuRkhwAhlGKDm8yfNMD
oPmUYShpZutbM8tn3PEUbT2FCGdlay8JF/9/oFI6et0fVfEr3b8/qR+74TbC2QKtTApygmeSv8vE
kQfOmXr+OBqCDdi2SyLUUtCOqlCYDfFG3HYD9iOs5z0S0eugryG+xaJD3jZ75iscnapkXv5dZedD
6amt+I+ygk5/z41cI5aMBcRzqvdR0VMINMVPFwMa1emMDUlx5DKDzVnC8ogMei1lPZ0W/PsIJX1Z
WLRZeZ2tXbpXCZxqNp1+0yTgP9LH2n9u6Y7lN8mdr6fXkr01aP8T4zF9HCC4puTHzzVxYUtVZSTX
HaAjZ9mV5cAdIaV527dg4TALZ1Rui424kmbJblOy7Bj293GMqh+t9lpTlGQH46y4bhLBMKrISttg
Ptsbylwkaljw9+3fAHSo4ZrRZDFPDk0LFAdkvwJr0Qm6FVi0k2UR2i3/s/9vLioik0poSA8yLhdO
Dh6stAnPMHoYinfKGnYvYcY+aj+tjLzlFt5hU5t/0VpasCVcrf2pDUy+2exNX99XNrx30pU/sQ+O
Q2so1874iZ9FFGhsijJsu+DucLd9l9mWFyBmym7MBzCozrLVHAh6xzOU9DyIRorNUo4cl9zppY54
Fbb+yoCtgMB1LKp0HxQ4sqsPDqu85X9uixbzEl+Fy1PKE2eA9lcNYRP8U6qRFhiObHciZDVpLaSx
83+QpL2aM+S4ZtfTWoiRudWytXAivjpQLOpuwB6LThIwxosp0gM9J5HmIdLnaVZU8Nb7AsY6MuzE
08VgNJ8FmIPT6p5W5P2VlUiVh21EY6A8/xnsn8oq8HRoGnM34LsmCDrc5ct8tBw7Tc8i/Az2OInc
r999g0jo7uvDL+zDWuytBaTBhGk3xQmE4RteQXNlD//4/M+4/j7xCUDhvMg/x+5uhZEYH/ibDR90
vX75/UtR3Ua/7AyaW5UEDXoSP15u+oojSkCmtUbEfbAOQmeMrAqZYvaNNn15k/JBfuYcTYqZ2h8p
LLIFX7+mPbnVNnIk0q6leyaavJRMsNStvsxtqzxmECByVl09+vHTFz72/mE2ZZNyWFCNU7rLTc+q
yQ881RhcVDIsvXkxOQXk+8gSutqXSoAvKn0iF4O/qeALII5QAphmffetGvRsFfui9Ks/kNctXo5p
Knhv1X7ngUtJGv2ALWn9aXrdr0mWkGN3o06DX1k6zMnknRP7jvG4n4A2BB+34dsau29dTDFNHOb/
GanQx8w1Zg1M8/L1z8ZCeJzatpRx6WmXfdxpGRYa9OqHbM8a1WyKUVG/CL2lkPNx6MBEtHNIKkNU
Bd85EWlcGKkmTDqXdpqGy9zEzfTAxTaQx4IL4EFYN/oczaouniIS0fdFI1xqidr5tXz8PgPvd9jL
4D0F4orbMWXXpHqX+4k2P4dFTbrmtCemz77V0ROHoZIR3FAzapYbp1peAZx3Bri/HzgH/XZ9EPYQ
/YL0JRP0w4LFhnemwYCjrVHUsqWM1DwVd1NbJpoEHcpyLKFdhnPTPoeGlRkK9HfONvRGGnjsZibo
Q5MSxxHxLy8/iAeOj/72MVQMMUxROpxteT0LBQ0cv4QEkq25rpniVsa9DgqexnI0iapxwAoTj0WW
NhmvJ641139FtlIuLiBhbPK+qw/tnTgTqh0Mkl/Mq200310pkMDBqJWwYj3eBPitJ1w7lkEcCixg
wsF3wXkNRJwvpz3XhFQoLULHIdM56lWMdKh8FWt51r66ToP4+NzFYNLLhezPMsCuZ3fbxdOgxlbq
8vJssQGSyrp55gHtHpxcOSkyGCmaRU8JXWp4ljrMFH/6Hv2nED01MqbRcpTYjUbcFJyGe48eNrwY
H08EjtsYHbH+gzypRE21nX01tnNoamfbGr+l9J5lPGtUQ+UNex97RaUa6l/xG4uPbTdVDbPChSDz
88u97DtJPAtCdtd4IZ2smBnLbk8O1WPfDXImr0fMrNAtL1a6KXeiz7Lo0gPy5JVF93PnG/Ui6clQ
RL/BdZIk5oF/glv06SgxBvIvajeTLq8sA5DerSo1dd+8R9DG4qj34o1rg77zWxiuLmnNf9XVL3Nj
47qSK0yzpu0HAxdPV50nu1u67PNOelDEFv0er4QI9U5zTb9nrJD9wQJsZIt6X2rkViNFVbAtl6qw
vy8se0oPvQZqRd47prBCs9y18BWGxjJFmdtE5m9JdEufmZtfpBlTGMsbJ2eEa1tbZH/hp5BuxWVm
D3Bf1MZfUzY2lGfQoF4Gwt8NgHyrs0J/v+7Khoo/OaEwzlHp4zZhYUaiSgXghCrffV5vQ3GcKdIp
WZpjcBYecqAMYbPkcRjryW5wm7ZZYhlhARVTkKxwEPOd20f3KadNYYHMu9Bqgc1boV8Ea3LgeYPL
r2I9jDJMomHvR2PYpxntcBh9hw0m5hRn7qoqMau/iSFZ1dkZuA7OZtK3mZnr6TBNc7ZZTE6z7I9T
aGO1gZpTQpK8QGCz8st4mf7d0R3sBaEnbDyyVXfTHZIBJU/mx1t1ym1I4eb8psw19GdDdhSKR5m1
5N955Q56MWhgrDNtQQQkTM7tTPou49eRNN5YkGANPvrfxHGXRMFUPIAcAGOgsbVohWqWYSV3uHna
+lFhCv8Rwf7LrLRzaWPt0DqtIY5rTzckSWiU3UZG7C/+ZPIjmlMZ7Y1AUTWgU7FCTjj4gmAjlE3h
ibwKIwZYYvqnS89easzR+RLcrjHA827PDQ9aMcMYMa9prcwLvpaUqRnA9d1Pul7dL1fpYfUKCaKO
k/htplNX29sZqMW/oswPllykWChb4F9Jk16KoTgI+xaKdQx8NJd0FjeW4rnkd4sVidKf6VCGaTgY
jIQJRfANnvQ+StXNUjyGwVgeaU6EzSiHH++upoaoPt0/JS6gyJgpsGBf3rnQfi+9b5QUahQvGVSY
nrG5nDNich9c2gyU9UVtOx6mjbJJh3AYAL0WvooLXYgqi9qD4B2EZNdgCWqwCOCzueut9U55/0ay
grydpXpTO/hZI8qetl6UdIGXjJU8BSDL9aYf+BTDnm6jUxJU7bwdlU2NbDHyKcuFXkFsk3CH0muA
ArNafYanfsR8rJWTd+qbQTZkLHBtErvuDgTLhOboOaVdkJ2CdsiGSa2CUTU/sIN5bSrOYLtQXJpm
DjI4URAfV4S3utdqub7dJ8L951gIrACyRhY1GOWLnra+YdhvB69+ih4vbTiv9FFh3STeCToM2IRS
uyvwTMoe/WnmJOWksK9nuD5cqHUZuXwK1LZtyZ0N6PW5gHYvLL9ctbkNmaKeX4PdTX2qEF9Rogbd
K1ESWICY/Zgn2Ws2Dm+eEEPrvexgytDSoKxeQHAnQggjs8NzjyEnP8go3JBoBkXxyP3MuBSk5qAM
aOowGHNU28Ret9QKPGz5L0U2+aK9G4sAaUQbbleaD8PfuuLXmFuKkOf7gLzDCE7Kko3BNRc+/VbF
dSLc+PXNpXqiY9svxgXf/QtNLU7BI1qSEbOCKSRPPIut6cjwG82it3LPU3FVWIKa/VOde+hAnU/9
2YLcrek87FG2Ofd2HIieJCTly5+UaGxKLdB1HHeL2dtvWfytLA/wLxqZKLHk4L+YRvQ1Sn+3CwKz
UMjvI2qWgo8ggARtN4nd5p99NCidO/IZ/EEpGsnLaBxXL/gRXbn4FOx4sz+xEvS12AKoER2aFy0Z
onh6GXhLcgdmpTf9ah7swVVkf0UmBMLkvanNGVs4BM3Y/4rKIxgbrLthD8YwvGC6unpYtvPKFBFf
din81S/m4fTcl+9FT7ltwyY3bLrHyOUZ+QMRMqQwSLEPy8dIKRuiXSXwNjLYzLIG0+jHrRJC+/nH
n2jg4idqcVlis6sutstKuxDYO3kFyBWpkQAuWGxXWZr3d2zab0NtnVXLprQRe5nOJ+rDPbSDwQBb
Jnz/gtT7qcPB5OCslYSN/CNp5Rz9sm7PbJTGHnKsta/hdh5GSQxbP6h1XDFeW3ntsbwwATUTxKwR
zfT+qQpaHVc2/ZDDnY8y8B8nx+kjgYbZVYxve1aIVu9n182zFnRIdnLtjks3xIp8gZNgItnHdEOX
LDal+w5J7trcMV5p3Vo+T/v48g2yDcCAJ2HGreXfVlYkLaeTwvwiCFm35RAqYEOpmw0qCVpBgIYr
eGPseGuIhrhLgHzfgvcywrm8w2MmMgvjt/8pF3nUF/Ymw5CgAjidtsucLyAGvM3AzXKd9zipCcaO
0mlvwgmjQ6y2JUYiNV9NNp+i5s0tsoU0w1ro42vxUj5rvhuJ5kdCNzYst8ymFJSkCsbUYzgevV1K
Bv1EmkYPgLCKjlpDqO1qL4bNdxjKuosY5tFy8UbTntVIiHqKmkV6MEyLosGonA2eXOT9S8RTYW5A
vFisNHF45zE0ocbKJPRPOBZUxTKiG5uA8QC1DgI1nsXCI+2CIJu+pUCRZY1N+h+h1fPOG1zXbb6N
o6W+UjNiM3vnsxV0+1jKxa5vFsXSApTDXVE6Vl3ybghfQXfApopFEyFGTNL9usULYzSgyO7WqofW
yZrxFs3ejFYP2K8XdZUUhWRdC4hyNsScf34MevSbRK7s8ZsO+S3zX1c9N17E1g9VCo1Td0pGa507
X5Go5owOquKjvxLejBZYdrVdvIIUvR8qHIgI7zILZJAsU23ufnjQczNdxJNh0UZrY3dq1dGnkrEQ
Jo8dE+cxXDkpf06g/xP7Uu7aiFZFTgukPNboNbcRDIg9zHnvbKMFhqulUyUm3sx5FmopbE51I6KP
/u1bToXSpbMi6hlLMqddfJfJ0YTbk2WgtmNzD/Sd+HDtHlDuOsfytd+cAGU/rMW580TM99R6ssvq
qdBNZuL1rLST9a4NpFGqdGRyycIzwjFV5xxgf+qnyRBggWb4mfrY6Fl+sNKWFMUvhq17VId7Vt4m
hwtd8YSnj9aqm0NPngmC7Ej8/P3+45Cewoljzl67fSfKrKy/tNU5qE4nPgvlyFWy+FMeEFOk7OhD
5lfYyn8uuF1Vm4xvZup2zMMD2lcZWfnrI9nnzGTFKDD0XOq1QQBEl9ZLSKvzGngOydPSp6QdX4Pn
vrsqog7PTFWnpp7hVmjiMBF4OkuEhZ38S3s0VfuLNKwRc3rgBGg/o89oOPWE2/NvQF/CuRpLnJgl
v1uQuaOx9f8Cg12iFzqhnRca0jbNCDFY7EX0/eEEtz2YOWv0mNCkDw08xgRrIcg8xTo0LIOFljI2
zPbqDOh6ItQ5AZmtyJOrTwJmAy1+mpo3wuHecNgU0fTpxqih6RUOXXETwJidZczRcnbAoJWWnGcz
1AX5RNIDkNtUVmhmNv4Olp4ZIqBOAaecjtxFgYhWO8lw/7nPX40hQw+RZgIyfjjC/Vmhn0zjApq4
USPJvfdN1QZa94dwHhL/+Kzq6EsGU9kAVEdMxjE634W63beTk6G5wFyUwKIZg6bbkXwSns0SVths
Alxfc0TIh9uOOcVLEbUyqW9N0f062uH2shpbe2k7E+GXxeg2oh8lXFJE+a+nHo0E9YFqJdf1FFTL
AiurHMwZYwJw3dEPrUGotU4em/CG+SlPdzoE3Xa9qa424n51zEHUl9sXXV6DGPJezL0mdVyLwgf1
Tesmfl/hTmI05dNjnC3Ok5nQLOEGF+itW1IPCkv04IY2hZtVswXxbyxRFAUzCCvWezTqHUiXU63E
7YDA3S9uVbF/heQSoWs20cpIo3ZQou7kiev9r3fMo1g5On3KY6rjPNoLPJJEtXksEq4m6BqdQ6Gj
QlUEz/qMYHAF9o2fJnfR5ZcZDK4YCqJy09WWZqphnhB1QLSmlCqb0thGbjd2mv9zHMN1/sLJU/gc
Wgv6okL3g0v+U9HlxPqlL7aRSqRXJqNPn+i6HPVNninGqvfuoUOVmG0rHEn+B27TP5RB6sSKIBOC
S1dLdJwkjtT/RDoE8D950QN6/HrMJZONNxKcECFLwPgbx88mLN76uMlrnmgMQo66Y/2fEYn+BIhn
Huauge4rbLwkAE2qN/lf8qU6g/BYOdG4Jnn4shgHfi9IGrkh2zQy7Eu+arIq5xWou/xgga6d8i2l
qBj2gkRO/OCzEocW2a6KWCLZ9MR+DEkvvQEg81BfgdHG27c8pTlTbNdqFFzoMiPtljOaDOCGARf+
Bx1Myy2zutPnGkCGK2pSmGcd7k4lYJR2h/d5w3ACMlP9NbsVqOXas8vPlw3I3GEK9MYcq54CbCl5
vBkQAPTE1+RAMW4MSPDAwXZCFV9re/c2wbRm8kHLbpFMQ2DTeCdxAowGm+IB4dxihyvgZnVXvxso
KZe9o/luQpZ2IDHTENOabWbv808ZsqFcjVjgIckuo2H1ndB86jLIaxJT6wophGWyUarcYPabaEjB
Klrl9bm7L2gWpWWY0oD9EjGBOh/u76xUnEV54vg5JXhClGa1HkwbhMK2d4lYq9YCSWfLa79FmD40
lxjB3HVUD2taZkfQHhg0+IAGj/1wBdQ8zDPfmBzntUYCiQ71KIeaaFLVdo2UWt3ZDeJbeQWYZcdp
S+sJnuQw1XCucUT4gVfUZNp14QpGSxm2lif/ri1FxdzWBb3PC6xBpv3sqzjD+wjEJC48cM2b2+zp
bEfjqWjRvuUE1a/u5tGgUx8QegLdlM9g9v94Oj5eTJpC5/OKGDd8oXViTB7lX4LKveOswk/veiXP
jJbc27VrgyRSRIhAhOUFi7KMmKfHW8PiQpgs6DxlWoOOXd5BeQ5rrjmYg/kANTEyy1SpdDkeux48
og7U0+T5uxg46JVnhOYyVbERpYgVFzSVamhFEYHkG4hxGHnZw46j0VJZ4W3bJy53wqiCJIMlH2mu
mtw7dDpjJBPgsckcK3GMxTLTBpVpg7eDU57qD57aSGVdcsKaIdcXDSHsyABf0XokVVCtXDGbS9+9
a58TwDzLl32xbHi9T3HP+laPcBIDxt4Y5LNLbKxLKsQCTheaay66mui6zOU0c13iXxAFvu9Me8Vy
0S6RGfAaqxZqHsLHjSX6tSO6fT+NkW5aPTS5/Lgt9uZxDectf2mFlBG7iR54/HxXq53UiOPM4pC7
0xmHdcUEEl1sL/Y8LxWDdCQAIDIxhA6YR8wamJ9J1H3TiTQL+fMAhCvWx2yQJIGkk35drwfQJB9B
204vEdJiH1q7OOO943oTTgCr7bg7auoMY6ED2TwerBj8PHI/I7tJE7ZZ8aiIYVPdltJ9YDfsYOnw
bPKBlQX10ua2r1RMjJWcLnJmk2rQ/7u+QxBeD7Xr5YXqDHQLYszMhNzhqzzNeRDZgVcEO9i1qcEZ
FLSnRMcIB3uQQ7SMzyzXQTdf2qlyzUiUOxHq3S0IMxbMeZIL+cAaAuJycBIBpLyaXBldbEuhITgO
kVATKCr/wI9mxMsr9hYWxR7i/WXnlvE9kDYxmn0QvnMk+Cwir25yeB6h4oUGh06pPM7PtMPJkg0U
iX8ezy6NPXOSZ40FdVzW3pY90sIW3ec4Ut2pkcR7IjQFnEbmQL+nsL+QDhr648jJPx0mJmYNYN/Y
cRzbs9/dZGwtNaMKcHeoTg/5V6qtVvsFxtXPXO2OvKpRlH/IHXaotI+kIU4nSrs6tki17m/GYkoh
MOyhHNcW3EimSUfTqEt/FTUCv2q8KRJ5qo5WzYazTflZKdvojd2RqxdhvzHbWrIOZg/3ovtWqWQk
akKzxJZofBvBUA4irtxMp5mbPdwOI+rsBrAhUNUbUNoEQ7sLOlr6yvY9EgSIp96m3i18/i69X4El
e6facQq1h77+PHxiN4wz89OBUl2iM0eiqAA0DjEN2kkNukgZ1JBfMpEA+3/lBKGXmbfxrG+buptO
GE2EzF7cfttNunYfy/5WezUeN4QR35bq10nixDtiXYjK3s2y58En4tjM9L7+nxeGbISW7dyQWTGv
K8DwRG6JdcmMVuL136JZ5jTk1LKeDIQQGgCUcNcI1F6beWQPNggEMtmW0iyfA8EuhZ2Fy1bB8qCv
fGgjNnwC8sQjztAaiRzFJ1UzcpezJvCWao+nfooYDFUS4cjgnt7bqzWsBKEbWruaxKuye5svBRWX
qQGMzmxB8zltViVL89Y19cSfyrNNjjOqBmBGpYBvEDj64U2aQdbI4u82RbPEnoN9/iW2++bpJOBh
mdrAJ8ikpHA+iWM5tjjrQc0a2KaM7BnEKj4Royc6QfW4vh9StvfNR/QAAFHby95oy5cjizgGpTvK
nDq6ayfUuVuG3akYmfg9DS00Lu4KQdUnFhigl+OiceZWMAHpjUItQIrj
`protect end_protected
