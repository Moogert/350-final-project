-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Vby2+2yL2TzYDTUmYPXG5Z9HJV4wv6M0KevDT6vdIBEzvwrUJEZOc4L7Ed65VoPuHgCa/jZzHcvH
UK8xIXrvLxJOHARtNdnSsQNr/pc52QnNvAe8RIxhokRdLI7HA3mWzuK8yUsRiLwGjrhFVje+viSd
l0IzEmjMKmPGpMPN2H9VImsZhYYfyCiGNjTidQA6pfTzk1BQ2lexAyLCuGvxGFRL7oGNuEZpbGWy
XQyD3vjJZhnZqyxhvFT8ZWOPPai+HVqPAP/h1X9S+uxWXYNDhbWHx/nwue4Kib3QuaMTBDcHWyu7
Dxjb+wHSKpvq/l1iABpvmLNFV6fXL4MyubT2qg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7536)
`protect data_block
f2/Y/yRoSIFdfZ7Z/+HXmE1DbxZTBTZagTTIop9d9sj9QQopnXcT3bjxh7hwrZGaKw8TPLZ87+NQ
HmOuwb4IF67HDWWIZtfozPqMqfYn7JPX/2rms4bn/f+nzLohM5QGPvzOVdxmhEiiUr1Gw5XcyI22
jsCSp2N/DolRPDcWRo23xp7YjReauCwkidFcb7w3dxAxu78x9bqRjZaf+QswRYfEF5GctEMbpsnU
ObcOFrlOYDlYaMq+npFOFf8DzeCYvUj/DZlp1ezPDd9f26jhTZGjh+h2fnEZHd/2tqx4OKq10t4N
MKOSHjLw7GFu9IYcu6zgqV2emkLpY5olw1rGinUtghxkdySgCeUB8E3WHImdph9YGPDqGjblzhQ7
dUpvPbgoltjtVpLNeeKy/5LgyTclKSxTUXfqRmgjeB2KaIeclHCx6FcvYRcGJNHKe7ChU6ne8jiv
hYO4/jsezQdpz16H8ynM3nH9B04CobXEH/rpDdv+UemsBhVmo+Zx0PwsRUoNtWbhqf1GriYtv6uU
H0sh8apvFYlxYVyQU1mSO2rqn1fKlNA92QpEvxPiTtMGKMw7aT/pVqvIOpbGiJO0UEyZcB5vFSWS
p25qH0HwADi4qM2uVRdMbSB8vIpzGguelLp6l4tNO84AGM6qcXMaxix6OMzShqbN488SiyRpMhQs
HGZzPvJVF2a8SdPdTkFqNAaQjvFcbgMmCjrsELPHwmJvHk2qmeQw9dJyORhP8d3OcgWrzNsrKayX
dWKD2GYZyzgwx1uapaB4ty5II4jkHaZOon+1KdM8V0OstO8UafpLlwzLtfVe+dvFLJjabu1OKszZ
2PQHnDWESQfZYpFECnJK+e/VpmNGspliAlZD1eq1/KScvC2yaFe+uO5eWqe1Fag/zqypUE+dcZz0
D96WDvxjMmXO9b8Iuqr19JpDosrhdIjjXn0CPRd/+NHrtCGf/ojaVsHvQiftLDtn4A9TpHjCMi73
HbTQJ5Eelp0HiWf46/WeYbX7aoU8dYDjVIpokK//85KFDrFDEvHqGOT7+/kRaOVFJNSccGbIKSkk
PqX/lq3Z53EdgRSNO9MUt4HPAMw7Fc+/LmrRe/cJFSc2W+lv5x4Oo6mkc0pk8R97g9+idH3etlR3
d+napOzFOC6iVA1Vo+pyIpeCdQLcK3zkb4onoflld0GAb2lJ+M3Z5JgkraGGe0rdoePaud9qYlFj
Kx05+CtOtdvkO/E0ETejYceGLg+g0Ems8afDRJlXCZ7IM1M1wBCFbDoBrJGilPYC/NMnKzbbLdsu
pNRFJh/k+ETKr9I7PQYuI8YKQXnTqpM0kiH0S4Zdp2IVr/WoEmpZjhVlleEk1NgTipmq6y5tKeLq
sIUrzHqP65+i7o5LJmv9niJEdvLUUfLzHWv3M8AkkqmN94Z3ib4Vso50kOHhqm0/bhoF392wvrtY
7/xUc4DOImLnSzYFg1B1tc4dkiJshZamHZUJh1TdIY56f0m4WbftSMcTVN27T3Ji/Mvl8t3sTRpM
evX2r1GALiDTBwDEvarG5bcUU6vy405A7S25Fpcr5J8cS2+fjPgJvRPPYG4V8dVeRbD9Q/my7R71
gZFmydE1AVW8rqfFrRldwYUUpsU3AmOMEzznUgAcgRH67s2cMyKMDOikDTmp8jPYy8BGyThOVBbA
xnz9DepfqbefpCYsthD8cKnqSOFdQws6UuRR8BkaHR4n2LZX7wU1p0QvTPKJF+VN3VAysknP6KNZ
nCA0fHAi62u6kUa0rN4uyNezxg3Ku3OIr3nmU/LtKFVKKllAopJqVm7ZLxSwoDpa96SzENhJ/014
kB+KFgTkbd0pX2gZLjGuKC+loAYWlQgjsdGox++639+/RyGlUv4CP2iTZf/7i7k46re7zD4T4bOl
febLHurfQP+OtPjjzuYSrkYIFQRaSZBSGQHoWbzJ+Sx3Q1pbZUgwe6tp18wR0P45Z5FgHxsmac50
TfQn5MYkuU4KvW963sjdd8Y3o+5ZkMnybWM93SuE2fuHGFcJdHXu/m6IU8tnRBiH4iZdTBX35u6k
BwuEeqVrc2ivOg45RrZbR0tBqaCF6hj3ELPgO+UBDn38yjh7Kfou6Qmr5BOh5RdkYcghXhLqVM9J
fl2h4CLyTZDbe3jaV92wuI5kODJowOTukZRLp28P2KSUqHw3inlETsprXZnAyZq0g3aYeu7TNYya
ImI6AWJ1S3KjfMMsj5O1Wio8pmdLQm/tcEH3Mls/s0p4ebv6B/Gid5Qi/rp2qRT0FbO8b1o1m7YV
r1UK4iyWTr+/rctbwExTwJIZW2Pcmfy1d0seoKF0tz11e6cc2Zy6VeuQCNODlpI47YRNVDbSzXc/
YN69tXDulNrKfk+tn7EVYmd2N6+ApwE4P1P6KlGM9bqH4az0JepWa+lHCZfm8Hxayrin7NJDaC8b
P1uYXs68Da5OfYfmp/IQGo5aRC+8TCYDSk3SblyB1BWelS+ZJ2DheJNGzPWD6fVFEU+OucxVBnla
AhiJr5UEmP8QLEGIB7GzXzB6M+SWlndFVyCyMdE2A1iMs70IB26iMuvrVVp9wnlpBuDmeTTAZh/6
3vvYmVgJWwEZQbjmLCF/5wFpp8UXkt3WxEJoY4p8m8ZUoClpMJgME7pLj+W6kZOOOahRst8ldIJT
RPmQ7Ff9ZRYQVA4a/vhWK4+adzzw8+V6jsOtw3kWSJyLU+OA4NrbijVzSmq39ZE96jtiHBaDptwr
ieiiOOc738HCkY0VLZzNIYXow/eNkf+2JvSkVbELwlhz+zhZ/T+f+nZK0c6kwPtnbegVfd7S0es3
uunPgD53MwsvURH+OFYq2+LDv1xb6gkI0AV3DLRu0AFVHwwTaN5swCiI+IDwLMuCoBMv8cdCAuts
+CPEkP9DBqidLVakNtNXF4urVHHcSUeIYCEz4m1p0It6PzBrKMi6m57Lpw3Okae3sTcO8pAhg0wT
nZpiNc40iI9SCBRu8EYrVS4qhRrjqRyrxsgI0VS0qsiTfjibxMG67b47FGKp/uwVi/L/oDqBm1SE
ROfWRH7JugyDzdu5Fmlbe17vrBX8lAyWRVaS+v0HeXV0pRBW8pEjm9qlG9T6R3+6qurg+DDPezX5
ASqVmpsNGap3o6tfRvCMIU76RlKRpQtHH6bgNrdXQZ0GdSs9gMyt3YnEvU0VvMih9THRBc2tI3Ye
o1agSlO4IuBUVr+hhPbC79lRi+L0zpXuyBH9KXuHTXVhIEMehePmlklA7jT8+sC69UaFZjFifHjh
w8VUxQy9vuPhw9hIBXVZthAZ+/wYeC5ctZLOqaz07nDpg8XADGwjlQMbEpb95rUoWNdz7z1hdA/3
CfOMaakK+OLPyfF4T0DD8sW53XCg7EHkIK2KSKuo88b4qIs4uqYdb/V6ofdvB3XjZaxMQ39J9jsf
ic7HFNxH1Ko7PfrYZKgSrOqQLdoeVjBE+0Kyyp7GMZTiMCknXy2d0JOcF7KofLqK7/OlXJEUm6JX
oSoDhsH666jIwA8Gwwfj62AKXoXp85eF75xpXIQvGOIaXXTefLuKVX0ABN55GAyxxe3gWuQmThWQ
ARsyeFeS9PXLJpVwXh4eEDAYFf2R48CjiMxbojEGl4bIju2F388EB3jAjQC56ERaRqF3qKF68FpO
Kd0B0Lki3jMtlVZzH4+zWK4iVWBSGrwUZ6zf+4IUAlvBT0ylLO6AvHMijMrnoSl8qZXXJ5eOImTx
cD+HFh4xOG4eQe+lT3RSGbswSPKHuZpdqIkOUcsQjMZohd9TdZM5pQIhRL4tdmsGBKvBXyXgRW9c
8+XWLlCXAMjCqzq5QyBL5oEim5kWBsKZ/mxrYaNBZLtry3xC95mi0Ai2gJqIDV1rB5cQQPMcsIN0
8JW2EZugAiQ8F8lRQ/0B903CnDjebYvxsOuS1PtnmNT7zXe7qrzbO70rOfZiZQ3KxoGjzwSgARGc
u6hz/kfJJu4enu8F+CK0oFVErZ63GdyRn5Ouxdu6TkXDXFr24oNu25v/WFgwchRpD1/V4K5Ug0zy
BPNcGGHaq3eLr0JTgx9a60+m1weGtzpi3VC0iD2wwa8DVLQClKBnye2/VH8xO42z/Sku+IwRWFG5
4M9iouQWDzK9GnBzvKqM8iv2czOqgO8rlSH8TLJ0zlgzMdgc0OqSCiHEyKpny/6IjTUiq6NzxqFE
TBC0LlMjdM/r60FFMitYfLtJTAxm0RHHSWMijyxT58glijcath225fonylqS1/QfSLogy6W6q2k9
ql0NyhCsCH97cKSfM9c93VqWBRRMVxXdvqS7irE+Is0eBk5zZPFY4ZizePzG1Kg/nWlpYnH8GWGO
oGCroRUn15K/YoI+iPevAc1UO7ZS0BXLfQ7KkN2F4oGX4sqIWOoL0noScnyYKxCeueEyt9Vuzxzr
oUn0cFsRVP7i65r56SzCCGPEAteCpG/DFXWHHe1Tm8baho8MbFFpit6kOb1i53Wu5r0gQmJwF+QB
Bu6q9ef1b+XxCy/0HucpjxeseT6i+LHIilw9dcQQeXHQkUGx/6DfZG+z7h/CLMNzBdgRqrztIC7S
N28ZT6gdQ0IctxyqRWhAIlK2sosbmwkl6KZkq/bvTJLcGnTdY8bnQzqAdT20iY6EZlVtjXVcrr/M
zbW8tjEmeVef64oPdyxaj/kb7DkCfYXiXX5z4rsNli+DLrhlV4hz6LfDESQaI5sMj/n5mjpehrdF
9QS0D4OYTO4u43ArRv3cd5xi6RvoSLQmbI93FvCkV09vFDEzLNccPkhABuDH1VNf+SOCv2LYb+j3
U3932DAzYBvrd2oxtCEA8hwh3y3Te/tZVfrJfxM5vCelUuVlLzZHCru+AgUdSEWF1a34MIW+zFRX
/Y6Tj21sm82cZtwfrGVg60nVvxmPPUKt7BhImmxLW3I6054DdPl7MXd+Gm0D1paifhQOphMNTtvH
QURI5foZsWflepXN0dnXqIrV5mUHCitNw0mETRvEjV2ZDfAUYMn81PPleVzhCQBvirj/XeJ+lUO/
SnTpP/LoxgLoValLGjwzBD+gLSHwG113AjTU6oQdfEQ0lTVBIofv6jMq/3HVxu2DrLbcrC0fU6bn
sxxaQotjJjIgYLX6u+UV66ag+xvQUl08sAajdXK/MdpId17uic5zJI1hLkx/XEYpXhK6Co8mPy9U
uxskCw//jadA34Xa6AWfKv4m7YooEtN6x/C0BfBPbT4HWHfAMcilGSVfuRvZc77T7x99juw5l/Yv
d8jiLIN0EqNgR3NZ5vrzg6zwuM34G19S7d15jUtZE/X7TOQxuUwr7gK+l+VWz+YVZexWCjg8p/kj
Rs68RNBoiEAoWCxfEy4MDjinY7VAX4+RyUvIxL7CIu83QdykvUakkuys/ZM1r+SvcrHKAN5HR+st
PhfyV4hNk14XAi6FksYzxIqu83hKAcJN3p3DDu475phqN0wzWQQ2S8kpkXvs8dcojM6BObK96WT7
SQO1z/wWNgeP7rlFDze/Ogto1mfpZ4Z9e0tKz/W/8cdRxOzOTf2njp/VD6W620QEDoh/75Flr3QP
AHGKqGOiV7Z+CJ+DWIRk3EfVP37TwvGn92HqFbGB0omekePUzfRr7RHcuCi6OfmKkCYYqABtbh12
CkEsgp5Em8VWoddcwZvrY3v5R1o+QTyv691FbLjkjVrduhQl15NB5kWOuy6daePbQJ/TAHEkZcSJ
jR7mI2CZT2qrzKbRyU+PVCV7CvyhhvCOzQ2qQX5wBCtu8UHss5t8ouLmXOZWzebMR/TuGVm9QDtl
lwEVhr0VSilYO4n7o4+UdQuqc/ifWky8nOgHHXeKQxn2tlnSh87dAX4tqIjgyatR4WITiJVmX87n
1EJBqpckNB7tweMBFwnob+dsaUFBs76wIq9oSe/HpF22BXDUK9XkZk7GRhBeFQAKclBOI1b0+hTg
bjGb26Aai0/wabDwH5YUXkv+K+cpCPeddsAi9D8Cpb1+zo9J5/CabYf5iE0hiQM3ZtAPYE79zieU
v70WMqwdxobrgD51N7M4LCO+uTonCp1l8XYITkqkvSZG7d4mMFIS4fQcbGDPIyPt8hLbSqC/uCrO
VYGQ7l+VFxunN4Tma/V/SLDopbkoSXGCxKxMA4F2gRaxkc62tPSK7aESnzkcjjUofTRI8U7AxV87
5+ct3Dx4GxrZwt5y7jHsRr4DL1sUGSHWP7hxCZ8RR7wRBlNndymsmbsq7MF+K1PxONHtHY0/BgTW
c3jEJR3teFFCsGIzaXiarkQhQXjljCagFU/2tA8uXrMVBuBXWlc+Hd9XLmd3xG4n86Q3q36X9wn1
Be2S0PRGbcVX0n0fXG+2s2dWcs7mvMVCRSD9wwGF2jpaJQyrbZVhehewaU7WpHodNPD/g0O5Vl+Y
rNoTFNMGsDSrPvCbeqMnBqlXDvg3V/MBKI+S4EOd3BcEKJnlcRwf1q0nIssDxFSnBcZh18cRrZYd
ybqnJMOFU7oezck3+xFH6TXPzqKBi+6j4M9REQVar17OvRag8WpUQwyYArWlIMLCaSZXtybkEG5G
vHWKY/pf3Osg9E0DxYpgp56gJcxqpQ9ldLchJv1YCbbgbxMpIjoSLUs3NIZ7D3UaUYLjNwuYsU+A
H0/r1F/Mr8oaB4YS6KCyU/cHKuS8R/6bN7C13pe2zJzSEralGZ4uUljg3vmk7+Q+nZZvlzQwfsXB
rqs0DH10PkHk80Wv/NFVlX/ouSdwbKwKn5WanavNK5n9qvrm2r2Ula/OCpa4iIFv99+XJ5X5xa7/
e3KvikSBr1MYsu3iPd4OLMxDFuDLzeiUsckkk3/XgIM+fYWalaUEHtGV73pq8j2JFpA6IH7rklpE
+K2rDYa29+P+HOE5JhepgSwgqq9sedruQ3hWJkMPk1SgjyBp1dGeTPOaMQnRGSf07H6jJHksb0Zi
BcStDh+SsKJeAsnBNVb0kiu7SKgm454S3xjGjPx28H7q6WUrAecFcTb6TI3ZImG+odU9h344eG7t
BT7TgJ8SnT8pNA9SMnIH+0NEDQK2p7HE5el2V9nhOQGBrv7zrk4j5PmftSN8pxfKAedGE/+LPwtf
zozemH0k5IIS8KMP50FgicRBJakGruuKCp94nUV63phAkUcRMVCcUgRnzSMpCuAT72Lv+aYChX0J
Sve2Oc+KA/89l+rkEKoewjnalBFJ3k/h5E8j3qbHYTz6gthIFjhT2DzvpSNk7uN9OyYTiZrqKZoh
bAJIWzIzKDn7rg0iNCa2Uj0uUq/b1hn5fFFvbX7NrlJ6Wdr0YMOOeWGMvNZf0c9m7S4KHljF8gdz
/JNM/wfISXzSgYJrTnAhGkiiH3ewOi7BVrN+jUvBQ5CsBe0RTxra+5RSMgTHCg4qS5qCRT77roqY
w7aPa7kEgOK9UMDaPD7GcqjYZe+aN3kDu3FrdftBJFu+3vsKXjVyRmOVwRSJpTPLdv+qEB3FTxFm
aOk40I2LvwWWSXhQdFFEsyuUYyp2NwMcWMaTc/GWjVNeNZR6Z705j+6y5qnDYjYmh6GkUzxylcjP
GsTUMaWiseYfC5iG//p/EmyE24K2BnNo8Ir5rOSPsHXWozo3oHVIkZr3u/Yla7aeEib2xHOit8gY
sXcSOU69Wraf5jwimNulOE/zYSnSMndmuWtl5QhT5P6LEI2blQxTjokMteGBOE9fUPtjOW01/byr
UYkienCy+pGuL/8yHCtyzoHpCWlKbUkwZcB9ZrLD7oOC1QuiqnPc4uU81ZSE8qqqwL1C+RoMsgYf
gmXI3zp1U59rDq1NMNOzKIwfvE0ZKY5ancxG8qEOuc3Pq/rlV/v3GtJDSQgGJcnACyHMQYXloVqg
HX6m9MR9sZmdQIg4ZSDFgC7tp2vEsoMMW/Q4YwkReyYJEi+bmF5pmQdsT76VITYztRpoQYe0dcfW
JBLV4r7mY2FRPRg/1oZDxYs5vp29m0AQBUKrQayG9aJg/uMXkNW9wnI12so36xYA7fKDQFUPjX5A
xTjMuoVFEArMADqnzsQuGtX36lOtcZ9enjTLxKhHR80cCZLzQ80bpuTLA1VKDm/t0+3v1c+IaIgq
aLwsFPo/s4Ly7pD11hAad++Mu2rsrWTQxQQ4o98wwJntNjxB/lZBMC32nHPmQ76qh9/81mpOauKn
uidOvTqZV5K+/vKSkEcP271DkGNz7LB7SW0OeWgoeWFVB1+oyyTdZDwlwbMzfNtUsfHSJqxsIYH4
Utx8KulG/3xxyr8E4v30QX3sP6sb8aBMCyHLJxbV83wC75/0XIoZaziCC5Uz907pQU+PMPx9uMh1
8ueaCJ/g097v0N/hCHZRd6Ln6F8gxiSocSqlGYjKlQPoZBJtWUvFk2YAoFwSvVQm+Gv5rZNgigQI
vupH3MzbhnuzdmZ3t8OaRldDYxHUaBNJTlaMj7dRc38P9mNOZTfeKW0QcVVsSO76y4ShE2nQpvP+
rZ4AZQpv9t5cuAdAHVWI6qEQevqfuBmfDPXz6nXuOlk0p22ILDpbfCHLdjsdySWfo46/PSlwL7U6
Ls/h2/yz06c22XoS34cPFZsJCfMwKQAxzIfZ5I/0gvGy7RglUXh0e7j6AGCqquDRUxhOOVqtfvCi
xlZ3UY0DQGP7JuVJNKRiFRsBOdAgtmHapvFpOn27YeSj5bFQjjYEqjGH+sUOaR21+z7g1boYbma2
eJErCP0GyM+MOpbm37SYlJecmuC17QbCaR4Bkg4ueN5SB2eDLM8rZWkFbEiF2HX7v0dHj6ljqCdl
z8klmnSP9yxVSqW6UOgxHqYhm2QKzqQ+/wnOfkLjVQRteV4BJpoFBJbeiMzXC3h+w8qi8CgPJjbL
99Ep12nQdt3uZrc1LKXFlmUc+IWYwd9b4bIVKdgSbKEyFa+Xz1uqU3LPYeCoerc+YYzZbdWD8gTc
Y/tXenZb/Ypxts9GxgTDjcqxGIMSsOjqShgMyquwsm6MAUL6OKa18g//icJW4bMMWpgO89WCBNE9
60e6kzSprt7lhzDjejZXxpX6XY+sM/cyvhhXUNGWbl4OaJzlmIFZ8ChPhuRkfgJnpLppDGFfdW6b
rVAEwX+rL0axfNB+AhOGZOBClCmEqpPX8ZdDtKHma1p6avdy/CE+u8v8XMXv7E+1T5T7RUBm+Ya8
W8X2pal5xsSRrIKBQhrUtzbpSrzUt+sJ9zNkycZnjqtQMjnTqGfwJVx/HTNtDf2yZHGTdBv5aiQW
UGQr5HU9LniUSOsHT6c0AUvKI6sZRtSlnr5rE7dzkJXdRF69BszRPor1iws/0ZzKnbU3EpK9z/LL
zF+kmCQDSmIkeVR8Jm1WgmIi3mHCJ6+ON2mkirro/pGfsPFPZhid8BRdFKnNydELy50lqN4ahUzP
zeQ2jhFRqdn9305Fd2ffAqQt7Hp+coc1/sWFE1rPpAzLxMDeucwoOcS6bljBCfRcy7oOFRDdwNPN
SGbbz5fM3PfKNruKOnJ3TITI1TlEIykdSAgAXHc3mS4FQnNzBthOS8XXjlKG4iqfh2UPAzAfK3VF
r7wuGL6aYQOWW/W24HJOwsmTmRBM+DbZ6R68PGEFLeUrVLIULwLHvUWqyfaSqopKpIrv4WwhXa0H
b9P+sD6joYVcwcMxkl0EBeo5dq527Pa/Ih82z/nDO9FHhg2N8DqBjphJXGaHcpPJldnG6YsITvDY
5cC0KAWpvSJHeliIsN/puDxBiM1YcIqV+i+vhY9T5cE9L90uqvpiS8Al6Xpj9o2J/BWAJjNrLePx
dvOQoEfUy3QHlMYGxiMel6ZRblF8bYtNLRI5Qsjl887je2gZgv/Gs6QT06KNDnKmAoH52uLo2Gkz
0RvvzZRHW9Hui2gAbyKJUaeI9rj4Uk8AgGvtpWF2GnzogJvmtLOs8iIUfNJ6zendM0Ir4fE20HSb
yPCw33+QUxkLdbnO+S8+u53P44A1bbKpFHjUBzpI7fd56UmoCvhdYopOnXq5U04Q8uTg7TbgO0Qw
gT614u/e1eVd0ZQW78YXv/EQYPW8KKocwrSD7PSlj9lJkDzUmAGNTloSoyCczFqZTtu1HKix9R0b
onTS1JMhJ2PTsyzq
`protect end_protected
