-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rsAmhwWUQYj1vctr6gtbdQZ17DBfxodlNYuFSPH4+OnCjlwT6jnLcZKGJfPchM+++z9f8ll2+uxX
MOw+TXUoGTonDRnPcz+0DBLpoTMrTDQkr17SEcsr6F+Uv8HaxXqL3sizBj4EwLplw2SLD0bmPqI1
dEVCLsPx+vGeROdeTlfDKRZaX3cB6nRGya+Bic2h9wUQ+Bju8jXXmUUcG7prIy+YipjB2Lqc6Tuk
pAinTPOVobsWKr2JBaf96KQftQk519VCC1lydSB05GzNhuYaoHErlSvWg7kkfrixybU911qHgyLT
zysn90EC3vMjpRTLOMlhTEh2RsDfigiulDMjrQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11968)
`protect data_block
6OrzAknjjb+iCSUzOxWQgKIBmmYvDp2ACuI2Kr6YMS14g41tq+rRdmJ4nkISV9fSvRhw+f+G774F
S2No1vfb6/7aic6Vw2QtBPF/DPbdAob/Wl8CC07BZU99NZm3DUHL61lsy2cmzU90Xr2L7w4/b0NX
u2IyFEufU1z17JBCnZfTu9IRE4CqufIJgqNBn3+P4FFtn2SF+CyA4bqecYRLBB1j37zc6iSdQiK7
LkrRUUWseT33e6c5kr/7DfYjkJVyfdYZ98euxdP734Y3Sq33fBDCT1ZBvkZOE3SIPQuN/k1xq2mQ
2hOMcmLmbNOqeY8zutG11goAoFdMXVBaX5Flz+AOOfODWmS5QuIFRGkENovU37c99AtudDaV6ETE
6JzoEw8kbt4d/AZUSXzAb198Lpr2SZ+w9Gt/Wke6fDul6Zv7G/ou79LI4yqeFtdNk8JS2dsccKZi
qZrYLbUy3qLL0c79kRPomICbZZybZLyEFECmppdlMnjM4Yc04MWA+T6u7+VJTgV4ZPvLtVzapiDK
sKE9mfjX7ZG97MakmcLcfVHpnVu3RiK0pAMETNKQnlrBVJbK28r+k5IaCPhgPN0yU6hOHx6kL/S3
iYKnmWFhY1bzPgiAp1tttyYxLvTnfy4I+EwQWuZG0y0yaUrEb6J544BtbW0xsJIOL54RTpgYWiFo
Ahec2xyOe2yUn7E87QmPKHuwN1hXIKRRmtDECW5IWWR1UuRRHdlkwO0H1QLs7M4Wc38iZY/jHttN
p1OZ+0gjc92hDvnd6yoiKW6WvPKG01lQby+O0bHGEsxTPNCYvzdtD41TRCrQif5RVy2JpesL5eC5
m1QaSu49DaF0eLcTTPYPkjiUKLFKJPIxLAJK1LI397CxjMTCuOa5LAh8hcIAepDQoBP3z1MnwKdq
oyVkBC4eDdrdQC3gUXrJQrFYQF4ts0sVlp1Nk/dscDBoex3A58lE4Ri76Rie8fW3fSBesrLqZmcX
lBzbC99WkXrM16kkfyuXGWZrxP96F4LLYoBl/OSDCEHs3LqPb1Yvs7ncBINT7qJVVuG0PYonuQ6m
M3nCfGl8EguMegdu9rfq9gcOHcWDlbydNsnj6wOOqEUYOvGfs8YyXEmn/6uq/8Ow63J1/zOAfxAG
0VKfnjCSr0FC0EqUl139OFDI6YFbCTvctnJM1r+sguhnYjLsO8en5jLJsC0BfmKqG3Z7jM0OJUXr
Ru4Os83d77+JB7imH94onEuEUOjAR9QLNmgCf4HQ0ZXoC4tClYMZvYqBlnXjxk28rbQg+COF9w1S
e61niPR7S6Fsj81HibrB8tOUrm+2uplJDtLTuIZ8tkOGomCiZZbT+4KryINwujwfztfokN1TgSX8
bVLP7grF03Bl9VgpKdW/tFttP9TfHkYNYhadddmtD3BpWF8zz4+zDbH+IP3Scu+7pV5DQCkKtPyo
KQKrajo529RnCObrDF+YGfNZfDP3XUusiGjvV6JiqNQb6ZuAg33VjzmdEDN+r09RdsneCLKFYCZ7
8lRASnkPUXVpFnbVMDOQYGPuwzwr/NTzZtZ+s+zWm8uZ0GdyClrOpicp8zqcikaKcesNZ/5EoIFJ
aorDS2WM+X9jbj6vcvujGa3nnV21JWLrkJ1NPquKjjznJkanRcn9ppAAAdugB4bjiINdz/tAswG6
3Z8DN/CwvnFzpk3bUWbE8VhLNYmzLvqbJta8B+/HUlfYisRcz7M5HNegXZzMvjXB+BZOFhfvPsqj
w6HgdOV5dNgo8ecJXKtDeF/ni8gdRhqwPICIE4Q7fdsSjhc97u1EZKrbn0pdLCUF2y3DcoNJ3efH
GP4b939FmAsbUVyvur+h8rN7ox3dVA0zmbFazpRPLP/tWeBxAjSR68n8IvRH/dQhbB5ZOamZC6/K
w/E26cXYsCS94HEDPm2BQ6aIeTcYI/vyItqPzJwtDZ9XrQ4EOT8PxlAc5CzEq30gB+/laTg/vUv4
Hu4zObo0QR8faCmL5BUaVQPJw/GUTbIHtDOMgvAsi7lBxbubu8TOczIM8q4lhOfhluHeZ4GPJwI2
fSfZ0Hg8QAV6z2CLLFq4DF/KAjhxYEnxhE2YeurmEB+Cec0eIfMAOZhppQX+sPZqGkWoG84hAonZ
NayfJW1RzWegreGeI44WoqKAYLKKZcwH+iaFJ8yj0PBofuawlLUC46LCkF6ICujZwdFZdtR55UJT
VgTUZviCWw2V9hQYECU2csmgyU5e2MSCknfEDrFc0CAtR6IJ05/mIH9qZwooLLv3kW8cr3sH5S46
q/ShHc6F2jusrzk6rXQPvFRsvjs74+I4CEX0jzeKTLWHFSN1GQ+4B2/Nwp+GJFSFUAaeFG90+BUN
V+4LpxIAY4E0TSrdtJGhfI6qVEtkJiuNenSITxfXzZU4L8boPCjpLZTkKdFMuMatMhhLBBcymT1a
IBzcYv+j9n3Qk/Xug0xDyOxeNF3cIIHm66BWCSpxC1gJ4R6VqBLwmAS9ImjoZJqysPTYcpHqwJ9L
MjCsImbUexsFYTx8GMXfUDe+h/SFN0hno9okRVXDYlggrKzQLDcsAIhWMpA+WEtwHRBopjDMirsR
4fxLbSH7ffpQPz0XHTfrElzBvdOBgAZP1/FD8ay7bpVUCGf1m37SHHAllLP4q8v/dQz9LmE5H6iO
4rV6jiLoJs9Yph6xnuORUKmZYIRahOa9bhQb2ish+4aPiGeadkCA+N4JsogUGcPnPbDHuq/IRemy
inYQB91jhULaMVQRIda0eyGetdOi/s5PMLYYfUpdeNkgY9Hhgmvu2NpY43YqSlcA8XL0BoxOxAKN
U3tmDjbhlHT/c8jWj9/PA+DiolUBqvGmxc1/7jBZqOpAbbZ6cZRfYTwtQhwakmdDiXQVgVnoWa8G
wTmTpSlgAnQ72TMG84OA3cu6edqII6LQZYvHiVMGYPJZ+SJzsz+zbbuPqDJNqls7K8PDW5KluNVr
OHRo55YqGw3yM90jTwroGtux+LvkMyk062dr0MR1tYI5eEX2IB8Wyo8TYT6esatPolbijqOiAkFL
EJQJJ7cxXA1HjySv0Iwb/ZT2u00p/lmfLf1njYFJHxeQITZRi3Z2n2OG2/wH31Ush3XpUOkTQA/N
7TKnq/B58YCaE7CFxDpJHlUTQRYviNnlvprN8dyJteT/qYBxtUaU9io1JSZwViuDYEsY03wbIDCj
HB0MQBRsCflPJPsx+uKtcPIq+8sZWXmiHksXbNmZFUF3m3xJqI2xdtbKcmKtiH3BSDZQtX6emGhl
8gyBCQZ4odg1LeXfP41Tb85aiDzbrBZkLzPUdLedpqwQ81xQfili8cmmf+tVMlcTkqFwpR7ZBNBi
5Zrua156Gl4asttXbeJIShyQBCek0buekexDo6MThyN3J2ZADklkjTAfDT2ZTMPrfLKAzlLJB0CY
+CaZDekYxiL6UasH/eQO1XPZwLuWgC3YhvjudLt62JU8iGT9m2fzmW7saXa69x6MYbTBUQbYbzlk
owbV6wygBSzU59XcDWtnUChLAw3PP0x6T2RU/BP0esgVgGrlH0Dm5heoH6+zXrgkFWvhy2K164v6
t6fGqeQEr5zPuraLsEwTQ0HmHPNyJ+K2UPBFyc7NyOVBVDeYuPEnD0I+ZD/gJzVouEklP3KnGKHK
eL/7K+BQKprzkUWb4k6t9FZahdsG4d4dAjBeMi6HfRMkGvY/xHWYHlQllh6T0w9kGVTdLnsKk3qV
JKHQgjyCcKViwmXQgx+/U5LXR/FnoMHOKPnpPOUvXl8kX/hgVTdrtWtla8tcYcQ0j+bB2jhkTfiO
2cxTEfZOMUFlc0rsfo9A7+PsBdrnyDT7KNJDE4TwaoOuf5rTMVndkS1L3lLTbHCoy/atS4Ojs3SG
LSNx+GTA7xeaiqFd4p3Hq+j4IDlVGuVvgDw92psCfcxjDLP+ykVILYI09H5orbRgmhKhN6PrM7yB
9TSFlYdnBYJvScDzRnhLuOBWi+mC/Z76jJw4F9aWCoBExvqJMb+ksY3E9HB94NhyNCfLhE6r8PMK
luh4crk475eqnbmlbZLbI0OKr/FTbY2Fv8M2WQL7a5WfyDC7OmRlJFoHbd8irIN3RPKsIRmJII+S
MQpEIb9Pqtc41E3kFpz8/0t/pdafAVeuberY36yAj4edJ4B4pU4lzNiqf4nfT008o9bAZhJpWj+6
QHZOwOnx9rLWPEMlrI4k7Rb6IWY0/lCLpJfWel4py78uhjujsj7hJSEmTu8jCHs7n9qZoEFdWpWY
TyFcrITdc+ucf+/UVVUiGkE8diiAYrTf8Gvotoc4wpN/3kIN5mK9ekhNGzmQaYO3yXEe7WEp8jev
MHPwZKs9KmwxGFNLnnSMGSiYFfccrG2NW58aTUxi2FAUM9YPvDUkdM++/cS3PmRy7SJdEHQEUdkg
SfTu7sL3wStfUvoISF4fLyOHR7cVtM15AbiF8icj7zZXskIGJKJE9KLkU5+C+XOTcQgO4nV0yIuj
9v6vL/xFCDg4BaYoFOK55/4eWTpkafagVz3yb3H64Bun6EvVN2pcyooL2NhkfLQp8NUqYYFT1Wse
clEXKh2EEtfRfJHuf6XpFZHQnQStJ4Y7FQZQulJCtTNJFhAnoqMXfoSsRo1lTb6Q46HsgO3WrH5f
zUjxrfj97nCK/0bDV9Myg1Ffc9bEmBsqsw++Bq7MNQt95cjTgIm735ds6TiDQOM06wRW6GtY/+7c
UfNp2ypiBwBqZ8DztpGVHZ0BaMXq+MDWsRQZOUZ8WiLq2a9XnlmyouKTQPU9e8ZLUrnFDfaoan6e
p8VUaqg5A9EMOYKzNXNd7PdGZ1JtHMz2zAH+CCv5oIyVlaEVakK2plXy0N6JBCbw9OBvYYwDpLcQ
CIsKik09PniE/F0Z9mTfy+QURTZQoVXRvcJFPcC4I9aR2zKy4sdaNUsM5xc3zmg1popH/QtWawJ3
0/noAva7kpkIRpJuSfdiqBbEaEy6R8nP3vieRKIoTlb+Ipi6+ILeE7WGZ0+5TbG75WeriFJvVZcy
yebOe6bkIy8rdMJrbUB60fKFLbK7RY2xbQh7L4wSV5ZxJehSvH504KK5tuM4N3FQ9qUNOE9KYtKQ
MWbPHpM6SqTGHXhmjkM4kMRHhhCmcrVD4iLBYG1yz4aLT9I16+8fBCvmNseq0fC7SN64aeRjoLm5
6SP+K544pPSvhaRjWsaOYUGLSabdSTeJETYv9qYO3t0u6cJe1x4EzHTAeEHcUJCL6iDviCQuad4K
J/6l8lVogxFnP7B2l8chwe9YO5hkF1PUiGfQ7lnefl3AzMUNPIGEZupgyDrNSCf08E+x+C4kQvTJ
6+tlAItz5JpMA1ckjLoGTySgKTkd9yMhH4xKVnYgWkrQPq+OjVUlYOxxia104uRREX/cGzxjVClU
+HbYguXND+B6iZFPXlEw8zR5ue5PZBcTwn0InfKZol1WfVDGMxpOE9bX1sMDGCzgMOWwmL00pygE
c9/dHXaD2vRfp7zomrK+RbJauEaCRl0g2l5RBMcixDgoEZbbD+Swa7SHCJADCb8pG2oaLybeWOrb
9BjIyLQVOXtiUmtcGrh+d8TVfAW7VoI61dkdXIWC7+dvXc02BQnZAQOJBYWhI/D855k14zSgs2Im
L26RxjHBcmZvYSjGn/e8tYNDe+PLFmREodqTdDrgqYbveaLSNPCHoE9t5p19sde4W4RVN6GKnKpi
Yek/HvkfvLHTU3OtDmxcmsauSFDxoSIixy3tnpfvDvBpZA5uGIGHjK5D710DQYmX+lImnOEuy6lC
aCamioTjaN7agZ6Ba/NsazYUSqDE9c/SyOgQUpvAqKCsOtswS9bIN2ZsvIFnG70XxHWQ27gGNrmz
d6Y4e/aBsrvDy5aKH0UmIyFNUET1iZmPKv9u6a0zPkYAxLD+w/Q7K+OvNDUA1yXO+B99rMb3yO91
7BG/HIYB/mcXU/JsmBviz9cdvtVqZp/WEHLhqdnaIzMtwObJgyA8X39mPj2e/mwvopwV80/NG/QH
csZM3nMNYsd/SsGQrbxTVTjV/1EUI/u55TV0zG0qiRHcy/yMH7ypj99opiYYtGzU6UZ2buK5D+Ca
jduL01u88+sVVcHhmEuUTsb8HhCP1Wox01ix1EMgxukmc8RHZsYRVUZVecYihEaBMgMoWjEtBxN9
P7kZ0DayILZh4Q4oBjmAcQohNDHjpnjww4G06bATqFEKlVDbasmPkHnvRR/JFdiLowC0cNdxmW7V
XcpX0/g7YNE7hPQfzcUiOrUWVJtsM6vvra23NutKinKceDpbFP6UZAmi730wdfPBFiz/CNwSJ08F
gzUV5CFnwtNZKlZgo+KpOlsaIB21b6GnvY2e0oRgtWI/nxkSUN96YdtO1qJqs1FKfE7jXM8V69y+
aBLytON9HSSFBSrdJmVVTMGFdm8KI8xurBwZpCec1xECw90OGmnkQhPYywiNnrBw8hc2i/I9Cug9
UEKQAhbgX4GzvcK/VqfsLoRN5kC6P444yHr2aiveL/f8U3ic2ieb4cwBqqPxo21Hvw7I4RDL7CxW
It8QG1BEl/Yh9W36TOrYGLkhFUE4WCUkhdq1Zh5p9StnR39An1QDub1LtYZWLKyEozZfmi6VXmab
bqoCmKwzogkBINqUv60NzlQRiH5QrY/C98oNHxVAHRkG8Kon7wH+4Qr/q6GxQLLbJeRGoKukq8Qf
s/I2gLY/Lchu336/0UQiVCM2lcrPmlwWay865zYB5xTDXTz9C1GeG/Io7CUgxt/5K03IxMzcxu72
1HZMLasfwus9tw+28JV973Nfe02kUWeJfW3/5/AsV7KwR77R/9GEENfiqtpXr/JNeIknGzbICN0D
RevlhjO40ty0KaYufGd93+YrcL1d01WZfjgqejqVSZtFgKqsTqFRKf6hClyPtVZDu+KlLdc14Ouq
JkGne96Ps3GEgs4dmTWcN6Y7y7uPoyqoomR7Z092H9x3f24OLvEy/fkWPvNR47g+6F/OzbWPeGLS
Mfq2pT84JBwIxhWDIVjHSYb8ncFbqsOn9uIwVJntQdmqmySvs+I2X472fus/2JFIoUDuUIZet76V
biDYFMBHc9+mb0JrJkSZH/kggjDAdDADEDi85E0KqCZWM016KdBTqDXfTjPGD9k0IMGlifLvd5AP
mhRvhYreGHEiO5i9ZIut1V9c5bk8/zNkBDAhAJkUsoRiMgGbRPLzzxG2u0F6llo1HsfevW7c55WE
/fxjeu8qmnA15vmI5dlzAPs/m3oqsDxMS+6eQneQPev8WlrUDYj4/1hozyTp8JgUr5QTZxhhY1nX
DiQgyXhp4MnHwpAQvBt3FXdaQcwtwVRAb3RkqSSZWa6/RZY3iasFshgpdYbHpHzJI7GTVYODE0o3
2g7oo3ky8I6TkvlpJGtHZsHZLD5J6p0mfDt+Nv7ap0NtVc4cLFHNV5b2Ec9NtO7ZlfVOT4iBdjdb
DJASpDg6rYhPETli4TqgiHcJE02CIdK16Ik1g9suBh2MCiIwg0jcD5LeEpx89ZReqejh9aa9bbiA
w2tnay+BIe1Ym/hxxMpw9C1d01THvMtmvQIuUBuiYtozCKa53zNlBHbHGkvs9THdQ3HSVs1ZzpeN
oFTiAKi348cc9HuQp0DHHqg1AOnWPylAXZykduucJM1/5+cEzeEGlq88MycmvlWLGrXIcqP154sR
OdLmoyzBMe43HsUq7LXkBTmrHlY7sMQULrrqqizjQe9kHWjTG6eErncMXF4oP5G1+I3E/jvs++IN
ee0vXpLmpOevo2xbJMU4J4nsF9tB656fTu/b/7HjWyqJJT2Yix6Lij9TPShKLX0OtGvZiWUM6WtD
PE549eK89ODjm0/XumgBVDEyutzy1COz8riOywhKKtxKQQds4wqFpPUQF9fufhcu/UFNgcBeM9Hg
062QWiyEnNv77mU8Goa29vusItIS9xmoZUUhY0eNEE2lnhwEppUq7fEpjCEHpM89q7Iy+BjBp9Vy
qePN96ivUWn1IjJC21siRTr1VsLXokIMJfCjQkVO/Xg6jqneSUECreBM2K2NZAX+ghUEfXs0pXG9
VphunRiprvDraQMIhYLYkfkNLlDVUdqsrk4qZA4WTOiVuMm2FNgK3a88o9MzYWVvdjx89GQzkSyU
8IcawIaDddPNPUSUjJ5AhNuu/2PoEvN4HakdeBxYdpMHD28xluEjyToMVQ5+EoUib2SmEHhrRCsM
Bo7asgiKnYTecToeyb6qF9STRj/NHXw0rsJY483RvUPNfwQFKY6dEQbgDXid4HGw4V5AwHNait5F
iQOlRtjlKHPzbyf4O9/caOTeYGBu1zD+5KGlBdRhdvZUeige86uHTZ/Lfg+7fgyOyfEUOLLgaX86
fGn2iLC1cTetmIsYg62LDeEPKCzwkT5SltM92kPUh1CfNssiRfhDSqQUd8OHNjbFJT9cJuXA/Y5M
zbZuwnMnOLyctEaPru7DfyKxttof6YrUKLd4HyeTd9oAmClXJF+P6CEFqNZiU/zlrAued4p9nUjy
fE+oB5WchK2i4yc6yHd5Tm6InYo1Wd5EYdU/Q27INuGSg11iT28po5fTongkYIgV3e0558wxwJM9
8+vBxmDtCr/FlASj/11R6ED2t24pIzyfdEEntiws63gjzTpHn4uHZPWyZpptevCleEtZ6Cq0ASCZ
o6kN0UQMpuwM7mgQwqLTA0Bt0N95nkz6OBLRYtZ1lDxmmD15Qatqp14YpirA82O9wvAfkccCsxgv
YBJHCb4Y5XYOTlOWP5qyaH/v8u1Ob28NwMXwzxBXtEh+VORzSg3HnetHq4Dhhz/zqv0NJkJxywtM
SzsGBjfXteeJZee5i5Rln/x288DMibUAqWmfTJdk8WB6es0lmvUGwz8C4khRA13lLduBk43CvVft
M6TF0CHo2i4D8zZeNkeWmxsqCUMwQl1cRilaKRkDnxWmjlzCBwNxj3WnbEjTnAJ88HEh74CyAjFt
XylhJe/itV0BOZHFayUYCiaXMUXGMiEUgyFtOuR72S9hOj42uWhbte+KyXQdhipro7T4MBE91Zmh
BxwiIczB7wQTx4oxo86k9wv5RpzGVxdIJ1AK5O6oMYvgePResCJNwK/LzKea3rP33CXyL3qjyyqt
c8BUrxEzvqLw30Ib4DO8vuAqSUkdjzAtm1eHXnL5HJQpxmp06znBeg5qZVgIUOOvow/DpAWg9uqv
NvP6HPkckkoXCg2OUwsCCVFy+V2Rdve8y3F+NdQ+NDc8rk8RYMJ0sz9YPjUzBjZ3vvdn/fWOKpvV
+DY52P4bcB9t9pnr4YEGam2AXD7KQQE1R+aozIlpbybxtvHZWIJCYd1cc668kesdS/Xe0/dOt2p+
w7NV2rHjgu+PCYB6JJrKV/ScsOvESsN+RbBF7CZ1pjWILpl5i9G0G/GYrNarfM6z1mbxj8E3NzeY
rWxjhgkJlk2pSLIEdhHdc++kdCjdmFWN5WbK9RiWeIYDwfHq/PP6dVpR4PzbhayNUCftdzx9lgHo
x7fikZanZgBR7yZc81OMKXaqGPcYTB4jD4hxrxDp+dvyJedWjfd/1/TXW2OiiHxEvlW/ARI8OV+h
3gd6Q2lx0LMvzKmqPkHsqysJDOr6tFw5aoiJ3PdKmGAAj6qVpetW/BHa0aKcp7hQamRp1TGD4JDa
b1wiJhqXg86RszKcD9q0xOZm482+NKsAj9Qrn2Cy3Sxuqz3lGAIkQeRI9QS2zoNFOmFt3he3lK2B
qqJjmraWHQ1HbWB8jJsDaiK6/oJrgaQAq+MNLVwnP7O2x3Wzg1i2WMg0Q3gMC5geUDLqifllkZCs
s+hSsXy3nKg5V2Lu34OKQeqjnnw8FP9tuf1N/GIQx1iAko1a2e6wmbb4nSJzEXZPdQVpjyrAvBmG
zthIwTbcjtDixBFBGgI8i8FB/Ua6XfyeFphxw9Ord/E2vXR12iYzKp8pLw20o1FOA2JzffEXkxw2
3mogJK+bDPzXlSrJvY3K9eJjl6ISRDccFzUSrJA28YkahzlONKdkfw+2z28Zz+cchi0M0VVPdUDI
Yr/6wUyFA51RlZOUjThnf5QQCP7qUvgO3v6t1LKkj5GioAyBrb2YKAIHnOn9R9bfg+uSG5hmYG3g
o+l0/0oCo3XTfYRsomCmUKbCjA17muBWEA8NBpOb3lTydLtGl7J/VwQvFXuVglbAp2ETeXlUJGKG
tTjh7ExEhNp1pXCNHDc88hDkC3FpCctBD/p4h6fqRJR8R/PdlyqPYHdAYT3Q+PRHMqJlh5qZuj3p
2/fryeEteYWwx9e7MeN9vTrUecWqvTWpKGX/wh12ADrAIedCobDatxOb2m1Um6JMFIL3vl8PxOtB
ksKdm5zkHLNLxUBbHEGEOFwfd7HcwhybT9pP+haYjW0kVi0GaYVNIZnDMvDEOMUKzhnjWXmK1Ayk
ZwJD9SV/ez76wZecWNSa7zujVFtY9OhDRUIRmMB0mYoRmpBpPpkWYI1wqT92LSx920TdzpG7Nt+W
j0frW79eE5XOwzgTp/HayQvQJxQa4IWr1BA1X2Ib/onLDenEAW2HblVMAGzsoPrr3wWJ3igbJ8Kj
twL5buBGFpbtBLzCoBHRRGS8gasvvd+VNF+FhDbglnE+Au8jPG9LnIRPBOqaXN2ynW8BBOe6oOgk
1DrUT4eRTGC3IeI/YtKFdL2psSNUv/eVMLv6DyCeA6BeSeWRvf5ScJ27m15rALNsTUNJbLwwDhkM
ZhlDRgYtcylbAImLMDIsd+rYcDsepT/hhjyrIt/mgVMwIH3hZ3UAUNKSPIDXcdepcuDxeL6HEgja
ACXhenDTjqdEb5oi3DDO/Xc5YjRm9tWz4NtAuTa7dtHzochPqfKDCuAlOYaoHw5QIE8KuvdNv8Fl
44m852ul344n+J1BGvWGigxJgcEZbxBMgNncFxK2/Pbk+kBQBASxfda4d44coABtAFkk7/bnxqA/
Mnl/pSt6jPnEu/njnfFCYMoGkDk/wuZK3GEv+HcLZ/JRSUqI9QH0AHePma66a9ffhoPxGfrQs2yc
FMvrEn/JfRvqz2jVwJ9ctV0jjt2Ua5/XCTUh33hv4rgTzAuCZfH2G3aQSIZDRYBJk5Xzwv5oCm7t
vw1OUEKeG0MlCWBUZJ+4EGh0HPZTbSyjX8xyf/5VE/hKbzbJi4fprAL9H40Bt4WYqifLgRfF+RgY
vAl2zYPjwP8Gf1BJ6a89q0ot+mpDvQcJw2eywfjYYWRduoFbKKX8oilUYTjWIHwu3x4p8TfRym0E
8X+CNgzD25pQgnv1WeVJ7AZp8MUbuJARJvV0YyYavyU61AvCQ5rWpwphlJYFOXWF7nZd1OgwshT3
Cx7mjVhHHn+P9gPqEDMHWR3hCt7hWTcd8TuhEH8FD/jzIe6DiNwut1F39TdmAcuBxvlWF+xJaUoD
44IZjE72AxPqKDEdn5o/87KamBa6AZzsUR2NE5sLkCwLUBW+1RA+zRlXDSD4jiK8l6dzZOkfvnA+
g1JuNbhBKFYtU7T3ESfrF54K2jjZMto009EWmHZYM/JP36WHU5CEaJEm+5vZVjSc5oOtbCAsT7Yi
RwNXDD5okZWxkCFXVEoUanDKulw4qZdbXEnUBEziNYGeQJYzUdqOaarbRfV9qkJFq54sX5xRVpPP
aThTnTv83OzZnx7wew4jSQL1pnvzwGQ5ldOu7C/RLNZbrurGPfE2+ZG/UbEQFdCmf9LpY4rNat5x
mVrsc2xbxotSNgq4vGwxsSNonbQqXrIUIwTVT0DZrF0iVkwTS5XVGnF8ZE6071iNGLxpHHx23ACZ
SucCqatL/2OBeBg98uNY6Na/8NucQnd45n1ctH3Ax3cOdSnpKSc8JYm17ZHZF5Moa42xMcNBE2Pp
T+TLdllPOCfyUe/etaTKm78Eru64fbDezjOUOM9iTH5BY4qDQbxAFp+Pyunixm6JEg2H/iCRnb0R
rDbms1TYep6NVovJOrk5LWXgTzoNwzm5R8DLJfEjIYRCBBFza6NckNJiv+8Mldl+tx/6brqVymie
pH6Ve2bRHM3iWYEFzFMQWnp+8dBYJzxxnbs+58/uHcWIogRWEwLXar7Am8HoeIrsKgQjhNeTX1aO
71wWPJ1DZRQH+spJz5LBj7pnL5MBBqGOvBhrUCKIcIVMU4RAFC5xpPPoxuvTxlvFDRwxgAaXdGf6
IDzO5gPTxh0uarXPASscs7pqSnXGUE6Sq1swcsa7Bpdi1a39Y2oh9rkdeEyVW1tFkYuunOf7ZvHF
Xhm5hz2UzXiOL/JJansyGlkrL5bkBRCEB0FugMNZRsdnU1Z+h0pdbODPvcCC9OnE4L+nKkaBKzx1
CjQuCZHWqQFYz+uLfa4tzH/pyCWpa4zM6ujehaIopo+JWYD+onFVz2US+RKdy21J0EkYpcC5KXyh
VRw1Lbn1zMbEsjvJvzfeCnLaRIq58OnRGPEesHiNw/57iRS8vxn7UTGffgN/KZEwkTGQgBtQ+gmY
xtnKbBSqFaspz2XtyALiffetdeim3Y27DgxxmcKaewuiLPUoOBPja/Z7M7wRb51G2iZYUNrT+c66
RZF5vLxEpVuEEFLQ5ChW0lHtl9CkL/2iKw228mVlXKexUDPPXduOhdKUrwD5tppdIr8BW+aqLvTZ
P/g/caAOC6CRTPhJVfS9mFqfD7ph2Aakch9FfHhFU1iX2KEApnG/oYlPkYb0LeRQ3T0tnzy+aNgo
ck9rWfbctBCB5ZTvDuHTLkKOj3+li8RcPZq0wFmY+S7VMwfgNQZvHlvAjj2+omIaykUumwOztepP
aK4YPh9KCbUxlf9BMBBU/6qTT+5bSMJV0dyIAmrE5+Bmr+FgdhyoZHlTEwqqsHaDQcfqtnwSrjHs
kuHpsDb5AnjQQnBKVoaeTOSJ79yOyeHYBQFZSJjZ3mAntrgRsLlElH1nupQ50jpRfvWKhhLE8KIH
DMI9OxdD33bnEfitEhejbqZpl9ya9l/t7D+OjkXA4iwF8KofRcVC5OtD131AL2OjbGtJqO0LnYhB
V2kTIRcmIfdL9v60N45FFSAt36OWdbpW4WcmQZMu2UcPs4VXS6beE7uDP3X/wSk/8+l3ZlCvdgMZ
n4bhVhXByE/QFAXgaINTf+PsI1xtTdxfRGtQXeHgcYy+ldu4RFabJexLfua4kzVjAfYCs1fV/cGz
22fFyTM28SxhRppp3AXrXU78vv2lEtW3hiYfMfMZnLdeOr64YlA3Gwncf3AOWzRUENOegPfpLwic
D0VbK8vhmoHhZTXZco+j15lFLhBIGe3kRtplmdUReo0+9k6WPz/i0fC8Cay3IfbgVJAYh/WP7KGQ
B9NRcfjFEaYf/prff5D8sKH35VBnE9/3K8pORcWXbDrI1wPkB6secJyqQ7CsvGPOh9KUIu7bo/qf
P8F0fXpM0rfUHE9nXs+WrjsygOi31a7/R8lMNzwwJVjUDmf1itKCoNzpk3bBYvSIWC3Xd2l6DBio
2KBIJkFhj0/Ua0NtMjJ7Lae6ohe8RklRNnl30L9Lm6qggTWhl9Ji4gCJ1g+Z1sDpG3ZcK8eIP8tn
pdR9pFxnScpamFNxGioDTYB0/hE7uJrDN65RIyr/UwH3o2xl8hfijfBH7VonL1SWSdtOVBwwd0H3
RMVTmFXc2Aa1ZxjoCWG/ZPhpJa+J/Yr6fFVyWQND5l6InteTTWlJLYoyFsiOQQAnw/prYj7o/OGA
5v9NgIZ2r6ho1Ndr9kbkFVztIUhT0DthFejVDiEIrcBpJREyLO9bwFXShxiSRtrL94k0jHoZYHND
ErHy/WsJhNGJ8kDSDSyaZ+Nm7sfDSOy2IObI9SSmctu2Cl2mfU73WrJ7C9t+lD/duygsBAETMvFe
FU4MaWGIvVF0wquA2bKfEOfjeYc/PIjVxyN3U5CC+yB6RJdtGcpePpV/nNSK9yPdt9ZV+0q26F5L
0YsRAekdQgJYi5MDH0vAbMaUH9rdkmhaWkYmEIAemdvIq4PXgBZWEJEyFtz8s2kxHLsFr0i/Nufm
DKdBjHr/85H1QgTpiyavzQXm8MYp1Hj9maKc3zWFMtT6Qly9Ty7YaC2RkP2dpO6TH4sky3iTpBWk
5XPq66bQRiG/xCWZ8fZ4yUJK+t2YlwDjvoHJLj1pKov3ufpAxxN1Jx9usxRKYaKJFQVoVHvI+BGY
nh+d6ITzrdyKLV7HOi7IsRigDRh/rliJYT32HrM4ysoZ4RmEFIw0r8ts8B5NA4ZPBhlN/RlIKjEm
cC0Q2NjbT1P+tMnyu3+ABlfstE7PYRXgHbBqxBqpQQslDWuUr4Ij+hvDASaonOCfIuYXbH0Urouq
3vuPjTHV8mW/1KWVi48lMRVN8eHHY0W4u2DDX6LuewNGnVTXVWvOO+QZLhVscYYkigga4eINir99
cYxo5JMo3FuWT3BzsZ2QrdG0Fz1U4u6j5AQNS4AF/DsPdKZmtLia24oXUo+bBVMMxtR3oKNA7tuh
Ue7gSDxTUEZflrzNIlQVci64OHvhgBDsI+fuVaE7uhB+xqw239mf9NYFIe6eEX1gwP0TW2rvnfKy
2W0427gXdnopmUmFdK/Lnwpu2sn8cIy33wYS1eF6K2raRcwXfEqkTu84XbBS1nLyWGPnE+oK8OtQ
mV85FmNh4V4SeXHLrFIlu7sMsJ8Vv8tSVD+JbiuO7RAfdvxyVvTPmfdA3mxdMkQqnBQO4ueW/HRm
GxqPsYgbWVEOHvPuiJKNelbk210UTNw3LIfWqCI0o+sA5ZCmAVp4tIj1LYa1nWnZoWuKyAGUecHS
fAm/8J8IKZCXnKBIHtJKCq4zf/oaRuLbnYtOOd/VRBzlM4m6321b0gosifJrvXGuxrD3MrGiXf3U
Mx+VOs6dwfxUF6M0y9v6y6hzwWQqVblBLniLaV1KvBToNOCFjdVz6f2Ou5xcEdY05IICjRwiKYJ+
JIwzBbL4usDhz75YWUyvPQHNpQY31f9FOICHIkR+0CimCuE8i/G7IEeZjORW1WhkE6R0SKii0ZOC
ITYSUsn2AOJ7tg+gK8yQQDK1MUeFMak90v3DuV94OoRPanwTqdIwfTcRCG096WLEoLb2AuRR/YG9
p0F5Gs+ptEvYJaDeIrwIvmmu+ljOchExDOm8g2Z2h+lHBnyJlrLBnUt3ZAqnVZv9ArQFxQU4W0dG
rcgXhsSKkVmWJQBq16zCDsjuEsbHR+2gPlT0D/ugX2LJWbRRhhEZSqQUprevuFdRrn0rrjRE0dn2
CjBGcEEw4I/LqE/mZKsORRap4kz5vV0Q+a6Vgo19onOU1GXS2pXiLdU84civ2600vC/vtXrHhDoX
t3jN9uXhiBHQ2wC0M61fFSXgGUoj5LMJwNqyLsdtKh4mFESpp9SyZVBmk3jLoWshRGtEeLwN4xPG
24JWKWPv/h4Itabm8h0O4hsJhAEp3mGj8ozuACYUQmlz8awUlptVPJBJBVz/rVCRDJddTJ2oJXf3
eC5u/GMKSYe3YUbHumX7F8++SaY0NyUF8MbyQU/58DolCE+1J4aT/22clHoizcGth6/9j68avt0m
q2gm+flwLhUMTRZPFJt4E8ok/eew5PO1w+GOhgY1HXyfICJAlwZ0SeqceOt46twb2IoKdJU8+5x0
pTZUSkW7hIZIx0swXZtUbtH/x7gBzYn3jbTxVgvCvFQinP9PvkoPMuwj7bpM2gX9+u/VNVpkmuQj
KEPxcX3kThcmqgCrP/4O6FjZYLmG++DtNvpOtDdH8LBuBmoDflZbU8DzjsT3rt/1KzARXnYn2cBp
gB0++tdVpR3Ru92lsNyNtKxa3gkHqk4/dfdiiF7jOomcFXdzkUVEZGqpEBpgI8y5HL5AR/lzeso1
1U+r+h634fIvQRHnRLIaJHpK8MPQD8slgm6guR/CeRzkXs9RtDiP1rC4O/kYXoCk581W5SiCzCoC
pVJ4ByPD9TcBPRf/tC1TC+glRGzm4slNFwE+zSO0xSH5DNSl0nNVXbAZEb53Rew3IYjs0BggOA==
`protect end_protected
