-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fQ0vZReXqpwdhTbz9y+Y10nv/wobHdYUij8b/WVD9XM6mBHrHc0MYeOevPNqCUsCyVw/5xN5jbpG
C4+tdoVoVys9lFfzlcQd1MYfdQQIhuFfvGqTg3/N+RsAzqw3as8G/jQ1SPnj3y2jlY1M+559MpTs
m49KCDudACSzSHL6NH5BiwP0AWBeHFSPH8/sfEbxurSpprnuIQKf0/RCYmg4S+C5byhWNVAES2T/
mO9UvIv+5oNdqDG50xxiRLyjKpQqMOhi1yt0oxFoh350+lsX0NqJO1c4aSkvkvld+/kq0QIGS84/
1P4iQ0ar+BkpIa8MDCdYW7iahsJ1X85Hl6iIDA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
tKiAIRQyPgscOjSOyra7DjgCzsMsKKIiwa2W7QF0tv8ors/aWOBKhS0Sf938odloYIEOAmltPSPi
MfY950b8AuSUNePZiHVcbkcQkj9oW2z1df+kpiiMBt/x97pc6W0wxmUnvHhJ+vhzpiZLYoS7mnAy
ePaLl64vejmA1EAj/WHJH01Sn2EE+NdjpPlOih0p/3wxHuI1o5W2kexxYCvO+pPzMNBykaQ7wszz
WQYpxGwI3286qND/5D/aV3DbjV6+HEZrrAuK0Dp9jzmV+/z7UwCKiyIZn7Cd2SVKfNTxdwHuN2O3
XkR7sMQg7HbmlXLjNBDLfggq6XuacQfnBe1+SPy0m7CEcWnXOMdhHXZ5CmHNY4VYOPfWYtPX7w2w
IjqhV5hnn75dBs+LT4v084JjbnQBsflFDc9UDsmQ+J9fuFT9vftmvAeMR+A/p8CmgOutzgjBcYVw
RK5BA9dZgINNE5qi3Tt1qCClJi5GyZH2JtY8IFUb0cgVw6627EX+x46Y+sXQ8LzkZxoVcWH5kdTS
eJa9cmpp44Rb0uVYDGmAND15aSlw9P8iO2BgFcr6qdZPwkhLByN23oxGINtwZMiLhLeA0fc/cs0F
Dq1kV8XsLNFpEyInH+091bm/+V+7xvvBA2inPvj4DTpnJ2QNj4pZhKe5seArnNTfrbU0Q3T4WHA0
ZSYrpw1JCklRO8lIgiYsL5Mts3EgjQPwHYQZAeI8GcDbJT+0sqkQqZb1FlimQCChGDPN4OQpdnE3
XrekaAad5mTAtAZ05iHObA98/bnJ3UJ5BRvg30WjC4d8d8JyxnGpkUP4Xvst7ZtbFpg4cjIOyB0v
BYwBCMp4ROiw53OeOBlW3GQaNaywwoMDJFoxKdj5XcWud68Ewe+LrXQm5mJQCnzzjJimb6izkSPj
aHHaYLgbkWeCPAZtwZKJy1kw3ianzuzxt5TkevRhl3T/+E2V8h5M0/cHY/bQnrGrmJSFctws0ZBI
rmVbAyCMGQ05nunC1qLP6c6PjyHHJu/g6XR+5xCeV6qndiY/7ZLkEym8IcGZmp2p4pBBlb+6KVv9
b/WbA0WsrGOcfqo5pSM7AWNgTzYvFmUjA+vvJgINZpjIIKhe1JA6sE/MB7N+Ry3c36PYx2eGfI+r
ycTTD90cs9c41JGoNO2IhmSfB9i+ORKHeXlgPGQmoT7nNs2GtUVuz7KjigrZ544CVW4wJYhSonHb
cywY4nFfMSwUbtEkRwQy6Jcl+IHUppX51lXa1FQJNoWloGNKZPC03LP4ypTjcAyGVUlN/cD/2vc+
W2vD5Z7a/8O7wDnhwAla88f+k4bQI+UbqFF4tQdRATwbWnf2B0WSfCHylmgQg4sPmJyLbiRT3rut
N6yB0QLGuTVw8G74EdYh/tneK8Xm6avo2Jg61y5b9GHH4wAtj5hAmyUnE97ythq7x9dZbE7zVeiR
DZ0k0W/5IYlRWi/TRadPebGqXXhAEv7Pk5ggKgAZeocSgS9aeHaj6dcGEN55bvbHC2e4t/QmVAom
gLf7P6dUoamo1N2jNulpWjkxjqhfA66GF/f0DVfrnNZnR8T3E+PkuI4IW6zF74u2zy+LaZCdLPQC
b/0IVIdewTH0Ffkn99O4Hk76N96gpr+6b0KXruzAhZqbUqvqi9WR1fkcE9Th4BzKqW7X+dU0DuSe
ygNy7sABSoY+YbPR69K+Fbaci4ktqGfccNuRA5t+rKHtHMiI3Dnd1l/1WXrnxuULCt7yq1x/pAFn
lQ/fPhBWzYWT5JgW+KC+2XIIAtucigsksjW38yLPQKYQL1IXXjAs9lfTXhH/lLpWV8WzV4t/E+Gf
ypJeoar2I9QXK7Gvyxhp2oRO5EgHU/4E1Ys4nwpRddXOe8KYNMlqjegVcc4Lv7Q11uiSYsHeAlh6
T866sGAuCJK187G01IYn/LPZ2e3xFDQ+kzQCJDsuef9LfyfEG+l5U00XiD/ll10XUZAFNOA4wOWl
8P5hO+WN07VAahJAQLx8QAzqNS7ilcjL619vXubPkmkS1f7Kdj1Hv8WZ2Nc9z/pgHPGWTehMxgOi
eAlZPC4kAW4KZbenVZHLzbK+ntc4+4czSElltceCNtnnnWEzl7XsG8Ptw/rNSZwuV6ZdrWW+aFkt
1uIX74Qfi2orF9W5asJwdltyv6KP7jr65GxVOYKTb71NC12qpc6USqPzUgtRl2DUhJ50+qiEb+Li
OQ2+1TVJu/lKELbpVuvAwp8Re/250Lvx2xGZ+vwDbjeGNf3zjr5xKsyjXJFujWnEc2veRyfeqYqB
fWHH8esDSuURTMrxk0/MKc/ksgDeAeXP+lXkfYQLyX7kwoNobJIDCH4vYS4JvgpVfMc36yQ6fI5n
iPoOBEMcna04zg6Ae2/dGkau9UMnHtriQ4dWIOT5oNR00Pt2RrMXr6Vx3A4UuwIYnzUmA7nX3+Cy
6gd7Sff+OrqbFs95x5oZUlayc7krausQO9JHo8tA0QfH7Ls20S/3QyijRNnocxohmJsRge52ddvb
QOyX72KYaIp6tOWw3IwFEr4kqOmgv7aQFtCErFrqlQOEVBa3a8sXW4w/oFFI4oc3NntnsSxE5yZx
FoHjut3u9tOwFOOynhKETDiZMTfD5chHCeNhlYf2Bu+xa1BdrVmrOWX3obYVhWExY5V7u3N13heH
JOsfGRIii6+VkBH62aGSsr/4X4FZ8I1z+dpRezphSFYNYHrNlnM+F5OAaUWAeFYzO4qONKujRTtB
O5E6Z9ItXFXwPhgtIPv7V8Ivf3neWyL8JI9tvt/osse92jn1YjlPtMRKFo/y5gdADjG3LRT90tEi
WlUl0dgeRQE/KihN2ZJTdQNb+HnnMXiob1al7XrtdSvXVtHe4d0ss9yUi3WeK7z0QLfv84CBU+N2
zyw/plsQcbDDAlx6kQyYMUHxkMhD0XcxClfYXE5z5IeBlk3mSxRifQ8gterLaZNLytu3Jg6xAJC6
lK6Uuq7lc6Pjj1BpyuDoC21lFN+YdfNT6NsA1XaHOWt40YM8+p/Yy3gd1poOwg/hgeBMzB2MV9Od
pA3yjKehKkTAtRglUPSabfJHjHauicvW13+oJBcMOx5PJo+EmIwomapLKPv720tMw2HzsLZgLwqe
Z3sCj9RKa493+pFcY/X9x4EGmoTvpbQFgtm/8bD9aLi1FtRKTfdX3z89gt+M9PuSs0ZT1sAjd42w
9ZpDSLBuymNmUZVMZWm1aTxQ+7K25gdeDmd0lzDnU0lTgIjxADebUUaKXZo8i9n+1BouwOBhMPna
CMveT0D0puUP91LiMIyoEoGXlAFrXySKciM7o9exYG5fM5jhmDmuXExKEKTx7qonxQh/sNz5HQPH
OdxJAoouS1EOla9lT/mULdGZ/ArveAPEoiifIybbyVtAcL+nfUYK5ntt1yXCo+qM5AMBP3kSDT3t
ShducKMmwPRmRNppeXa/BQCVp2AsUF8Jf9jp+JI6KVL+1DdWAJsxAieg2DFMoeKwqPKXU9rvmo7H
jAOu/WQI2/poy62BFnN5MsP4bF5OZG5UjWcUx9o1kmBTTPtiiUUGY3eJgtQKeeqZIAZ0Jae+uBl8
bfQpSX27sIc5pBqP+aapoJLtqMBTAP72J004GCTX3jxy12kUf7EakQM2RU4LHzSnPxGD+HoaQGXG
yBpeTES5nPvq7qwRg923wHRmPlPdg1Dq8hnr5tN9wyTXbNEIU4ql2VkAuZdarsogyevcF+J69TMK
2bLKMHGYdmXYHVVF0HwrfhNUWm91H0KQaF53jc0pgwOZ3+ripUnl0os7IXrcv3y7jgtU3m4ikvbO
uVG65b4sfJJvpp1VRtWpKx1pTujyEkMCrWTHBF6omk/eJCK9MgQQA/exY38EzU6+x0M415LQh3Q/
yKOm3QXACcVkvDfQbS/rdeIBpDLeVj7x9+6TvlsGDsT91pR+9cojqCANQjTd9yZ5gijr7gM1u4D3
eiFQQEJRyXsaA7NIlu/deIxenh2lCWTSeI9nh6saAgFTJkkK49KTzebLq0SwH56tIhihEEj4UMeT
zPDIBc4Ep6KtJK5JogG2osa7JPbDSKpZ9AnXTAqHss4LD81Kpx/hRxayfipcpJ/ASE97G4hwivau
67R6iipSr5M0HYT7/4LctrYwHNJbmXi42BuaIHOLi57ZMH6sGCiNzoi3oc545GtRdkF2MCcv5RGh
mYkKMtziI5ZJpoo97TrYRZIsPwAOokD03Dq8S1SShQ87NDcnOjIouWV++Hw/f2Tmr5Bd78S3iolg
Ck5X1nqQNXpXuY8dJmtyyJR7Z1lK7B/Mlr17FK/ocD7oixJRv0S1PZ/KwoKcS2uMvPUMOE9c+wyk
jChxSmWzzwtB7W2u/+4eOWNRpcziqEVHgHcSzvyF4EkZPINMcoqtJ3TexUiHVfrG/WVGC1kgqO8A
4ZDBjEe+1UAOQ4YW+89YdyA7zqELqyp/IsAWQe64xBRNeKoTBGUoUfBNu5jhHHi5zQrY+Sawfe2h
gFz3HYEaytnHXXiQiaAlpXgbaG6FJzx/o0PlOARLpbt+fL9V+4GqNujb9/9oRHz8FeK508Dc5e8Q
qq/M3rrLIroz9MwCnPwl37hf+UDgrym02qSo+sLmh8vykBuhv8bcwsRGFFrPEebr/ERqMjjb0MXD
GJmUwLSffnyT2UiZpiknLMgjdyCtmz67z4/PH8gjZOnPYOdQikmOHR1E9wWMkJ4yeZWneVAxcW26
vH4NnZJjM6Y08VdHhUagMUpbfanNC/mB7HdSUjG8j/HhHXI2w8oypFxyBXeZp3b2MLCWLBfauhOj
ppt4D19s2zeKAiBcuHaSeqmdmnCelC5EJSelDZYC6dtVJtHU4wJ6Iv+uLmUBU3igh8GmYtf9OTja
iA56B5fqp1dgfmGl0ZBUtqArH1ID/VHhpwzF25TQ4Obs1XKPjFBPoH6D/zK07fIURingAxAqN02h
Yv7eMtgOmssZbqQQ2PY7iy9W//DFUjCnsOO+Vo/IhVlJzLUx7ntU+jRW57MpAwZK0cOJKufn7gMN
hBZNDA0pHqyMls7zNkn0D9nhJyOJKOZu1VIlHIMXOGUddtiOzOJZer2BGnkhsQQJzfAwbvXpwWMe
vMZKybFNooT4XXslkCqbUYKw1QxdmWBHzuYFIDrUJrrt85QSgo4s8Jx4ZP2kz4tQEkapAFmqWctl
lAj2ZfxxCPaYI42avs9W1Qt8LPOQrCgP2bAzZpP9nUNqwfHyUDHau++vaZ/LLYnOpVmaq0QB/grT
N93ZNhhs9l68BlG8+vOBXxOSG7ebHWcGhnAoARVphycTZwvfaHZj29UWMyfsXJhSFgodR5VAChtx
whxHH7xOkdp9cSeBGYYQwQ9KIDXBs4Np6Hhkf90WYIrnA1EEYqSwlW+ynZc3xSNzd3xw/3kIXZez
jFIDqG2eDsZXlR2LGBro86BCleMDRgSp9/H2P3/QapDakdVBGwD2CMu3zYItx5qje+pz+Hi8ur6h
jfrkkxTd+ghlvzUmvO6sgDYmlQ6K1rWqwQyEKc34tOnIfzFsb7/2rKpRhAbYVJ0BTYviLaOxIrmU
qtA0qk8ahVklJo2fpHZt6xh6DlYhZ/9CLxJYt6iVDuY3ZF6XX0GXKi0MKOEB2DtHi/mvzsxx4Xeu
e1cO8VLTnyBXrm95spW6HS31hY+WJHjMGoxn1iXf14RX2GuEda0WaJLytDbiVCUa1i+Nozuuvmj6
X46GVXm16LN3sHf4OYHIp+C8y/nnJGjgfQ1I/z2P+9vauOhJ9QYv1lSTXD9JMMRWNAgkro0gkQ4s
75yfRn1zYEZIE3rLnFrjbdb81QoGb4PIA6D19m/I94TXVuw+TYNtSjraX33h049fPWEHb5+6q/wo
noZAVM2qkHF4U15qtnfdjhPp4rO9Upe5Agm/XPb6AxnAJjUp+xM4+88cNAcSYZnheKl+G/t6H7yM
WTsEVIseUu5SeGY6FFFZHbKXSkjFpXKTOhzLlIRHOd5es3q3ZhW1PYxlMPLjuJ5O4hKL8IKRhJCu
9HR/gDaQeMQgt/SYvjjmN3x1rMjvzOmvaqJr0kPr44xq9wcpTIeOUgLN3yyvNFY89/cdd6IUukvS
IWxXGvQP80VHFpuFEsc8tQPCgTUqr1XEDEAuSpd6HDXsNUaQ1sekJxrPY5bN3utYBZIkPEMcQDlX
nH7agEdyvzz50lRgYaEAOtFhJvjwW/hQOAt10aOdr1aYuscCjM0mW8vSy3fT8iP+0m9dbLXMZ9fl
IdSEJP6kXOoJwT6C2dSz++AF/ErjShsZ7tN8loVQYvCvKkIee/VNqj7S1oIfw+Jg9OLVeL3OlHN1
No3jRUEP/tAflVo466wz8qmg5IYua566uw6N1ErOQDnnVFTtH9Fz++ggulw4PInJEsA0O0DUR8jx
aE+VSZOXIQMKUb/kjCpTzPCvzLJv69xVJT96uus+XO+VjEKwo+LVjtiOTrUogjC/Hm6XWnE0UtkT
Ult1tZn6Q0hvdq6itR3vcD633+alz3pLzpt+xt73sHVwb2QMb5GbHC4qMKUQ91kByKdVU7Q9A4kV
tgn7U/SaX7BAEhjm3yp5wgQKL3+S1Xu0DuJ5FeHhFWf1eO4f0MGqhiFnGnlFUGlm1/ZnOSVxN6xb
SO5Y+KaM2YR0WgUtLjBkI6njHhjm5ITTlsYJBI1jaKKsl56vbWq3i+zUdGUhBjgTnxfRtq5hvTSY
kbJU4WwcGxy+54SKz+pGi83LEiZPBxdqrYnMTN038DyMDEo+IW8MvsuvBRlXD3b+6CvLqhMPoSr0
SGn4F5YItor9kSA27LJVWX9Hs9QXvOe1FNSJX7O6PndarfVK2dxJOkCtZCaIaKpc6cmccRg3cDiG
Ydxz2L7StArqElBIuaL969fFxU2xk9G6bfFDBzq17MFxnkmmXnmV6RinIVlzAlvo9MsKdGuL/veI
hLE9y/YILKemWzpbDC83eIei6JTkQlybU8DMse+Ew8j3eKRdZgrbS97iq3R6i8HYmrzFpMjUHDHg
/G/zdlBEbLyKXkvzxaHuFUr6IQtij0ATpeJ6gR8JVp1NAQicjz5BAGiKPdoWhzHg38twgMVDRFR5
yUCpGkrIm+3HVo2YJfwa7DzDOJOKaXfxywewUSlWQpuAX2qFxaR6VXcO8HJA2Qo1Xrno7InGa7zz
sF44/uPf0k8nG+ciyINkfvXG8j72c1lYO3/H2WxdkeSpcK0NnP2u7tlWHfNSxEsiKvqjiYWQoDbQ
jt4A9sRDawBpwh0vrYz7l3lH7gpSz1U0V8AOGkWy8TVs/LD6+C2lrnyFaMjVAOFLa0d3zgsgVTvB
Ip6a2la6N1aO3KK43WCBfyvvdcDwmJdGWrx+JfWvuKZ2kanxNaLnRLYOmxzzq5AZxiFALiQ7UvNm
Jm3uUW6bxwmXUuRWZ5fdQpzoGPNytocd3josMjp5TAIGLNheIxlFMEGboaHZCyGNc2R9naZPIKeS
mCoaeOsvsNlOgguaePzaHnso00uXuGBqnwfMyM2RG3zlZ/y4g8YF6JAyxeib0cCJc776eWidKG5r
c6D8zaWRGuEQcQJcNZcT/EbLCGxAUvLLYjVVm6RSd54NzaeebPVXt6lAb8hFtciiuWtJfYaRn51V
xfhTXj49Hnr/GGCo3WkqQs+VS9oYQlQQNiwoXejfNYQEm98J18/T6GrBbUKrkG8jc0kCJJ3kuYBW
cqZKEVdeNQIpoCGDiPkIrnwMUHRUd9ELr62nLGWaOtW1LB+LCZcDeURGihRqldWy3WRhWURE9QUb
U8+fvDYnKM0HQJlY1g/BmBCcOJAvEIHXVU5okfiXo9LOWWr+7B+wEto4tVPswN7gNweg5ktpReA6
qcuWSZSZOrRJQkqpPL+1cNu3M0JdGKe6WSY3hAt8S56qEuOWtavXbd6ajNRVA+T0AGT+UN9pV+R6
jGVu4GKTdZF9D6eahmDHxiC9lCukk6srGzGFezmGAl8PpiGrs7tsfJPffjqTuuItFcQoT7YFfZge
faKY6g177kSTRxt2DHo4cyHzddcHVQD8VGsmZEDbUP8j2DaffvE6GAqskc44vxAM/mx3TV0RL7SR
As99RqE4ZzPT8aDgzwwjlyJtnAZKLIVoXYlQtmtG0q4B9bfe7ovaSwuXNdekFKr3sM0zwZVCBqUl
GNlNNuK6pQzRnx29dtfjXAMds6nETNW0eXujWkdgDGJigCp4y30NvPX05k2vKvn67oZFo9mFo00f
cn6Kirb7RBF4Y/BO3JpWyhSgHJUd7TB12OFFn9VflBbTICl5g4qkGGvG99w4Cb7BIOKJMU8sJDnI
HG+XNvxnNj6aKizCBdBx4k2llqQ0HwqhR0n6aBuBbrlWa94kWOinmQ/nJ4ut+C1rMgU/HXxWoEWf
8kYSiP11LU8zGg4G+BrvsVMJSs6VLCb0O4JXvD2Lf5Nkx4p4aTAZJCBAnQrSn+xg4IK5MFoIhlqP
DCETBxWtKfCCM/8Hk7wfWJRpaolHmFRZcTKR8N/oku4dgwpEn9JYqKJ6/2oYmZZ4160ul/IbCc2+
I+9b+fu+hnZEuFgtvi3sSfUJGLsDTY3x0nZ/xhbxEDokRMbaS1Uz4/fcQfckRdAEwPINz8A6UZrF
ustIVjlr9sP3IiVSY3gWvm1UaKTCTcn/Efdj6vVMQB7Xr4KXJLw322c6ZUsBsUicemy7GNU5MeFW
A0T0v4m+Vk8wvBqn4Qx5YS1M9fxuc6ZKONPji1gk06a2dysYbqhzuH9gO/5TVkIO5T423SEsU5xW
5AfSH83R2U1RKSNOcywshlRSs34Yb1Kno1ReSP7PyCBZhYCEt+FNx4Nl8DQeXdm1HAluFvOVPTL+
R8VWQVHgVOVNmqQ4hQjjWpftHyrnRZHimx33pMNK/E7xRHvAWTBrcP2SMWvJdRvon8baLOLDexU8
9yfv7OkgLZ/oIoapkQ3mPtQMnc+Y+boO/vRwmPIGmvxW5NvpTx+ryGyvchXwhjcX9aZQuakq4Qx1
n8/2bRu5mCqsWt0P9Ajm10kQMF58KUQb9kwiPIlv71rkbk39+zNrVUqlfkWGKJ08x3S5SL8EDtsG
SroodsbuchdbNoQGm6K8BgiSO4Ucke4gg2D+5F6y+/be1dOtg5i3Qxzh7iHRX0XyHPo+kwypb9fr
icZa2u/ldcgZwzhP4rE7qvrp/y7f8ppBtYGWLRM+eTh1att7HSWGlojrwV5b7uR4Tw8yBVILP9pT
Ud6ZQ+1UW1laBIfBxxhpEWAQ9nom136Ib2sejk0HiZ4Ak1AD5xxS8Xys3g3f0Q0Tes8MTy+3P7Lm
DnevN0m6gOADFP7RaPKcBuQEocCgJMszfmSuEzesAU6mrxswWheYofvvX44XA79a4JeIDtihbIs3
vhAr6jWb+ttXg+KI0QzMI9kL37TX3ej73LnuXgjp5cxD0P2/71st3WYDTeeHbewNIT1jVHk76Q43
9ZPYryy4sVDVdzOwpxoogKodODk7wY/rgdJtHy4zlIbOxEyKepyMfia9ZXu8bbI3nmAueVxaJ72j
r4pSoCaFoo3AA+wRIJR5Gp+rM10WIcU1HkvGtXdtn6Eso+vGPBMJq3/T0SbOq54y7u3jnanF1Y/f
VCRj1sMLwjc95GmyKirSNXO4BFto6/c3Y5Hge2cLXJdq2AWNN5NgEUFfpmETmbvpjEhtutu3f7Rf
cKqXZyASxGIe1g4LL+ndQrdy467fvt/qVEAPt8xTOYQtlXQrIvx+lDBTeyI6z8pSYvY1m7+FsM0D
eD1bPFuB7iZeF25yEAJPv50rqcrJl1uWWn+3NeyzL72cTOEQNLZWiEOl5IuPQWoxTWyIoiBsGnDj
dwxb2fz78t6NykP4Ouusu2qbvO85bDxCk9hKAalxNm/Zks02z5zodbURTpUR60XtI1N0YSKX7Ljx
9OJBoOEG/cRCy47i6fUgaQgiPOSquIZ3EkdecyAm5DHHeFeWDwDDLjXJaLTnoaXhNJxQmmqI4dU0
bjzoIOhtEiYrPJ9L852wCYOudA/j95rdmRrOaoOje2EDntMvld8p6GI7PijEvRBOVGs429ET3FvE
oRnnfJhUfLOx/wi7yU/Y0FEWWUwf8s5QfE33o+/qaB9i3BXRF2sg/piHwqvAHRvr5N58zpOvZvh5
1ScvrZtnf/2Tq08EEAtu7YovtphBdNwNOvqWoS64bhsW7RR+PQCp0GkY2zicnpJ0D2d7bQN6V3iu
xj/1Z6QeWb6OoqR3UX0fL+Jf6p4AlBi3O8GXP0Fw4iZ+GQrx+HXQrkedpahtnA7WPXpnNsSUctb0
7E3Ww9cqSGl/A/FMUUTFOhwsUsFTnoToze8Zpl2wVhfx1/usNM6FD4j2KWskDzPGUau/S4Z7P/iT
wti3yC5eb/NQQDQ0otlBnbyNB9KPuSj/H4mWH9wlpr4DihlB3XtPI+RZXgtgVfqyBTYUu4PoPq8t
MyMYoCKnKDlsbZ1zJ1IepJgUqma/4PGe2ecuNIWKlP/FfKA3J1tsP/p3kzR2n3slh/a24QWqSR44
KYxm09B4tWS1gowG8Q4DdLvP/4+CcKcSHsNXPQBRK/TKqHhzW+oW7FouWTmHkmyDnq38QPUNprCW
S3WibliJg24iwX2ekifXVGzCqJysfz4k7FtEs6lyaFWu+0Uk0SBTwo5yq8dMF9YCZFusM4rewi+E
ZbiBf9QljQSKWGIzdHOuTSNhoubXOLMHimdKTYtmZ9lp3L3j8+KLRsCqQH9smIyKGKNmcO52oaOS
A1VRSwSa+9xjr/gzJdlFvvcnNo1cHbA/U0ZJ0S5TOaUGnbX6RlMEG94F62xOA+KT2VqF7GhGjeQy
5ZkviLFfcrXOaKyxhpdytauws2AUhIN61LvWSmSRuiGTKrb71vVtfVC2DhqGEED625q6NKbYhs5x
3Gt1ubLqn1ohMK9pHUvTCSZ4rZdBOTJB2JMSPvSKzDdD/qOz2D7eJVvYJ6n1ufc4OTmEdF6CfaOm
K+9VAM52jF+jIsLVuk5xhZ51TCy2V5EYAZk6Z9RZmy6I2tN9OifYkzlzZEYWhbi6sGdD0z4MJjMh
CQ8IG10agQl/jF8cNdCqCmHt7IqpWaNVK6RreUdGCKl4yiIVx0/kLSY6YWYfz2dGNJ9J6W0kbiFA
EuxAnc4D5Z3+wE6pmKTnrjY1zINmD1L2vb13sbk4OW0vbnvwcxHsJsik2GFxcjOqMoS+eMqDAl4h
uLQ4sS5tkidVTW+h1u5tMX/66maKRiFrG0UwXqecBbDwWBwzV5QGewinyfeZyaS0coJEvBWx4vat
rnn5RayjeVCPRcObW6d3mSo7aC1RTqauxtg3NtuUTHpnyjEt3xTXHvQKF6KxIzOdAULST4fJiUN9
X4hhka0ca3Cp7oadfotzuWf3gigUStYJogMWWIGWp+5O+p+qxJKtkRVTLUcmot6kifykgp4Lw9hj
TKnpEUACC3tyX+w+HLb4isjmhekoAkrOgDTdLX92SW4GFRjBtouiL2o0b4MkrF2xZgvKcEfEqlCw
LDoreLEhFrRpA3SSpWeiDuXKUgoFaDwZEE/cyG9td4H4+nWyCkUz6naNazadhf5cIVOO1Rm7YdIx
hucApQWAZl5J3UO2KSvOR4Shi2KGXeZWv1bCYQCL4aRrqyc0vs+8bm6WwNoTrXRk3Cd0kfOxPBHb
tyyixoVv88V2rk7o+RWFtTdRYRtQPgjf5JELQ/4OCiIomNXfrv2MNteZN1opZidiB1NaAGoFSYx4
584aOPJd+E/4c8odL7LcgdeUplb2rockLv8o+dnc/lSAAarBgHnOdfdBIprhF28imMpNAX1NZjse
DB/uphKJymogQ1pFIxTfS1qvESup4WCfj2TOduUQUCoC5L0P7m5TgLklj0YZlrbxrMb6TdlSMmB+
HOzbmACxaAgT9jntZoL2BV4Tx6ZYW0FqCtmiFeP71bQhOg4f+RL/gusJM017EUJaiDg8KJzIvam+
//LpPYrjo8HD0rZfCoi3ZYqau+FrL9YX3PkxPPfmwhyBmQsxGfCCe/JJ1MIuLPKEgHBeuJ8oSMlB
07WB82N7JSNIjWLFwsRWngQkYRHPlWVHvfFmzmSeK9iFnwrc0l4Nu4qcRBg+/vrql68zIiGegLac
uymBuqA6CMuujDUSssoJdZV6w6K1ubnQuvHUH0iCw4h6nMxdnUvNVYbz3Oqec038Evq7mCGqvSv6
deBShT9ulHdqGih603b53aRX6Y2P/AQ907YJDa3Jf3o7BuRVLTkleVubhmD9bJ7C/Ef9PnAebuFA
5r0cmfo9AzrGxTAhN/FL9UgiKp+smdfvTqob7mZx0lKYEhaiENdMUjc2oGQTXRbk519TBV+iQ9HA
78G76c9rAGFHTpB8W1XqSWI4iMkyGdWcz4jXpvi30SorJhyYimpt8OF9YNPhPsHTTkHm/LFZ4a2e
JYMf1slf/f8ute/5i6tbr6mFOuzfRswspepQLmYeeEjYu+mHdR6eo2nRGOYuGAP9GepHMZamvG5r
c0ldu351yNn4D5ZE1qJWl+y+KzXYsqj+g8z/vTXW3ZTDXBQr6pu09nUbULaPiUUiSkjwVKa+wJFW
6QWHwyBDNjOrLssPpdaz7wYgHscPozJqHfEfwwYx4u2LBZnyJ+oj+UuCpjnJwOzxnrUhhQ0mwVWb
I5WTDoOWoTp5FhJqI0eg+k1YCOjdfNUNMr8YNgzhy9bRD+2LOLuGhpDpSalvgVa4GZSMLZDDj7QJ
eu+V8uHj3cF7NFf0d0E90poM1vOX6yBMbNc971poiqoY1S7XxUMkpUsW2qmIO8sWM0MWIKkS53Sf
fPagTRoVbYH4+rKbrjL399tXPFL5jUpTbPNESJVeY5ZE6NZ7Dc60zvx9Rn2z+CViKoZi9RmChfIH
6JyiTXqwuAb2rZVmGloMpIECJ8s2eipIclhFpYHHadnUDLPJPd1RA8KxOgzj1hezkHnbPIRCmAI0
DwOrhvRnfgKAurV5YwH4S5bXAlNLuGbbumI98YC1MERioWSxq2GnAFvLjw+FYQbb/8Ah5HcsnrIO
zHr/ltMm+NGO9ozNw6pQxUXR/OspUgii7iJG9ftdLoCFvgtDU4KgVhVV/wSUvG1GZY0UXzoOECny
iv5tYe4K9mMqBLGTUPBmbME9K9HB0Ra/JONlDw9h7+yHEWra5QF7h6Wpjxu/y9uGTT49dHI0KJZf
O/O0ylcQE0nopNko6ezs/vioBQilnTeux4ZN0s2LPh41q04mwjbpxw7ORRTB/3igd7FkuozN0Mb/
nqpuatN0B1p1fblw/FqWNxlCBcjq5rSSqmyG64t3jvVtLVp1j0c+vhvkEf/Sexs0TL9G+6vRh2p/
YANIPipQrs/keaBVbYMbINg8HcMr9fFUbrUByU1w5Pw/IDngQzm6Jlbmy3EZuw4gcm2NK4zuw1cR
J7wWN37p5ffQe6ndvNc4QdgYcP6FlLIj0Y1WJDNAb5FQsDLF3A8jOsXh2LzoKz5vPOFcUUZyAZLE
KrRSUhyymIqNyFG6sJs/NRaCuHKRk4EE8EnzbTzQkCnmmAIsFVzmqO6eoqpteUQoi949i2gCYOlf
rfmTG9u3q7Ew39L9/P7euJxjGTCqMoAzftgFBG3wg2IiklgmMHLK313FdinVheJsteIx2iQK2jdX
0kvj6rQ4rulM9xp4izm4sMCJyY0j+i9MN1z2pRJsA5xCk26IiEL4nTnLVhvVbUuvARCidKA+DEHe
cJLjPFGZvNBFoj9YLgjuYSTlAt09xsH6CAWHkHrdMkpQiwiPPy13Z3DuKQ9ZgRX6i1RpF6VZ3WX9
3mKVi14JDqWBxVUAXpJnDzzIKJo612mEzo9X0ZeZ0vHqcdBJs85Y6tf0ru0r8LUoLIfVSHLCm47e
6svWsRob1RtiyNcz7vyYAT3PeSUSuw2hiBEZujnqKPnvvGqOh25kgDXjpyyrktmHzG2upaX9Frdj
NvieQD0DfM+sN7WA6n7MS5uBOG44d1J20OfC0YHNgDbJkXaJ5wTFLyyBx/+jypUTcMsVwys4lSL3
qKDPZSQzR4vOfunFGI388i5Zkyu1IeA1YvNtxTXdbLVB89lpNLXRCx7vpzHloTVs0Hywa34t6+aT
G2OJpsqxozHlM+qc1sWphd1By652SneTXoEx7CUK++MVfl7NBGeSYvU3k7/12Uy3r9mKmNJa9v0J
jAcZbPkdvS/Ce7UW5JHnQ70QJH37fcuEl80aTuP2Z6O7j/qCtcJ0wrD47JEggIUB4g7u0yVihbfr
/xg/EY2cuGU/1kqX460CU38yJLOMPBCbJnWe4tHpCnZmxAe7NW8I+c5Bl+UNn1xbqiPyKxcivnXK
cAjxNYIOi7hWP5RnE0GU9Sv2r6rHQQpJYbA1MGTdB8fQM8Gk8C6Y9Y3Ssar+gg9QHfT82DSNGHvh
0wAIh/6owSEr1YptTsS1Z2cvlS9ddJ6ruak4Sz62Z/JlWdKdC5N5RQrBJQL7LfJxFEB07+tq8GdN
b7FfQcNgiAb8m//qOPY4VVB+sggU8C3w6+hyehlWjPQIWUZZ0RJ5IqeapTFED0k9cBSahrlx6xH2
iW9ROndwUE982FtVoRZZS9aSBrmDpW2+eiOzmbFkX7+ChfQV4y+W72vkasPSjFoo4MW5nEvYuLeY
FuVLUCXmUpxhWo4spIE7kojyJyYiggMcbGm3NXRNxP+WmrOoI5E0LmnDz9Rj/cM5NXo2GrBrktxH
YDhh0rbtaWgGc6iLzPkF6ARdVxm2I3j+Y7uxIgmK8RPwNmMyGv6VArTA/KvK/bZFXDtsrWx+arjy
7cejRj4CMFZxk0N/ia8YsvzNiUZPJWPJrRJMUsQtjYVbkNF1WEeCjKgrR6L56NiW8zYzgfeIibYn
NnnPsNz1IooEMJ5AJJ9QImt2okUnUiUhxIvibxJjMKBliPdvuxsjJyhevgGhx1ymx7l56NbdgmGD
hB9bTpWeAkzF0Qozx7RtpHjQyGKYVQUKDDV2YDfbhnZ212KYb5nJ6sBZf7J0xRxJlDgxTY+BaR8L
q95cSN6Y+jkDvv15nM45LAwOuL8FCl8QUTuipAYc650AnwUjxcXVFCJopVu+YaqfF4WdrDup3nqz
0VAtBAcebqcjhNByI+7MjKP1Ggg2JYdf1ueHxsj+UJbBJjF4J7FwzUuM6UZKPfJGQpE9LrSR+M7q
5pfZPX5k92qpoLf3tS41NKERtuU8cm7C4I32FtnJyQBTE4nmFH3nAc2xnr33KT4+eckjobnklQoq
uPoFERcgpWjgc4ja1B3uFJMzwjBnHQYnzF2CZZI9oScpTSRV+KvDsmhPVh86qKQChxAQ/L3SF265
7/pmVc61sOUCDwwXmj0BGiyiiTNNWY03FFQmM/3j2jkXt7fhhhLFHT40HpoNo6d1RgoeVxRKqrwg
eAd30b9IEmRRWORHhUWnzA/nbKY3BvQn6ERMK/hbHDZxy6hWKzubuZIUd5j5WOBwdemQPsqxCJwe
BdHdWihe3xcVIjBbxbTXzFd+ivPV7/IjVcLqn7FsogflLvS/tXiOy6SHmdqDW0Yti77jnVJSePUd
ApgiY4+daVPx/tA7KRvDNjA+y0Pb2B8BK5VZ8eQ1RPk6BUYdSBrIE+ifKSx1ZT9ER9wCjggaweOm
Nruyk94WAtJ/6mHEmmeI6vRzvu3rqUfEGtZsa2mhKsKaDW1Z3NEoT9XUF41865Pn1rKT/e3a6eFK
NeMnsPDVfHRCROl4peq5CrIPzpoL+A+w2XMPOT4+r6lhwqv8NccYvlWN2OeSmtnYryeP8ORnzMx1
pSPldxHlh6SlQA3psyLT4vUix7wTewa+5xRsLQcCm3Y+bVuy9o/QaBpGZKFs4dJGNFCuoePlHSkZ
AABjXaxZQEtqa2klfVvvTc4kH+RRQ/NIHKOaf3nqWkxh0JMGpkXh1CjAKs9gUWA7FIBgDqHmkwYv
Kp+Cpx9HCrH4fdTdfyGxabFfrA3Ih54YokBN5IsO1w/otqtXF1RqDLkhJfMFtL53DnTI61Ka7eXN
pCkdENlSQa39mUJqfSR5HvEitnwEsSikYh979fpR7juRiApmIf15p41l30RVkGRL1+Sh8NWDWpsG
cW7d0PkRdtb5CGg62NfmE8cQiU0HyTM3NGOxjQBPGgm9GDJ/CpgwLaGc4XtbDSx+2g1QNxz3EU11
5zJPQG8+UUAcZ2Ey9PBhRICZBphQXVagWIjx+7xirTJh+XeoFxmzls4Y17Ow9GpPncn2kab6KsKa
sNjcNzFyQv+FtnNfyWsbycBv/UTquBgD17zCTHsBRsaplGS+PpyUI/Rmzb1ZjJ2BYaEShHE5Pmqu
YVDiB7czcGVe4B0g4rdnbef/Dx8m8jgV+5vVuEvhm73P5RpGZCQVZTsS11yyKHYQCHh7hJMUb0R5
Wu4qN1iv7u2trBqi8RJ8XjTN61Tjd8tlEB4lxs+0U6FKH+EiFF/YZgXCQe8mdnw3biirMDzHnPhd
dvyMtSCrS/j0YjAuVc6GuHjjyaNe63VPYjTGGLKSCbbrhQq5HyCLYB7X/xM7c1rz3Defqt5o6qyK
d0VaB3pF90dr7eYr1D9mVSSFAdlUXW2X0bEd5Axz8w2SLlapXpk6LQgM/BdwjPWf6XBXypaOXaZ7
5s341WBAzsKnMdhizu5+29HrxGuea914GYzYOgiP1gg60FHQ/IW4NCueEM0sw+whcMOr+YhVHiys
uk18i+Yk1a1ymbFvbILLTVtjNxf3IYz5/l6VaRigGdCuPUDQZZyFQAFLNdBgPCXAUsEOmiJMWPV4
VEWU+phlmqyWZSOEshUnrsQzhKrYVoebKJa0yolWJjJuhqG8p8vxLQWuaorIOmAAlERtCMT427ta
TtPRE+8/KCFWrt+aBRP3tszy/KWgJF5akovOWZD2mg6IcLlNaQtoFTwnXiyCJsCLoqJ9t/54sXmF
SE+OJqCBl5m5rBVgE23ptYZpdnyfRURO21aWu5xws0DY4c1Da0GS8M/7xtzZmro/bK5q3lQ7o0yF
sWigoN6dEJ1Q7/qdwzX/9FhCevBv0msYRKIXLBAHP3LwU6rL+0ETSkbS4qQNsYeE6e8Nx+yCOcJ4
gE4ebNTRb55jeMdCvFmsq+6FJhhWbAo1mYaQAUgPNjZzyhkSDphlbYYkzwuckO6Gcsf+wn3NeH65
w7x+Er6NrOQMiTjwsx7IM2ka3QnfkfXf2m+ZJQEsP+5Ok1Rr3Vjnk2byhx+ePl26cPGx82zGNA1u
LeYA7b6izCBdShZC0xx1SWKoxQHHm5EhaE6jrYcHwjnTtT8WcAVSB1yfQeCONq2mjXPByBzVmLf2
qRMglj8Bh7qnt138k8SCeGvmsIk8FBJ1Eowhhm4Zsu6BDd3iWC5WmC4lU6azg06d+W7r9ZegZNKF
uUtsFgBvW9OYvZgj4/5g4QmQCzgVOR0Vh9GXgzzo3rolYK7IqoQCMGqsMXA1ZCLPUpItsR10twMi
CUQhHPGiXRhZGAEfBHD8R+PiQefu6VesP5OZTSlYa/yKKWc/Ez1BNAciOkBYlFU2FaGPRX3DWnsc
yMnQK1JP42MmcSHgQLI1ipA58aSofHvz0flUT20D50HemnC6W791cwYRHWej+uoyhdyGfEnn/oDe
tf71ZCB4vh3ChGcNv167CskD+nTgukN9dTheU6ZOuMh+l14UbriJvVtIB9t9g+3UpqcMNlQRaDhk
ZRadQW7SXcD/9OwTLPYY55hvDc9lblA6Y9WleaWcTQ3IPBE42PF04LdEFegffv50nUsOfhL4P+xK
dRqsgteKL4KE0ZpvITmtMsngT/rZQeBugfGYFNN+ioo6XssGTvzZaJdPDnSR/4NdPqjimB+5ez1o
6QxEeq27yWdO41MFDL0LrdD0L6NDTcrARm+w/xF8/xsigR1eVJ+XH1yTEdhyETJ1J9GxUk27gAkG
AFkUc67JCb4xwBF5wD+cpfG8cyHpuhR3d5Pzz8Fz4Xx+CePinx/wvEWn/IdPMype7JN/XZDxSSsX
CckYdDubX9915KTGHLCGv/Fatdmn4RuUpXFEHQ0uLtgOjZdAY2479PwhVSQA45b7o32EhWMAiU7L
1w6MEUSRkf+JacARhDmI8Ayy1a24TEeHJ4/CMe9SgOAbHEXmqwAD/y5mHwuUYt1qget0U1VQwOr8
yKQVd7YITjsL39l3zsazyx1Rq4SHpGNCjA7kZYykJQ+bcqhg2j/l7q5nqHx2RBfDIEW3uIoFNmi/
FOnuhF/YiOuzzqav+0P868QW1YL+sR9mlMVIpF6jUkZH2x4OKRwRtc0zuV7tIdIzqlGTKAPtSHHt
Tu4vvuNRUaE98iJJIymb3DwPxBBgeOf2sx+fjkRKEdGQaWb7QnBzC9sFh72ln7r2mfoYPKB578tR
i/tE+r412N3q4bj1cz+w8mMu6+pvyjdjBPklcZKhlXi719+sC7eFBmrK5odvG3iKGCVXZIiMQwa0
LTYyx/L8enbAcTubImQ63vSrJDqMNd7KwO2zrBWCbwpJwKh0d7KQHEwM8EifmCGrah/J7Plk+H6z
K3t766ORJ5PVrjUHYcVqfGN3lqgqwtaD9cU8ygbpCbkmdq3i0SWT2pHmjg227KCM80/FpRDLkKEe
eAE5dzvSxZVVWjGDOW3KXs/KoEdOJ8mFqp/WX6dRK9uPtclh4bgPpqCw/4PebGcXnTZ9GiuiVf+D
4LCEFGyZYoo42TjAIJZz0sXYj5kFTn/thJNBTbDdMQ1+vIYAZga0PepVzSZwZBZFeJKIo12cVbHt
2eYslZdOh/7KB820BS8ocI2soXvidZUmwjxrbL5/uB0/9NiDWpyxKvlBkHMCgKujtfLDR80KCGeW
2LmZzO5nycvGrvgOfCOvmr4zpr7Uzm5fT0pDud3j0luo0zGaMxidQAf1jNzOsPUnvUtMpp81EqWO
wIjEzQRsCsQBBBs49VAvifaTtloZpdZHqs+cIck88cjAc+gRZzBc/pcoipGrp7RDmnjZks/eF0kD
psKaC7Gr0mRdOwpcyUX14ZNCRnOclybgCJYJlcL/1VlEtTUWn+Nx7httugLE3j9nbold74qEBm7C
lvvgSVST+PnSRvl8NP9//G0co4IFNobko3XlTqBRd1Nxbew5uNUJPRhNJfB+hBGg28vSAmgQykeR
hUgfKZVQsHKOt2cvaUpwZ1JvbkH3fOt4KqC8mArgdEWOCs44OFw3uzopy4bJMB3L1nLNPVU6TZjr
aEFhhmplj0p/rGWEwhKli4mLyXjDyk3+IotVItQXoMhjp7Q/MgDIQo5K3zYXG7iehYTOSqp5yijy
GxUGbaE6f2c/DOS+Y/1gm6GrPc4qy3Kc2tmaqvEUKe0szaDOXD3kI+OcCDzbsLAa794481FkBAXH
7BNj1beuJf4d1RRcpVaGY1Ye7uHA5EaqXbp7nBQgNhsnxVJ+VKOSscjfwNiX4Thya0Q4K/qiYk51
+jEupB2BOTcEYXV1hv5u/mRq9HzTQMSG6R3CyUtyit0rlxTitD4mdlXXw85QoU9oFbxI/c2Eg+2m
perWEzl9Z20ANyhTwTiXGyztrFjRkd2L7S8HMzNXJ1l7NebxoUe9kMwmauxvYGqNfu1LA90798T8
YBS74sS3l6STuFtX524qH0OBprPiZ+o/wxltiEVUIwAILWGBu7dqqsluoRJMAw7+P+c4AVYprhfi
c4iGlu6eN1HRaqaWW8vmxhXFdM8O94LIHglK3rgwIAsjlaqR0imHbdOb0Q+bzxBn9m8dn6zRc+VG
p0ZkrBcM7Uqbh7eyctA7wkNflRpL9BOsfuXUkgeYLlH4WjLAwAtZ6htqG7kfPUXSgzLnricqk0YQ
zZ/5YNxr1vx+Tt+yzEGkU7/W69rx6hbokVWwUy7XldFpVULb87swnypJdJoEAmiHKVJ5OKa1J/l7
/mSWiHddrA3aPGTSn519Bx48MVBIzN3n2nXINv40TkwlmZmhRWZt80vJ8OZAtQS2BIL/ZlPV9vew
Nn2xVYdeUOszYhh+BtcT6udQTSxr5iRLv/enU1taj7zUhPGn2XGlUb6VA17UezJZbM4inQ/jkHHn
pNMLCHsLuIOwRQUU3n38JD02FViZfRB8vrKmAevuDTQnkEgjAXrdhTSySE31AdNPWjgbjuYZXMVM
uV+mvokEL2UbmHscdimrV5fAiMDED2AIgT7WkC41r3rNUop9OS0aaBdZWCDt98yqmUIOBXDeLKii
gygZVTWKc8JrvN7F5ygI1zQSpUjuKHx2pZOresSdJQ1mpFD1J1eXzdYLuINyRMYujNjMhYW4OpZD
WZ4RZL6jn9kbG4+HwLYEZUAnTQGeX+EBMbURwOkl646H3vMLFnMDbuqIj5un1WinAFtNg6BSjVGY
Sv/7220JTPmLxbJZRiQQKdNq+oTp/L8m3Q3eZEDBqg0me3m9jB+6oIL7zu/hARkCZCUgMy94hkuj
9bdqEN+aoSwwUB205pmyA+oBrDu48KawzwP8OqTjqNzGuZWjF654uV8An9ZpDyGAZ03/pUYWKnlu
1VeMGIfq25p8k6B+79ml0Bag1z5oqpzFsj6TltncpRnGASvdYr4lsq5aGJhV3/TnQ9DN9624kBVC
ECIIXM6uwf1dNQbI8nS4cxJohDoJ4TwZEavkV8jY++M6bKwz2hLaQZLVFAkRfyWY7O+xxezzDdlR
0LvSpUt9W3Z2XqUHv2V4pr85jkLKSHHGGWNVXFoYPtz/09I/hnRSbVKGdMu/qHpmAQE0KdtHFmND
0k4R0vN/P2zjXRCaym9AfAO6jQOgmR+ZMR/VGQRlvRh8/B0B3mPz1LyHc9hUohMtD8Jp8sJbt90J
kFSyB+N26a2ATHETfpGQBY1Ia7CCdPXN7nbNJqGgRJMQKu2Ykc4+CzNfy7zI/V4LitexDtJzySAS
au5mQfWqjNAafxVYNs1OeAf3xZxXr9qgjvHrVhtub4B0ZPbMQ5KldFENB8JVzQ59+diVAu9PRrgJ
zoH9SOc68KND2Hw+PjTqFM/ypEvqpRNARyyDhz7qGj4PcZGhPKJDVviwVeZReT8+xE8pZtyI7crv
1F11ECA1bLloNE7e7j/mak+x/t/z2aSYnEeRe888lDND1MrUHRLsADyHPyFQV4bVz/sN4SQokLrq
grlbORWVz4rB6BayEgx1h8ZFFHoYdB9OuQRa1h/861iNOWDjICE+DnDYkGNyrs+NYDBiyvVuc/lC
+n3PGyLhu6xXzpByH7kUNs7ScwmHBZa/4wT8FV3nLMh61Z6WVD8YbVHKNk1xFyf79E8AdvTdYP6c
v0Lk59/dYQP2ZP+HlXVejivBOy/VEuy9IIq3QJ0LxKn6Pv82oxXv2AxZrfP4I9js/FN7Kg6Om4is
654s9pz3yX903jOOJIbP569uXVXN6uNQkx9oyNtxzbJdUs4rg/Mzev+8Jgy0aNoKteeldHNu1dcv
xfFfgHZZ3YP2Mjg6KCh7qdDxJE7YKZXeTRbjwn76otYctS41uaDG/2fgbHe5c2fV/1qCZdrCY4XE
s070PT/r3WtPsSaUsimu07KMZxTydCucOS521p+Jz2vz3Cat8vhAR8GxlZqg1PKo+fEIbMtTnkl/
Yz1H8l2RpLcRGTwNhRZ8AHGiZLms8d+rXyWDv5ZK7TPGBe8lTYBHyQPJl+1Fqt+Z6L5yQlK1wK97
giejFMUTvznXx8ypl+QOBbZuqn7JnMW1jWyTZC2KEtQptmH5TcR7tGN6Z2p3KXGcuP9acHwp+vN8
ikPu0SPPTioUc93pDvj1d5g9bSIh1f3nDtnz40wcNfRUpPMAGt7BeBpv2q0PETqBpvLbLIO4RAgu
//XN1iKd6cLdTGgCuLyPsBErLbGU1baqtZEnbL9zbFbOxlAC7J7tOrZ+W8yB1e+D8VcDPYWAildF
J60pRzhV+1xMQjqqCcPQhsn3VieDlet8ZwOWFYIe+qaVE/tSkYnkKbJP9SJuw1t1du6wGF3yI0ny
B6IdVW7FbsYf9HPr00Utv9JO3jKT3kq/ZCLSkuZoR2ZDkjhLbqzz0v/QvGokmFTqT93fB2QyeFKK
4DhddAAWg+5xixJs3xoJLbVEoIEty44r6Tu7ALovfVEfbDCZ2JdUDXqanM5k9+P7BleRQFSON0S7
orQNsk5ip5uLCAoFJ0/F1aoV74QjG9igALvy3bRDNUjuoN++jxsQMUz4lJKPRFHTO9AT1H/r4/Ae
9McB9ryobJfvTE1Ue25m4TJkFw0z3oJkNkTciVchiCy7FZwbgtNtPNpbJaY0TjTP6T0uSmv4a4tk
uq7jzgR9mrjDlnCMcOc3CoPhSRn2a+Jtw9jXDZjE+j/TmGVvR0IH4e6jpJ88pDjkTZeucWikk9gW
8lQZu5JRdSwfK82azByh7JVxxM22SiUIGSUkwA8qj5RQ2BDvXXpmEw2mrYwWwsd8Hezrcpe3Byrw
+s5GiJbUWEwywd0D1Q6DhNutSt4thr/1cFRpMmZ0CzNkEa0lCsTMhdqtPsV8cQ1+z7U+Tg7a3YRE
ElklBt43clGjeGI49TJMzO8XdN8I2PEoS14cHk9/6aLrTmskXu5r6//j2HJ9TMHJCGOoTi5QIRvI
Hs6kyiAexq3S/BiESNF4MUH5KqHsDsVnNXyDQvyX06QEvItPQIccVUeRVrh9IJ0g8vx/QaYatVRr
hRGrkcMRjrAtjb5KR29pNMMUDfLqZCrIglzuK0jitKP8gnsTCM4k22tc0fNAY1Gzg+PPgaQg9BXW
eAIZppbrYXAe3asLZyDZ/5wYQnW22ijwvW/a5htVkp1jsBW7j90CXm2c+pN25rn/l5Wm53zWohY+
0duOd+ThR54iSD+3RyOE3K74NeHd4AkQ0vP9GEPokRs3Xr5QD6x5QmYKXm9jiUQkhB/KyQh93W4g
zFxH5iRA7laToRyTt6CFDzAOrneSwKNAqkPTG1xGf0k/wDUhRJBkdoIebzZaiVSI1vqiGCk/jn2q
sRXYh1QY25l/oUxPOhD7LbHNSFV9K4wCUE8W9KFaslwTSqUwWKAWcb6tfiqLv7IL3Whcldx8o006
6bVJCeSh7cC8bxyrT48xo2goeBtmc9xPLs7edu2l2SprkhrrzLFuFdwUUSImBEvDRu2aEHnXKXWj
ZOU5YkRRLhQF1Rso0u90R+NR5Jlzx56iKnwp/SPkuwdgKNtMOPzyYHN/wFW01yH5zZWEqDiU9HIr
WRHhZsEGdRAKAmC2INwOk4nRAojpYbbkhe6tK8kvES16s1YPbJFRTywKtItxfrqa2kMiSZVHfRLV
dMdDHUF17B28KT7LeZl6LDO7o78OzYA4L7YFFhduYeHx3eGXkB2Ug2jng9gEIJ1nfFxFujAzvT15
b/H/kKahhTTsNZanR1K0ABU9dkqml20knsZu/hiefn323EHYqTXgTLRRB+1hg6V1hIiJAn1CZ1U1
98RAHADEjwIHQ2Ssa+EgzcQlsZHsjaIoy6vIh3unFEg8qbzsbDiw74NBCVYZPxv6mjwsegednaq9
2xVQQxHEEzF6qqmgAqDSiTIzt5bUyR9asfQMGxqkrIInj8daGvOklr0apsFw2Gvzk/8lGUhf2Id5
5J+QW5a7sYFfnIy+g4V5drVuKSY/kgneFfn9V+JTITZpSUs8qrnziSWJ+a+yA1KvZaPo7EdGjNne
i19oO+TD6NMlIWXhq/9SFxt/it+CnuF8t0ZACcoEt1ZLgiMUL6WQR/+jdAyoKqjebL/6Vvq8Dbn1
HDvAXOrcSCl11UDt+9pnGHlILB2AZCDwx/7zMBptKpQQaIaDBrWXCKsOtrpri1t0zqtzrZ6uqT38
2EvyNvnleepXrZAgMP7V1QbAz2m1jpxhq8Et0Cxm8h5Y7bq9jUgJuoBHNHdL+7Z5ZoAAu43S9P5C
SVlw0rKezW+UO1Z+VZH8JfRrxoJE//cwd3D9klxdTLdlLNg1mDfnglvdSMtXMjlGUE9VlafTraZl
ig58uXu+8Fd45/03Wda0lPzsfaEatpJ/n0N0JEvf0A2CmZ25BzCjKs+pANtPMzTZcBybgh90aVGv
dHfxYe7cScv7x4/aiCeyaovsct1e7KvurhJLhPhMe3I93jZRRnz2PKd/EbPmFuKsMl9XmWFXjOwA
t5EJSFaR55zl5GMqvpsQdhH9LZ6R9/H7ZopeRwlLcE4m+PvlC5DiWMc0Ssy2QNC826gqiOGlQTTT
xwbTiaGCDRbMgP9T2PtnTuw1wg3VbgepyN3PPQLZrbMi4AWs3q4DA7tO4YWFs0cNzo1C/JzKzpV2
rVQ5WyvKxTOYP9BmldUbVNH95SQQ1AGAdLlJnFwTeVtQdoygrpG+AwwtOtzx2Alj1RtdsYBgOicU
McwY7VrOz+8es+XmZuKCbWvKEljN01TDnuRYvem780dx7PNRFb1KcybIx/oUKBfw0fB65Id52Web
R0VmglUoJws9VezDXBC8+TDjyK1xlySg62T8PwACMbPFZokHQq9JslHVGzpnZ8Sm2jWUmqxstnQD
COOd9gKeBqDgCjF3czvOJdGG2zn4qdWbc+CxSdqkWFENmskF46jJdgZnMdlbezhdXckhq0JtjrG+
DIZvBbO864sNFHo7+48lHkSM1jsi/HxUTSdSp2VlO2LJxiG3PuZgsNpRH8+oi1dX7mt20GLLIhoS
Zw4zcpub+R3bl/RC05dtXYiiXwJXR1TFmwFOVtwUGNxQ7dg5bx+52c/D4PrTXy2s+1daDSqtw2V3
WB7c/PiaA1G7RlBmFWfJtEepG/1LW6k6bEm2TJz5+3f3ap+IOLmNITGo+anOWsYauOIak8o7Wy5f
gsqLk9Pi2GyC0YVjOmvqJGc66QVms+k3qpx1zVq+VDGF0MqjVYJ0FpPdbXpK/p47Lbdqee1R/pic
WomvKKIpARLegzr/axiH9zUvdR9uaHZrUfAoQZf+LF7e+zk9iB/NHzLLPaULmlpKCHj8gYErWtlW
tgxBEvuTS5/zq04Y5JyE5gwhH6oEzTmMQYW3rXUiQhz4RqpOkZnu/B/D6+5tek8p/OKpb5fpeLPW
u9hZLSof1Q2XC8L0T9S3YgiAkl+GtGIPwQGKhN+C5nFurwT8ziHxyKsLL2y5zaQIWFzgXMCOXPDJ
sE3sqLFQ+gP19vEpDwWkfDDBQo0PRr8BICfB0t8kKLxjPvs13kHZBZ2zDbI+uU+xuFFMeEPIULkb
3TyQye+gbxavBeyV9/8JiCTlpJCINOozc2gnruZXPIx+B/qZsru5m1Hrr9D9hEPE+EcdUVBafWNt
VrtYuYpENg8wFGomKmy4+ZyzADgwrN0v/l2Ay6WdtV+thdoS/PLr6vOJueVhv4rerIByp97TgzL+
6nhQwOqTkGDS2mX4nz8mK+78fNKYAlAKwwGfTxofHdicgHyCRThnQ0uGLT0yO+GIVkA1JwdGaku1
foGFnbqIBhnpfHZbt3Gp3N/b0o0dqdmc/I2sG/epHtwQ3hAUECfG5Qi5Q/8ZMms9g7gtGrsVqtrj
/9gGq4WsfUe772bGGuaGKlcYvZ0mcDM4HeuJAlAkdhfq7UDMlql4IE3r3s+TGl964C2NxMcXFkRU
fN+taWgBHa9D8YiceGF5JvrX2tMDJ8vBdO/ZWCu06/Z4SbxM0HP2n/W0CYhlWz//Ix5CwNjRYpps
OXuoNDd561N6ZA8nz/c/GJPntwglUux825rvGxnUdX4vAnMwK8w4JVwX1IuFbaPbqdY40Ueldr3e
+XnsqyqWzdqlprA6kWli2RLVlsC1zOkJm4kLWnlaBkSt54dSu7EI6gVQ0lwTauzzfoT0Yc4oUaon
9D2fUlbkwEbCeE7lbucoTimiZxCWO93e0m2xcIxpJI+rO/RNcJrqZU/xlROxJO3tyLA/iF6UuebI
cBYCAdZRHoJgUSIEOi0rRgofit7VBjodiTF5mTGHb0B0BjdCshSbpwPWH217UTkEcSnTvEtNu6nU
/7Q2dF4ekAyv0OKlO2qedrea4W3O99vRa4eLKHsXJ7nP7v9iPL3G0mTlB6zfSvMU0wdAwXZRgMcl
swYNe8/iM7wv6ssyTz6P1kfAJXopxrFQ5fOGyIFePKPwCZFX7DXGQBMbEuwmp6QECdMYMW1Z5Sc7
cFFCO7Eu4ZrXOkn0J7URK9UZON1yy2KrlsNR5dNEbhXBJU3T+D306Tg+pX4w8Ea3gV2sLlQRqd5C
853U9yD/+08EeaPG0i9TfooyIGikD+TvEtA4wA7GaDtFhX8usShqQclvyCjo2S1xQ/lu1xTK9bze
Kfk4j6TCgXOMmkFfdmiiWsf0b2NLInIGBMyJvkg8Flle8BouhVSEyRohJkSRCihnmKXAtuWgWMOA
lzi/yxhLUAp2Tb5rZ2Ptur49HEiSnTMljtmv/n2RizPkiXNUGzyKpKrqgH+i+X5a87rEULoo4/8T
/ypuMt+5rlSVSD/RP3FCnffY4sx5SdNwE5lzeEp/t6hBB9k+rvhtG/erPBF7DQBEqxSBaitEvqRQ
rUaxH9AfwTADw8Yq8pJ0tlD6Vq34N0lDUVajEtSwCbCzsJKe6Gg+tI8t7pmkdWOjQ4mY5F+fBAPu
DGShBQRAVL3EDe4O63aw9+FQjUIEfnsmL5G54jfdSzY4J3FbFLgRzoqakg2U/Fo7rv5CENhH4xGI
ZxQpMjFzMMoiIClBTZU+k3bqWupLgiDtaF8PDfYRIqYWTJjLq0njWBM8bTC+8BAwyklYjCIXkRtK
WRpZgT+RDq0avO83wH1NIyOkzSOzZF6p43v8dZMWL5taGtvkdcl8zkyhD3bP8StZbeuVKI3NeXtS
gudjE+dZnaRs1R5+1Wiuji+JLoPxc9uXwXCBxzJwzGq+HBT7oG0D2DwAKFCAw8Q5dI53f/2CPZfT
l65CtGRMoR8drLrlknhZXaD4OTs4V8mIfLjI2IRQGoE9rakfQoBE4maaqCissJoSvMwo52huw60s
r4qLmUW4bvlfyjVh5icrB01iRidvvGuTA/lGvZLH/hGPlCfLH70Z/cyK1uyONSn9KqIJZko+Kuzz
HH4XVf4o0AmBzHIISGeED6YrBiQsZ/Crqkw+nvJ143JV0HbtpjVWlGj81ddog/mhGYhINmEtWyGY
gQnXx2M4lgt48dqpH0kDeDCWjLi1uMCgSZAOqeRVOflz256WoXt3o1DYIwCTxBdsNSOWOyd0zm70
i+PMAPvfmvEK5B0B/i7FJUrYinEr3XF2mgejBhwnFv3toL97K8yFvmuZrU4gfsGw60NZktgqkk2E
hFoCj4nna8CFyWLS0/mxE532RLFcjFiFH/TkdN13Qgp2tBwylcvrS9NijF7gEGwq3Ir6C1Ak9xct
xjGykpZNJ1dCBmUZVaRp44mxXvtisHaTLwokIrNWFxHe2b5uF6GJlSxPd9NmzvCJfErLRxBm2oKh
TLJnr8IQ8PPek29dcSrCtY2SrW8lZTg6v5sqi01yow4DMxLmjoDyhkVPV0F8EvPt4brWnTxUnb8A
L8zROG3Ehh28nMyWWItMtl3UB6fYEpe76QlBacj2467j1NN/kvOJJjKfFEF/saCtYAFhuTEkcOP1
jSJ+dXCPGVyLHFUMKFQEx8MMtHDBhnexzT57XyAlt+lulom/GKdguCXEYx6L7quGB0+jRVYpsbX6
dTWcH6RkMvsDfm3CRZrGzqNoM9r5QuvFrEtsmN8z31+DkcL6jjbOVKyLfQkUs1ER8rIkSPUI5C5i
m0JCD9PqANY3wli2gGcuddz6hfjQ7kagX/3TKH/16fyAd3Vn5Fq3u34WVOuuOK0h+rSgHncZbQh5
DVS4FUif7dYmN/pCxEyS4NHfzfmWpyyJQP/brR66OoytdU+YDK4/t7yfCXwUXbYHqQoBLaUjlNzV
Bp2Y++uq/avO4XfztN1+R57IUOR15/mGurgPeHEtgT/BkssdEP3o6uRrDVJz+4xYh3WO2tCBv4Jo
TBmbcsCz2gQTRVLO61utHa8eZiMj3eiF6ZZR/fXXOkxcHAgwPVD9KsHTv/R8F/kG4Zp74fjZTXWa
Ce7S//vQkPsvImyiOAR5JlGDZiQHemmuldzuIrxEzkeCVwS0lLFMylQN1Zr8+MVu+a6/nCsSE1ee
XHhlZQayANufM3mliKTsEEXnpgkvOP65fkQqUqbjGdfpJF+dmBzGTs7St/xdWKkPCJYxol5shHKw
QJAIFkqXD6bT7iT0jKynFDYN28SrdkNkR5g/OwZ2GoIYV7MLP3aHVmcxP/GL8G+k7y3o1yOGa1ks
OEJk2AvC9x3fJZ0JkwF+KF6u5ZwQ+PgonVngggnbeJkiHbxgmVxqCSp6vX+9KXDRqXlCxSNXwayt
/qf000Z90jEmVsq49Ro1MAVrLSkWelLhnoxFI7+Gu0QnVkq5IiJIrrvb/hxVVU9KQPuqgELElkci
7v+W/jnAzahxdDfEXZEgSF/gOXR+byQzrdr7E/b+6KChPZPObYeZEVnlWBcNslj5RIgAWrUC4FS3
HtYJMOqsohQ3OlxSUluEtCyq47uViNoeZTerheCoEKL/fODksUfIdsTETAFD7uwxaHkXUQNIOa9t
UPdrlZzuiirDjPGm0pNh3A4dao8naW8qY/KWPTJYmxcrt8gQ1qgfyFA+18ElaAlNdUsLWnr6B11a
bfjDswlcgoBk1tFP3dfSi2XS/Kc3+bpAhzxBd7ySInzEzdF9PXUGUTyWZofBqPTy8dUlBzUWGyQ5
UGLJ2M/y0GdE7Hz5jtQv9rqQdRa5UhbBgFIYagAB5GPjubjS+wc7sH3RYhoNBojZgs305+xG+1uP
tivY1Ss85plShUSG44oN95VLWoEnRLHqX2NZmtaFmnCfcI3uzcnpIV12fBD8jLuihJE3clFcemcx
DLmfhJ00XspOlRSLW5MbQTxjU+kMcQXvw00YqaoXjpQAHmQ6Hc+9LjzE9/4Q68OCUk/ShtfW4k2A
e/ws4NDCo9f2rUMZVK6m06qtH2yONRQWVaWaJLa50G/pcxz77bCrONcjTHgzpGrd81nHRvz05GaN
W4Z8N+UG1V8qZhGVKfV+ru3TQZvIbnUha5FIki2qjdsPxy5QIt/do/R0vsoUpzPlDgSXk5NiYAqB
YruS8Y45GDz9mhob95ebc5naE91wyl53p4ZbvtI5y70LPM3RwbqFl+kC7AS3934rlIMsrI37XHUg
GDvO5AtGjN8g+M7ETO+LalhAnG4QC5555maPiNdr/4Dny0drxteVPusxplbzjfpgSga3MdYYDkf6
zngIUTivGqJDrRzrvIFPZCoHiUUzmWiKS9x70/+GFFfN04sUsdyQZmOSaAvyKMowMGyK6U23tnHG
+yolgT39CuS5wKZE2sGYl7zjqNC8sWmUHvglXDkT4NCdyIxG+uQUna3K3Y0I05Ez9i8tmjk/VkiQ
mAh1mdT8HrNJQfjXEgKinvxt1QKsimp+wRwjfjvktmpxEJKm4tfm1sFBxVRBP0utArFDH6FKml4Z
Pp58MFLR72nwJHYy0st6XqqSysHfaEg51HYcNCJdBdc14Rpl6rSQQTTi0vODvctLJahjz4nJPERy
qIb4yxsKHs/vCauJrlWQWt8uXaCjpbkC2LoPAfgf6rAXjo6VAwOgJaNRpEZxaiz4UmjHIYU53DP+
x6MC/ZoAnpBI6O/+6lJS89dUPxwDcUjRpeNbtHBFpApyB7JMIL8P1m+dhAZiXwqhmQvg+NGUBdnm
4CIZqcXYx/0sqvQaZrgovwEmiE/fAtA0yWDQRPZQgbRHHk9WFJFTmx5rZVvslaXezM02mz4UmwuO
/aAB1uA0jSjjKgSo0UdflQKYmNR4V6IJlPZ4Ndpy/Rx+sTaIW54uvnrugGZElADqYmPvSlCQW5ck
yc2aygNBWBQ+1gpMrjPON3AxFokJKzcZ07Ip3cQY10PK7tGf9C1vZv+0jUDYMakvMwZa9mz9sXdP
vGHZ++rcZku5xJxPnFJ4EKIy1J52H2i5MJvNro+ztNcAh6A9oBT8g607vgZKZPI+y8Zoq7MfdFLx
uRrewCuEqlPrPVdYcn8S/+Run9SYmVbccn++n3Z/nntn40Gbe//+JMzfsMMHoOrGAGgzNe69aRZk
5sgLXHNr0+3URbxW45U7ZV5xhI0Z/iHULM1p4sgxiGTsf+nBhgO50UX/Rc6x5LvZRipoqKtGa3wS
g+DByfycS028zTDiGKNZUQme8tz2XBD1xlOZH86b2Xb38iu0CwYHZ6WvXFHc4dO9wtc+ik4mQg73
ugSD4E/V5vpo+qAvF/H1D/orOl3AxcE6tENt4yJslO1T55S8IfVq5yWVOMITcFO/vyVEr7QKvppJ
TzUacmGrTg0yooHmCoJp6RYGQPoHKqLDUnDQXhEPTZP3jXNNhiGRrdQbnwkWLWCdKTPYoxtrZGtf
PH/R8h+vIoTVML1htj8RXwnbEmayfJfLdXT7kaS2wv9II/tH7XvK1I4Wbh5j7TKxHw7GEBVqjPTV
vuAkYc0bX95Zhd7lAlkERwlqS2L6XQXZX7RX8EozS4xF1tsS0jQM4SBuuSXiKrI5tPjvgcWvskWp
i45tY9/7iHEiaD08ARoCj0STgEE4Ub1iO0zQaH31IgtltJ8m2i7k1YRN98rdQoZTt39iORM4jqJp
9fZiP6XdG65JwlTsISXzwVRG3zTGSLQJZrpUgl7G3HA9ulDdr1n2kxo6KH1bOBR8/8bWB1vE949l
hO2lAbWFnQYqvpx51TWleJpmPxY2rluC2a6FANulx4PggM40izBG+PL8Kl+hP3NA3ih1ZEsJHIXi
O5ALnmA611Uc6IkbN0mOWb+2skBcOc3M/QwoqCPZmbQiJYCei64aufSAuWq8mNNiulaPHgGvFL+9
Umr4aWfh0LqbASEES064uARWQM0MppFEOZWsKnzkLP3AEepOia0X8YsVXVJdDNuf9zkveiv+pEXE
WC/+UqaEBJSllBWMCBkY0APleEDVtvys1m72Jc9rdqr9mg+suG5umuuiCWtUw711SmtyjrvkaYUN
tLPP4WMitGsi2KQUnPLdZGc05W9z4mE5ySr1nYgyZQJLrztLxVHcl6xcGF2jDqb619+KdQPpopLF
KCZUeVwoApMHPCuSxZu6XFNghbkl+wx40wcF+eH9STnYeQxla3UnjURHZNAO8gr0xnGBHfI8lN1n
TFt7nYarOekaejXqI2UjIc61AO/C9SvKRGhk8/yJellIPUEpkY2SgRXafIl3T3U3MujQ1P92A2Ac
PiGUcgwgEWMN/F2SjmeoTChyYL98/XPxgLpg5V1CG5AGQx6+KJfDTnE4Z10FbnyHpuxFnD0WlCFs
kZifg/IAO3CcIMJZzxe/cV7D5+cbDBZGJknSnuuvvUSgiDA7tL8J9EnauIuJXGyDnKiTDMgxsCjJ
Y0i9CT744nyKEn2kzVLGvVd40NAFy1oTyiP+Xh00HGIVy8MTUV95zdAPAHzTN9a5xhc3fIbsMZF/
AjtlghvVyFgr5Z5cMq1C9mfmH2BnhTnMYKM0QHAYcaQFgegbvgRbni9BNzWU5CcwtoUM/tvpOoUL
ONU37kdVTbEw2XJN700iDAqnwB+lsX3lmEidY7GUJM3HRx+H1dAas9/17eTD7V+JdbtQ8mfDadxB
NzCbDrEIua5Bf2OAcxMh876TN8B0Na0VqxYUMpJ7sfUsvl44nq6SKRxfNbAkA6eZCYXrXn/GTvft
RLHsB0b4vrVt4BbE/q8zj+N/6bEZY+KP9TuH3AkYrF8ZHXWkeCleGXvpTDJUKwEN0/VBgdZESOSW
UtJKFuziT5lzi6rMqgv2taXjeUu96tGFrtqHnhSrN6Ywnnr42/wXlJoRlNl9dtg56RtyeqH6Xdan
I0/z7MDXiTpaCXQHYd79FHsOBVeIO0fQFYuzSk+y5ePYZNm/ueRVbAKdgva1Q/NFPwMFBBkOUP01
ccxGiW/RYmN6jhvnC5V7ZnNErj16L7iA/2A0yorw80WanZ//N1HUwYyB4qliHT3lwd0YQ7ROBXxc
ntfLkFT0O804i3+ElwvAuDwfbq2gM8zzgtJE80/hIWOFAbTFmfJYAHJ8DxxpKWVknNu8UKMrEq65
t5EehzEJKU0dIoHIUfI/6sTq1U2npZBmqTR+KT293UZVtB+JXTrX0Iz1tQHVIlE44a9b84gIPmDu
5fp5PVmbafFaCGNtHPsme/ED9iKpIxzQHQawgrVbfsJWzq8eyjGV/OODuM+uEOked2f08DI5++QM
5UFG+nbQUtOqamvkFP/TEiMtGty44wIPG25V6k8y9r6+xYMR0UU2t+Memhwnwf0mSk4MwR42ZoGd
14DG/v2beLVXDbE0WBMVMhQ437O9ncPIH3B+HxtyzlB+ZE4p4N7l2gy+H/fB29FicB7BLkFVZlbP
Cyct0r9i/Mi19oApfUiPLvGMdmLfl9afqrhz1hr3nVaLQg4i8X6yQ1n3IjSwEoFwagPap6q99uNA
Ohk6gWadYHSyccdpu1QJJpy/jhPKu4kgd10zwmS9R3ysNpcKUS0yAi4DLbXbDYMlI18TdY683s52
QpdkqqrXq0foINMxSIIQ8Iig7JiQVjZLLopYcO8npZn7wCMf+ks0NZlkTde9ze/wxnbzcST4G15E
QhfnTpMqX8nikJ/y4nJf2e032Ctv9bOKGtnWau1PszcekLlgEdxfijs8iHtLeIaxREra1O9hW/BU
zjADPZPioFdyUC6y4pXB25VIEb6GFWSeuJnQPjzAgEWN55poOry+PxxwyzgZ9tOz2pXy54bDVerl
VcdAT1tT6Oer4fRBnvSMYZkWE/dPuvclXq1NcAa9rGvDrfWjg4N52PXTrU1uh7P3FQx17IXXSexk
enkfu0Z0233HzZlhcKdbZfwqc23UiN+8wtCFEEacEaC47Vbd6e6yfBStZeH+IuppP0cZjRseUjTf
Rx4GX66gVxU0IXXrsVaZCmzJNUzGOv4tbet12/eJQhMOnYS4hJWXo1g936/Ve14aQQQzB2PlBXIb
VvwdhZl0S0TGcfpqUk4lOBjUQjiMoIGL0CE5+xjDDZWryCuh3O7nWICtIUx9nqUIoqMClBmtuYRd
MZJuLytZTug1fzeK8HguuAUFKv/tzHpEMr4tYNsh3J8l7DmfSGddj41pfFQh1Ml3Vmc+kapUPEfz
AyptWd8nMz+yjiCKyO6gOG7inacoGb5/z0OkDUQCgpe4EobCib6tuDgPfcmLRxQ++kWlleHiIShD
pcwsz4CdfSGsESd2hEn6V7xZZyqX1K2YAQJDM8NAZae4xl1BKpJcvvDMjQy7g5FqDWfODUCq7G4G
31RtFNtYCQ5r3aUzURc0mCpB1kEiTqJwb1/kCo2n/fJq2JlBVdCzIcmpOGUpZvAPPsepRVKX/WBH
Dptl5vhSbuTxVefGBozaAucgwDiVdppM+wTYT/b9ZKMHARGgNUN/0Wc8gwDeT1jLxVz/j2UwgDPF
gm9dG8rZna+d01d7ysmG1sHWO26SvN6kSebkZ7Ur9ePAoy9cHaWxcROR9yK7OMvC2PsahkPn4XQS
HBvWLs5Db3Izzwh2MvmabmM8pcREqJwNZuQtNMiec3u+1g/t6q6zbeKVYSELzqVFbWvr2+B/jb17
luqwgyOavDnXOvnRNKyKcS6Pbw+P3F4mpCxDJE7amEKDwlWi1dA5VrwV8lIRsZwo2sAF5hQUb+3B
s8v8PGbIEkjazO8esmoUI3+2xYkYU8poH4++y3z8Sqe411kwSg1c5KK9sTU7pkpKZmFm4QiT1EBK
fAzz1RIIVtmNhkl4S9E6Ufegksj4JfAY9q8NUA9i+vh/0+g7SbVV8h0cPlWoF6y6uMw/rpgmrcaU
a5c/2AYC01/7JpbzO6bYA8sKFOKV6LqSQJNqgLbfgcSNfPiOzj4eWKjQ9kaB41YckknpPp55ME4o
gKS8+L8Q9W5A2npxOc8MLRg2RLQRd7GAxharg7b/lghmm+9qmSznRtUATyNMLRNtWOJYnzr6OFiV
PRybRSqqwYiDiBczhlgKrZmZJI1rlfQA29/XkpM5wlA7MUYQZOYRUwdsT3p4a4FicqeGINtsJMcJ
6/zB9y2I1IXjb0bA/jhZ6J+6J2NGO4RRirGhO4vU78vGbE9qd09lzG28ZKtetM516+sdy3sLSb7V
gpUpUzMWDXmHu5LC7rS2EdlDaiRRSZlCSCI1lGkLNciGFiYBoawjWA8ehmtNwm5A3bLQoFEvM/4J
hu7bpz10I25Nx8uYdw0x687GmggWP5X3NAltESpPgi2tzmobWhFnV/8KKMyrwLtawOCYRxBzyl6O
WoSxw51Gap/1RCWarOjlvOJV/Sel8ELcHz0oSWqw6A6hQrkpuY5g8SHbK+/jWIjmHldTA1w0vvBJ
8o1GrAUZ3Hp4ri5SIRZH952MA2fHprQae3PMVz7QL6ktcLClTa/uVCIzn2Ej/bndvSh4CDwmtBzc
yzSBj6ZigdZI78erRxFs/SBnxCASAqug/n92r2BOm+XUCH/sQABlPmsjAmc9Ht4wycixdz/7IaBW
CEZCTXZ/PX7lrQirOEZ/pP2EQuHVWZp9lEP0kMaBy3u4k5TRs/GLU5lkM/LmohXuNFQ3v1mlghJn
/7qcS6Ka2ci4CyI4TA74VbZKH7+rea+zatal6BD8c26hNg6Oj9SiV+x/5lBI2spEaWjqvbRKhUIp
MsZLx3+uBM4DRYxNGQKoyEfeBIYsBzUh3iQeXX6FECtqrQGDUcCYT+Y3yWUdGCmwdKYJMiqnKCGt
CIiP5INzcOtRR0UKVdNXMWMwBsIv907GbIUC8OhUpwr7hlnxxUDCddtbKmuRrjr2AQTAiwaGxc38
d0PZyGwhTnvhXed5Vxgc1ke71YXB2wyN/JkRH0kV94YXcsTJw5QQzz74RGwFhmidJVr7cCnWv+If
63dMA/T9MWpr/60DY9HvvEAFr+MMn+spUIaAjZctFHrcXD622GCrhzHOMpRnWtWVgoI4XdecO10l
MtObLw7JJWa7A0701JqT4iZYYgwfBl3+hnZt9uF/BN150OQI9MGXIbcEcghaELVhJvvcIRe5CWNp
pJWm+zvrfFF6oo5q2Vm8cI2vGun8ScQpOSwLFClrhTMLKjNxSQj3244OpFxCh8bzxLb+KcZG+72T
yR2s6lU+Ra66aMD4Bkju5IGRglS9U2ZVub1njWvgm1GHBJeQJG9Hyc9QRPmjmUH4VKPcDhw3mbwM
F7rFroxw+CulQrqz1ollXWuw4arLyIRCHDvInUnqfHf0qSy05aehGIKZ4jaFRn7zT3NEAVQsAAvR
cmuVTLJ4V4Ag1C3fWwozys6mMLmkz8ExwZ3C7pj7P2KRnpptmAVSr9hdoOrScBkDWj8YMsT8OtE0
TjbANKd+nfAjMj0FFZQx0X1w3YplsM+dRy3UeBFu9K19CE8mgHnnP/bEXLgy5uV/kGQ1fZakyMwg
V8k0PNRkAW81FHo/PUycnqZWr/nvdUBqmb0Y9/kDf5jq4XrToCZHtEXbmhAAZBtT76nI+EqOsDqf
AAtNEtVSJgSbFZcTlqCxMoh27mG9yAY62k3MLKB+4WhT7xOJA+RaZ16+D7up9TdKDz4t5i76HK0a
9CPaBop+x/zsKgU215aE5sztOL3s8iTWLjNsmyfnxnf7QCNiFcUmJDyJ0jBffiOEoeLqoGdc1MuL
aoKQeIakLa6AhCfRTQQkMmYrKE7uPE4vE1A1+DDknPIZQz0JIbnWZeSPLpcA333P7Ytl8elewRzP
P9vQAPT211zXbbbyyBM97a9dCuMn7LfTmwi7hNhPkVHua3PeY6DSoNL/BBLjqfwXBXvJUS1ZdSnU
8WyoQzsbLf20yTelv2bcvuAWlgGNB7mOFBp4LWx/QYUiYLb1TPDaVF1OmdgZnwJ/HRCoS8c13xX0
YH1lcPHFB++uczToMuzb73m3ouAFYGPl45HyXvrU22fahaairPKv56ezk03eBJnygpxcVWK2a0BG
hDFT7ZzsUpEBI2egZLStzZWhE/o9f2m0bQ05czlXTNEALHDM52/9bq0mB5uoS7cHmvSsKGWhRTMW
gh8obl45DZvUdQyxyHLFe66ShXT4VUeDBah3I13VQR7zTgGaxIlOex0WnoX8ubAZ8xUEu7NQyeWK
ebr3Y12X3Ad5EyfFS9b4bEwdy37rG8vYVwBv0tQIctZOrKJEq5dCauPYv/Q4x87wH3dNkCkiif2k
UIbDxio9sNQuhDeHqBh58jGqrQ+z+v+h+H/3MIOOhFkEpf5hi06k+6+D5FmqayZ3pXdPShhAo/h8
X6HwkTLi+4JZUztgrfVHTIL3DZdiJIZEQwCpiuov5qCYuzFJJnIx01h7YvsWwSaQoTaIh4zLdtlJ
tLamIXnMdN1lcdKNhwR3quuHSD2cDbUvgipwufkkusht/9dnAqkMB09UFOfHD/mdMjYKxOGRxtY1
4WG1BEV4glYhZ8dccDutOkc6YLM2Eqqy+/r9OjYU0aNda+jQW+bQOF3nOzkgI+qGpIZ/l6izc2Po
jT8EgnUV5TLU3aJcR7hk4+MiqdoBN4FQxHtlR+o4Q//DPTohzet779ue4r5oBtUU63BciOLM2crS
o+ykZ9Ih6vQnX2vYxLgB9Ldg1KKa988Rl/GtgFQkzMKB5O2CEVYGvShe2CvECVMHJwl+IUBun2ZU
MF+MSnNHJ+6EwcNk7GdD/YY8yhoRhyt1vrtKmAeKb+ZFxPFulxBjlkzL4M1S8bxp2xNoON7cEkas
PN1XkRs8eqe1fW+Iq8jRQyQ0pksveNX2UwBO+YzXZwTAnhxPpSUSChjL/iCw/kkmC1PcdNvs9W0n
aSi43duC0wULn9yBPXHJRpOKUcGbIRaoFz4uoqGsR9+p0y+Y6fkBYs83lcj7MoWb6gdmhcU6eYeY
uQjkc5h7v8r+RrX92oYeEENrqLe5hyBNBWiRQdrKF5kIGCDDw1BFwIRTzSGJK+6SwDveab+Oa3wQ
jSpGgk1lHIXfRzpc5GVLhBERgvvjxYVY5S7CSeUuQ2m+IMbTkO4004JndQTOXuhj/8xNK7V8suIk
10XcmWfUU4p+eaI+HwXYDMJLPgFJCmuwMZ4HBSlFkdrtj1kTtO2EMdbhM/qbC0XTPsm8z504hj7v
fehRdqdUkS5N+GvrFdgFAs28UKVS1cZGCoy/Jpg8J4T8r7+0Gti3ft+kfkzaFER8Ud/FMBrQK9i4
KH3gGOO7o4daQQ6V/rZ1j3SkYFIvmjZUxOxLWHCe791UQELfgu3zqK9AIgEtVJw/sX8IkNq6vffM
cc14gDGdFDAymmUM8Tv8mn3qnP7utBrVjUe7+BncfrqxfL2dC81VP+EjxnZnTCb/Tm7uuKBBla/j
U7W1Tm1pjS6KSzf5Dsf096sQmWr18HtKtgsjsCA21+l+B3RDvnBtKbdZSnXplPwydhwAvQTbC2iC
6U7FEgyOkBQ9xnvTZHg7OM2QrgkwJikMbrg3X7B0Mxz4fX1rq9VLoxtPGTP9OW8jQ4SZQGTcoq5J
iBZBkVxUy78vW35nbJMDliHNPV4GsdURGRumRYvoEkMZZfPcZOZNlq5FA0/aC5bK9BD61Tf+uzBb
F288HvOEiAwfeu02iB4R2RRK97VZhjeqbXsAiuALV+jfcNTgO3ubGzKyhClyx2bfuQ9+tTeLCd5+
xFIJ8tCFO0eddvpcFSc4dmBwAGU67sl5G4MU+sO7kcK6zgGdmCqGR/Amf8JxTJHVAw4c/uBcRZ+2
GQaIWYz5AJxfevuT26lfDe65UPYY1wFvArgY9/iQrRcN8jY/jAi4jpBf+lrpLwpn3INXAmBlTOt4
6rh3JoJbqhlWFjCxW7q66wV3957vscshIDD9L5pu5Bt4xeWNDTLDTJlMwsc0wUYcyAe4XSePA0bB
AgUuW2zVrSD7Bv1pPqgwuMuwkipbIyncn1ojjhEIF1RwGQu9z0bjw+ggDC1tJ44Hs6RFH4Likjeq
OPVXRNPTwJjCk9nMW7TaMtxsA2U28mCAkVAZWZairmwKdXpTHl5QlXVXejPzuVjQ0D69sO73s737
ulbbLpk8wMLNMtT8+D2s2zAta3I/9LM+45aNMuKpZIfmVq6c0Pf5BpaGpCSDMhUSI938CetgqAHW
ebg0zqNj7GioZOs3BUpb4FCEcDbqmtfYffkqt6jiSFKOg3yOKhGUEpNYpGjGkytPAJFBjNyswk7h
PbjqsdwvUEdX6MhlyAMREcX6461QzFGBBdcKgvxBdv+EWW+m12KjgfQ7MkqF3k9LjIStr2Kkh7uv
shV5ApRW+mzreryGEn83eMn6TyHpIvALjcuzTUHSbipiYM+fNjT84i28WGPYYIkNt8+/V7z8RsQU
7LsyGEdL24UxBL0+GL4ZWxI54EFsUbhMbwc7Zl1aEyAn2rS0OCrR++3zQHdF+b7W5n7LV94cdYnB
vtIazvok2x8i/WlcEJ4Ctvygp9KHZbsOMyu6rN2bUKY91+wv8+/U++Tku533q66/o9GPjNcdrjrS
cagjVOGCz2PG4iMdhJtNzxK/N1qVlbKwAxfYkgdwTCBOdssiBfff7J5SaHXVURsP/3XlVV9ay+bM
nTtJFgmL3rZ98O+35QeerqgEJ8HHvcWjr7tClv0sX9tVv2/7YLSEuV+ahPdrvO0dPxv8E/Wwrpxq
axtemFKYgm9NcrQlMP+p65dQ777iQBqqHMyH4QQvqro3ngGiMBkal0fb/ja+f6UZc1KReDdcjpOE
/kxStMhO3j30B2HEP4DX13Hc+wrda8Uzu/RSvRUE/qVw4j0KBmqRKsubGMzrm5fn6AJp5aVXHo+C
eVy3HMmOw690Cr8lZ/2U6P0EFE0aYr5ORwocDATfUUqP9KER1OXQW4L9DybWkRnpPlHGO5dlmGjN
kgbcgyjxUCAtpV3xQIUTj7HZmBOImGF4hvTvufpiKUisdR/Rnif1rk/YrwyNZoCjU55idscJsba6
xnRy/8oDwrUdBRdgO3xcuyoD5+m5VXaLodwF0gIyl2zvMfl5Q3LLNwPynz0AGtFC1DS3LtZMge7E
21hBb4Fu1j7LB95Z+WMssZyg+HN/VQcoO1drSphFBn48j3x7ojNV56Yx9DZ8pkTZFqGf0SgVv+CM
Xx1BuFtqt26Gnpao3wKDSP7WyjX3BmFIyZ9s1UpYJ/npdbdfMTah7Dlor6S0O3eneoc3fV2dv6fA
DY8zzrxKbe0WbEZQRADhjW+Mluw1El5WIqHt8yHhnUJyf6cLGVBRaVLV7T+eZYV5aGCLgChKZV2r
s0JHYCQs/vH1Okm2pOIsR7cOOjVPCcCI7Zv4nvfPtgWxo+oqpG3CAhYB7BjytrZIgXDxq3x/em5P
jGsqPcxh1HAW8/y1JCuzlH8r2apGhNwbMhvBrSItQnOeDveEki9MpZVZzxs6VXCni57zToOvdOhS
TmUWKPwpf5HfsBLLFG/pnOvq/MNfF60j4RC4L3uskZfjngMqhDDUKS+rJGfj/0OFFZ3Sc8YAbwuM
t7wjFTErx3cDnrxpD3Hz+Ki08JHe1P43S7pQByW1C5vOqx+e2ng3GHj98CBzWFBsPqZNAoqThdns
gQ8lCj4bNxkRrRKpeqgQLL/EZjFJ+V5h12o+L6CEDT22voNLO2dOXOtSTYBORnOxngo7YKiBuxDP
bSi0R3qdPA4zdaF/jBLTGyt/IPmxzaD8dSclmGN1viBLkrzUoptKqhkXiQXl6HbPSQxnLA0mK39F
g1NRkskTIA1Thtw0W+pCMnsIZLe5pdv4KSnXZSiwKsexvhnCAYF11D7fowsqvmGIyzml9G5qqkaU
EtrUx8YRT/StKtxqowbUwSAVUYA2eI++UiVnR/b81qNra4KqK4oDfnFxtcIb0Fes5wGocNP93+im
UNb3W3thvv6jJUHBB7nmwuT9IlsNl2o9LyxamyW6npBctSSde61pkF+oImNOhYvO/hcJ+UcSdt+D
X/U0mEYWPuFAP4WiLBYz81wtbMVLJD9co400v8wRYQbpvhTaGjqtnB3QX9GlxSK+KCuUfIgwZGKU
UprjKC+9MLuI6IBDtsoPN649jOQOrXqEnskrF37IJTI+HzM4Mo/BQlCg9EyfnaFK73QcF73GvCw2
IaN2NYcJ6d2A0oOQ1ix+HrE00ksYxl9sb0JLgMKnT54NuaarY2mUrIsHQ4PLsJvdgcUjyLb7zojF
FPCdkmE8E2WPTHleSynBLCyQt4WA6giYx4+bIBBbXLfse/MazwU6YoqYKd6zXvwNPxRQE6ZYl2FF
wIrnKDxo7W6WaNvz4I4nheMKGL/tbPPoe/MT7mzjocOTD5AQsYXJlLgXnC3TvzdKIBdrERtmmwJ6
HiK4J85iUiWAd1HEamSy4iH3eWke2Eo+1x+fgWjq8abTVn6tb/VkzIVC67cCmEFWf+zGiSBTwki9
Z+fDWWoVlWhTfBzNjVLe5ChfjnOgiMzTX0tXB//QRQep1sd4zrBHk5vQtJms6Ck3rTrvgL3YfXji
0PA1FLQqlQas2Tr+S3EvBftwbt7jyYzaNlSMJpT0kzUqeVg8aatlG4bd7sQx0vccdjlnmx/77vnC
bowdBscJWK+T1HopLrOoupE/KAe0RHXI+qkoel7Hq8GFObRKsDeeKsWbM0OWxFKmlZkA6SJpe8ya
RtJCLrqq9I3myVwxh0zzLRJOsKqGEYaXmwQcrE03UZoU+2uRLvKGp9mahFkoVywkDKy17PMN0YlJ
T/KK6Vs3xDC25Ep/gDCx/rAboRSDY9Zmf+pPvmD5XVg1dleK98IK63GRAkkyEMotYLRdmVpNoDUO
NTKBJzjhjhxwjr/KCbtsg3i0MwO9VcaThHC9L6VT5POGv0oi3Et0RhKn8OIs6EfUn70XEejvSg8s
sqRZLYyUpTPvQ+r+Bhrz6KpfFIeeazZXDteOYe4I4CjL303qi64MUdK1gSoA0c9V/DdW26mrUXCR
WliGfoveDGGbrh2qM8DdwkqR4jI3PpgaMF/iGYjGMiFUAm2U+Rm9jNnaHgazXLPk5jE52j7Wrr8j
Mv1SVSFxeyGzkrEoeyWZf3lgCsLVrzKY6gou560PrpIj0prnDSbDyHs4RTnDzByXPtSNBByPu6Tt
ORHQBXBh+Q1oiTrtuAezwIqcmSuSYn9L/Mhl4S8kVZmoyTtJnB+5n+7PP4EUbjvZ4QODyrgrcIJv
JYw/K4ACBO24ptqw1Z+5npnBcAVtg9dJePEvg3wsQNOYzu8+O1uEjMiGojN2C8Rnecui9w2CqVd+
a+W1WAMRctFZ843LnAO4DDyav2oHerrcjLElxZCNXgZ7lv7QLYNHZg7BzuhXRxT/5OjUZd6BoUHD
8jAJACBT3E6Ss0yg5Iyxz0svXm2Bpv6xD9jXOnQ3UUpw2f8wnoiqj0EHfavvgYvKRr/2wBgd0DM2
EfMxSNSN1Wybrj9B3RW0gP7MsjiPAwHZp/EV9V+ZcOZK5wZV2yyO5GYx5kYizxAJJ1779rA28FhP
sH08LbJpGWg1V5dEYK3JvmjuZm4wkuIPyl6GnXBPLamvvj7konzuqPah6FFSw4HLBhjIPbHeNyGv
4QQxx/ubTYq3MAb6tddL+HPGHtFii7rfjZ8D2U7gawzlszR57uJjUmwx1m2GWgqx+MwWLk0uhbJz
A6hbkGVWDchDZXjaT4lo5FdJ+SVll7JFSSCH6bA57/xTMD2a50NDfSztBB1vUxluCgHRKPArRWRy
L74mtCfg5fffe5lh0QewH2vsYA3kKRxnVJHo42mGKq4ojMmI9dHj7rLSSe/iblImpcEUb/fQdraT
yFhTMZyu4sHwPczyrt0qaqSaKS0tXCtsBy9kaQTdGBtShjX58EZAmhFcwiCOYbh/YccjY6OpCeCR
CyR07v97NoS7W6R079bnRd1RrXTdPw6mK+mg8tBShkFJ/11XUrKpIDUiYTCPQf4MhkjInXoLRROZ
tMKnmmQ5TpemZCRx4oHX3ioTp/RP+OOwREzLRvKtYUeyfH4wfqqe+CqH8NL8Kf0oJG5SqdSqQWOX
1a/wYCqhL1SV+EPwm/CaVhd/1JztYTC4P+LWTv/PHngr/2ofCZyx260eg6p2f4xTvsA1wmzdw2eA
zobrIgQGGpZcHzwYuccmw6ch9GG/4gHz876y/cPJrYFDI7D9q5nLJVTbWY1Gxke9kC5fy34WCNAI
tK/waGNENRaGTrslVXzGEmKn0oxkAFAZAQKd+kp0rASIzW7X+9qXkiF0J4tAKrB1xz4TQ6ErouHI
R1yKTLjhFxxvjWMvojVoqlQDFBveMeobzzmXuCUJFh0QACcsq4WQ+/gsGPnvs3y81dS1Aj4HzG0N
xAkLAYqeVVcUgXEqCBB0cpwlr4ubczXLO86bg7EMBd8GOuq+tF9Qh7/HR0nU0+7MfPqRscxaxt7g
l/06XavhBJOViXNcnr0NWAEDkeyZuVCk6XZkn00gPGsl2TLorNNskNDnbed1oNstu0b4jpRWv9Tj
gBeHd41wcjhbnodhcvrgpGmPBoQh1eowHinh5swLHSEkm4iFVaspVBlJ5QpO9hUjl4JDOVIU9DAs
h8gyvewydg3DlwyLTOrbGKKxeBJx/aFBkTRIR6aAOg8689CiimaCSeSyEMGfNIq8SKLJFzvlna9p
dydHXcvFTp6w0roKEZrssOPBUUeI+rvU4cEsiW/PCt6hgwP9gIimldNeAfeOL5MBcjiNDtZVBULo
hh5sbXJ38zk2BqbwMn2ZzGoEOynieBzEtDQ1b23I8SPRrDATpRN7AfsPF1QPImrleXVTKrCIJkLk
R3oJI/F5QQQAx6UFmelr+T9HJQ9XzdmxQzQxZQwgLiKMrtvpfgt1F0Z9b34UUSxi5rQKPoQUQcAF
+xOgyavLZW1LwpKzpZslMWcA1nXPsCXRktgvvBde9CNEqnXfXYDeIaGqqGHrc3PwnyJrvf54j5EG
z/P+vPVa/w9dnJ6hQ6YemWhmQDbx2/3SdbrhqDFLxvUKORBLXnPWXv7J4axar2JWg9UvovfJEb+p
DRsAvBi/8Xhjg3vG82hhAGuMN8yhVBgUMKy71e8aiyrrp8cPONeg0srDm3jpv5ZPVk9G5iGs6Utx
c/hX62ucw6oXjEWP4LI04ag5/5OhOQailn/ZK6zDsQ+IdoteQ5EMD38al9la9lCY7DaqWtllSQ0u
FEPsge3B8r6Kab0iYbpR1TEv0fK8kPm3dlYUAubfmYInX/XlO/ube+0pFRCB6I0nQ3CGSLMNjrQr
LjK+xx3NXYNMjwOLvB+bLNgyqLhphmFw2Qyng+kmMRfk21ybAckF+6hUt7vJ2eN7SyfaisUkFVcb
XiOWpOelHhQ6tM+/PcpzmLhjsTCpo2O+OZgXns7uBXgO+LxfNHzIZmT4FRKJMp+OSRtY7Dtgafwi
ElbjM2r1X2EeR6D/VwW8CwfkJdTJFw7iwTf2Llp/+SQnNSWWkQaKP7gs8yjOe9iRbQUZwQXmCF+H
L7eENMiFBqQoSPUQ8zYXwYn2854IVTA89b+XsJd2vACYhJiDZdLeG0B0hqAl8fH/qv8rkxz8pzok
bLezwja5EOT0NJUdl8WPKsP4c/b+0DIS86G0Y7feruWJjZXHIVDUfY+NOPbJZgBmjOihyOgSKbx7
NbWN93bM+SUalqbDnsy61YYM1nulJbSpX78en4tJhieiiZVGeRncNr7nA+/0vdkz5wAFqilOafw0
z31fo5rCTgtZXpYVtuK4XW+F9rsFSlZfagMU57/EGRQ0t3i3kgTB12CVrO7zp4kyPNEtHS6TYKaz
hEERdba6imxFHzhc6HLulgaF2IAUUL6DnSKLwb+RKfHPUHK6QrynhS3m7XCwxAAFnRPleTuPoB+5
1WFHrh6QHbviYUJkkW4aiq10AZvxbir49EmhTdLTXFCM/cXj6JMKS+tn1rdtBWfbEsj5t36UIfEh
KyNjEqhNDENqeWgGXwuRnb63a+orFgoRDUFDJBOGcdO92cDPkGAoMQ64oU7/1c77R2dvhiULxAPT
ZDcNB6CfeN/DYjWXh36tEEzUPahTLm+8rtU6uf5weQhEDEmNkWVVgm4JN8Rf5jHBwDAbHNFTSRhd
Cy/PydKSkDNQKImntGQaxLUdd5KeW0/1rngj9v1MHml5A11jzsOnY1hEq8B59hJGGZc8T2jx9h58
z7r3vsAPG43tqjFwwgNLh5Htv6Tn7pYz/nV+dHU4kZQkdGp06t+CztwVhZLnKG5TctDrA90V3aU1
gsTmzSuRR+Co6jcdp1ksQiXko37/R7WwydaG84K/+4AP43Te3yp6ZCCOZfgIMbwKZ0MqWEfM/bNC
O3Pp/caGcGoP68DyLqP3crTmmkxmnEMVwbOIiivKfhsAXhg/hqubV+66+33JwMwzrB7xn1YhQngZ
Hi2akFFmgAvgXj3dUfiTtEgCVjPxezs4ebYRO/BI5hEKV5uWCTdanQy6Qc5Rcg5CQBUv7xMoRjvi
nNYJxgxWph2baSfLU1hSSbeee6W9cY3L0QD+/HbAGa7kcEOATPWDPGBfJK/sQ+7PNWJC/PH2HIMb
P1d01cH5l8pk075RT5YsGy8c23xU4tHvWMot8Jtast4qmjMqGCqi6hVRAi++9slcq9B5Mb1sMpTB
1eI+m5HKxOK4E0XCzK1B9vWhF++0c60cpm8cd99jy2skiyk656fqT+GSXG3kgHf8Wz5UOFNk+VGX
KSCO1LW4a6LaG7VrIv2kbl25ckwauvUidfKx6nv1i8JnuEWnRhazBziqOl6Mex3sF/nwTnkSi/50
aqI/sVQyU9wALxKRgXQ3QQHkljBkyO0q0nq7if82K9OBk8hGyM+OBdeYCQRh19pIDjXVDlXnGnOz
04jNcPvxHYF40yI000tC7554fglny/9+8+kcl4HOEQckhvaJOPDJHGEo3psjaC49zmdUC/ip9QCv
w95MhoGCsfNDkrAEiYGcH5zrC8yiOsNc3UDoY8gIsEVgXMkgHfIF5IB7WPdxCy7AYunUmg6O82ZF
ZUDL9NVl2OQztc4EBNgVa318FfmpXRugK7olycf7An50wGxvu6UtOU/rmOhM2A55OoQUlOc3ko8n
qwjWqw9GcIqRhOCiNnsM8fmFUwCXFLwHfIt625uRZwn2rFRNXA/MmWH9C49juFBMbbHCTCxiOqVm
6oYM0TwlmQ9GdPpETlhpMpqDCXTKsFQovqp9o08I2R56CcW59UuSR7nND3qIE/zh1P1XV5qTYczV
RPnaOwcVaZLhGSlucqY6EAsbgPOjKti+BafH3BWg0I12E8PpUkN8NNFDq14NO6XWS/v3216leOdJ
f3bSdFcWR0IOE4bg7qOZhdMQhjDTQOifVXsQ7BBCWotZPTzwQJTIu8/bMRkSiLi7UgvIE/MWe2os
QI7tqnmotgeCaJB9O1x3WL1tg6cbUPgoKcPcNSFaTiOTDGqVOA0JEqPDKH/I98Y3chjf4FBfcklA
t2Vt7VCHpAn9QvMP5oiAXZC0k/Yskm8LbkBdPmPV3J33UI6BSyo3bBl7UgBaKDtUDdBXFRHwnW1n
I0R8IZPX/bIo5nqBaXUcxl9TUEvNbBANPivKMNML+uyIEfFOOY0PBnTNHcIPDg9eRRr1jX5QIIkg
jHRrZ9JdZeseEVILhZbRSgYKnArzHaxyqDNyF4IpV9LKD5ek6DyC85X2qDyhUm10LVnLbRNFMcdq
7lcggIT11Oyjsjk/a2ao8v9orVWyCAAVJjVa9jWY298KJ3GeMXbanqbrlJXivq1GG3NyTJBjXjDg
APbXTN1o+TPz3cFRuu9fBUoW2w4tuN62xisU4bvPS5ICcpIEkWM/vQNi5hpxMyoO5wCzjCPcqSSH
k05asHO1rE0nhY6X5xY6UaaFcAbf4vTBpZdWqenUe3qO2LjRh1tAxkJZ+ij+hTMcAfrPeubKNgA9
tCtg31Es95vkGkh1LOc7Hbx0h2skI2pawcDi2VmsRvNyplAgZcKZI89rZMnLbjNdMUwYrtdH4Mvx
bdToaXxbY7ChxH7XQ+mizIe5nUxKcSle3uELszEuEmYux8PxQs+tGphuH/8+b1ZMyAlHAYRxjVlY
9Le+6WE5OWMtyIYi+/Es21tq67iqCfkyGEKIjignKjyPu1ogY8kQhukvyfMOJ6l1c2Im0l++7rpd
C9Gro8J/Ypq1Mg52Wb8HKF/zql3sNroulcnRDAEjhskdLTK1dXH74lomcpEliNJaJp40rwLnF1OB
oxaMLO/LkMLskcDDbC6BbIFaiTQ2WwlVw1PAnzyJH1OuOtK9UD70zAEjKDXPP3nliEtQmuxAc/N7
/1kA6E9LiMQnavrCo3hEUB7XIk6Q9h48VZf24j5aODv75DPqYnCrruxABvIdnXu8MbFIr4Ydlh7v
s7HwbT2tB7pKqfLrgOhZYNXQAajcQub1gFHumg7PeN9vSRNg+wIQ4Lggcg7wyzLsouVVPcUNeNk+
A+XAA/FGwukM4nWew6ZmUcrUHwG7CrjH6YX3lahNEIBdAmmSDtWe3kjvX72aBDckH6o+ygyO8iFh
dk0fkOtk13Lr5WCRaZzqzYcIoYMC6Cc5ur4jjXnFcXdkP9tHVMtcwe3LEEVYCQ/UxclpLBJ29SMJ
jtmlfBmpyQ+zo4h8+yf6XdOOL244QeICwy0+83wVUZvo9EHCc9XLaqMBL9GR2Tl+ql19OrClMyRp
khgoU1OSKknbtLJpjDGB1zVcsquGKA0P8ZPHKOPYn98IMulgXxxKGqY/kKfBr0UkFES+a00LjfYG
bfHgTioCaj14JCnZYnnAwobMARHF1G/kqP3O8nN4/A8ybkdQichGGnQQK4n6xXA2cYf+dxMWT+9V
g84USv082e2G7qwxHT+Mw1bL3//bddtJBKxWCzN3vFd61/Xo6UiccFW/BnC0Q/P87SrACUzjLQF2
iknZCMlwtwhHIYr0SzZ9TMaSlhX7hXrM66VFxp6wKhXTg4d0m1K+FWHnQfPLgMH0uuy9j0CTlPOq
Ze7RjTh/qVTbRRl2gjsmjmCgipaFFib2Q+LRYWxC9phBsdm24DbHuoqoIp32gXOYl7J9wmLx20ho
69kcneaUQ6sa2XSzhVaBFJtqg2AHz2LBMnRiuBp5PET/zZzD8027UyNESCJ0rm4QQAJ7nMaXkd9J
hVQ9EQ0wRf7Xz6UsKjQ/zbsh5CJPE6gOuKxKS6ZwS6ITgVCXF8gaqRoWSBQ8xjNZW5sE5VJmEOdj
NO13mLr6kTEjp1T45WcqiSWszfqbntQr5ENH6J/YIWstzAOxAD2Q8lU/lbjLqVbLLL0eRbTSej3X
HJNtNU6tq/FHe5wTtB+vFM8X6fdWvHhT+Qd2ErbFoRb9cEXdETznrWpQLGdi3ja2yj+2H65c0MZL
/F7Kk7eriD+8aD4dCD52/MqHxc0vYv+NGwa2lBUC7TwenRwrrdXBGdp3grINES91PWwiqVdNPwl2
0jwNW9c8A4H9CqG5GdLqczPqHksjY8ylEDpkWJ2KMwK+PXjeprOjSsJ6krLZX1PefFca+f0aSn/Q
MWyGmUC4Gz/CNksqZ9yyl9XcMdov5uUcx5HqvdzCxT9eJqLrFfMonw8PEWcE+xjRthj9vHo9A0XB
buhmMXR/IIjl/uw6w9a+YxI9AhFMR+dVSR5oYx5Jno4yIc6fgjOjrw0tuq0xYkMew6zSBTM/YAly
klmLwvJTPZz6pqd++YcmI08sRC+WkpRX0YexjCQh6J3Kwic6zgYqTy6WFhqrarGZZicBqKTaXM6T
uyRRsAxMyqEl/itA45X24HvFjcuq3Cj2NBI0dJDvhdAdCGR7vmAel0UtRIblYyCGdPjVFsjOeYwk
CdQLgdTL+RFngFjp7ONkDN8HMhdkoY/ye2F5zkHMJ9GB0ElBdlvW+kr6zC14EcjfEmaxV+jz/4xY
5I88CopUk7FdjfpBL26Jcz4G4+iu5glXxLvaqMATEjSB8YRfoPrNmyvRtuHdMhoO9ITkeZOWdPx2
Kjv/25HIuXHVAqYs3bpEmg0zR6ao1tMIVQ17+4kX8PuMPFwx92nwH9JWLd/t/iQHhyPPJJgTs/K/
b43ueFpr/QZoRLGWcMEGtRbCPFS+OgFK885odqxEmQkT9IcEz00VnL1OotR5rHDNTin9fXueLJLo
pCAZ0VcktMJOTEB2xcY1K+lX/LHFDwUM/B5yuu0gxge/62QiHSVm5hYifUy04T/ucMXpyW8UOziP
E+f1TTtDfYToGyIBrNHIcJhJBkpKW59RsFWSVv7iYcrUE/p2DLk/M/xRZphJ0mxbUYV0maIwdCh1
h3Hw2auxBNKGi6g7BenJBWuXlyX53JA4I3yj6zORsoWhuFDoDAd1qhBTNyATsWXjo5Pa9v4Xfmxw
Wdb0UgZb3KvrL6+VmZl0nJxpV162HmMA/G81cUeo2z8T7b2nN/LXFyByGfLkpyzTEXa/zF/idc7P
LOYiCUgKICyMrihDLS0tmFWV7/jcmgfJWAPpDsc7/pWXsHH0Ww3gV400Amv/QkR+Av6q0UAxHlcO
nN9BGwNLq/6yrQtzYsMXYzxhHnI5D/Ym0wzJuGfYNUOLGuyjwf4h+4hblXdjQHLCnXbHxE5gEByg
DcaCxtHUdU2GF5YE5PE4gAX8UeQQRrcbNKPtlz70N7g9XN6hFGkLNOkzJy+OLru2Gnmc5bPaATkR
OMzN4rJGPLJ/vshBS/QelT5ahqkvnuYT0R1/OT0B4Q3VVFWxL1b9ty0V90iL8zLf+Z5Gb+6P92xJ
GP+wai8ac5oJQpm7IfI0jsAMuIPAy9ai0qLWKMurbpoJFYVTUxfpSUXd7OvXsIstD63cIXS/ZeQD
oR06TpwgfEKClGbqOc396plMBJ0wWBr/qkzD+NoNNIuO/nHiynR+2nVZgkjBu7EijM9vgo5EnFfZ
KsJCBTmV/zW+rEQP1Y3Da7hPGu3SW0tukQwtXHzWvvYtCPX9yaJvFkePujl+VE70pHX7TAdKuTBQ
OvAB4gzm9SXDGiOSGgCAWZI0NTDiQuyC50S4QsDmJ4wy9+thpNMdbJokbgL/YnsLw77llFl6tFO9
c6A66X/+JXCcsAlH8DMTvk2XRjl2VN426SeBq3bL2s+EfrwVj1KCK9Oo/jHR9Mpgnf8uUILgr0Qx
TgNrsQOyWscmM6nVJ5eaGSM8FdWgk8z4IgCCYY/Tm4/YTAuKaGGYFntXQttp24sN1dZkL6IoelgI
EbaZHLArcCOkCumunckiZzI266VOQW7mdByNsbKPS1uetO5W60BQk4Xj5TAg8d/Az2zvY30i6gk2
YullqhURMwpLKmKnsaLb4oEpz05vJjusJ/mC5gGfMTvSVlJY8AhmmLWye4zmghH0mWrGlX7y/OSw
GnzULV+BxGip47riGkjNIvqYUKnHWZir6du5eCmhBd7d555zdyVk1KGK7iJorgjtaIKjQ2Vlzut3
GkWIHcU/iN2dOAjxOhYr1594VrjDe1IWL6eC6+nI367KiRmugkez8jua5gkFmWkoyzazOmFsGolS
akVmX9Y2KBpS+9gg2EMADI7Mj2qmuOxkfGUndCCctpMQ3qnDnfv/0mn+vbT9vdUBbhUYib3XpTt3
gzE2RPHHJKWurOG+eOGHkef9X6zjLUq9DFiF+yI8RBdr+Odj2CwGjlwHXSp8smkzjDgP4otW3Dni
yDx+Awx89zNNUKHHZ5pe6/4MqKnmblC8qZDRk5Aio0D/zX0nuHMTq4nd2f+lqR30//L8LvgQcqXg
Y0I/bDTk89QYO5aZXwMhxEBab8ECy5xkeaaBV65tw76LLrtf4OG64cbvycMsM2TGNg+f6jkb/ILQ
7zMZWz6u6fBDdsTaM9aGeA0cm7EVvnIkXrCYf4GqJRRHvb5Jh0hEZcOcAqtLL6vyqUHmFvF5dIoB
n64Jq+aNXylLkYd+m6Oiuvjg1Y3WkzIS2XUsN5/5zCXU/wFTBnYb8tdKdW9Mhpoc2t9+51a3I1w6
1N4d35/NySf9YZc/b1sXQJkC8E7PWHFd8MAH7TursTcnuBxXaFFVfLSqz6TrySpsZ5GS2jm7mP4J
cX3gWFZ94Ue8TdgDkv6UsbwebXt1ZOBAiAfF97S0HT25TmWIuGyexKbcIOzGR0nAeBN/E/+DP8x2
k97ITR+0w5bpEo6jwPzjIM9LJXQxtJFICoZudxy3OQy/BoslkuSC7ghBmbyHNGqILVjZ7/CJlFHy
7/OgZct2phucjlkdfMbhjw2cR5L34bFFqM35pCjOLoBSktOlBt+h4Tay8ML+xnY37BNBV8yFrTMi
3c+vLq/w940UkyKXepI06cqNOP63xkzc/hhiggxW67+74DCbwnqdgcyDj6VeOlx+6ws03d7xvkED
V9HJG1X6bbPY/DVPBd30pAyM0yrpSLxPdxR4EdUR1waQqwcG6mH3pa/ILdflukh0UG5VX+BH+IZr
+2Xmvv3MhVm6c1qRaDNQ1zw34AWXKejE2Vz2ieZ3pyoTCa5VHDg58TGMIL1D+jHGUag4Vm1X9C4w
Htoak2TQwN0vo42ER502y+AvFBX81+5bW+0Ar514H3YQpcI9RUgGJUxteypuBmoD68+xubah32+m
bt3YF9leGGLtG7njKziIVbSCshI9THfOlzgawhZWPO6JTc2VP0bn4DYUfwkKgyuEJkL3O3tpsDGW
p1zukuHB885F7PARJihJoQC7KNaWAjZmmtza52rG/WCKjNLuVa9L9J4IKeTTEuz8r6KTu47uegBN
cRg7Y/9+2AmHKl9578dGxaTcnZPaC5llN8Fto6umPwVhlXliwSsqdUbtyU00x1FpKoFBL7sgE+6w
mQuBCHxkYSx/BZ5Ji+SUF85gBWYEfap5jOXnCRcGIWwAp0VER1HYA6UDzdTuYaVUK2D47Z3VMiWO
WsA+ROmUpr+9fS/qE0nLf1+pgc7ImO0EpASMiQElSVNToolQBkJHUa15np2VV1UQXBMnRN/TGzq4
rGy3hYyJm49cYhMTx6SltfsVPgrQDQKDK4Tw6A1X/2Z0vcegS2Q8W7hUFPw+EsvFGOo09eqEf3yw
Df1tTEjdI0g1/8it7nyQ1sXJYjaMsSW/avCGA+MmEWrXiuZWNvPMAnGHkuF26CE3rUJt6V6ZEzNB
KakTI+R0BKA3BcLw5inNlEZOegkDOjmqqwmUbe43esJ6Orf0wNbuO2Ma6nR0WEw/PiZfjZE/9tae
PeFdRUh96FrQlMMXei9sDNZA0VdaaFMlQqeB6PFZfWZzZZafxvjKE6nGT6X9Gunq2Ma7zS+pGB6x
dyhJczcgZS24AU+IW4qmEOvp8gGUlvtk0OGq7FFL3Tb2wqB6AF8SR9x3BOXAVRTHZwJotzqo1EDa
QN3IN8nTAgWfjdbzmb+dK8HCuKsxJyxHWgiyQaExlOESQNTC7vNeiGCPJuiPvswGj1CPnT6jd69+
ktX6AZmipZOefLMVWCeQdLIKDV38/VdxgLl8zZaclmWR9SOt0Wm41caF9aZc2hDpat0h5mGzMVbR
EWiWHw2xJbV6k+7axoZBCaOKieTUfVPUzcHKQ9+IWpW5ktWKaktYGy6AMURz3i8J4Q3qn8I6mhAk
u+hXf5g4uOjp8wBlZ6HesJcDPdf6NavjWNbsF2bewtXFBIqTrSH2ZfAKTKLrqVHPfCvgcSBbeN8/
dhpEwR8Lu4MU915D6KmDVy52lkO6TLso84/FOP+Yo5l7373vqUjliIILpSPJ7pAxWVtKmdOy7EuZ
9IK5G4cJbA7xPMrH5QX8DOSj5Z5nCDeiyDU7vRcXdjsjeb9GwJRuCQxLG1W6N/3vxHiO622tO9p1
oqnZiEZwKBgR6VuBlMx37yyB1IG7PBUQZ0D9sApqP43dAsXPB2Aj88N64mV9UZhRUQKC3zxiECZd
ec2LoAmDEXT91gkXxTGfDQb0anIhU7Zj1OWnWx0at2G3t7ryiYgoWY63FOe37kd48dPVScd/ZCHa
454T/y3atVlxyJiWNqAHAmrlvuxrxW+Ov0tKOdhYzo5PNOSHCh0huVSqE/9waje/aVzSUXN3j39+
LVx1yiSssKLSLibDyMynNT6DPCxCI/0kiqbTEZGBH6pssjQJnSSNVFDUKgLiB/HV0arEE455lkKv
KxjNAlLJpwlUHU+Hm48oGKKO9CokQ0pbCwP38wEs4Hx+UWeQeL4R7KCnUSG5SfpVMIJO+kGsOTX7
FB2pipJTIG9AGZrZV8va9U5bmxOtDs9y5ZkqVMsR3HEi3Osj/IezI0lCZ4dD6VpIbn1T2Dys8Gjf
IqY+hdGGYDAsZRCOR8vHj9/Cuz/4MmtRl3+/rwpmjgLGix/6T013i+cuD0vnHCpNFJLsbmeNQWEN
HsESNBppJU5FpHv0EBFV1MoaHDorig0SK+ZGvFbIdZAUcpp1nvBYNQZqewHu7ag2g2pUD076GlyA
UKXvtU/kiPTjJRR6WqJVt1mzQPl80suJwnfLOo8gDAFMvIItpuCWoqddSqyHho4OpRMbL+XT3F0D
CezURiyhgt6Ht+aywOMGh/cx7gviHgsFPnIQaeTs5JwbOxGw7wsbRYnAmX1Tc57JIrgnTqE3knaJ
LfqtAvzlhUFgOvBz57dokKr6ipjjq9BZogX7QW97QA+NhUEd3wGLn+sUhIsKSmZ72eGQWcw51kJT
dvqWqSASeeGlPTgucry++DFFDNkff/vDKLKiURkP0fvqh2RgYyBp97X3HG01EDudl2nr+WwHF3/0
DERodeVWfGFuJ9Q2UdQ6PNYeV70jCzlxoXlPXTlvEqMJ3rQ2k/rNYN3bAuDNNprV0NQsgRHpE7sm
mnJ1XmjGoBJpmuwVLoG0QGm7TkcP+L3KZXtdFl1fk9WYOwbZyZTyt1lN2WS8BTfzJ2wJFzr2J87w
e4DodAMOyol5cXX3p+TqFj7qWRoAi59Xq1Z916tJvMRXqJesve9EMjjVDwfcoIE/8bqNtifz5o+V
Wo+5u6zoLP55bgPWAN6Dt72+RRWtMFnzjEagUChJvFWkVgFmMdTqB3af3155FNj43GZy+MZ8UJ4J
srVGcYiVWCENLCy0yetJBGIVJpewCfJs2zgxtUH5styHGdtBp/BopYRZ9lPT9eEn2ciht8NRAKeY
mmwe+tWVVZ77ZinbgJVN8wseHnkjs0Xel+DnifpIRr5t8Ij8SCS9QI4DB7i0aBSrMb+wCJRHy/i6
6bjMsKHg9mCY47bfSKsJrMHEZ1aShGgDEYwOcII2DUGmQ8Josn3Tb0dGUyDO3wjD1m5HoZ9JRrNJ
lcOtzGcDGPI8+v2OTA6qrnDe/kyqJGloDYWrW7DJlTg9ObilzHAz2eH0gdtaFftaQsoGtqjMBmR+
Nog6ZBXuywxkC8qzRrzV7bq+BNTGWKLzE5GiX8+UKz8touuyTwHDQ/A8y+PfdrPIttneyB8Rgitp
H53RFt9ZYYUq0K1v6qmrfVBeSKxoIqGC0khvKzgxtoTKs+9QLfIfoyPbVTy8+rKifMjvIw2Yot8R
59krx/iNEdFSnmRELMm4a58ki9Qxjasu0wZA963aAOfMx9yhSOP/OyzTvkB8nyxpYp9whvSbBgpH
RXDMmtbOlLBDpSUon2CvHHS9r8781CHxpxzV+AySCwYKv5EiHMM37CPCZAmI66wWb10yKxFEB+yM
u6gN2MFxQ4KgfSvlvoqeEU+07yd47jCj+4dHOFYn0V6CSdvZ2SAPb3YkA8Nxjtze/QJGx5pXvW7o
gsImxNklBGQeBPaCMWLWr9kBabAMz/YhjApuKk4m7iYhPCYXWfjFhd+HgSmO8CN5Y1YpiHQnJmT/
iCLa4BxSvsnroys+1Ay9y0CoV8kHUWwnUHFpr6WCEe4gKnzNoYM27FZfjw66qz4mQF2r5E/dsX5h
Twi9x4HbzP3DxY3rEfvMNIDKEuXKZU6C/ZTG6jmrZJiteAmqYPWBBPGzHdzQ6SQ2j4BEc8h2FDwL
r4VTawkvDKSU2Ua0vXVtfqa+yHxv+50OCt2Tgn2CQsZWae4dYzTUeT7F9h425f3oYH96RmwwenLk
0xmA1AKjOpoltiAdAtxEIBEFCPEbmnsPxd+LRiuevkHfKdeyIVePhcNvjoQZv76Bcxr6tFMj7yL+
jWH4h/9aLgV0Vba/5q0u+zbhUAOSeEPfMQzt9uzefZ7oeEj7omo1+36N0UpZfs6/DU4cAWfMKVz7
8Ead3VhXOGzD2bhmE2uY0H1H2sR06iK4HYWXxT6iiQRQlOdPq+abhVSBlPqgF6u25Hlt+ybbk3s0
jXn/OisgZ3lfYZ2n15exUzdc4RfyUcLjirwo/1pnEEtept25gI2V3w+SRrLhY3i0a9iF9OT/2xK+
nr3Fv52mEhEDCgvHxf25BZ3VsgV2+gLXspLySjA4xRCCiiWj8X+Bj1m7N/KvYM92WkOEknB6NiDJ
ezx8uKdvpgX9THqkcUj2cL7YMwK2rITPObNLwI4Qe9u9b0w/R5fPaXFbHzqtQwEOhQ/5E3Aj5n08
90c2fkdw3k3FuwO1zWPq2MPxYmns5QqiN3Uez9EaMNDJNFi3hnZMb26Sq/UI3lTxZUfBDz5TEIk9
oth84wgpeJAj8WsK2h0eeE+LDYhGJcuKHoyIyPVAu47iZQrZIMaBOCy7p9r+yQZq0iMm/pm0jzYE
yFcZgzeWpPg6KMrAy19BlCIcATwXQQmyCWpl3bivjl3ts+wIY610hU7im1yJXT1Ex6vq3JqHMuuc
VkAaPa7BN6M8UD2SIKV0ieFrPvnq4Ukzfc2u7vD2JNql5b6Wm90WOgclq0bJ6bzOiwozvPtgHQe5
C0o3K8NAPj6vKoq6s7z6qP1F71x+rWxOseRgj/Jye+sMKfzju+jZ8j2mYh9KSy7anuh8ot2HRRuY
aJruTSKprJpNklmMsekVoUyMhmf9TF+gk5oM4NfUc69IVghJbDTkgLCgumtKNjarjz4TgwOzD/uD
yqh1xtied2LHFEjo4lZZf2V7pDgwE9sVD+4g5+SFYJiVfaeC42j7DWRdO6A8Z/1qzM6nANpl6nhh
8pdEYfHorvQsckgVzip/RW9+lDYu44lw8uP7yMTcganxq2Cb8/+sG8TQNBLN/Pc8xtZoKHFc4w1V
GlHbPjr3Qd38UqYcBnhG13LL2RbPoMyGaBthzf2wVLXSH1NnvZlLGVWAjj8pGhIY5tlXhMEby1vi
VhwLJ/Z2n1NNUimqikVILTOgnAv4qB5k/+FeT6PSX5SDEiIMUUhTaJwF2IUuLAuU7My+RhEAkzTh
CQeMvL0HXEGqnggEs6K9NVCCLLWHtVIxt7yj2r4aVN/dlkiP2ZHbAqsPvEXJyJY0IA8Wbw52JBGX
XKaelfEF4P16rhCZ2hJ4jsG6Kf2Xoeq+dLA3QsX4GCisaB9XYMwlcH8rGBsvw4MyIkmazxYF9nqa
trApTAfsL/a6VC7d4ZidU7yTPQnMM2cTF1kQo69/Lrm936NVgazkjqIEGmELw90aQUD8Wf07xRxf
6Th1C/tKTcNrc3+SC0RQhsQqIfehnyoppZXV8r9dHJICVWLg61dhMHkKaXQPJk7a+u5wv//fCkqT
cTMdB5XpkyiKUjqrNskmlrPyqN5q9riLK9PI9RSxRro0PZCn1G/8wWXHcbxS4tQKNFvSxbOmo50U
m0DYS3KQJSxMbfk4zO54P2Sj4y8xEuzk9iaR7Rk6v0pq14hbe0WcpcySsh8xqTIcdK/GpBFWHKQJ
s1Y2WVXvIUwiWDF8OOIwccERa3bFYFyI3tNhdUjTxwyIoHzdHNAcoCL57RSNK+N7prpmpZapdP7b
mQaMhliBpYbQ0oa0j35NPVld6pWDbCoKJE0BT2Pi23yiaEHbiZQNA2jFduYxw2k32ivbMJpPXYPw
bcsNdTyeyafIjrqdyhPhXOe2lpkC3JxfnWnTPOpf37L+MCx7rQS8HoPT94dRr86wvSnrs/OssFGr
iypuVrQAei8vTKyPYvJjZuuZN9bmglUKs1IwztD3va25gMj8jvCddDGAsbS3JLt1k1J4kb7Xs1nh
2pcqJHSLjlLS/m7N9ouiQB6Cn/euJy5iEKmiEpnaXw9q99JftapyzSUVtxqsZay4scFWuiUw3jd3
LSK93qj0UMyXsGyfs9YwMmnlvkbiOEoA8lB+q8ADHrCiTDxOuiGFlJvIfOuDEpSj2JJWpfincaiz
BAKekSoaqdwHqYBPTB6+yNGbK/WVreYyQ1VxKHsyjm95gF1PRZsbdb6SpSAGYAwFpVZ6UhI0OjXc
i1/1HPz+i34BiZV068V/3I8nF18CfVHpbA4g+sYPX5/2cqNyVmg7mkWO1NcvLzum2ti7PzTOjGJT
WcUABpN26ZxzdgkHPN3ztxiaNQ3F4KPWcOU7mmDKK98B0xLytuUflWbfBX5ciMWlctrcdoCmBHN0
pxdTBXwGqQcn4IPw18LoADTEq1BYDHSLSw3twdVY34v7/q1miY0TamE769F/9C9GKgzF+aUUGlM6
zptj6Hhl0PpFFnIMcEEb9EnA4Glmhg1/m5xOJOJVxM+kfodQObyJGgTH6yUX7RhhkKc6jKtbBBKx
j2ATPjgW6fDssXBU1973mGpHEjHaza23YaYt0YkorVKnitMBMcSx4928LmMryTJ/opNIBSM7tUdy
RWPObrf5uBDuF6l/ybz3ElbQNjvmfkgrywwUlCr1Hhlp8ZUbMpVB1DfMov3DO8E8Q4SivGTnf1Du
zKWkakBeUaHANARM48F6vJGdJcmWIl4pAmQDmi4AbMh7jwkBN+9B+b6jlSF1x1/OSs0uBYq5IG1r
c+FpG1p1WLjwO3y1Xq2guIQOb4mia7zIL6ZiyiOT20zBMkQ8bVVfSNu/GZPGy7Are4RET2xJKZbM
Vyl/CcHFqwqDtCPlc6g1cYLKTd6jBi3vJ2krCD1vdjiox8sIUEWjrqXFg685+bzWKBeDuOb1A7/e
oE4LBpvh0OBkPWo+xqHdsZukSHXdZoUjpnkoomp113bDy0H/swDOaJRn67RDmLu/cZhblgG28pBG
GjNjMSjiwst8Hos6y0hJX/U91078zVUWsXqkqOWW5FsywPXFWnBL/ChfDee0Ci6kaX9jTLzCJdJm
qR483Z6e/GYxehQM+RVZtKWqx+OJ+hke8sxNhuKjz3GHypDvl1rFVF4tBssiLgZC47A1hRcua9Wg
MRwcrf8fblnP2qEGzzXzkeWkE/e/oSfwLTYpHuSSTvJ5ObL7of21bMG7VwdNz60VkIQRoG9eNa6X
k/Y6tmd46/waJ9Y3y35vAqwEcutrGJvbQCv+g+3WhB9YhwKQ8E287Uj45Ou9li5Yrpvh4Kqn1hgG
+xYq2A4jIolDRU5CFPz8gNb0zC3uEI1VlJWM7RToCvlK+egOEMKiKew50/OHw0GvveepqaT794iq
a4tjcg9BCCX9FQtic6Yrdobkl6FiY/pIAPEe3NIUWurlub6tFXGcrVf85eAF0Cwpokrx9S4OmM9E
vgM4SPC8L6GWwWNx2eXqM1SRjSF++DPLREW4+fZX+Vva55ViThhqWWS8tuVS7JxOLG1c7tObeEzj
11xYLTZBwl5w0fcy1da1LibQRvmT2eBlZIFIQHR/61spfpjF6+7MfHEggcAXLOsKPGk135XbRk6e
IwWnKeJqotULHnpApd8wIhUV9hL0iGrKLePqzJOuiAo1ArmrmbiT+1zW7LCazB7wGKw1FnTpE+t9
qjbD/O31RhUaU/f4YsxvnjKSGH5XmUMoV9N350GwpLTC4nyc4ZiR9z7qLfiDF1MNlHDbA5R7emAW
2OTwsI7upaXWZit+6R6XRKrkoRsqYCAmSWRFYZ7ddtml4APDEJZyIDa55PoDAWO0V7KlO0551Zqm
UodZ8/EgjsddT4Xu9mpJPpvyHklfwMXpPGpj8iuBn9uwVH8NzEunxou4bHSnA2reiQxMD2laAHLE
zAnm4A30F93OUKeY6kwIeRKX7gacZprtz9UArx9ZGfmpI4Aiu/E66ijm4Jt1SPjFO2oqfcNVj64x
xgYR2EWrnnPSAA3dLIT/VipWxx3uYUjRDAxu+w37TQsLlZ9l7NwAoDEFd561N9INznBCuDeFY79r
grTeT8kbeYpPAHO6ETXaV84By4he8XnZe3RT3Ujfr/rcsKQf3Hm7UTFQWgt4ADPtLkCdwasM4pVh
TkX7UhfAinr0CdlSPhquZ0t1dt5ndo2RYtGikXkIravXjvoUNvRYaAB3FR6GlXIIaDoy9LalnC5T
NzqmOCyz8nElrv8hk0pso/Wp3lTJSt2Cvx0WLRvv4YwgaUu6ty9gCcHUXXQIIHsiNRkQ9lFiJVTi
h0I9pDp4mQRX2oCzz7WZOg1pJTksMsdSN2gGu/M3BY8IoKoCkx3MzWBHlFFpj2AYWAQwuMajYQ5J
GA7gGetx72Em9JbSLRHiMes/IYwQbV8uKe3lniCQQ8zZQGwdFELo8GcHe3FtxhrwonCbYtDwcets
Q8rtCPz9YJI8kIRz4YGYZuOQW24oxYAoLmNTrqN+gd/MgdFDo8RD6cqCmx6+AGpa1gQYT07O59Qn
MELYOVPOvhwOeRU/aQvALsXaW82Lc7JkshL7ssDD0l60Ql3HIlsFMHsaLh19szBRU4a1EuwSrFqs
xupvChP6ta3HQHsYbVxM6BVF87SfmZseGkynkT8SOWjt8Jx2UoE5lgNBJqiowMP1PUSwqS4INalS
E1y1Tk89yHTtLpsLLghZk6uHIvCM0zYCGvftF7FdlsXhvSV6O+zKWZtj1OF5iraXoT4/i5fzTIx5
5dpUrizcC2Qm33aR4odR/2+tQ3S45TyTgnU9CazLx2dH0ha9fxmkjBX910HZbKtJv1BziimIM5Zb
1UOg5ukmWA9wLf/HmWahY0vF+pLA8FnSv1CsDrF0JWinA+hcXIFBFgIYbggQvEtr/GKHmUu5M2yf
DAoOWvU7Ao5oesvLvFsTIf4SNDHxdX93/Jobw6Rzuzmm2cht8yY4mFKnab94JBRRbssr4ujd5uIK
OjM5AtLyy9gkzAOunDgbngnUDB5CPdIxoQddsqLIqPsWXq43HRTPvRLvVeOp8cq+9QhXVVhV+otJ
WEAFHuO3owfEnsHO41h+GHZjXch3txZysbj21BPX6RfHyY1B4A/yMsWIvG+ewl4v8cmi9rBGOXFr
Jce2igmrW+HsX+GjEyOZFM8qyYJBUmdflfhSWojkX6WMN0nc5wzA1issu/UlzsGOWzHparwppSDu
kXM1YQz5uw2ky0eJpprTHqsQAPq1hKAFeROZbX/tpNTLi82Swq4Jcrug2RFc8ahs8k7tYXcksCEZ
WVd7YuHoMSiXpQb2b8Djc1TiC88KYPjqrhVPo6ob8PbwdHUASstRvLISmmPMe22scQhp6i8Jjsoi
taOgop8npJEC7BmCQjgTr54OLN4iHUWeSnvh0Fi+aFj5DlXs7TOpBr+bk9TdswptKdzCsL6+Sacw
093amwcVLDf6GE3R7SMxwPOn+D5bdx5MhYCw7po+UD1G+3XhrqrCockPgAnQcumd9ajvUTkRRiHM
3xvDcUHRlGxAvlSM8IqBnCbE49s4luuwBXVykMtNleWtFRlXZqbF/qpccpCQA92QUPTbDTS1v0zo
KQ880c+CtQW/ErBO/ST4Ge+iRsO5D4kUMwRx4yTs1hz3HR6OPYu1N6zHufEOs9RJ//PnKrj0fG/7
RrbrCPZFxAKEGsQ5O2X4KPyeDqGw080uEZ+YXhdeVSrGetAubm2XcJG9WTYzFhPwA84H1IsKjNej
+VhArVBlw4GfzqhibnE3C5NOVVOuPSBbeTtys8rO/3GZPCi/a5yYnqe9Z+VuScp2L8+c/G0dTfMZ
YXIoR/yJsqd8ei1qYnnsYxf3C7StilOi5t2XyyfrGDl0cTrDKYAbQJG1Cvk3uELAk3LMBdnjo2Oe
7/EQPiym1mppKiMF3rhm5xNDjsOiD5yu2zDz1urdnCuJkVgeEH6O+qTG3l7MeotFfjWFPZOmjMf+
KAtHQPvi6a2x32mp5S+P5M95UljQANqVh+BO0g/BV98pqxBatE/JuWlJWWI9KLkftKeUtS00nptk
oe8oVHTQKKrAvrQ/9A3Dy7ghPKykrcizRj87cjudS0EwIGl0dcputXF2fji9vO6nzVKV93BO+2vy
MRPTXop3pUvvKIq1Y2TLd/dZBWYR5ATD6RKLZ8A8iQBtnFsBsTKanMkydnAu0Uzly4gaQeD8NPtQ
iMJOVL/44H86408tcEenpYejB1ZFrYtel3FP+dsphfDWCz9zUGvqPBBZW6vMrBGjWJpa1g9RQ4p9
SRmb6IO/na2s+pjOaXRatcYkMgITXl48z8II0olvmV/ox7x/EuR7AaWY3TX4EZAJCmlCSE2zD1tw
5HDscyFfiXw9Si9D2f8Rgj5uz+aKpQKxIm70jZu5DRfbxxLc/MVyIb8bJjLVMI07thDZIfcqUCZq
wPAcSdsAkvs7iu9ffhfs5fLI18aTHkFADy/4p/6sDOX4i9d2E5e2JwuXgQtQJY2HxZhvVmpgMZP7
rLrvBBwD7Kg5KOXDSd/5YuZ6SXR7PYA6bf+lJXPqwgxK/JvNs9rnFthjgoJpwk747XFZXYRpriHG
4rITfO2op9i7TsFWPklB76mhFy6JUP+Mqf2/i39QQPNCUQC5iCI2Bx3X7BNUk5/KGfUf3Xgk/SIZ
L7kCKBiWXt3zBqunnOPgnj8IjAVRmYnj6OhCK134W5JXbp9rgNpu8t2TxPDC4nNN8IPtE0GgW+Sn
3/D0jSsdIN7BB060vs+ehNEhPpYxiEvZnWoZwCX+V9BrIrk3Ia/rElN5GgFiDnBMMeTug5KeiY83
uR9IcuG9UbpWss6KfBjhuK4BQAaPOfsN35LXiWJXP4NtPPbiqbHrP6qJPjFWz8jhTVl45IemNfjB
AOje0t6rM+RyckaIuGk6MnWEEqQnwDXudPpnp8ItGxy8d3IwnmXkGgQ/cW3zYC+6mjssm+iOwPpf
cLyV/PEENSXQ99WTIHA/+oJwh1DoPBCktwuQ/ve0XaYDCrornVbfvAbd5U18PiqS0Gg0gOLK3Xbz
Bukzw7ogOuICNu6YvWqqwmN0SPLjEBrWbLSamn9y2ehZDW0xbc2x1CzXtMTOruazDbRwqTT+G/XC
AhiOLFsTXjKLJeBqif/i4U09ySU9vCT9PVRqrqJhyt0o/aigFkYHzs0RNfof2TP4wTHFHs3ez7oP
UPK+7iQSMY47LpMBnos6tO+xW/TUlsok/zU2REy2Sc0eQ05QANGVou5toutUTcnoDujxjHS/6hUv
10WGOyxCEt4bVfmRM301ysdK0XpGucWejQZLAPd0pKgoFfOlVbRvsh1m9d1sHRMf28Mxfv5wPT+Z
+aa2OUk3OOqIfGdEeGZqkXhByLG18cInARXKWJEMraazEmaCm+1fOqMS4MWrPJmEzfPogaYbyIFi
NjUQqR3Fyh11vzJ8to+udFJZbrfFUTmAuL6GdkMAd+Vw4J/iucqh3kXNgQbdQhQOBEOe4KLbbpzl
aA9vyUpsS2EEQfJDYtnOJA1C8Xjz9y9pT+38mEo+EKLTH7Nw72ScQ89FQlsY1Lj+dtj1Brsvyroh
F29Wbj9HHl5qGbKIoWkE70m7IgKme13eVr59MDtQMOii9f1J2sAArVs2pZV6il3jEla19c2Njysn
h0gia0wOs9J9PsHCAcWEdKY6PHyt9BSQPtc+ml845X7Oy4hOvWPnI6uVBuQlwi8B0bLbDB9QPar7
bHz63l7ZplonnsnXd57+Z+pKH3HPmrlmhASapZrYjTKFuRuoX4B7SG73R6wC0RDEqKszkwHIfB3S
b7iu9L4CFf5K2IsNJGJqDes4kZ0yRqicESU6IYUz731uwXeJxKm2KdURNv6SzmVLpB0iuUPovqgi
bk6NVgqiFnFe5k75kNJG+EhxzB5FKDaj6DC9D2l45YNQWRT+DqMDcMBW2ZCCnKz75SOSg8OCj1AZ
Lazh49OU7qEE7pRR8oxOHtNDbxGCx9uYppw4YA1hznkOrf61/a95thegnibax2MZUqk5ZpRg21hR
K+FjzR5Fz1HSJAAVnUHm2vsuXhCoAm5A9LQ9P6QrGq49qwLObdQWQXSPzAsOQs23zyK+8jSPZOtb
CVWjPQCymfkkTLrF0vSJ037bi83SixO+mz8hn3vqRV4ZM65ieslJe/gGD+vu3qF+snX3hHEPmjlv
jWbHv6Drskss2oaeoVuJS87KVeLDkcZ4FOhtWwp0KsUY+rlp0zLq75AU2FmAoFCuGkqtlLeKgpFa
uXAX5Ll8AwNtw8HP8K/Yv2CtRehwsqwH8eM7z6k3lns07kbXs1OHHzAR12rFp+2Qh2+j0LBQm85X
CQ4k7nKySKrhB2XLtTtvfa3jl9bZO8zKTk/lslPkQ+qDv1MGCMgK8ufQ7gbUWZbMqKmUL1T0olDU
fUVjcX9eG0674rRsfWOi7RMqb94k+zA503s8lXY4FrwB5cju6wiF9z+8j0ovj5bAny0j12iua6E5
KG1Jnqi31fK3GDPu7sNJbur8GDk8r8kLEP1XhXH886t1hyq9KDxUDSSREg3W8QUjHdx9FPIKd0Z1
MIWq8M/H4qGvJNjfDzjqj2Eo4u6XcqdMaWpbsf04iuAEQRxJD65ZEUH3+62iCqgWJP35lv9J00UA
P3Rt0Y5RWF6vbVi+ge+AATPjllL+C3qrm82/+qs1l5nD4DKoYKYnfVuobJzhIICX1akOxqh45nNU
Odg12cei8nRy7h5sHU591WNvADXm9KxMNt4DFiZq/gmBw+2pnZfF/oGTmgVewDSfTYvJwfPdYC2u
uRWT6GIZaIJJY5ywPB3LSnHTJ5smKXbDT/vGfpXW1olLPT3Blw0z0n9hnP5qz9Scxf+6/ktcR+Hq
Pw89oKNOCmakXw2zaaLImDMVpiMMTR6+mzctbQKTl29ImQXPfeDAx2iSmk5MhfljIIxoc/Z0RoCw
t6lFAaCSETQzj9UExnLYt05TzpOq0BiTcoM3G15w+UWqivwkFn2iZvxjQZPux6KrjMz8jFanJFFi
y33PtxvSPnSE4+rfHOFeMkKmnH4bRMZjVWqJoiiRy+cTnL0ATx2HmrjXbdibyeiY+6Ybtvtd38IY
8H+qQmxxClvPvObgKIXLZnjzY6Uyz5jfavb7SF/ZBXFvB+NnDHM9SaCJQUObBcva9QHN8ExGt4zL
hz6D8tXNCCrwzrf+jGQdLV7CWa48EeoO11k+jhC/5NR2DpdnVg9X9zl1eOU3sqpkoT86n3+k9l9d
Ggnq9uJnI95Xti3wE8eQfuO/ETX0P9MpcNcE1aQkSzvoB2kzUaCnPE92MoFz8F62VKr9E5FGoHGW
5Ip6R1yRoN86jK8Qm8s38iyRRwDCNmuOxBPGOHMxuFICXyuzbDIM7nN+ofmSz1/+S7iapnwDAEU2
M0RXZsu5BVw/8bk6Oqfed6sqUAtCLOHP5BZeojI614PO/JCuMhdZqpD3H8vAC6PwE4WMGj5M182t
ex+0NhAPFFs1YNOg8r92rxaix10zk96+0lIQuULCp4ybbrJfv92xjPRlZL8QF/K0WXMLBDc0/ymN
iFl+fAy5NW1lfqb0BIqST9Y9f/cV/nqyqSCseWOsXVAFv8K5viIZaOlgmb0fLyk5kvVpNDE1cj64
EELr6k2uPLycjYHunB8eilOP+Da5FuFvOKOZcX7uYp7LY140VeKYj2q9mJvBfebyTtmUmSFbT9wc
uqKJb0IA3LVKk2reUb5j7gLaF/2kvkdfNl6RwHi01VjKQLViDWWkhAMXvqLlfXr+B5Ig4eiHuZyZ
b5W3dQ8BxIPQY/yy7wV3tpfgEUYpwlD1WNpf5j835sa4cSaLxzJZyS2iWSDLJqDJbCP/7lRbZP9B
Mb6PofFeNOA9SMXAWdOOdC2rq+ERuvcXLjoCduOpGoJSSjmpunbcosk8ydPHOOapUnEwnirLXA6r
zpbcBU6e8AQqi0hDnhVxTzgltAmFI6IO3k27+mNwxokTkT49bn+2jAo7SdL5pXxhn7t3o9oBj3cT
6S1945ctrLqJGjV/JlICEf/Pkh2BE2dvcjoxvmMAW1n8U8WbzUy6iset0MMU6Ezv8x7/uSxgF1yt
mS+j/AwaoBUVUMiuZTRHOn5yyKxBZxnkh7DXuKCT1qcqOWfVbZ7bE9H6wqxP3SmYK3dQUxCH3nI2
bJGgqN4vM8W5Rz0BK19OD0+v13JmJ74D9zrHNmUEJcIF1VIFj3YUI/uMwOVbO3haae7Tr7DjUyQU
w8SxLNyOCe23atG0gGSP7yX9BkLoF7cCdCNIjvOLOoinAiwewpTqkyxgL1GnIWhDt9Cs/B8KNfSS
RgTZlO4UKxzVGnBg71INw1mCWSo7BJZXYLePHXYqs2GX6EIOg+fVQyECKhq34z3E0z/CAtNyggvL
8dWJXB7mPHhFkpT3V/+Sz1i4FQrqwJjdzwZH5zUNksTi0+bIObOz5h/i9U/DTH3F+oXRDYmJkNcc
cuRMfyYAy3fbOjrHR2RgZXvDZrLF70LBmzIPmElr8mut4nkHw+SVvbR0D6YWSNA7iC/NeXhja5Pc
8ugN4mjWpVqISCYJex2YaoCrXKtcqezzSewc8WK/hmvAO7DQlA35R8sZtoKtVn81FGzySnMrlciO
TK8ICBcGYGX+LkmTbQEtEKdbpc8GeydwdT2pwR1FeTdHQtG0i5KdNsUDY/vUrMGudAObRK3tR22Z
/0prF7diJe8BS5chWE2JZTLHvuhnAvqCz57xSj4Qh/ueeKsghuO0yM+ectU3NuEuyL/MJ+NtjNlq
osgQN+T5v2D+4clWI6EQ7wOmm3VbatEHZ1dwaPfpeyx8WWh/q7PJ5DUn7aEQjajjCC1y9mj0hNsn
Bhm0PtbYW6rrKX7bdTHO63vTZ+qv8hnQF8KPyrflMmHKRCA5/c+xI+lA7ylwz0NBhvX1WWvkVr61
3mirYhZE8mg66NkAge8DnKv2v/QsIive9CRx3yfQ/twqrAL3EDQBGcliYk3keEUvx3EA5jZoJPib
jtwkxWF8uwuLPEYh/+5cCCot+alLNqlFuntVm4uXrTNNncZsXyJYgFPYVhI6HwHl0hFOIF8lq9RY
i8sSv81kiWTpPYRDHw6cTmZCch8RqUBq/QxfVAAwGpeFrlhT1gq0nKNmF/Kzz49I3IJ+VNq9qd6p
77m/Lp4d9BV6MDqO+ReOHakiYsB+Dn46TvQfA37THXwdzk1xz4Bos4xdZw46/p+1cybcuGQmG7XT
SLc0N2MoHvTG7BEWVKPf2ZEd59we+j0m/OD7oiNg+mmXVem/lV5MFLvnZe4GBEKEm7Ee6zFMKLBQ
D507YbTU2JFgwzdYh565hXnUaBENmfw9KLYWIfsyFou0DKnxc/o3YdWYYO70ZPs2MnceK7o0CSE1
uz5245fehAYK7p5JXqXrvb5Ei1QpHlRhlxFmvq34ZU0bigMvJl4tkvDFnFuEIsxEOHejx7F/AcA6
NEwZBsPYtij9Nz3LgCzivR1C/imlhRfH3b80hMoBoPIrxYlPyduoDic4LTrV8r0wzMgQ4W9XI52s
QcPSK64OaYAqWuofv6bgEQ7rbZp24eWZyDrqVCWriMJf4qS0+oJ16mjrLE3o3GwoEWaW86bPGcnb
xDlc6eQ48lHrB/MKzKmw9WZZUrh0v0E0vMKjpIi8VLUByTYWF7HzVowRRsQXDeBlNMnzaLTXv4N/
n3a9E8Gji1kHjsZj3mZ55FyXbXLouvqU9idp+OkefDyv/V9oZPsTzzDb8GB5qQYmaJJ2SFwvMZYD
NhtDbT7vyrKjLGZTuKA4SnQlBY8ZL8wo66KRE3kU5zwS6MMJ+F4vvg2h7NyMTN5tGdaToCPiunWJ
sKFIwEIAEtStb8o9e/mcTTLSJAPoB9CxtaNW6mKQy2UwKbAtAJ5iRRwJPWuNOpADs53y9TB9Lebo
LsIVkUpdfr8SA+U5qzukAh94uojicvmPr6pBN4w66Ikth9rOpLVFYLRG01+TUE8akArx4axgG9dM
+Zb/jf/MCpukjg0yz1c2yyBjS2kifquTdhhEt4gz3rvwbJC9QuH+GnP6c1fbfoLZVclzsZ0ypAFX
BrOJKxSJ2k99dwz2Zwi2XVg7vhpxLACMsCeFMn5qCftBd/5tA5ZwBeUW7cNfj0m7poPY/l3A6YMG
1shvkls29r0W0uyaDm23ZmfU7qIhrJoJELfditWskQ3QtSuiclQaWoSnAKl/yEpmOzRNtOSD2/Kx
xLI8qk8viYdradU/Qx9dBnxlEwjp9j3YWuDwovbPYgFgHzFEq+OtPOScasBTnAtYbHNVxAn1toqw
kbldCIMuMhZLv36I6ErBc4P7zKj4k59NsCG4JeKdu7QKzAcyl1pYDR2UFkYA6bJMC/aiPGzPqPFI
s8TWJjHtH7MxrO8xPjULKmjOAON/OGqp1CE1Rk8TmPShrE7mAHGtv8nTifzX1QmGRVZJBGV9Erb0
/fGJP9XjJPgwXGu5XZOKSuswJv8ldlNpg24MDPsrfn5W9E8aV/aBc8adft3EtBnH2irV/6G3lXga
9VTCol3hIyLCMrhlWc5hJ7wZeHxOBEpkw7WN8dbKEk7kSD2EoxfJQjd1/lCT62/K3wF+lCVoLIYj
uUsqTHayXUbI4DC/9gezwwi9E6H4hqdJxeZXNzoqYyNL7GB9uIxpCo7hpvKsZG5jWYPgzGHl4Ikw
coKH46d/khD9KU/lZDSSZMJDBth1ql+YOjE10ha59zK4HPzlj7hUzr1jjVnvgm8FZek4+ZJpl/X/
wCg7/dfSQDHH4zzwb4ftR+qed3QjFrMgPK1CCXEuAYCRh9Wfp0Iyma0CGHt+uGUIoffx8Ms8piFj
IQeHa45rgGGZ+Dw9HPZQjnyS+mCH7ErKFV3Fx1UvuXXbpIrABbtdWzUddOW31/UTC4+MnbfDRwNs
q8RpVTzVhU3u5f+NOmAnKfDoHMYGQt8hOrvTvPr4EFqjvKz7wk4/66pnAimkU6QZHrK06BceTF7k
E27W2/B0LURmjf+AkTslNdSNAUfsbRhF2dTwSwRO/wGRp5aE939tI0AvPGhIkuMP+dEsrddI0iNf
h+ALGiNMIIaL6CkX5l1MJNHtVcmQmqzwAcu6wh9V+G2E8ECZBIBNKmB8VazzXLbP2LMAjQqsKgFb
9Z3hVbWRXzPzBwhZkyi/Jd9kv6lLSjmExrw1eXbqoO3yqh74NYJepsb5YujL1dCfjdG8SX0GuG04
hBPpLCW6N6PLhhAfnk7H7qjTfawrHuh3+VeDYZTL54WI+D44HDAkn0IpRxReiXYLHFWjGUyxtmJA
MFzCPB1/SzMwceTgtyZaSrduNSl7rBdAaals7hEOIpuIDNETTJzi5oSUzHEbLr5CXYnolImdUXRk
khYPNP0TC6UQlyKsBCvzQ3tfs8oWSzaCE1L8Ktoj/fKAWKlOtHdwAHyEcUNChPl01CowGf7ItNn9
lYMNzmZVfbY1XXOYxxa1OsihKVKcnG4LuLSQZo+SeETOsxaRJVetHmdmXd0ewHQtMGQcXbjAEcly
HlyzSjwgURa0gsdBA20obNv9/zJuHJIUtuyY2I6CphoGFn5yGYJDFdw3Z8Ckxw00cfVqL8+cT5CL
3PlcvpR2v3XOzJi2+sNq1W6OmRocx8bodXKB3sE6f+x4J4VYzC4jvmSBe3avFeAa0Ve4tSybiaIV
IsnXr5sfCAEzMeEyyKQocsaTJB2XGaTuPnjNww1e/69+XAeFslxzc97Wsmu9Ba2F/dyemr0J0iun
yDAZSXitW/P049ZCn87NXY4b2vKH7Yt1uZuevbnG8TMlXoSyow4d+rZixF1i8nLm6mRWkEh3PqZs
Q/P+IGBtd0ftPsqPViQ385pwoK0tcJ9BqYbtYzAyXAUaIGaiJjLxL17IJ0hFbA7TdWMqqNIaynil
XjTMtzsUlsbtXp9UtSxxIz0t8V8QhcnybOQYG8qL8Qpj4RKApRDOfGS5vpi/MlJSC5MJ9GSGmJDl
bkaj+yIuMIqqb5yem9oyiiV08yIa1Fe3xYtDNDKpTtZDOxE6YPcN5GDKZAqh9e37ZMEI0L0RIFQT
MbWGKaXX65m/n05UoL2bSDA+HKMzQZmezHK1p9YQidqLYMfsnYSybuQNA/7jvhKG7Ol5y03WZOsw
Y7lnQ+XOcq3BrC1f9Xkr5teq1XMBUaIcXAbIZ9IBbi2LwymgYh59h/IP/3AMYxH+DBF10p+hSuhh
0+hZLu8qX/PATvuj3tbCkbX+nkQhd45cNzk/QGkp2374ARkJfxIEw4SeD+4Xt7HdyLLkgqSRoWGe
HbPsmnEmIFy6R+FFMqscpEq+eaxPVYZGvmGlmRmDKGFVU9ZhlhRokmJ72GapFq3A6Q3Y5RGH8AQu
T/4TSRqEMp5cEqq9QDvkzPLIxPPhq4A8GEKVTDaV/z2Upqd5QOCBlr1MUPH+CcBFR+DW1EIqsVI+
5pR+yjcMsRG6aRXckmbFzIguEA3hGJ1z3Fea1pW538tyvX8l4tJFF6jywFTUhmxutxNiT1PpVU3Y
ZBH6aB9/svm80tPP67xl/FFhxdxqhCFBfnoUqO9xEieaXGgQP0BPWxO6ngzrw//JBLs9eRVHqdnZ
Lfej+hFsbKQZoOd3IIhbGm1ikwm837JV1Knli6SY+GiUfUoVbSgVFzAthMXMaTh1Kx/PuDidYMI/
lZ+z7dW+2DtrE2J4mrx5R8irst5bw8JOELVFXp3n3OeTjGH1it1iaCl4WBEdxakNBm6+3zXKrTbT
3lk09JsMbmLvrXCuEmRODajyGwUYI0B3L0dg9ZjlBeUisISOxHexAi4olf08goig4me+lGvdAWR3
pu9tJ9bAlO7l3e1wArVBrGIYII5562eEQPDmoLOBd0xYmaKQNqzBugvUS5whkmxQSyVL7m627LCh
ImPCvKuIcDeE6fLI5QhXGs/aB2iSiAT0H6qm/UAlR30q1YUXOlCdwtEeZMcdbS+Q5lbOk0uzTQEE
PEsv/9CEOUJCNbQsZwN0HKuvBHKRxnossvrGYVkse0M2HSJUl5fdkN3ryBjNe3I4NfEH7uWyemIA
NfEgxv09A6Hj42l3ASAg8wxGTGMZi9LCbOlX4R59i17yJUROTyIz1JtVwtp2QaWMflrvYJeP66jq
QOcXk8XGKnT7G1UgiqHO8Gftu/qhsW7dbxtTvrNkF8IZgn3cGWJZWRvWEwHY/BF6UbKgdc14UATP
9R9A8QX2J6OPkWpA5b66tHEw1ivClMyxFV7aM1BwOBIVtrqMVWevxR+TLDAYco3ll5Dn8aaNPjFC
Nko7jnhn8CmRtqNMF0sjX+uyd96K4ckhQycbz2AMfTzzsFD4N2TYuZIF1CA5q4HJsZxdmc8NVDgg
non/fQdkaV8BtBnfq0RVZskIRRWqvGBFlG/pkfNnLQ8uvAoU77W2jK4nHedwdSZrfTYCpIzpsxDT
aLvDGrGJNFRBzRP0mRYzXLLubZUXauTxXhS87aqCqn7sgogjZ5Q02UEf1OvSaw3h3I900VMMqs/n
q1iad6PhWOZo273McvugMVtI4GDOri761YgXBa3vZIr0QbtmRBvghLz+BSmO73ZLEFJBoCJTDa7W
Glk5KlLuIgXuHOv0SXf1Sa3hX0mPnyT27hfd8kmQUWR/DRM+cb+gNgaX/QabVWUi42J8jfrLtXlh
q5cPi5BVaYO5IK18Ix7n0sb9OzJy6K9kTEEPm7/+LwrbAjdaCiPbhklCVRxJEpyVQFOtUiUcaSXV
/hYpFHzmSw6ypXBdCIvLwcoFyZXDUG/sTiSfIfrlyMbv4qpbvQPjoQ6T1Z/AGmm9hFdLeBekI3QB
uIWkLv05T+OW3O3mUqSIirifrD28yVUapSPdTxchyXWLxPe1xdhGUnV50NRsBiFJIbjA987HYPio
GUOoICm3mZc1mAlnvFBRTwU6xKvfeUdIs4wZaLIRmK3y5euzWxja5OEji48SYLDj/9CmamJgKXWT
yw4f9cIc9ZKuFNiAWvh8VbJ9+BT6fLKu9zWXQPPrqSEWweeG5H9v5dkzOWKVp9UPT9IovfFhlrj3
Zu3n2xjKmI3lxdbjzjXqCzuRlVxZ9eQwNYOvCP5YIQu09IDdXjSjUDzTZ/rnkOUzlZ2y26+xFnO8
cwTLXs/QTYHwVGgAtWPaOasnCN/bvSCsNCJpNeaQvsmLILxs4YS0ojDz+5fjeC0+uho0POQ6Kz9L
0ZtF7ejWqyDNdjSRtreGOYNKCejU3OSkEYtoFcp8AdoGbaDNBdpRG1JLvN6tIZqmRCxaYi9ta7Tx
HInNYyTG8O5+Tz08j8Po5eiu9wRwrn0rpfzHl/Yg47aT/ZXJPwD/kcPTGYeoUpN0TJtix7cud2YQ
e+b7mp/tmId2nP7soelmIhreETo6njTp0BIU4D+yHD8AYu6z2fKCPvj9NuaspcAJM4GGystGvRTR
QedBtcD9lIqy1I7X7BJpyZGhAppzpaaLKB3sxsKgFyDHjLj6EVh5vbYqvpudEWC4w5L8Cc+/KHFE
RR0BLUxYddDTxYVI5n/E4xsXMxXFivZ2yNTnt2MMDHCpbyGTfYj+y5KkAodya8ifoOJ5jUPj2GBQ
9lJEQMmfqVsv+ndjx6pVyeS1iAj34XINgA1QS3jVUMGTeYR1dMdHvkGFVmZiPpmCYbBzPSYBoXTy
Leyk65BD1CBoiBNRcu3Us+uBubiKtHX3rD6PcYwO9DZuUxXHg3+4WWu/2iTbEDmURITWXjGz8+yg
Ysf7+BW2Uy+GoMb9rbL/OIdxtGHd4rj52oXRL5z1cpuiw7GpWFQzdorYNo6gn2hbE5rgGOsLwIZA
LFWi8cw85eC2B9TMLc3HASfxnac7ZKXRHwnpZDOS/cRJqU3uJBceKmJZHZVcVVQs2t8g9t11aZv5
xr4I4E/q6J5e+ud+5Eo0VsobpyVWIhnYsV0g2X7CVg35Z6s3aV3RWjg828fgsm+6peADpWqCSIgm
kFoKLZZOBy4a91APFovyisZ0neJGwok2TMGI38YkwvuiJASqWSTOtEWuLiod9CMRLz73JhPj3Hqz
bGMbjUJQR3S8MDrKXGFEY5F8YwEsWFOyH9uiCMnYOJaokaM89/NS5uC9jSizUVRJgcrW85LRlvBD
dxt6XBYdEjBC+/giZL+dK6UV3u3QiqzR/ZYYLLqqno/NkvT5jZAOfXMnQGoff9fibv3eM++5shEg
5/pbyvDf9Q5jLLC7bXMsRuVdgPsTE6DIfVHRlkohgY7vuK5ZQ6K1c1TCMIyouDer8UU5UOmrpq+K
3eZIwvNVREGL2BulQOUB78D6A2ol5rfrR3uoR47PPgv/cfo/dDzGmTTfCY7gKyEJiS5l+tbuOmmZ
JyixloxK1p+Ee1jglntSb332SsFQ5/J6VLxnVxvdhdXpTZMIxZA/6SR/eXXb/GHPjESmJWBb/uJs
a0HVFXvYj9y1KVIehXsfMJLNc9CTuTiRGvtYdDQ8/oqwJC08GsUCR82KKme9MGSMDPedBkrWgkTR
SbOnWYhubbAfVkfa3gJYoKJSWi3RRk86eJ0+Ou9zuXN+ro5+6Gwvy3p4UbqHmz5uRCJ16KrKFsYn
jM8ECrQu4RMIasm6CyN7+D2nmVMiXekdFdI3j0vCbyO2zwVSUdEA0rxzSuAl6ablRaIQAI4TYtNv
IpGZUHxj3Y+fXpCWQfVQizVlTNgamjyWc+mY7uZJHeT5/cwenODL+ahm/ogvZvExi2AGiDFliwYz
Mh55/btA1aC3I5Zj+T4jPbaC02enOc1Qh6huahbGCuKLP2TL6CpFUVfv7qnVl03Jjum8TXgPKMQa
OnJm5n0/6GTXJ+b8UzdUnfOtu/vveVqXskeeTqwtJqwHYiWZnvref7y8wNLQc96+SIZ4xlpsvhPI
W4EUexmuIHP8GP4txeFFCgy4SYu5koaCBrbIkqX4C4UROSk89iUySEkpbbqSk/+GCsPq5qeB9xAg
iBKgj1qIVxcocMQLv8Iybh+r6rSa5c8w+EOv6DgG/LQiWJYFzGyugm7/MmVEX4ks+BlNR0E8VAyl
8aISfBxZ5xxCjTJKtsfr8BD2RZ0IpcOyI/ngJiXnNLtzWWMzAtQjtq+dLjjF/R415eUbtpMLcsLN
WED7SIhDputbuLxQYybbvDzqwu1Uk9ZKvQfDKfofZpIdtYk5vPcwF5pfl9u0yBsV9GTQv0rcYbd5
rCsdHMXok2ZTJxdTvtM/ND/omubW1rs5AAba0oqkIw97/MWrBdYW/Z24mMwKxoT376j7Qj91WDAm
0XYPlrSwJyZn3Bh8g5xefnhazv1gQ5mSh0WbZZk52ZfuH6YoToQZfed5wvGQ5UZVnDbWSP5n3i0X
lWVm0vjvl099ZKtXjREOZsERU5JLujFOjIw7T7C6cIu6UPyF5r/4QyJsuWPUULGZ3rZZC2F4rzYc
w6B7uE7BZF6ldb6pIqr9xsW3tqtt0mwXwLEBXIRIL1k42dG3q12zi7G+vDvjleM/1FmI4MhetrUp
f7LWylja9RFIgqbLTyw8EXMb3GBjUq3tX9EXs7P3aBRri1lLSjzvUageEkc3KdCP/LETvpwK/fIF
L3t3Ck2RoMOIos0rVyZYTHYT0nNsF1FyBHtLfp3EurXuKyIU8rqp1jYMu4xnHzVJ02E5KvEPR/qE
JZXn8+TcEzwd2QWKMc8hGT0pnt/CRDnsJgJ7b1LWk7rZPDDN1eMnls4y98HywRWyGdxHgm/HePvd
9IDCa1W1zD2VwUtH5Pmhz7a2ioSZ3tHJmY2W7CkwsEYFEPFfLA9uBf4oFs0I7HBpq8wajMCfaAAh
vLNiWoU8GN/oGd+EFtPeUiZTaLWGfuiIxoxEtPtmalR8gcA0FWoL6vuypQUGo/U60T/wY3H6ptU4
uACb72Zgsk1GSNjnlhSAIYf1jLiUpRtJQrTYqqAzZqK5Zt30/zg969gE96fK3kGNZNSZexeMcaLQ
/PtN2qm8TwWmLj2sBvoJjhPdgKMdjyDdreod3ao0kRR8FU0BqHhHTgM91W6MLMV0BwRuqZk8pR04
fMCPtjSAcJqlpvHMiB/qsbujh8m1Oj8eOgDMCkkQ7VsDA9o9w1MfG59uALIhRQDw1reTsDNsJzVk
WXUhEpvbsurx6423H/pJX7BPoSVTkoO1HDPvs+B2LwFRrxsLKEd1Syy73btpcJ4FgCK05Mve6QY3
FImtyON4fq/F72lBFknxWXMCsl98zVQyMtD8rAxwNxcKwE7L5EaLXBRo4in8lwFWq5iRJdnSdv+D
cMR/LGmE+Nvfe6wbRNTmx+707GEUF/1dE16/asiOE5yNfpxSR9jqT2Q5eKY3CLAGFSRbXHy+H27V
2cuqyvitFw9gfHTcKTWD4SBp9t9MFFsB4bICrcWox9dp6goSO1GnsvKjh8j4b5LDwnWZAGn/yo/w
xLDkZdoxRU6PVVQpDS0Feg3Q7e0PF/pd7dzqdFNwVk02txvTiDyD/vOs6kfhcFvU0M6sz86QF+gv
S4Htx94fElceEVSylzoXqymTSn7xOmaFWz1R6289rMMt9cTMlL2J91cuPyXZhY/lj1O4csvxoj3e
M9r2VOeuBW/6u1Z4pleRnjUj5k0YXz7PG5Al7bXDZAGqY5WvvggmqKo/+TEWAsVBJLXkjttmrisK
xtgoDNwHAEdvuEG6QXThZH1rmkq/T+0paTWfrckBs/7Ipni/DZG3gN4EUuv1nh1Zxh6XWgJInx8A
wiCCcIp5CaBznZfPIk+Fi1P82niZTN0xNyw3PgWTTzkp14JAX7YN+zAfGJU82mIp6Y71tPPXL3u2
tzF61meN6KEVquZ+XkHoRPFipGBtzgrsCkWzQb+5TDocWCYzU0Zybl2zIJHxfFs1GCvyS9eIaVUj
t85j2k8z6OrGLSEVD6YdvcPFiCHLOvqNu+FkGTNh192FjedHHpysN4hUTZUUoEQxU/1YHQXUiaPA
XrSc+21KndPXBfhvfAyW29N0l/Vsapu80Pfco+z0uDLwbVop2v0XzntyY0rp54eH70zhjxKa3avR
783/X4fjoL7dXk5dShW0HUGN+Rz217kgPK5gwB1yikKang/Wsrb8+YC6x4wqL9BtobHu62orJpeq
iBthWKN9QrmaZ8MgBCdlatKHkVtPpUo2Q4vNvtfESgFpSx9pwVTmNi6BE6yyz7zL2nrGtYu6F03S
vW1VtSNSo4wtiSlLT2mdKYIv7Se0SHrY76dAwuoR7BGNqpokt8qZxBCHc/YYp4uy/rS7aG+zaW6M
BbHUNbLFvIp9axEjFzUHAN32HmFyUU0IT47zovAfCQ2nTkcu1/SH1G9z74LwTw8jDgfMjZ29KdQ/
kNUPtTRINjAz1XbLxdR497rsOkY0rTvqj/302swIGlBvHoVyFesqKhImQGpVoXxgmYwFHmfY5YT5
DTdmj3VWgvWmacagSRDjKEBO/GoaXTDRiYXrinwESOBEK4CrncfHVMxQfOtudO+pFOXeMCYX1n43
0A22XlAJgemNPzB38hhkUbHoCcPbSUe4rlhBqGSKyq3sveLSBkfKL63ZdjldcjF5jbzZWE+BDrq7
x8gSr2ObfdzhiuGWCZqZBKlTCTPLf2KUzG+E2Y+961zM8wjkZ1jv9GtIEhkZTzTGsXrqzhUQOlUF
IYxBqKWZ/3iklO0SjZE3SXP8xwJHAbLf/Gg9Nsiqbq9Y6cszjxFVzqwWPZg0cz8sI6Wj7jmeB+Ch
XY8lCP1sOnArMOc7Mj3YXIkOuHwtBgjnFf9xcTM6LKvdlYuRT5TtYYakQ/ZdD1A5fzmGp90a+2tU
rIgV0QdBMPPrxDhAJ+79OufmlIbgPDkxuQHbeLHUYB0cRm7kKrfk6tzAOVqL52wHQ6woMczjJWhs
kGx28HNL7R91Sh5hav9uCHGNaixY5scFSy8nPTCnNXcvx82BKX87nJy2gcUNtm73mVoDHZhI8Cwl
myorDuL6J2kHIMTp3vg+phsIyr+KdJQ78O3vJF0WZFBv+BwRPTztRobihyHc8O0sULtqyhCY5DOc
sXVPgehCbI0WLG+foqTDNyg/kaQm06VB50vLaNKMrWvVJhLa7scC4yjbTQyG+1WJXaJA8jIkhC3R
qILRQ7cykDANhO8cnUAOjlf35Tq7A4ZSG8r+uRPHbTtPJpwHd2xqxXbvHu9F/I726lok5oDGY5kr
lFoVWubQ2zciW/Qh04gLu/Px9giz6v9XkHGuFgEfwaGtCXmaFmGq+l3ZFSJ4h0+RtE4+qXRR08TG
afwkt2VmNfPADSEk0q5JLTrGB5M+f2DOUaRx9LX4Xbo433BGCY7Gbf5iY3u4bUpjmsJPr4PfZfnS
Uxlf/gX5YJP/Jrzu4wHiJg8Jz3z27IqY7oH2eXgbNX0zR1BlY07VLKYK91qdfcltR2Uo6IZVrxQU
nl+rASePtxhmgrmP45fbDHtycWj/Zq9Oi+IARutiMg8Qwy+PPu5IOiDTasNXk9JkzqHq0HgaHAP+
Mg74yvmLhjgSaO/VM4JQGPmcyNZ1xzd8daoht7B0jH8oWR+kln3NNPKh9gKpzaaP9/6xftYMtRuN
SLi3lknmkOS8KswpsY87Bof0Nlmz13CZu6A1dCAFRjqGWnHa//hs3aipS2qVaAh4+2cTYIVLp7gy
M6NTm22BTjb/wR6+5f8T9I+jqFmzOUIN1X3q1yHcgamsBj0gnBWRiuu+uUXpiBIa4obwIElyYlih
pNboDsLPFm9w8w8+UdIRh8z774S0vm6CIBH027U2T3vItv1vYOldNr2dnw3xCr0mmSMvshuLNgB9
YyXuPHSuSy6M/JNS5BTwuY0VGGDrdAvLycjH1qXdvibKqTNWxF5wJjYpTcUKZADJkTld3C3DpcNj
FcwlpB2LtM0XYKdtiyi2y6WDs627jNXI+ar0gSYHe3tDV8RE6+sCHD/96b+corymS77yzFLIcWeR
JvJjYemT1eyBhG2MhptAc9lPNB39cTPFJKpQhjCSoJLsWH1nwU7tPfuIi656YueQ2S0pW0jCtSn/
FyxtkitBPoCI7RkbbkgEpFKqpn0D/PMfEhrlwDmJFyv08rOkHDiw8PgqsPQTLmAPllk1fWzZjb6M
kcpO1Yph1Os0CVhow471NPWzspMMwJiikCOMyU3Gtglm+Pp9RJ+ODHjIFW+C+9Zkx27Qhcz+mD2T
n6MetqADZVBAuTKBFZTeJYA6M7eOYogBV2NdDOUaOam+rCY+z0aZo5z7w5afSB+CNiIFMj8ai1Ma
Gl4xBtpN463BSbS0ciMrMzJpgftpy2Y2j2cG9x0ipIgkg56vseYeT2qvOapRkaDeEup5Ikp5szac
1IQ+KYG0eTvFUq1fCf0NQSKvu+RvhVKtrj2chqOEsdbEBihkMsPn12uu9ASoCDeXuz/arBnNNaGP
PScXj4Er6dXsWaoW5c0ItDWq/hflrotGz5Cg1qShfP8UNA37GEqNY7q11KL8S6XAFAl6DPBM3QCF
6rGHo0n1EfIutsxdySkOGbD6h6K/nSJd2JDaTcz1qNa2x1W19KlhAlNXXWohpCfWallXWYOH10Bn
eGhx5GZOR2ZY4xdSQf/H+A1SbUWPMF6MCxLD4VRxS7lggNyI9deDBiHQ+OI44h9c32R0G9TfTgoK
tj1x//wyyUXZ6QiR5dCVyaCN51wV/+/P7YI4ZlsxnDI7D1hEGl8PrS6rURvg9A8h2pIpwWBrqvqF
ucrbgoLy6YFDQn3nqCpdExBZXSbGZ1aVI/PGoEBVXwb0fQyWR5XYxj8WE+C3io9ngdOeiH6FOLNF
gZV/P+neYG9D6klOyRJgQWxqohAM3WE9smXolpuEiqLYb8LHNovd0S+GnsksF0gBqN+QLTr/a3dz
fms0CdukDqZoHWBnBWa+oHXMR7wo6V+lPAAL4H8yIHcyYwNjDAvovvCbEnzzwY0aaCSwg7bY69eh
7xxuD6fgSQDxfFMJk+hyen87iCbxDiSyDuPoGoEXevlEmNzOskT6MZ3Pr0qE1C7xX/0hQaArb3tj
R1VkOGwubjH6q3rLM9s3+DlldxpkzLPRd/pHIpRVKy8Whma/UPnX/17WcJEf+Pu0p5jLo4rxIwT/
rxgkxF9xaOJVDeGmkoMbNep8MRSWHemsoUzK9fyJifqCehKi4Z4TakwlEudPEMPhcSt4xsTzQ4DZ
EPapTCW0q3PUUxMGZ/CiPBoSWn2EXflidJktHtKNl/ttQzup3D/qllCMFpEEzjxp03GBfrL3SKTF
KVjEVW3pasLil0aUBKgsT+AQVNj12slQosz4AgmmbgInhX1yn3xGrBt3zPrdYp95w0ELKJ8lv5mo
fzeMs06zXIa65TF4QA3D1rJzmQyF5KxAR3pqiwffNuf8SJUTcXiG1nHudPoKie2zzEE/QqSQK6mY
4K4SVNkQvuPgRb7bLcBoOKsqgSt6hLZM+BklDPLPaXY5Ia2uYVW0azg/S4TektTGyNVHBmVIjNTU
y3PGYrnMZQ3dzxP81ikgJ+YM5gkeWXQ/OC3yr2qq9C6jjjkLGANdd5/VRJSGraoWgmHcg36MbSWj
9RsyDm6P31mTgY+MiVYqoelGuwFIN+ubQ+h17nlZ28d61rzOkEs/2rA9wYY9NI6YYLyNCp0nKZYd
YSbMjka16up87grHi26xBhw6k/HXJbsSYvq1RkTFL9x8sNVshpT3+ekq0xUrGsRQqSn6GtENjl5v
+xFQP5SxACSKOOkMsOX69rPaz242EuXS/1BJWnO71ChQt7E62eOt3/cQ+IMbqk4u4sEN9hlvO5+H
fzRKnfz1+X6RHCgtQD2wuHepXVcsULTmGULbprbgBZHLqRlBsSJ3Kt8KCvz8wgQt0373CyGTpGj5
jLXmoVXjmMEaEUwr5lJyxT6zJa46aeSZngfxCZlWFPsetQNWTApyPmukIAFklP/g82UOiv2YVor5
0vxqiMYmmZPo1Woxzp4T3mavjajXvcTguJBDh5gTqaVaJnduaRGaXpTQVdFrC/7sWEKCrebenIlR
eIQHAIRsGLtqvSNiDHD4ZTXN82vL3Gv6jko4QMz/sLmOZgNyBwmK2ojUKMiZTgzAXOORNX2TX1pt
wiOZ6UxiIW9h7gMx+AAmc+FduGpW6Gxzet+Q91SyPd3RWLXTe5vVHqSuKF4edLTCuOT452bsMyFC
F32FhzT2oGsEN31Qp1upLkgkhC/f0Tu2qGHo2jVEkxLFV0MxwcQl7Tm2bd4XMfRG/HcDhrMI3ulX
ORqQiC85VUAf0bePjx/LLVLCT1tbMoOyMc1Lt7DOI2mZwQocyPmWAn039iOpMNRZBFOsVs6PmqXV
9ct6xEBUhMvmjry0cDGMiDiC93dDtRl2X4mOPD8B+MS8kfA8qm5/TMrJEHHgJu2LDwwE7EsnvDEA
UwM1t+Bmg0JynVr2cEjiVXT4qk/zt/Dm4dcg3QZTyUP9b6VKAsNmJ/6FJDDuyFEoFK2QSpIS104q
ldcSx8MefjMCrUjVjgDSVe4EiMCe2npdXSQhbJ7E9I+Eiz3LbAjT686L34BoTRe61RVr7q6RcQ2n
wi/rEkAAZx1soni6T3ctyn6PHc12klraX/9PSAYrJtfI4YqMdGAv2bIgESGZxJUuH16kcu20kJKa
jp6S7Som3W8zuL+wts2oi42apzYp5AKFZwJyn5+NmbfJVBNq4Sp3SrlrXdZMe07gJZT4zXbT5MoM
m0rGoP2ng0CJvUB4tYpzDrC/c8rQkwow3TD7kRTLvptpKN6RtGCRqC76CpHKXDUCQ+5Qdyt79snl
9yy5eNpMmCQiOJR/u2EE4nwm8DG5rRfZX9QoqxlB0VM1pcsquoTTuWJq3hAzPTDc9QxBz1gi7sxY
7ezOekQn4xIACbr/jGpov7IZDTj8AhLKeu+5XcfIcHjq3X7VQicGcYVy5wDBAe05gYrqQ7wEX+RZ
axEXz8/hQcV3HTPjwCpL7iGROveaniKIkJgXRiKIQtWhdusafQ92xfMPYPbt4qPFEvZI9VYTCvDm
gXtpNq+aGC5HnNz8xekEgtka4aCepqXX9JXD20YzlKYNY8WWdP32GrzVPqFM8aF5iZTNUFucpdrQ
bNeKV19LgqpUCIO06IxFRvPKCh25L5O9YI6iZl8tAmdWBouz9E95FVddxrETifihCDVXVJn5lbll
Qo08ZCO3+ud/DJUN4HVMwyKghtk9rVrR+Zc637yykhMvPjgFGK5/uAn/bGznh9XdvuDg2alJTsoO
37ryYQwJiN5qt+Wdpz18CFBOOCFe8LTHpCAe9PWtJOEneyzffuhWwD/tPRdqw9+JEj3EeF4RWu41
flyV0g/Y3pn8UUqzbwsCeBhdzhs8jYAa947DrAadYtJJY5prSR6QCba0xxt+C75ZLcfbpn+h2cfZ
rlOxywMFIDHN0Tthle2HpWbmFqFuRupAvAcF/38Q8NvPDecxI6Dk199Kb0hkOQW4JlaiAm+M3bVW
HOGG4KetpbsQg8e2mhnOinWEAwn9JeutiW+KlW7AZaGVSYF9ce2X+q4Ld19fO/X23NX65mlE68/W
B/glBzM0IbO0ftG9jZF9GkCBB1sGawff/hDmlXOueqaaEn7lEYOJ2HFlY/1KkJhyzt0pnOofEUkB
VRyWvTi3xcZoIYOpxttusV6G8rcSapRLjvx7AX73WWRMzctjMRkdkAtdSzuV7wiGnSMVOEJaL5sa
mm4+m7oz7eC/4wogUH0eyrQVNk5cz2DIo1EZm5BRGgnE+NpPfzJ+F4ZyPgHHFs9vlShFinufe7LT
jBSB3NClAlMByGUHI27iGHdRUiH36186cX0QjNiAmaYcWsId5R6m3Jx/uPImwD73fEpFFEJLc3dd
/xhlgB/FzcPKZiVcE65pffBTh+Y8PBM0rYoG0qM/4Urw+STMvAIPZKNPIiawhynxusMHo5b0w0rA
DbFxx0zIsMgQ+izrzhYwZGB/6/eh7ZxMoJM3v0l5hzlebLinCIGubnjIgDqxo3ND33z3WhvhzIQl
BHxo7zaIYBLQH9XMnKifxLJALhxerMplU5iTI3025KUanrG2sT2hHgh0c4umxmHdULZ5JrUweVAn
UELckQC8PvhtQ9gRdHI92aONsED4bnApM5jr5IfCvyTc8SVtSyY1SMY6mS5puEOw9gsfKujeLd5Z
Tx5eGDNpVLFwflfc3LnsYpCNShYoheNSiH6ngbpP8xHtaB7bMSXKajYhT1gVnTA+8xIb2jgI/dB8
oPBGUnL0/JgX2eTyGWY2QA0/H9jtwJQ5rtmCtTGpxOQ1lU19BAlsdDWAKze0VKFzcXvXPL3cOnEh
QpbihfeJufo0IE6U7C10KoSsYVN4xORQpbBUs7SVoqwZ7+vuNAgfYA6EYixZFxrf/eN44g1K5Pnh
WYXbsx293JwMathdQM2Wd826bEU9Yh+9hQRgLANlwFb+EeSG2jWPwAirg/mEkJbqMJBeO6NQE0BV
ZFwSFPYdMlBLUeiwBZusKMK6s8yn4sIdA76GiHxJbIYWhi3SBu+GlW4D7XAV0k7kj0Qj8Nt6zMge
cQEUoB9bknlhhMIvWiFId/JoKbUHUzL264wrsnUOoD0S1BJIGiFPF1RNEK2x8KQTEEtwtX4Nj/vx
W6Gwj4P2pVpUTHcMUj58DapnczKGr+c/YyWVMwvEupYAy1gUEQWvBDzu8Bloaw1N0IUdOFD8AaBZ
NXew8Ix6+gUgyfmqNwV82HO9U3LwOKK0kvGwBnYtq5q8bE/+zs2vfCWiz/uA2ocO0mLvshegj25W
V1gTmueTxbh5N3MMG2KXmE6Db2pou4xKISC5GlbF/+ueUlO4/JvjH3VlD7Wh4WAgtDTW+HOog2i0
WePeEptA1lXFXPbTQzNP0uwTpps+Trs9kHu5ac1lkElLDNqViC7ojRWXHb+aVq7+fpHcWf4rhEBv
rMqv+ahOXSHQGbmL57Wt+p1NwvqZcxSsfMKapuJjmn7Gf6Tvx+nI50Ykh6lvvFpAjYSJOJmXL9Fa
m39jpdDw0C05QM2cApbEzw8hJfRWBqOIid4c7K8KiPjtDbp14uGNrvNKFm+H7Y6LOeHsX7MJgwvj
7nFSPe1cgkjtDQJ8pFITX8cT2qLLqN8aASvAhhgdgNbjWCZgrfqeJfG5h0JiOQk2SsQOJjZ/J13R
f+gimyAcAt1ra1DACby3S71dt/St3DrjbikQIpXN+EhIQ10EVO9R/kagoGeRDU5MynRUedgUFj2R
f8zEQcMaEt9Iu0c1ieoovWdccibP4G0V+mtBWC9LUuHzXh19wEYvOED467nNvPx9GBgUFjGoMlaL
+d5RmcZuqtC6klNZ0Vfgcmya+91epr4QKRO2pt1U26XB4Q3PQ1465sJGfOeaWCPSUH20tgb5uc7n
6Ny9gcHqSFGgXcjGGsB+b3I+Obkyi/xU5mIgr2+aAJH8eMgsXKzknJ90hcowX8WylVYtMwX44Ayy
fEjl5uFDDkA77DEku/VhTNh2AWMqXTSFzckCniFEYb2158HQrddiRNcv0ueAHIrklzPKT+fEjyNe
fEx5O+cgQhlDuYgJc6j3H5MtsV1qUoxxcMvtiwZf/Hy23h5/2L2ZsH4Fiou3fBXUdprJPyFMebz0
LZm9+/4rfGghjVSsTxhBtXNU67Ty8mGs50JN7Y3DnM0FqpJHksLtot/uOJ1YHyxKjjoRAQABriC0
xWRTmjoklcwstgs9BeJDBQFCI4+UGztOZi8Y9y76RlLZbV1hbT71JYmF92bRFvE64hrlxvPZy9vn
eWryBWsftnFXEKQBzh6wyUkP1DW7RWqId2twYQlpNzFEPIMRqJpsquajL/OzBQvvlRZytsDRSSGB
T1RjH/vaBpG2SoSw0FVllC17E5l92RXDJT3VzogRPyesuHV3eUFd328cH7LUmlpVM3iJMkirr3iA
MxP+PWZdpnmu4v8LDouzhXQ0kfwCtpRkW/AYGNUv1NoIdf4LxQcKrPS228kZaPOCXSofW2m8zfVa
Z+Cz18rg8v6sLsqz5YFrNn1otLwEP2fOaCez0wfkuqXDgx/+vungeV9VtzL8J+twg4qYLgXiu0Ok
hoDowVuTEU1fQ69w4krJB3Rjuo8de4Vj6EDhsX7CfSt9SJ3DgwhcrFTs3uROi2aptZT31iVmIHzt
NgJtBT219lnLGyQPzCdoDeBy3UN2MkzWshqSe+r6K2tAlNg8Ufs4s657YNQn0uZyC3KnS+u7Dn34
VEOYBXATXGqxzly81G5y3rH4386BkCaZCbPUk33sXylghqfJ/u/dwUMy/lIHOugN9XZlpp/fLpTd
0XmU4B1J725IA7XwHJcMpIe8vy7v00PBhy9gV0AjB2bTMlMPUnKBZUzr56EBup3y+x7zkkJuvS/Q
FPj8nsxV0NcVxTZS5eEPIdn2szrpxciX7ZFEDNrXJOWaiSWoVn0QqySnoTrKlcNYNkpm0yISEjAI
tNwfmpppZR1KU/AWZviPryRwVYSejIp/vb2SAfQN/DXXDKfCavKWNWQcwvdBlKB+DCMVtXlfMPSL
EHjZ+Fz20aES8sYN94bVkJ7bgWe/925DByly8+qnJiw0jHmP9aSnRjwjlbWSc2og5lBrn6mfFB2j
EKz3ajv31UPEyBj5GmNRjmD14YveoN8IBs96qK0bxw25tAGz0agtgC3qjCNlseHbe8H1brlAx3Td
ZXbzkC6P9a+RAVSQ1HOtUQL3CASFCPsd00PFqT408iZopAK1QYeOzn8+Qfvg8WAp0KnecfsFUtg+
iYo1tHdD+XIvFz9TercMlRn6pvNpLQl0grtJQdIyVMTGcRD5oZOAQkh8zuldZSpJtmJxUMpovckj
6qCL0QMgL1E9r/T9dOEQrd0QV/99EQQ7CcL3D9mXdjeFpetLH+N1QN1jLh7kp55ibgPsChhKxHj7
ykeoEMiS107QhwGgMbgJaX3eTMmt6m+psGIaE2xo/6KzAiqR2t6PfbrJljDGxi5KLKDSoEoWqD/V
Ld809IHUzdVew8Fv7SwnDYxKOugZ/TUsqgqlhye2frL4eDf497c0RB6Ptq5C1iUVmU2+eF5DOVsI
5TcmJw/yBMr8nmjEdXjkhE7+fzaOTyRiQGMLATupZtKcA0D2RFCxtvL27ElPQJpn2rD8Lm6QZoth
hZ7K4N8mcBRsNARSBtrjMjcGauNUWUzUVxYYPKcoxz3MB44pBxSeUURMMDTODkHRmtEbeDfWkS4r
/Z/j0NUUa6rAwB4Zn/gIEk4DJMcf4Fi472JMM9hkuWC8iEJ2owLWuBzOhq/GjrzOeVstJ+0SMKHT
DImNKCFNTjfZCgeHouffUcUDVAEFtweJO1DUMw+hXLdO29COBJxbmyaL21Ofvw8DRp4ExI5WQQMs
MC0mW6B1DyQkLh8u3Hi2nWjNVzIx2YhnfQFDi45MBp86+veyHCAVdt2A1glJJMcybVRN6riS9uMZ
9H/tjquBJi6zfsYaZ2eGtN8IYacukC+zqKGdfV2IWjz3wK5Ek4ASb/4x+s96pXOJeCsg2qw/eawP
SiHPmRE+kidZTlDjOguk3d9lg3wzg3RZm4ETTfji57sZxGTb4fcXyspr/gHMlWlVno5lGIOW1H1B
5ejOO3It7BjxJW6KHul/Suwh8h4qu/8RaBgAknycxjxw+SoRKU7CBAjh37LTsuD8/V9sAGK9DPKU
bOQMmbDPx9DCw6gu5jwvtlxrDI8hAH5UcrJpwosc5IUe78fZmjZeKENhigv/e8izH/sx1IysHzjm
aiU2xOEsOzVQi9+O22sgCScAZa5YFpDxOc5Tx+Eluv54pNwvPGxUuH8ggIdoqt7gwLh2qdm/OTqq
DhfV79NkHTcVCkvAhFuMIgolxxGCPiwsbxnA6bpU57Le8YNGDqQsKOFUOqmj8/2GCAGy1wbjjC0u
Eejx/N7aO/06+diuLD5fiYpChQnI0r7PdC8inD1vDmhgPRclrinNXEfIEth76XXA2OZJDk2gpUKb
j8TUCtl8fjGMrRmt0vuo+JNtzphVfIX6U74BHIm+cViE6PraG90eK8STNEIPnatUWk6C6sXKAg/k
ew3L9Jue+bxFzUIB5Q398hAFCiHhwWQhkjNuPS39dZ3Qvx2np9+bCAnQ7tF0QEhB2oT4PR4r4H9c
v7TYkzvOVmCKHhRGnhWBX5FAMgOolAFQgFcU4iUOVuTQ/GQOTCOthXAAURdpeFA9+0CcUwUO6GgP
wFcOiTGn+yEgDdSl5Pr4AfaEGrQzWgcpTjxAPjD3WCzOGG9xlB1Av3/jC5ks3/xQNTKBq6PJIajl
JtB0n/pXTViJSGf0tbmqx6iwIU46lrHeeupnGvvvg4Eg8bltNuLHaZhNdpiWL0Fd04Io88ry4eBM
ULNszBqrso9f6W85m81dwnI4K6Y8b4IYBgKfwhZYIwcxzGSh2kNquFP8NYYd200C4QYWSpq5rniE
ni0X1RMg5Cblo8Q5tMRIcO2+Pgf1c3xGQYImXpSgWD1ht0p+Xk+RvbLjGWOLoKY713lLd8rgqtBi
VrdDkFU8/buXXMm+BOVPf29v7OSLANpsUP08MpJoIES71dESVLdzemmjbYpw4j41STqUAi3gqvSf
0rSHr9rigmXwvjDGTks4259hQW3U32fCBjar1OXruoKMSIP85uT03JwMROtG6/kPAdQQ6zO3C+Wf
vQ7s0/Cg6gTzDCVlnP30lZMp377k7UqA0favCnT/K2FEHJT3fa3Co8hFGe8EcX+acTsyko4q6S6/
SW0zIXvdlt5m6hAPJkXsboWTFP+1cqXwtOdZgrMtBCGK0ss+pYLwuNWHLxCnElCFzC+F7ZIKMuh4
ahh5yGGDcNDKmhppkRs79slNAGrB9XvJ8RhssF9+ajhu0yqQ4KRnzzvtgkar816mvtSvf24Od9Et
fQk1JWZ9Jkz6EjQ780WCodB+s9e0nhb4FM43DzV5bKp+oTS8gHu11JFF/4/9JJ4zC93K9GYjUzrp
haEr5WuQvOxGOVuDf5fsGgZKVwjuewTpCMVL5sSmKlTYPId//sIwms67XiYStAzr5WaO76aM+UKr
ZhRqpEIryTrm28RNi1afefT1x3cLvckiXYxocHCZdEc3McFphp1MfK/ZaDf5Wyr4HBQDS7Awaki8
+uhB9mWypRU3OJBmEhCJ2kxkUOwq/UQacrsu/eWADCOqcE4p6ZH4QYcl34bJS0MvGB5ihpw54dFt
DmF99Tuf0Logu8x1EbXHBSZOhE6rr+xG6qyvX9Es3KDDbziklfjs5141IEeIoZoJNrthdxYoifXk
pNkI3Cj2HpnwpBLX2hT3r4YKKjrvPX49Xx/bbpwx32NgnKjdJPxUmADCK+6TZpVypKCxPXmWSxss
Dfq03Eo09SrIqduHxLZkoNuDplDOhzYXRdZkPWunA7RiHJagLaToYQcjiBq9IOYw/IP5tZf1lrMm
P20L+yyvQifyP83IloIhFjwAEOx4iCYizn2W4RetuT7dwEGFCb94Mo8BrKOnmftzz3FaNrWE42Ua
u3yfUb6LzzXpulu5GOkmDG91gd6iLmgWs09vLI+daZoPlBkyXc0TTbelHqWbTTlZWW3BcWffUdJy
vkmdXGF6AqzHHT7fsuy48K5D8dNT3Cyaui1NhVrhLKyPAW8xEUzifK52c1TTI+h5EoIGsL22qhyY
XOYmx692D85xwOOaeuNh/G5eXXO6Vw65Dlcb11zbnpI0Dmw0Rdk25agEq9O8jRoxhDQIqOIuixOw
ucbxnUU2Pei9cyP1aDha1LTJ2RHmoYV8rB1GpHxgvreOd8CnFG1SQVCs5iVtn8dUz9HBYaSw9KEK
rCZQfe5UNEY9CCpAiaQgEwx5ZK/Mg4ffk9uw7zW9RTqEhMiQ8xPV4ceyxMXfXyOb8TZMZ/IRU3Mr
oqa+zB7tvfSghhdFLkJQG2K44z8i6k3fCOQfK1gPpeTkJONcTFHDz7Wz5US7tvw5GzzJpZ1Q+rij
2gAIy8UCTk84wcm3bZVFzhpg2+D5hU23ovfE4xK95ePEjnFy2rLt0qq/Z7V6gkynB4JlHPo/+WFU
Gvb5OMG5ZmzGNaA9xyaaaSVReAbcIxKu+h5AC7dGfvzlN5I1hp5/G3lDI2EeJrnsYGgJzzoF3Jly
4BlUZ2Dqq3MjJtKTjWSsGxOL4rw46RKWS3J1bxVnPRjnnbpOKRvvbO86lhMmMKWKcf8B9k1BfSho
ifZlsusjMIH7tqP98ICEIrULEaerIGe9ZxjzXCoY0b967HYc8r2QmWZQr62IKJ7CEal52TslDLoN
g7BHNmw2BbewUrGTvFmnow7dAh9w8IWjKoZAu1xRFKfs72oxCnGtOLanp1NqSDkvzaEvzSZcji00
ZVteh8gFo4qYZawEmRfqgNfh2/KC/3mJ9slKmH1tfjLlsanl2s6Oa69fMuOumlRDtSY8MQJ6H+NK
MGTcWSgaoArYB5VrZa9FesW2qJCyqWpX+FiE2n9vht7EpTRrVkhEONRm+5r68jv2+6VMk/JdV+2i
JNd0fEPmyG4FaevljHL/4d3kf9b+YHIwyYK2MZC3djLaqmoqWUHC/oXyFd7tIN8Ge3wuh33gvzCh
H9ULq2qJqBSprkjBrBrX749IEK8n5NeHQd13u6VWb8pRI5iPuV1ILFfwe8dU2jnhvKSCFKfjnafp
Y+wBPac4DaIYY3hL6BI25gmYmwibL4/yzjT1hvvnj1cr5/sv5ROUmmraY0Q47eLyKCIQ2F06yUAK
kCI+zYVsxtj96vtZ5KrHJoTlGx1BjV+pxG+aoF1IWMPvYWXs3THszYgQJ/d+P0IOsmjz4DDaAW2l
Im45UKwYGbP+7E2UrrwMUrxzJQpD1D90g3iwfuKvGeRNlNArEIESzqFXWxq9MyjD1jzv2inZKRF7
nFGVFgC5ezuPwzX/g1zdDiNg2OlQsx2k58W5DHXszZUSw3FcDiaTEkB7hL51Z4MqevYTakR0BRYY
uLo9NR8WblHwk1HRqxg0gGMbRintLil5JKW3H0pakN9cpALoXJ9aYgLyhuwvkK+Z7sLe0Na4FVO4
7ljeVv/EVeJ9Icm1UIXX8wxlhLh00ujWFCtNeLeZmDFhSG7V2vBAaBd8xVioguKsYtUcKtLKjZF2
T3lcUgsgEFgahD3UcYAKRTenRwmh3sJ36NIDA3EIpS2yJlu/ugqiFZxBcs24RDhgGS85Q8sV1H2v
SMR0dSbJtKsHqIWg2F2zySD/jTkOVgCaWpgOsJ8pqxN+cyNVHH3SjC6lhvlk9/muXGfE1fIgdNFt
hzsArRk7RZSehbeULwUm1dJ4gqMa+unGu1dD+IbfSdXjjTJvAWNrn+GWeyWLHzVWaW3oeYRC3h9E
oXKRUn0nTBdw5tKLmg9MBc2F4J/LvuXGtUagTKxaaGGgobgS8celHiZVX7XDeKW8TRGie9kBtESA
yCKifCPGFfiqljXjX3I2EGGFnNL+RUmxKiIL9yGlWmk6H13lifLX+ONibl0+VwSXvH0xz9mpdYKO
Mt0Qcci+i7dMZLwukkvOjpESvzZ0v0oqKiQEB59J+pvQc5Cd+pwzufc98lB4OHAZtqeoodGFrk7H
5Olbc/ITZTDLJRbmsMwx2QLYXnp3QJXQERQcbCw3Wwsj0CGZxQFeJ/Cg52xiiA8A/UrhTXyrkAja
ByP+RC/eMoy8u0u5RJF7SuXPoSN6xqW858CJ/t4SvPTInhsy9pBAx1HksSaT2BnTOtj8pjsnaQbn
2McaOnvl/HfHZ1ziP2olCx2W2B+VW6xkZgKz5UCkNry7nqXQwM4C4XdanfscfvqgpEJuQwovwjZh
DcFt3JJObXobUrWOc49pXMlQ6zOFbZ5z9Sx9ud24MumjJzy4orACgaoZOA2ijoTF2fngL2egXpy3
G6Y1iIuCn4eAyxH74VFkfoRUs14ZIe8ESkXgB6kUdAqSoi5jewHZ5C9PEAfQUOnMvSQiZL8u8DCh
Su/38bz6nUgTSA1zg8v1rZeUAWDPEErLeWnrg3F6WiBRDpFL/RPpEtIko3/5A33BV9mfQotVnW5G
IgGoZ0sMdINGWpUgZ8gr1jOaOqFwNGGlNY64GAtVU04tepmMW4w3gVa28CgeLrojfv4CPlrO0kz2
VChj+ofaXK8L8Bq1ipq+WtUnv+D1kmyjW/PnrcmMQT+BkmVuVrunnjJAAsG9854iYoOElhgFq9TP
4ORzdXDb87kT4W0KQ22dQE++CxE4S/S5uS0s4A+GU/ebwflUj5376mA8ZnfNQKYHM+K8xaEeFB/h
rXfIpq/XBbjgTthia18iQPnrRJk6a1tN8UxutywFrZW6KBP9B6L1HJjuZ6iHbKrYvUgKsOqb4LWN
2x12OhMEelepUq36t94AodIybwVQ70sgixPCKrpzY50XJWJJrz76mBB7/y2B/syMqErxobfedqkA
22VQ9H/w1SYExOlksFAPtclGHb9RsGlhb8645OoMNfRrHGGKMrmw3OlTJLaCGKwNZetzYwveeVdB
DIITqZPdM1lpvLJKbxabwJ1BwhDDus1cjk+PII5rM9QFRfmIY4sWBCoUbfExRSAKmxb3TGQ14sEw
WS9qJmwTxDtxIayIlome9BRqLiAnZevVpg0X65QTGncoAaaf77+hIoUp96CwKu7zgC3GNyR7c5fB
HtYv9KKQShcNxdd+uiYEVoSfmMCwNGWqBNTNEacq7UfMOLlr7z3gu8PKxlXxzqfp1hMjFOSKTZD9
SofBv32qaex32wldUlOUbRcGWmEGq8FHN2kUTiCa+tbeooZFHXAJcy/oFWW44mWS6b4XaPCZy78i
ZF5hANL0cp25NiFMySBRMx/NNdjUlw25Goo4pLjrHcKGlas3oLa2xD6cMs+mP65HUsoPeakLhcUl
oRfb8nZBr8oPKd+pk5NCvLrNjbCC+Nm7GjGwZuj5FP80BIBJxlc0wZx7qCORPcnCN4Z0d5EJjWKi
P8WdRwo1s3CUtlxIsK6Ls1MiqFCV0p6w8Mr3R5ROJvOw0cn38+14QX/EtPe+EKhd3E/zjqNvN9/G
r6q9QRf3JpwB17wVkueg2/7zg7Dz380xM4kIKk7m4b3sVFkitJY+TjE3rp6sVJS+t43PnMssXMiz
DjTx9BM0CJx4PJz76Uwh2tyLWVnbPwsd5ATUsa93l31+QjRolZhLRaFI2UHKTZTLLEV2jxXUau+b
PEIep0zotR1XxVwEhnT9wez/D98NDqlTo+iXZbmiDA/4peNPkn6Tqi3zXFf7gJSL/KUue1qAdO21
8Dfh6763N91LkmsTjryy7AU2F6tCr4+BQZH0EVIhIlI3zsEWq1fch5pnmB2PciWnWwn/wvv6btQP
uZmHxEHbUxwAAuLZxeEjHb/MEOCYatwjvKFYDgXvvXVzGuX4fyMu8Bemq1q2UnqI6oZMQK5SKMSY
kOv8M+LkgPid8vjT4700Pb7aTFhRaBFL/TleKwPh1jK0ZXhGt7cLq3RNrLQLJlL9WGZ3U1NtD/3l
G/uFDcFef4vRonKooOvllgTPs5ltmqFTMQAKTYoprLRcOJb6Tpyau/NO0vXhjjB8Zk2hw0P3l6Y5
G4EeFb8fASSCllcY45MQrIjvPmtN30U0IIGXUObb+Pj9bGXFhg1jgrXfGyiKDaYevgw4CQuGOaXG
ikwvF30ilW/eHJbwe2ISzjHScwQvEgM4sjuib/6qdfPUr4n3IeYUohDbvfLAryofNDTbBdLuiGWw
IB6YZ/vYZOsYHcjyubQzsm2Z1eDQVzWP8+mmDflZvDzi3/Yg9kkA134yeQAHhK2IF6XhBQYyH/Ym
9IcedYbiQklMnh262L8rnb/qpRvxmGjpcEm+qu6QySg49GvYweif1TVFC3CgiByLTlXcSfsd/bW/
xwlaG762iL1n0Z9mBfaTmM0mjO0GlCq8rq9Vp/yoP1Ivl5DmYYPwHTjRCu/VF9NsgUTLGwMWMF4u
a6/tkzBTGqUA6gd/4tYnkIrSAtJWpvuNr6ksU1ijiTxwAqWslYRuBi5yn5vdcPGGgJqZMpPdGzMs
UB67K6FlRwPQNbQKIzcNkgTmz5fOUAxnRQoaVC6XILi2wpHdPYRFLQ1vJgtCCh87Ut/ckY5IwFYj
sWktjv+YoaTbijsvJjqJ+NncX2BJjfG/NMXZRx6ff1o9v6URaOGzLGO11CgJ8VuXGR2UyFqxDSQH
Hmd6EgKjnKfOd7SlBp/8dqTTe4ehc2VG3u4FS2ssLcjVo++jWwsV1ue/z46auXLVk67ZcAjgn+QO
9rPXkxwZ+5CGIMODoUN1k9hIn9gUyMflISKAnhyjV0OyE9jMhIROokACJIFUJDz2aXWP5sCcH53k
ghv++qs8CZynJulIMT+qCERQOGROuUsERuug7MN6iiDcmuoHoQhZiCR/p6abVZw82i9R9Xx9gPME
tqS3k/+yw8b40CB+9Umojz0lRuwXIGl9xc8ou2VzyKbSQy9/mvPPJTdYetgWVwdVQOs1RLonMlKp
wkT/U1hCVuQjkp4+sJyEnk3j1LQ+ZY0mGGK/gsuOav3FBN+4m5wGeYy14RaCLUAFc82q5rd5XldV
QRvFfD4SocaKfj/IyXCXum8KwUnOFbcbC+ztchJyOKx3VRJkkSrLXQpjlNuIXGLaGYqbD6xtCe6x
NhhuIr5qo4VERIBCWpkGW2LBnWiIcQ8JcOFwhfVl+9no8rWG5M3sYCmzyc2jxo21y1vfAW3H0C52
o8RtPgEOxyU7GdAGaYV6lQNxFglI05l6iqHQk1nMagxPxnbDWsM3anFogIa195FygaAlRpLX5fAb
N9HaPvDqPe4rUYDN65VBuEo17i2zN+gVO3j5dSWSznUdt9cCvW3AioIWD/1xG0MxVZ2pOcJ69nbr
vr5IOA03EJpMhvBl65B4ppAbtP+JrJrTdJUJ2LaS4NvxBz9+nLXD0oGIPAUizntHD3lO9pDYWiEK
tVk6qVtPic8tVbeb6xR0htlCJHdkIBqa3jGRCIE11YeBGIUAC6TtAJSNNhrftsMyA6hC0z0SaN8r
JUBwQ0NSukAFL47u6WSufTAA/4BYvAxmKwOG8+8zZkoDDNl7YaepVeWL/jUG9zaQoMsKpOfjOdx7
k08kQrcH+3Dm4K5jdtThxwM/6fLhnOIzmKe6ZtlT5f4vD1E/Hp43VU8CxLbJmGHAJRgKZRJsOiSt
VVocm4xX5O97sn201sUCE4bji8hVePz+m1u/SwJetivfx+LVIO2YLoMwr36VEF/b91KmXC4aFtyU
KYTuZzrleD1CBTzZQVC8sRWOSHlesDDflI8dMUuDRK23OmRx7an8WJzAMUr1yzt73IzJz7rxKZfz
iaTIEgTMH50PQdLhddVOxaKwXTvJSJ8GfLQ/BaFd9jG7rM1Curo5i4fKNtmwFdEVLotjXXoUsjcX
OL900JVUvt6U8VqunGRwtsi+QZ0lvuD9BtkfUIW1SsDEYFjL3GcGsL+Ssv7YBnz1690mnFXrppTv
hglJ1dht+fqDE18N1FxU9kd9GIjIgp9qpeJ4uBMiC8tzj1dKJyx6HPxggN4JZ+8WZ7wAFu4Rglan
p3mBcYyji+MlNvapl8OYAbB41S5ZwQgPtG8++ySiV3cOxULHwXHK4jLkLNkENkX+3OLZy8LsbWg8
Y4ryyQGdsNL2LEZz4F+1vZaBYFqwhA0UmXIUXxCLDUKSibhn9m51KSld8nPW1qx5Exekn3ESTpXC
SgJ5XvB1Mvl0jlraHyVbmpcAzHY+U2qPb4m3mw8tXEemZzECUm1CwiE7xdcV94cmmT8d0CuchgdF
0bKTFdJU79b4qJa5aPFKr1K5NmUQ/WUQSUooXFzgw157e4wc/SG8CJtBh/d7kUXNp+fY0ZimiIJr
w2Yx3DMb45BmjvnKievNljk2tRnmoJAf3mdVGTkWh1CYMmiBAU5BoA9a0JSexhIGaNqnv+pwMYKj
sJipWyzPPm6KKywHk9AKnaEa9Xpq3qn24d+H1zOxUqdnZXh+fjc6lgvHSqvO6npaAfWGiqT40vjR
u5QoBsmbiAhjOqX7jH309Iami0LOMLSWFRZQWpLYRCfz+hfaM+5ezcmP6jNqm3OvuGOWDGexz2tz
a9tQnwuLnaWfA2Dzu3EaTtfg2rC6Q7CIhecPXPW+Jw7m+HfCHOFNfn5z8vcyLFrgL5+ODYpbaftz
eKfDAj+lEwUdIEat6ZWvufyVvNO+P+KJcwfxyrJ979EiGtsNpPBiKg1UW8JyIaABRhHHIH7QdR+W
plNn1hljY6sSKVBQLW7+dwlaVG4jdqNBaYfhcMafBC92RSFkcLPtZS/LmxI08CpdUtRYCcVUT8YV
2ZFiGaR2QyAZuok7pNDO2hDPyVJb+6i8nM7+R4RHBmaSL9BN1jU89rlVRq0oCjnSzw86CKObFoMn
Oj0c60EQaVk8rXfTVKPSGjXFwrTUwpWO2FAeZBimHyvu+xT9D0gjqxQzHAw3WyMwWm4KeOvfE5fG
7sImw3jDkGGVsLqSpag+jL5f36VGDHTRG6pwRMU1YI2YIOctndlkH+zoYqjtQTUN5HxKWhDOO1UC
LVNXjwBPQnDtp37yPbkciapgqtk1/riNCk+fyjJL9N2a28YSTi8/07Z2RiwTQ4csQKBQ2pmKSXTp
B4CXyRNlP6DOHZTRAx6NPtJipNjWff2yuAmuC6bpKq6lDp+7/cZpA/EQ7rXx0Bn2U1pvBrP2ha18
7eTmv0+IPjugWfS9JGKOM/I4grVN35375KaIYO4ulrkriHwYASDXo4IWgsAR8c/ngwnrGfWuUTGa
ckQrZSeryZMjxRrdVISan3+ZMDVp2jdkHKoj1P05rnLKFe2ZooS50w2wVUrbjRGw3j1HMcg3fmBs
SWGaNJSLT2ixDWfGCzgug5En/0usdynKyMx94ig22hCigG4wVWXOPg1FGGD1hjw3nkAq4jyEHZt+
WxvPe0vjO1CWqwXVxNuqk0b/ZHo6Y9OuXunshS1zzrT2Le/P6Rqoms8J8AJcQpE+/Tedo3VwYjP/
KDoXBTVLq9JmNqGC7eFwiR+99iWXzFkFccrRBQ0C9f2xfOTQTksH5+G/pRhUXOlSYSYrGOIhxXNq
WXojnP00FWCRBm4wZb005Akalgjq28/Mzjptk0UPefyy1MDRo1rUHqe6cd+o+ih0Eac8Cx7fyR7j
nWv89SN60Im4ru/l8WYOtNXWrU1mZL15yVmin5afpi9JzMcpskFBEmEP0SQIRCVdNqlcypkyWPj6
fXEJhHh4okEYmyYrRsxclJVdHVVwDtYHbEdVxgB9prnUAtlLbz0HQPDmlSqh7TWHq7dndrgrF1F0
SfeTu2XLkPkcPoMJVh6iWOIee/AqNWQvk17+3Rsx3LqIdJKH/2snqC4Ajk7DwNUBIMIKIRi7oRH9
MxQCD1CDIuPnvBvxlfqrF2NCyTHv/gqKdUy9FaQg16GBCBFoB4Eoig2RWGlf9YwEWjlXmQjtH5+K
/wHmzY7pFXkM79DM7KviOjjbVtHS+TnrsyqFI5Mp68WButCfOSZIWr1fg6VrF+kHC/g4OTaTcgJ6
F0+eIPqLCK+2cCkeyh3gV+P3KXRV71Qfzv7LHBiIkhFUQwCnAzp4b+6RpFR4rCKro3WuOumVFCrh
6HtvvtfHdZ9gB2kDI7POYsTE/IrlGQsKAjCIC4UaExtTrmeXOrDkB4hRYhGqj0G7ULbpmrbu+H0R
rFUoVjXFsRzSvUlErzrC7oa09bU+f1Acph8mNqLTK+vYPXblBuxR+WxG5xzhxFSGHnLcykva0oaj
Z6FJmTRGxpB5+GIXuhiOM5zfoYVRnBak4EoifmKaMMr+xdCU3P3KpAR6vsI8Mp7nfTNPw1YHgshk
ESQBISpimhHIt+io2unEEdWv7O8Ol/bCtbyeqMI8BRppO0QtC8IBB3y0v1b87eC4j28pDH/zfY9E
XCqER2ysvzifuA0jh4zygiVKQi0P5KYG4hhAptq82tdzn/j++jf94X2KjaaassN/DTcpVA+ZoH8x
uUFdiG2SkjolSBe91nom5PmZzEYmHvq+Dek6MKZgcx8eBXMMdZjthb0ODfinHBuRYL70tyw7vdTH
QEqlM8YluAUdCXUvAzlyuqSHxPQhwBoQhAWUvCV95sKRpw7Rhe59EkQXPugBmlQVDQxJ08NhH1LP
hwc2Z5M4egEe2CgMiljZP3PaccRNJ/BkvjKWjB+gxjfLXdSdjE9rg/5qbr8dQesqQkgsrLe7CS16
9nzDHOIeAz57hVUVnH8he0XfOAm/Mv1AQexUkyHbS3DmjZezd5ENa8Oxsi8VL7GMtWX4vZzzp7Nw
N2ghatmKBy7SRoFaja/yMSIvxLhVwRBfv0OeA46j+sP9Xx/wN6mIGfAtS+aIebu7vILTZ6AES2es
uCGabUvY+c4EK3XtS109rN/bDkQcIBYF/4GBUGfIuaHEDLXnWkeaVYc9WRKsqz1Lz+1ZAiefI1WE
nN7sXC3+vC6mqMVBCr+obksJm+mG7vvkBqRhwEWaTBeQ9v8sMvtKC6O4QZ5LlNfbbVhpK6anTSYL
BHV3vvQDR4f/b4zjtqv24wTIFOPwgUQXhRfO2Srif/Voqz2E3UdxNtbtbOi8Xm2Vbtv82OgDEwCV
gjl4q0P4Jli+859dJz3CYtDEMB4VQeqnIi/PdNUyGEhAMCrfX00s6CwJ/Lv6pH94kpVTDo4E6W5c
wnk4yk6w270yWxNYg+UTGocL7u9QM7jvLTBIyAZgeasN8h1QJaXMek17pY8/6q97roxPAGD3DZN2
JCcR3r2GVCpKtKEnm3LUs/MWkV87s5piEnh31kUbLXXBCZdxv+H5DxAyDi1V2VP7xvn6Zkqnfqx7
ABWXqpmTAHtbFXcMIHgmYhC2ijJYsUAvsnJSH3K+7CtWe1M+jHMVm8xNnQ11jccxTcTGnrHDjlPY
OGJ7RW9F+XkNh/rzNAp77XThw+MPd3sIWTg5NZIk8sHpXl/xuOWldB7hetp2IMuA2+6vkvTylhZW
lu3SB456Naxs3Sc4wZRLPHRQgYVnmgwHMVzHB7C/+GP3vq7a5GbaHUASHovBYKTfV87Aj30GQbDi
3rHaA267v3jJECLiJWdonBrblqNRnZQ/pcZ5c1ZrLlRYNGOCWZFFb4BqIIoedjNQBiXgyRaq8gR4
jNGa/m5x4rBZNwJ7UrRl9u4LxhObLwos/cNMPeIOo+qBDBDMvXSQ/iAw8QG5JenMpMHE6huAM/d5
VBfMaw+sbQlzyzM3nM6RO/cf7tcNdj48iCJrxfdiC95xd0Z2kDU6XqEv6sibZY9op8Z06HoS+wIS
NSgUcC0S9W9bU0Wb9WJsPUw6iXf5tFhln58R9fFFynomHq4hOBCHjQRK2c0yqEPQpRzaORz/dgnK
vnUqLn5kkIN8Dd/YIkXvijg/g/h+JbyqW/smoozAEz225oC5R/lCxtmoKtnFgLyf04965Yavom+x
39I85hwFijoSRWOl9fDL5xDJ4CDXG2qB4SOgrVbhh6D8TYVBFSJk9tqs1Q3Ob/PbEySHAL658RoZ
Mo8rnUkguRtNde4FJ2VnykIGNe87dxlFoeftSosAOeFnsdctE/ShIqvWokBvNsZ83zN9CmP2MSiO
ApFsIjTI0qWGLOk+3JHydYBVbtnI/nusY37Kjjn9Ly78cQyfAYhu9ZOgWolPky4rTLJGnGE5kuO7
PrZdwSEVZ+fp/a7/42czY2kTqKJmlWOSM70CKWWlgUnv9W6UEfZeaClAScJqJTgtFGRa9ynKUarS
IXjPldC7XKmTkeVEeJoSvSv0X2LJRicjQZbmieJ2iudmRGD9g68g5RQXUJkWzl6PXZcw/idjYOYX
MJqlZg+ZSXYSU8PxmBkC68PyR7Amk4TVZMxXkfX3UUdYfxImQHysFhbViHOVVQo0LoPRwloe6K0o
07lyIGktaKBgskcYh3jjSK3MK1l52OxayNiH5nhD7tT2CBRCwR7R1Yj+nfLz1tN4U91QKtcrs6tC
o1Y0BXgvVcgzabh1mdkdanCKMNUOIk50Ia43dUeP86JTyiG4qwonGnT4bW4eVX55l7WsHObRDL1R
eC2ZTFu3uSqyI5/TUk54e44yzpXcrAnPbfPP4pHYs4s2KaBqPcqeb2f3SgcQ+4bpun8sx4ouqEsT
fx+tsZZ9jfXXwNZRbYzOHNmQcWFDTBfOpNFSAAaSoOY+KKMLlAqb/j/N5gdqqFwJKPEXHI0bbriv
+lUcOG1LPEPxCC3nATBfYOaLY1TFy4kllHP/qlvnRyyccjFSrAntIhU/y6b99hbR+FEfmyDpdG3E
2INhPXPbiXYwGMZC6tZ05YXllYJTG48/7jg0Bx5QUUDq+blPoxvIqyuIu+Z9qVsmVZMnRvg8dj3x
XPNqmaXvzGzSr1h25AsOjOJgD5E4MOzSNlxl5lIvEzvYYBeVxChsEDsGupfBY1IygGgFZvD2b1xy
tCcFYrdClQXi2oJcvefRpS38gSEknK2nfLzzb/2uMeDw5i/kIJ+k/wN9WIJs9VauRZS47eGYtbPl
+cXdqMVrppc4ITvjN0KGOfCJc5ToGohIh0VgDYKqAkHXLlfob5jpuXzOfSHNUbcFaob33FWhjtdC
nQdGs3uODiN4YblndI0msylrhGKng3qtEUGAlcl6s2tZSk8G9bZFg4ietAtVIO/zJyknFLvWK5J9
NgD33NXR6WPcDUy/hbzVcs5fbu0MZWgZyQW4/EgpyMH7Ao3lxygm3ziMKzdPG4qQHNi10Rnj6R1D
PdUsbmrW669G/C5IkDEYxofXtePyff1JVqsNDkBGYnvOo/JYPEilE1kgJKx792dSaB/r5AonVu86
hI4wAvzFKCz2uSnu33T20vskFlA6im83UnUz2FC9KRqbSGhnzBNQG/uW8BeuNHwn6qF/BVa0t8Ur
AdR8b8RYLaK4ueiCoPwYgP1OWnyatDj4R+fnIOcy116NGpEzZFfMwZtbujZaXdPMDIEhhvxuVWcd
QSb5yF6m5o1FOnl/WVaj3mKkbkZzny4UdOTQkMfVkJSNGwWMJ8rhV1MJth55pt1tj6k+NrINkUs6
tgj9qKpwTY6vUD/BACqu+bBP54+ViCEmWXhB3vwRikAYFBbOlvhmvudOsBOlBTmqK0T/uk6wAqyv
AUe1FXlq1+ZTjbNlvNdJ3Q+2txxkwB4bD9H7l7SuPUIiQIii8saxIN1Ur+XevNBBxBkJ1khYA0cG
mC4FIk5HProgkE0t7oXgqEOsBqBZeKCTqCkHHY9ys+/q+gaTodyvvqgK/Lpg9Dtk661ObBo1knBn
rTw1rWoXc6t/9tHB0jjvKitIE77g8SBuLgoV9IASF03HodnHF39WPyrcN8QbLBp/ArmBOViqfoRN
YQIxOts71KXRQ76SsmDlj/lEpcVHTuSgEf7F/dDSiH3SEvJ+BdtiztYEkLUN2WKGMLbWF3JqLEoM
O5uPtT+zX1xfuv3Q2TU0cs5Put81cnoE7fb0mWLQ6SlRNYqV3BKGv1d5ag1WE5XWH3bGetDpGZkm
gHdoVLwGLPdAjBv0fZsBnHNIhl1War/fO1LpBH9A4bUptgpmpcDbrhTE970JCI3ynzsw5+Ncdtur
Y/9tteApl2WzEX7HYBuVi87rpOeiNNApsA3KDOhsdb4DGG3mPb+I48rlfR418ZHxB/u7iarJgk2T
PfIo7DAW8sTLYcIrI3hsYp8nKDvCePqFqNS+mQ6mTVsAKaoWQkEf120uzERslRsbV9uYI44ocQfm
VfGzDdbTwyjIbEUCDOEtlSc3Syy7FISsaQjOXnmurBHKy6WisgoV//7a4ImhMJiQ11Xc2f4BQIZh
dfJpGoZbRPsD15LCuBQ3FbvMkeec8tifXDevF8j7kasPvAlTeuq3mZdWbi+aIxZY4toNkQNvkAYk
5RPTbq7YLwdye0T+/wGSwrUzxid6xTGTbeJEflSoS44qVlPSKkOc8WGIdceercIwyulW6Gx4bLRA
8LPrSxLAaWWiQ/Sz9trcmCOyMs7BxQleJHbSQQXqYWtEWwUYvuKeGJcxFbkO5fucCNdow4fHvxsT
tjvJTEN7EaxzeNLknc1usQhfrnb7J4w9Bp/nY0r2faBDiYQWvmMSbSx13MUUNHfdzkv2HP9s4CZM
+TM/4RFJXWEweQoD6Jf6BTjA+0wPwPzhNYuKgh0OyI5MOb1A7NmxSgeZ5/94IrHMmAuHSvY7qPWJ
QXpEtNVQiZWQ/muSafH8CXv0MRme8CLRdkHzhDpkWBYY6akUQ+CT28m2KPVqHn2ywM4pSw3KDQCD
KEfPtuRliu7X9HZfWkC7/8go21dzsjbyVZpk5awhcQdgloV9K9v6ep6eI6zVgjNnPkYZGCLopBf3
Sxu9jERywdc4lalQeIRpFlLO76YwyMi12mKuNse+z75qVh74knUqxYaeUrlQEHHHYJ/+AVUl3Dsi
gZBta4AvyJXWofi25lB5ndPSd3M0FWp1AQzOKZkWTHCc+uZ18AF0U6SSkgIeGr7dtKfPYFI5hICS
2kkx35LdjsoqlorM0P/3mo1TIApJhn93msr+0Fub77Nc9xgfg3kcMFX3fzYQj2e0StvWxf0mbjxH
QBnMMpBGyNFJV+BX9sWL3p/+aYK1fI+jFCBaYjCRq1RvIiS7NvzoKiLGOYYcv9yvZDn4OIyETMSt
Kah304WOHqVD8xMrtPQ1x6D+gaJngYV1x+kPZ18nH3baAVlbKuxo1BIE8OTwTXgVVKWN7EB3j/Xs
OuQxVnRur0S28wBPgLlFoQFwzxImn1F8dPTAP9x2g2StnHMO6dH1omWlOgZw+4aySVEQc5O2uBzR
FbBfSYQ8IWJYZws66cqriWbLpjb9e3bF5tDPArG+IGdtvCgl3WEWRLIoosIeoBLcKql9FNXk4k04
uZbdRjmoyiSg4cfXSQ0ReN0SnXY+aEm2/U8AVCq16ualAWlh1Aiq9sNFZhDoevsTjnPI7x9YO7Gi
1N4ObVVqYVSgA0XfdvEESCw6b0848R3m8PJrwcdM+fXsWl2qfH01IdThk6E/wvvhs4wZ95nMq1Rr
DDm2U8ONNLxGAcq0183baFCyyIHBQglsYgTwFV2S684v/3IILpzzFeC1kzVsJXbOAqDpQzDS5rpp
0stNPIs3WJGXb33EJFhAj3UKgXGIK77jC3DljH2n+Cwbrq0sRUOoS3f229phe6HRgCmOsifQAvVN
33NulOttoNX8cw/XUep/N28ebcGoj+E1sUvXd/L8nZIJLUQ6SRQhDpcYQmzdm4Xnt6O2V9FYOdJ1
oxzLr32VnDWMzBvUCNTfGmKcZcKmGGZPr6V7v55LJ2X2RrzdYDeIat0ViE7wbPuK+HcP9d2lY9ba
V5H8KP5arsjfx3ub6/ZU3r9qLszrf1SK50OiYKgx/PjMfo0hk0te5yb7YKvk8fspaAhhogH9V1rd
ggpPG8QHvv/dGRNi6A2qb4HumfRHEhxomkweQ8MQcWjIXTmrNgG0TMwZFNTjGBOGL8fln+nWRVIB
IRLru/qOxB4Wc61jtcFjvKystxRu/9hNRFco8b+IjWxqc+lE+8HpWWrVb32g8C1LBYVl+N+8xNUY
94xD2w7kybb+6w3N2mMz7INLYvzz18nsTONBYAKtRUq/dDNmgejKiGU2vNiFu4tRxe+Fm37p2XJ0
NXHK/XMIL8n2JaEPp0XyqlgkfK9ivg6fIG96070vDmxUrp5EKGoZA+cRuU0PyM9R3vd9+kJCuyvu
2eAPAngCi1dNbGbjPvbT0EkyADlWbT+2j3rQfMBvozjpuDh5NrpuFWHPOE3gB19RAV2A8Isbg8ST
z8ENvYNZxrVc/OCQZIzaPqZb8EWB66bxOMFAfK5gD+oiTLpdOYwjTwbAv6M/wfNROzit6zXy38LN
tDe+jmzK7PdiFh6B0rgBiQLo5GXR/namtke7FGIPZV3hJkn8XQcJSHFcUTQSIwdPFMzDMaQcSwiW
t6Fa/cBizb92i98sonib1BjpdzVu/64ZeXnWrEVwrXrHXyZmpKZ95xqYMiNTLIzO4/hwCR+MVBo6
l7EZ5Inhb5/TnMIhZm5iNc+doMCf8hcpAPawdZfe1HH/m8FDN7fI2muKdoOeaEQ3vLaMefiog9TJ
uW4M4wRR543hZymFis5Vmt4o7vMe0lGnL4ODCRls7hEOOG5ql1EwBFfLk1cG6Xo0poqrQNfmj1SX
Ga5quMsVAgQ6S567PtK5Z/IhfwYEl2IupTxnRfCftfd6zNKw0PfXoYMQR+3DYzer2aPc+tL73YfV
wXVnb5GTIvHZ18P23F11rUlTAlkeL9+OsbSaxmaDuYkTzeuddqXcgp2QJkVX2pqjwSJkjQb93Y2x
l4bdYEhDgvZ0raIDfdInUUXbtKpAKgMz4j/IohHTZY2u0naAFqxqEOufkW1bAEZZr78GGBCzAVbu
/yDi0s3FrQNWO5ZRoRSL5DPPsjMIofWPrHlXjMQiZVWfy2n4fXps2+xW3MWyJYs+GtMnFlSN6B4f
vzaJr34/YNXQPv7G/Fb3RE0VHc8fsbtZow5aswJrjkSYeCFCWNLqUL4H1cVFnPx4xlbW1dOSZnES
vtKb0MTcN4eAiLEy+Eznzc1gu7htvwOOs/iQGrVNuiugSKolUSNbp7C7ecyBzmy4tIPPsrVp3q+L
5Ss/H1B/X+kFVoxX0gKeGqhI0WtCQpxzLLtjasAPNmJr2ziGMAgX732laeANEUT2OHh6T/42gR19
89+K/F2xPmR2RUOKfKoZgNDarl6NUSO3377DqfVHsx6Jv6WJ6zyH69F1WbC9yZc+J4Ti6J0qnNE3
Nyty0HzDkTfI+ZH+2R2Tc8xOat7TpjH4lk+tPWl82RVHd8Q/UJ7qyRojXpNQFPxuOIeXhfhwgN8d
LevcdWIijLOLYTUlJJhCDgARH+GfXY8ekQVR/MFOKXQTw2PSu9L5GkRb5+RRRc//Xx2kWc0JENf4
2vgZZ/W6aZxEAR1rRKzfEHb24M3OmYmFlg3pO+72OYBBHtfea3hOU/NIQ5DE5Wq1k0OXwqDCtG1D
b829yBy1H8KvL0+NGO0UX09fRgDug7eRen2K1GmuXo0/+uArgdaels+AdkvuPuaUqOIOvUPvRNFD
mm7nY4JSTWf+52r/FJzdeUAV/ToFqJDli2ONxkq3d2VMN9UNjdp8Dmzvl8YDtpUcBcLaPT+36sj6
/aL6QukstT9hZHx5ykLbCdF5ZCnkLAGyuZ187qfepPxJ0gNr7ck7X57LXb5Sq/ssiDqAHrx3bsuR
74RcPF80FPoe1J6QHRfbknrFiVyi4xu5O91O2mxFuPTtSsLGIHi7J2E55+hhVuNCfOJREtuh4t9B
YCA49b2TVjTTSjPENOSuj6km6LbYeEW0Nh3heUjtaZOjCH+IPbFpfbC1bwTtKSkgvDeUUUg/o0NE
1GWWzxoERxkd2XaK1gVs7D58YKJpv287FvrqfmAsIWvbC1KNCLleJCz0ot4hNNcWTrEkQkI80I8i
WqaWJFIuHofrol3NieTrOepWrs4HfWGJbS5ZgBQY7J4qiCRNMRsA6CXWE+QUAcH2oEq5fl5RuEi+
cPeuo35u5AQVceBelnS15QZKvXCiOh9vEbFafJBzNDloJiguyk5rGruI1qGJNFpYf/IAdOAYv0kv
OuUj4sSXC7uGbEPt6qI7zQ1AoU5OoZAp0A/OipUrUGjoKI8nir/GbHyD3qFDJp3UUWmXB8Puv+Lg
xdb3lHFeQzFB9ZclOojTndlGdl3dcVF6BR/6aNxEXtLY+kMSKawRFmRY0TWv8l7uTERh1ictyl+Z
NZZ7sgTImCC4s1V7zuiZroWQwe28dq2JguDmdDfbdiund+JfrUh0G154721ooTIIvwi97LvVJUA0
jNmzaPq44LiOyJZqtvZmXC+fw/z8dDJXUt8J9+r7leedcqpRcYr5inKMBKRpQ9TjXg1eXcxTX0En
nylP5r247blylaFWO3/zeHmyeKM94Dc5syQWFdAQs63nnFSrv6PWW5A93L8BcedQ/g1bMMEZuQuk
UmzFZbKRxMXoZz+rC558ngtcaZUUsBPm0FdWPnC9YGUPKrNsAtPUKN2a/lAzj2Rri0/ki7ckY/Kh
9jYdqK3B/omtg7GWiMhu+vuv46BtE7ciahlQTx0fii31bX+QA82Nhkp0OSxtLMFqrPKXv6zDUkjR
ju78YrA87/2tlaR98+MCCcKQ+UJEsH1quyMkqfGDbF3HXtyy0dDRZjEcIwJOBKqpiAYyUgU5xJpy
ACflSSZyDLQJJFL7N9p0BPnEVdcZuaOnUL+/E6Kq4JjtILVptesb3Wm4IY1hohJy6Cb9JZaZ8tJZ
YIzfzaZHajPIOEcckC2Oo0sYtHoqc09PeEPZctp4dvbB6wmAQ3V4QYfIsFhlIdnEP8cbU5SXPe5b
w/q9SKw+Cm6DwRGAXXfXjX79sGCpwbZvaPMd7PTcSfAvkuK+hf4vXm6V2GNtf6hkLJbyMsjUHqFZ
vaPP8yK4g1iaisDvZZl9owsP9sJdsQuG5Vft7ua5rZHFK3Kdy7AG1aQw756ZM9GNHLprNE0LWQiF
cgmgwCmLjWvT1PR6OEux3sHdrmHDUiRLWyGRVO3PHWDHEdf/wtc9p9xv73P9PWGuQjlB+DYDD/EX
P02Uqbcfj/aK+x7p/1dDSmuRu84lpV9kNsz9rRJULQOvOfpUYN7Oc+0dEK/6zTzhCJvq8EYf9ubA
DWrfDGkqqFx4l6V/D7l1Pi41FUAt0vFXFUWblHU89nHg38yVphVUFN6jSXeJC3K16brvp6OPIVDn
g95nbBUb9j48dSqZ5KzWTL/PZw/psB/g+P3/woNZ6aVK+2+YL4XvVzoaaC4HKO2Lcr6Tys6CpxcN
VvPTK5ulOmAhSQG7eUR6aRH5EMzldIulKjLf8nlLr+KqUzp4aPVDpEc/MaNz2MGqK/7jt0FyEpcM
xVAzvTZnDYyKMEeQPSYxr27c+9gTe5zP0RTzm/23HhRyVZ8C51tUGL+kJQAMEqVkkRmyuLQXsvd8
9Z/UABxL48SqAuy/1A6Cu2+9JzwiZvK6Mlp7ERFKE+VAHjJ8e08KzC7OZgfhkbhLHh46CFj2RxXV
S3r9NjyYzyZRsMJVP824si3Xxq5CgdYgPn6DXaxT/uIx7m9P2imyKraNOFdgj/NwORbzTYPDorFz
TouikmGyqGqT0pvrAa7IEtERMqyc/JOdhp29rFbJiGABIrb84L25E8KB84f9H3dSbgaMAzJsBoXs
xxW62GpX1U77Vntvk2W7kt6DsXee2XOamTWLS+2DJZ10ulBRjPX4hm+VhJ4x1ulOQ8/V3kT6PrDp
rnNDeKj7ZNRQ9WUPuctnZJ+0gC7b9PM1Xsc76rd700We+zFe1+r/DZCcxE1iT5F2dLqVJcYFyGio
bnUSsVikED7IvYDpu5EW+TmTALE8K2k74WAZky1FtW0Ulk34MyMw0r2ddEvlbCIFkADsm6V1eGet
/R+V6ekJef+C61TwEON3OkmGaU9l6pxmaBdXD2smttnnWXwMfg9QOoow1HixnzYpnttdIKwBxhR+
vkjBY8VIC8UE/DPjS2v1CT2TSd3f3OzhdSO7ukjWOJkLsp93k9vri+b1N+svqSMwa0FhUwmyQTrR
3md6ApoOi3JCI5l5do2jG7t2AD9J8p1avEYyydzkWuAlM4Txk3TKTgQdRLUDpv2RZLExW1+MxmNr
AQKPYJOzs74WG70HXPbEhgrtA1TxlPIvQ9BP6h6RRwNva4CBmgRaDYcCy4kUtrlxzgwJQTE0bRoK
7Pbjl1Nb24VjFtjFHRd0zxe26jwVNj5KmGvEfQwe4251MVegTj2nNHtyUbkXlQcQoe1950ksKrbL
sSP73Cs84LGZ2cOXG+BCnyg7u41VThx6R9YytV8NSvUtza+U7nDTXXGwpcTIduL8k7mYpW3p5u7B
HUjCBzkv8eNrcBkjwLogyzFOGS+R+zKYTU0s9x8xZ4y8cgFjmwntZMR/h9OrZ5GmzJML5/IROWul
bYzBNqwQ3ExdF7wr96Yf9KiHXriTJwyAkrrc3nJd2vm75c4RJXGAs6m6imDgg1L3oRNX8HARgsno
Tn0amj1KW6YaZqH/kNYnL8eMQi7f/YrurfbQpXi5mvjrP2q2Eg+xpVr5BSycOUW4dXCn5SaDAdVP
xOSpgIDKiD0lh+7f1l6C1kG0lOVpcMGslzcfuHSsnRPL/wg9H+JCdtWWyil59uf78qq9JbZVv4bQ
2Eho4Tdv7N1ZOt86C6hvRs9fToctz7HM2uyRI9w3PJStwDpcwPoby11NatKMvIjDeEV5CyBL6Kxd
pzL6b7Nlk2ryoD5NVTJCnapiwYDOCnLgg4gT20ZUK/7qGK6rpncjEPG7gmAzFNsEoQ97sZQH7nA7
iEHUkWVblXcZlU5StlbIv5Socp2Hgpbz5GbJx/dCjYWtW+/WJH0wHXYgPxXTj3KXmnydkLaRih+9
tIqPIkCoIyXsA5qxL1ANOWaYrXuwPfbFUxgTFZGr66iMEk8ZXhScUoF87wLJGURBjrnqoq2VTWjE
bgSXtaX4mKMyIexS3ekyF3+NlkVQ2aQ5cK/PDPgImfMirtlISLtMPtWQ5aR1mJZV7tVaQ8Xc5TOC
cC+9ZY77kXc3RAdlZOaRCWWFSlOW7J7d+e8YeDRz/GtyynIraB2SknMGfbZS3BZUWZv3Edpd25f0
z8HxLAEPOpfnoJfiNI8lsngyowrOEk3nw3+LnJX4oMhOJOpvFVET9TMJ+bBXEVYRxeYs7YqBZTT4
qOve/3QNFDHXTTZIRFubO1+GslWwvSH/EtFmz9Nm5PvC0GbjgqPA3/OPQspgH67KVE6zH0FQ6Fjp
jJGIvm1vu3X+e/lWzvr120KhK5x+nYqB5clnbMD3HZxb3AxZ4rD/MPa3LfGlrJ2txyQu+HCj64v4
CJBIgs87cxWH28Q/xv3IEeSAPDuxxTx0whIPSUEmOj1uIqMf5txIsv8ziHn6o9qiKqBJcTYUowXV
O9Rg67obq4mDRIo6cmtYviejQCF7N1Zw88cfdtuG+4Agbc4b/V+M6H1R3Gg78Z3GNTpRD5eSrydf
U+TZZ0kz0sHaUVzVxolGTora2DCf/9jPJm3YT8AtKS3XefEuk54dpYnt0jf+VQIq/MxvIRtDlERb
58FBPpl8PCptUyN5ibf2HTdwxZxPqFZ8xuNZIEpKlHIZxZ4USCzULXvP3/eh+EZ4/WsV0WjO718+
t45c0s03My94U1zsF92NPmk7vafDsUPuNPGDWqXadVlTQHiSKazWKRZQouIEQBLU1xKtw//vBLpc
WIOIxzrPZ7LMXRCTJABI6Z3WMoXcvtU/MnW5BgiTB4yzcKzK1NYOKzfXujz04e4TzZRIyI2J59lr
b98nShxR1p1TIh9KBNRU8/VAjlcHFk5CRIeMx60SfbzCe1q9qOyeWjw/4V4HxP1/P+pVdzHRHtcL
qtIsc4sqPyNncaNpxpigPhRbCMoMMXEqsy0z10msUdIY1BU2SxBuZFbzNDBxXVfgb3Zbx0Bflh60
WQKzMBpH2juQqh8ecW6FMWO8QyzjfwgfDlu9DA165t6e8jZt4DbvdT5G5S8d11u0c6xosO3VkEh2
72Yb9Nn+GHEZw1cvNB9ysN0cI3NLU9xk56Lo0Y0NxFNr3qAnUTjzkPOcX28dPuMIJAQU2WwrbYEI
1RR9FRhVjh9N8V+CFOvN4ppp/9TMBB76JVkaixcdAPRAAr4zdg0TtdJHvWxo4KtVh9/R6uYrCDGt
YCM9HNC3/8vVjJ9Ad/khcbToTBnR45gD02rKtn1mUqUrjgEhybw0nbfnV05DxTiDooKxD+zFfLIS
KnM8pCQaL7szUq0qx0DXMHoR68tXfy9TnXSneOZmLcrPFUOKe+QOyKUdc0d/eSvOZ4BZhtzONdzW
eJgnPYy2+LKhP2HesBfpCY8tcH+9i5Pr3h6OnX60WoGMcI5oQBD7DtOBk2gWbXxlMTOhTQJyWOiV
uugF6Dmk8YalxQq09fV0p37h760owjzKdlYV77GBhBXUNryoMzBc/j3GmGMpng+oShVdJrx5kIaq
ckodqME818cEnNd1a92unQufbwfHfSGyB4isOrPD7Q+DnvQdXlH0Uoh4chW06ju6txt2lmHvQK03
kB9fXzrWyQtdSszUmO5k8Wds/gQoP6FS62zGu1FBhL1V4HTSBCqNY8J+3RNy2i5H/rnDZCp6Rgjj
POPsV5XbKzCXnwz/XVUYaQEXx+H4L8En+iWooxg9WkTqux6zHSw+Yir6xfBUlM9MaEbfQT5kHD6f
cnuAviFvbMx/TaK7pGNlof6cP9onYaYn14KXDMk9YFV0S+2f48NwMZ0f4YigSYcUw8wQJQoeKuLk
gxsR3T/SaQKqO6KM6i/aK98JYADaeUy1qEr8yLgtqhSpq0QapeoE3lUDE+qmx1F1HtwPtYGSukmV
ttqyzRD3G7VPamwUYYgoVtqTSWHHyHhEWM4MQ9UNbetCx2zY99pibuF3I/0ZurUCT8eWSI+HuiGW
LjYYXWRq0OYYkEaVmQAVZTwzRH0JIaVDnbwXgXLbBkPfTIvkt5KuiT/rLeE2rIziSPlSx2wRxhjX
EIBCsFM4CgK4DBbY7qP4tljiNATkzXkw2VHNH0sVViNNq8v2BajRRNf0QKX7tk36Hb1hQOXmUkm6
TXBCnbcXcmp9f/1UZaaR/Y8OrxuAngkIKSfJO+A6lQrl79bjyHlUJzbOLZHMfuiWTxXHiFduffGg
+krqVSrdB6a3L2SdAFtsS+DQEzPsn/teQ8MoW6Bp//4maLA3QUOWs1+kcoTBIgZGAzRHu3xfXK9H
Wg3b8nOroYmHOdgqRTFHSdIZfqyFXzUvwB5HFbDDHlb2sr/5p1hplgweCII9kyKNe9R8e4mddYWt
4OqJT2IHDAPOEjrzuerW6x1RN48s90jnEV3+rWNMSjbwCOOFqoBxkZ8qu91qwi4E3q79tLORnPl+
Fh3gjKg4kNzhkn96cCzt8ZInpiT92WdTwqHNhlBpzhxv1dA6PtzlJrIsGH4fy23DxKw/TMlqdtqp
tZ5PFzY5WAqCVVMDl+r+CdyhRm+yr2nIn+LB66CxHu5ZkJUbqHa1/vr6JsvMSoqYZHtergI5iC4/
X6oPqSr7wJ0f7gDLRbZ77TNkLauevecZMEuSObYbJ/91NkowUjcRYsv6eHpfM7u5MUkOSFjNbYqT
Oo5ajdD/npXKvKMD/OnU+y7Z0QwoYkTMJusob1AT/vyrwLiQesoTLsq7RekJGd/EXu1BgLB1Fs26
AcpkEgaWn9Sch8slyGeae1xhDp1ZkP+y3EC4fYJbNbH/cbS0+sBG4wEaT9XU0SH8kFomzsX1DsNz
+3tSdTMD6W8zZQV8KYcoVvtzfQKzWPKmAHCxjXGFU8Cx4Tc1pOtKVf937M83LPIAH04aH74+bYUc
gVTImGUXtjgI7Dzb2BfyBdwAl5bV90V64/0LkEAWNG8M+b/1yYcoZp29BwYaugAwof0XPX+WrVnr
yB9MsCOZ1TaltJ2dv8y3WofzzrY6cPBaJvzxmSWarXreT3BorwS1btQze89XOVeHxdYuM8l2qL1I
LmtQ/Cc0Eh+QNrm+RcTgOu8uSrR1YHzvIU48YNjEdbfNAnd5b3Z17pFdS12YabmE8uLj2j8FMM9Q
1lfMHPGR5wKWM2bpipenvWxPUUKYSloEoJ95v5aeQpaLEEdQQFSqxTt8KJUicGLXEUyMe9DCXIUK
hZkrrV+k9t5O7FQAqDiCWveEfTW0t+3M3YzaT2X2bkN9YSSEKHHlT1J7X13ntijtHkF8ENwCVl8F
S7stXnkl7bFmKu39VdbIgah8niDRBfLCqvyxpJA8D2lRYroCx+EYtdY0ITZd9Iidoz6gcKQKNXCI
+JxYVM9MOHD+IuwB/L2nZmj3uX+tYlacp9O5SR5ykbaNWdpmtiu8vGc2Yvm5VHCEKewPE+19A3Um
Jmz7p9SQpTWfQUbhkkDq8oD2BQEmRNoqyVZelSAakwdKqjN9oNlBmqp9/9/4GpzH9PVGkVcYIHp8
dlA5qPMQ16/3BXTOQg9+8rt5GELjmzrDIsuo9DUEaC+9usN+AtNx5WzbfC0iIhRcAK98I592gdZH
muPSDPRJKhFQqp3glhemJWPA9hujFwTWoIhh0NiVh3r1GqFFMVhOUxHrC2CTB/WkBZEQozHDjVsW
Q7ROHIWpD9qdHzrxdUAS1+ity+5RKHM0AFu78VTXqefJ+66pS17NjxnDnVozRmgEHt/ChSdisrr8
fjCU+RA/x+AW4qI6B0ABrHLpPaCs+RQBHFi4Bc9dnKvOTatcln/lgb6dI1iGZ5VG7oT6E+l5K5eX
caOy+8pEIzzIjxtvpUDM0gkEgJW1sPhKjl3mbzeCB3+IDstzK88wyF++IdNg/30MPBCQVlZu+iwc
T07VUr3+mULyTgo9NG5hbejvxZX5/2nfD1Meu566N3FUew05598x3BTJiX5nbfF+FiBOGoVPFkAA
SD7KXpIX0cPrK7d7VIHoX2Pc5KxHKK4slYk8m2UoXLsGCLX5D+L92IIE544cRhazVZ1UzQ+nDj2W
2Y/AvYNM6r7Ms1j6daIMemh7RWJB+CGUjdJJvFVjhJ7Vp3wupGewoU+QipVLPGTTXasEOlnSBtLF
9W5x91H6zfHdLvodFddCMOKO1Cshi3WPmr8bbPcGo677Co2Fd9/s7cJVXQbnfFCRgOYCugOkg86/
TdmYqaRhdxMrbdSGhg2urIj5aY22wuuqLkfUcKrjV1iZ5g+QJ3726EmxB2cB6vPfNWWHSGj5SJ4V
4VJ5KLylXYNSzKfpFWYvuCjVcEkqJcbVcwFEo6dRw8IE8kqbcJPs9j7gewg5Zy1BRTfvMeiJzDZl
zX2vZZUwu+EWXnjgBap4BXGoqrqfLJS8yG0oLqnzjiEJRE5Q1Cfvb8xEG50VV1QP0cm0fxzOdDVW
KEk/mpnBtE3bHfGrx0URua5ga8BxLJXPnIuLIyBNTgRiXPEK6TTF0wNOV+Ura2GfY4eQRyrIiz85
PW5Mf5h7LNFT9gTCyMnnNvlAIkpDW05OYgskpSKyZv82iBuRiayOY/g4K9f1704YUrSQjb7SqQ7K
jgzXz6RIv8/PMYBt6llg2Xupvq1dbLR/Loz5FvIHhuw0LDMgW4uw6aR3kp7dYuSkgNEiHs5l+GZl
buDpOOOZ2Z1J91thFqroc8b8IgokOtd1PlV4L08Ag8s0MzlZyGzCkeEYORd2weFnwYWys2YNCKub
XjvTSQgCBjoizR+MHTFhBfRQyt6+UAWh4zXz4OoyUqkOpzHlnzCxMlM2vyd1kMDofyUGLZOgAFv3
4wWVcRc1V4D19tIo/PjkuYYf3CxXkSKFWIlNgBuGjyq3FVETcsoXws00iXtxB6g7VI6cZ+ITQo+u
CRWvLPnCs+eAJJtLyA/keFd7MLgUR7ELN19fSt0LWFSjso9BVtrFqGzhHaOiwvZM0ziG7pd2d2Zj
icCeoZEtyYCne9roluqPufqyA7tAclwPDVTTrdPeh+K8yjJn7zoKxRKRy02mIGfR2IJcg/N0NECa
in/gFxCsALbXO/wsP7VTFiuhzGvULZ4UwYi9T+AIYXyYlhorxEkcagFvM7GzeXYvj8F1SOAQ3qma
CJhD4jn0TD92VOHNlGPV2PwjBgVNbcVN8Hl2GRPXv/lmDqxZVxO9npDVriGOQeBg6sVG5YhXkJa4
g8uaH/VtFgDA9OXrsaoxak0clk21MWv/MjGcyLlEmaNP4YGsXWoXVwFiDp05zpSon9gdQ1q4JDo5
DJEG5PEwg1zkN0CS9bqXCW1FANtYHcfL22DkpzwnLnc+MicSCgo9QjZolKQnWFWPTICOyW+1YoCV
EdZLrSn9JU8vf/Yns9BRjbII0LemwptAo9BVMDumzP/OnLCGSzq8GfwaYnZKlRj0+XUa01RZVkOG
ntWz5icvwNZKbza9Pnc6cTVPnenwWrnk3Q==
`protect end_protected
