-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
g5EMx86vS7RFgKy8YmKsXALTZ0foofnNMSzRDhhsDl1Rslg1JV/4pp74aJkNWEgtPuXcLac+cW6s
oz0i4/EEq1BZBZrSOa7s91LthngtDzHsfnv/QfEB7zblqatZrdrkGNgHkCWDlWM4owGFH7Vxloov
rA32Ru9S2DJ/xfpPK91Sx6rgNNC+ohEa5Ln31/bGNqovZQaL1uwz58PWCC2eraXhPIgXkZVMtpzz
acvrFnQU8jkAE2YLNpOjncbWkIYio4wxvwEWKbKQrkmCkCYVj7r0XKW1+vsF3SeikLrbW7WKKc8T
LsJpQ7FZPkJwqRLYbwvyx0NvXFh7IcHNjg7hMg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
MjQ2fR67XN/pD3eZsWV1Ly7iOdrqI9HuUkObsJMg3ld8EI9ztuzjm5YYM857z6PP/dq47dLd8jWf
92bLr6e2gBXpRjH+QBKss9yVAArxW6K2xVrc6u4BFPQhb5zI3yFO2/W1lz2YlgYUCfvgVQLRM+D1
a7ysZK4aPX+b6J71wTa5FTqEBZcBnezIa+6BpcIKnohFKIeuQVuqGBSPGgLTQciqFanGgMHcXOWt
X0kpIf4hsyVVQJERPMXAypPMH66U+XimGLWru3F2/EHG+QP4cwwVGS2MPUKKXdSxDY65vY329LW7
c10MjFmvXnR0DfLkHmisJan6NlE7AH88N/EVLgTVI33KPOHjKxay1B4OCvnSjtAZEdzNNGDwfa3J
kpdLarCmFPGKD+TeOMGtYS1NMDMsrHck29/vHYuVrFVUCXoweJ4/qkYiviCndtQ3S1AaeNvh58QT
jsVmANQqhLfGO8q34MZB8TgtzBswF5L8Hwb9T0ChPFr2Usj85DzYrDlAdDWkDVmwG28KReA1ajwG
3eU1u3ud66NNKfzTtAERsGExkmAWbjeD1mN3nuIHSs046jkzYOzpfEViCvfWLZYBfsbbeeiPYRKw
IgEGPgn8/aTvpYZTtB3sYoWmka5dXGTcOgKGopAVi0x5CWEXF/nhyQvmeDYQ5Gps6sB5bBJlp8Zq
wtjxICKB53E+O8avgim8YHuiJG/xeW1En/GG/G7Dbx9dJLDtJPSYoCC5kdV4lbeqIyYCbrXlGpkD
o2UktBBhpGEt1QK0wXsNUD1vp95tgH1gbveDCfmw3CbnPJeSnqoic24rpJQZvvVNkwJ06Xh7DzzS
728EjrRxYUsbmrF5MJke+JRKpGpVeF7BFSIZ1VElsQPSByjE8D2vXsz385SY9JdCKLMWHyVKSKZO
4rjPknO+5ZCVMmDIK5cI0PUsJDk1nHHoY/hun3sTZ7PXV98Drq5kROmyVuf5zjyAmTTRJJwE+T72
J8kBUMA5tuWg4MF6+pwdYZJCBs8tnoMVtjNGZ5xISOJvBOZ0YPnevsCfW3a2Jslc0RH0omM9sVai
B/MfE/ssnpmf2whgDgMw1V8R9eXxab9fDFhQVRNULhVHomwGWWnYIL6GQUoXxoh/N0CEwVaACMGU
IN+m/505wFh3NvRjLOTqZYdMdz2dunDF2W+jYyGQ+fBGn5fCpwICP+ecZ0EM8e4SCF3z1zDaZTcv
2iSOzuwXKTJSgOcWAQFdLtdm0KyEjRX2VSWKPOPx2oIt6P5tOxXh67TIbWtwu8AmCzBUCf5bv45P
9/K6AZXf6W0pS20CesfHcGo5v/ThD/dbbVoY5rCMRTdgCUrI98pTulwh49SGyEqARc7AO1RFuwCt
Drv2ESRLjZMwlwgx8TUwnCE6pRi0DXwIjcsNVvaSLC4O4H7KcHhrxiVSUuCE5WO90qpFgVljto61
eR61Hwyz4y8eS5o8f5S54Cxphn1K0jZVL+Sx0OGeDIwIX2TwGZK3X7jMvyzwuZSxD55B+mJxSTmr
BuftoDmSRRhHZqZWD+KBhIWqQMNW2oC0J20euLsx84AZFzKzzU4LBUXJPyeOxIFM26rMAtLnCVJP
fhL6036T43oEN3HAxFU59COcAhvYQzm073r30Sb530TFuRJvaWBDKHvnaaoSM8jkzVW9tYIAh7A8
svA0b5cnuetCLb7gQwsiojM8W/oyzRJIJa96UCVZCdjIjvYE1XZFSlxpZJnLdo3x4CYUaHv9yh5s
v/0Fuid1tETMKvbctj87tPdpVfgdoHCEdFwnpi2ZWN2bFp1xmilZCTIX/fBA6vKZpF1na47oUZP+
5Te7F4pjHVfeRsBN64Wnr5e1Nobo76fj/EQoqrfAB1MWcYCAiCUfHTjgXzB74r8tPw3nHhkggEJD
4Lj/mYpa0/jT1JoFo0WGdTZfeGhQEH+8Lc9yEqREDq26PZZH08xQVB9dIUTPwBNFKbdia4YRSKO+
qshHwYFN8Qn8ApfF51J5lfH5XYpUj/dJPwZy1bY8xUIxEd8OZkXkQgVqtvegdxehAvtebCd1DZE7
Kny7kh3nxEdYp+u21WwksQ8yzc2jb0FSJMOTghY68LWO4iu3UYjEm1wHPnH9RMYb92uC1Jzol6gr
vnTFapcd+IgNBxTk5Q6Z2n4vzbUYTxQ75CWzdK3aW1xolmIJLWXYFdX6v06+MuhJfRZTQ9CGpJ1V
G7YwdusD+NyHgDAsoGPLJ7QN3HrB/r/IhIi4kIVyjvwa9ZUudr59PKtiVCNUWWi+1uCdqwpBEjpG
ioeNRQD8po8m+kJQQ0NRtTlaptmkTCwWl0I6czJD4c+fF3HKwUPL8MBx2medt/Uy5O8m9eChJrNw
7WpPEvfLajLBw0GSy/4JEiqvxmgEqmXbOebnuC/nBvq0zF2Ba5lwViFpHKcNNDilw1X/y3tOBRAV
tE8SnCA3aXRXBL01tYUiGS2wogTKV29lDnsofBmTXCZFQyDJ4Nx/zVknBNBNJRXHEDS+Irnn6Q0H
bJZLvk5+ozRC+ARG56fR1AEsJoPuqd9PET7D0ic4fZuAWCZQJJ0+KdXTv2GcGky4dYRFRhm3qroY
5tqvHJ1grQ30a/hA2ODG445ntTyNNJd992krXrVnSQfWfRkbFsuB4HKBkEQbINhbRgu8SPSXN3Bl
UAbUTkdOhoIoPcvR+D/q/9q65/n9GVTt9kVFDCNAUYciE8HZWns6kkZeL5ed+CkMV7rgiLWEwtAS
pd83fdUGeQo9S8J0GHeO/5kUSKm2Yhl7/toXNfG0PNCbTIDLlipfJhWmn2TxOylWPWbKL7+ha06V
CiB2tr9VXbfMVaABMjOqxpgdSbZdaB96vH4HxxzP5PsdEhKwOWj90I0lYGpf+0uLpBU5sSD6lvQi
+PcwTkRGryGEmIY9lAI5TqnTcM/mpAB40Jes/NyGiKAgrw6IcAnI0Vw6sAkKw/csibsZJuTOHS6T
OxBqZtRM64+lsD/kDZrsn8OyM7gUu4Z8B02dY5MqVZhgsXqXKe67Fha18FmbbL7nFEs8pwdi1NF4
4E45l9xM/apF+B/tZxHomBrVqgLsHgfwBasAG9DsNOwPPAyPYARInnHg3NGfKzTQe48z4Xh2yWOm
ejbFeSQ+DL/zzTPKs12PT0BU5CdWj18cmcLYs1KknFmt5FME7JtiHeQH+vtvqD6xT3BodIRUyFWR
ztOw408iFMcE4xjC9urdbZnd3Li4bsj+PxxFP9md5bY8HDDYi3Q4nNcJULaRYipej+t1M2UXp42g
iBz9FVnafHWshxB/s0aiOYQkxauCaZz+Bc6bh0aIDSaNYhL6aJpNM7mFohOmD8f3MVELUe6jaYUL
0HZ951FMXjLBlwY+bimc67lSj4u7wOH0c71Jv/DRdZzlJTiaQyUtRaUoEQj2rA/umi0eoKrixdZl
Ct7PyVhBQuKAt1g1tfYIpN+RmtKanLIuYrzsei4xzE8yrKnSj5DKAlN4UCjpoe84r2GGXL6ALdhO
mscHPKI01hkC4P4cf26JwK34rru+jvDdajbTrBIybZLvnCf2DRnV49JJlnrnVKj5xq2K6opPVRHs
MkkY5oqAN0BBUOmi4OSQFodgQQpPqxy4MVKj0NrM8SyXNbOrk9klwhQisHrGExcrzC4HWLs28PN0
PrVUXF4Fw4ADw64RyWNxBg2eK9bykzwjExAbO3tNIAjJWSb/MEgOOKvdSv2qkqOaZuCBbHi3AlOB
cSKIjL3i7dunIuY55XyzrDRgjtUJvNtK3/dwWSiG1s75zO9MiYKyN8aSHIOVFuMQSG5NDy5fJZrI
L8Yi1CKtgOaKsRvnCihlKVn8ZrRHrCEuV4sEO4A3Y6gcXxHJQoSEXXcXYhz8yCSMLCbXeMIg7RjN
ckBWnXAXHkK7eMZSsTrJk3TR+M254ydx494COPd2c5Bfc7dfvWozycnMtEvFznIaP8VQu98TJ0wK
N36DyqMz6P7Hm/39VuEeBgqkTdwBgsHJFs3vqKag+JVnCb0QMLEF2y/PSkUMcdbp8y3aWlwESTCT
/0wLKjLwH/XV/TjaPJaXmtlbkUaokq+9wArgcNJTWEpSVnaTuWetsA8+mEG+TFMM8eW/wki5N+dH
i2RHC7vJylQayguuTkbf0w9LrHjgkW7kkkwbNHIgRZNgzncuKxY92Q5zQKjSrmf4O7xlH7GV9aou
Ps5c/wgC7+I8XujrF3uUEdQLf8EC9k9zRuIeoxRzq4g1cKAbj3RxbklAi66psIMkhlmISbSIQ3Ty
m8xRCISpE/56QnPy2SC6an7UBouBmI5FdAlUEP+EBFn/2Jc8XhUk/Ee0gh3O19Zg4Qar686Qa4Bg
fTNxLu7P+qKrl4a5Xc4r4aolCPdI0PWCSdbZzgrMvVESPxCLiQot5i+z++BzjR8xYSQ4mvqpCeja
RG74m/UdQEKcTotYuUhDNLkXi+BbFlGw1fWllRVyo+Ce3UpOVV/d5GuQV4tPT+s23p2mrp3jQCph
6rnBxLjp40BSO8RvcaVfpf+t+Eud161wG6tS2ZgMelhas4susj6RiSQqGALSQT7ZeLboK5AUVAai
frqH7tvH5ZXujdn+0pgi8zTro4be8LbHGr2vU02IvxMwlgO1q7FEThn3mcJJaZWZyACBGvJ4wlZ3
/mj3/c+mMREmLqQOPWYN7p0+a8MU/GRugfF+5yPdlUSTGyigohA2CCFziBiQi5OA37O0n13f0LTV
zD7pwIIlmU2PD2Hn0kPhgLWz9FYl+InMlqroRRg39hNSqgtmnB9HCH03M6hnQ9yAd1gf7WUmpFg0
3JuHUawG3usqf/27zixxzQpJK7Gb3hfcmdfS8z9c7XbG6N4VLY18t572qYRp08woEQayfOMQhwvi
eJiacq3Iwpz2iSzDTSzRUh9/igA0MwULpoCYhcJnX47IuPGkCK4qdvfRCKHCPWNNei8Inh/Z3WGD
dC94Lt41hNfd5pBTVYDLC2rjrelLqrXbCbHMPZRKsJoB2JhvzZ+pt/Sim1krUgwIe+0eMeVUHn0G
GaGrHez0T+bzKKlUWBWcBwztZtC02x62G/BBH8XQeICqYucyz7ZiFbMXNu8q0kkgtgUopPphG30S
dU2j3gmhj57c4CBUf4MS5OXcUhmpvWmlw1jYWUkQwsUoOLdA6SzLfCBv+WyOr7nc7WauSexJV9y0
rxf3+1YMexOv4t4F19QNwdhwphB1skqflTi56OWCa2kX6gXiffMmSYLU3l1039fLh1Y5tOT+ldvJ
ePxb/4ZbXX7/RW8TyvqEfnYAQH9ewwQ9oZLVWYkvAWEWJBfeqSNmY+YzfzPqS3bhdZGeGw2WyiPd
HxuQRMH3Hx9ljAs3ZraG9yR3QCAsks2Pb5PZNSfTX2gAWWLnb3SnM4A7PNcRfT/MnrT8uImFQ5Ez
kfewbj4clQRFh7tQxi1UDzVV97Y2c59/ez1Pxitrf94JT1WahIh4Vf65tbx5ifI83z5wV+ktBPsv
KsLtwjT2cEf95j/TbEKN2rr1i8Iq88/89nZvUGX645BkoEEgC1mqMBUaR2RDQbS/JXeb31TZh75t
wg8RzyFPYpVxfUf5yHoECUkQodkKV2NEo2Vp6c7yLFiR6EaKAHKyGNgeC/XsAijj/B+2iuXwvhPT
ftFNjw4D0ZUn2y8MgmL4UVrv/1QN0UTPEcoTVFY3OOZGx3RxAfo4u0YmxC70YEHCihH1/H3Cr04V
/jXkrD35fIAXvfAUdjbi0yc4fb9KwG7/Iuf+eqlHumMOECIa+eIqG1HIfrGOGdHG2B9gzg+y4Bdp
x5213Vm7m10oCKjx/6T8Y/FqFgVDRa4nCxDeSifhyb0MP4EhrTGyCph96AS737GVi6NYsnfKl7HO
dDFTwsScrgSuPobJf/I4soejyi7XEHF8Yz5NNPnpCkQHWUso5MJYq/C1ZYmNEmZpboA3RUiLhDJV
xT4ddFLXGieuiqHVcD8XPpfZrHH2FmrPFdhNCaGobiEiD43hAtBeQi4Whlr92l5IoU0MxWxNSyFl
a+rhqEvme1Q7ioHnLoK1PvpcZiMQ/psG0iuE7F1bT1pG7A41BYl61YvTBi71VbRG1iZhEJ3GQreM
jV4fWE1apQSmHWNQ8CUJA4ReDr638OMhpQcEciMaaYxUg/U4NkvYDjFGPmEVqNqU7fNw5BtETurp
iR/prlqopGA42zvzWjCvB+qdKfBvDJBxzYwSZfR32s11ihh+UxdSmk9y/OtVePiJRUgWhPgYShMm
ELhCir5OvNUKclny71K5iTzs6kr8NMNLApX0Jb0RtfHZUKffhJvRYfT9QThXG1mxiKwGy6O91qSG
g+iJseRdkN/iRFgTsIlUCVkywtO4kjlJeBC/zuqvJkne6Rn6K++fn/ZAzH9IT+t3Y5pdHhN5839U
+ycC1hntFoa6MzsMHpHuUZMqLvmziMLS5TZIQcegLZGL1rBYWq1StiDGvHuytSzH6hF2xV5yzbM2
o45IEPBdw3RTu85VcVf+5tWVwpQGaeMJsbqywjBM5/gY+6zbwgAJqTzvSSIq3yHRDylrTmgY7gDJ
6RinLCPrlEEDCMFlaT2QYXXejL847mPRwyrN+luiXfi0jSbkfG+ZTTsKuzehXLAF6i9CJMyqP6Ww
Fc3KKsA7g4WSomOWBXF6ZPDbkgb1+3atcYmr5Pe0TQqO8Uv3MvOSJfLxhJlWjIhC5Hv7aJL2x8Bx
wNY5mkemAw6ybcaqGJ7ed0UYCQ1dXnAO6Kcen+xLhS1NElit0Ek/dyUgdhnqJ6CzSeVRNT68hX9g
zBnZFX24ymfjNftNmAzSlS8C2AzQyPOusXUAaW5pKwSVkSQcCBydTeT8K4RJyMG8m5YF249cLxmL
r/D3XudkaIXb28+rhgxyFMhkh03m2DDXU6PjmMFiIwQs1GBQ+sAVuAoRw/Dq4/ODGHQLEjY+D5T4
dqmkL021qSMOCzOGaToclyALVlkPrNncnm+Nl8Sm9hX9Z1fgeg6Ktix0CjGhnzw0Z5Pood0jca7V
lEMyA6uMacpciWYxuUBxq9RUb0WeEVr7bXkqv+8wC7LeVpOQniLthNod4Zvi+VDmC1UITqlXqY+f
N6aMqY9JhpdxpD3g7wMHRcO4U7ad2OkeI0pqcq5X1B434xqasW2T2FalK0ewaCNEaokbBWrQjppS
JpY6PAOPZauXjSF8S+IJ0Q5DGJXa8j4M0UjNfZqMupp2lvQdn8BhK7B4aeyv0qUrXDtjzPIzARQe
/H+pfX0mJQKkfgb2ScDbKGIwDdEX+DK9Ijzb0F0ARd1HhhUq78Y55n4uDdMU3d+tRnU/35yxu4HV
eluxbMkyk1rrMscGa35Dak77DeYKzy1Dg6Lq3b+TkV+aDHWVye27XktTKfneBYVvy9CbhugRamJy
Z9grmr0k0jZYQYrCWwVawkS39oudoi8b1YiPb1j0IUYTPij2nZy0mjk3eAbOkWJwn3KY9O/n7PkE
K16XrQxLBW0vW7jwbtUwV2D/kfnAm7t5CHXnIWgFwOWXCElfmKYzI+xjxmNEJ1/vV7tcpKS1PRLZ
Kti7pbcSWtVZwrbOzfg5RZvTjfflYQQQ4g5N8lOouq0LYS32soUSpF4HNYf45QW8KRKMUx/Ieg9d
2UW/JxnczcdogfeM3LoRtVMaM1q5AeI6XgXcwgnp43O2Nk2RLGcknCev5ybAn/F4dE4i97znWl/h
k299RyZ23HBE4P7rD6/O//qHL2UT442e6SWtTHyjyKyxtBVUIgsaGNiNwNBfgES8tGJdhmwuhcNI
RwDwNXwGqppZzumpbncBFDX1lRakLF/oaKoAYbGCXlg3SJzdgAvaDVFbTcdj/6RGkPpScU1AxcwP
5sGE3Be/ZJODpxQ0AIGVY3LLeFqUOcOy9FAKAeOHtUTGO7szAAWfvhiEVjXz4ikdvv83yt+oLPv9
4fJfCMOJXR9gLMC4k6Fc2jNdtHDhUE7XiXrdbvu8UGn83jbG4nvvU1ZYYUwT3AgLpo7Y/P6s0Pkg
+9fe64zOsQGqKfLodkFImid/H+U8aUSoetuxOVwyYsrVczDUC6+hPv7t6J/6/MAoUU+IYAGTomJN
ZtsypxcTeOhIvGC1H0SMvJ9aXNls1zZgOxcHGE6JZGoh3iCsVIp9Oziotl8lvKgDmQk/+ciTQ6ah
QS9ZkVT4JQtc9IHdZvPN7lgqhH/LiXLEtDP3eADIcmYt8Ii1sF1oeV74eZkyqtXYFEOzxsheNsn4
dU6b4Uqp3tt/bdhogXTF2+bAxlxue+UOaNXSR+HMOcreO1EsAvObtet0zFM7jkTY6xeE8UGVvkJo
Keu/pVOU9d9bo9YQJsOqaw6YlsJtFf1QBPnSBbndcGxUPD2Tj6z7ylDRrdPY8UOvwbBPDuwNaDo/
WtHeMu6Jcj1I7xMjJWNSxf0Qtrjou0GzHLuDfT+IIK/mwFzYhnWdIM5uDWi0MZMXO4eA9aqzcEDc
ha53u+HoH/iqqptET8PobXzSo5t7mMCFxqhO+NDN7ilsYimHa301T/cN3zN4kb0w9Ic6iCJOwA4c
hX2AbscMWuGDu6FOyqDmjN5WNz7nvJBD9IL0vixnG2DPwQoLH0kGLjjfJqJievaxbgPF9TyFb7lh
m3NcHcYu5cttLPaoY6odJ7Lc0elBFd6DlNzFd3VEj6q9mqqOgvLt2V8XFlUItUX+VPZLLKDC/kQE
fULIMqHwnykkHrinK+3K5bldBv2gYmJ51L0/kB+ADQll1W/fxY86nxJeU7d76UfWytq9QKphS3qI
OgmRqNMzur13iKbpbYiT5MPeZP9NKzMMW0CEtZsCshUCkDWUzBtjiIvHl5CbbEZcv1N6uAk6wOYC
xWIdATls5selhkS/mBnguMwyTaO6AKApLO2XYhHU+9yHDNMD5iwLlZJaV8cFsOJaMYjKFWuDC8FX
4iszlbZ+67WYZkYMMBbe98bFNEnFR/Z0uZi81WAXB82GW9s06kFBa78FtoCg2iB3RGtcOHvLKZWe
r8Mv0tec+dQpO/IQmc3IfWT1V9pri8rKBjRe+qsMoUEeDsgOncOHXS5xxu6lcN1uDFwJhbfrmxVk
QpW5fAVzOs/2+9FilBFRwHemOvNviT38qBVKJ9xLQX7cvVd7iolQ/nGYWsY7iSbuRnCfOKa8aaTh
OYEIC9mF0E+k9spopqw8rU9o71gZsYZCgeXMxUiqofLxumlRp1KHQUaWphbKT1tZZ/3cGHnI6BZM
wGSZ7a1gfx0jNOPq3gl6Ns1lLFQlf756xZM1VMevoZ7l8K6lujQYdGRgJ/RT+TL/VDV/jfzBeDwn
4S0rDvI6z0HNs6qoyDg5E1FuyVPNJG2FtigSXlPdT0PwzTI+Ki9T2/J4RiVW9Aupzmxscqd+W6ie
+5wUFJ6ezoDc7/A9mS61dh2Ve1q/MKRpA+kobm17HjvW28XFHGLrVwflLfUUxH2WUAsuYljsBir5
hjs/xQWvCOP1SKxZOoIgHFr3D2t7psoa3sQViYAYoSqn7h+G8Z4hc3/Clv5vg3oLpqv6qF5IukH9
LRYpq9s77ScY2lBav0YLVSn6aCGZx3UrCIsgJK5It4bcAbtBz816+QtmvMeG+YSvephzrB3N/eZv
QIouExgczTvd5TE9LvflO+njSEx40HhjzqvogFb7y7thuBAOLwk7waEeBu2BiTY2x2Kj2YxitDZW
I0IwPUTtrlSV/6aVXzSECEiFXMMWjszTHQlfD0TqcZi8um8B+mD1AV+9FxVbuNTrUp68XxoVQjmD
i9x9OBxTh2eQQjwxzt29iJ9vEzwe8mjJDAcsjc9yhMzgmIlSRq/Rx0xm/dZdvLI++jwS4akCIV3I
kKCNJcUUdVYLHeUYidEVrZixo2mH9RmwqaUWy9JJImgZxpIzopJ+MHu+O/jZ/3Yp+M8E0fnxzY41
mNNI/jfQQP3nYlViQebAPhqRPsrV6WhKBEq1qHbwamVqVP/xxhAvJasc14J0Ji40i54foyryjts5
TBFCFEikCZnj/oDyD3n5rmJbU1HkVH0w3J2GfOPifoVZTLuyzI4uGexnZ3xeeCVKKxFDgMUuern0
MOjvo+/DRn9XZgdPEWk76SyPiMbC+PEq9d2gUWrFfn92J+UGo+H8W548bMnZe+MnxkM0plsKyxl+
AjcpH9panRfJU/F88Bprtj+XoWOl6oyD5AvWCl+5KEfQYaFL/QTzpjP8cfvEuKFn/h1mF2JVpIcX
Vs9Ft7Vw/5oH5guPbzTXX3fvW3yKi9j6ErqFH5gUV0yPxR8++vm61SNRSmZpvK3APd0/JTZwNFFS
InNG42R19B7X6XvMLFU4tN+j1Lj82OX/Ti6gTp+4A98+cTBPY3jhlcDACjwJRzt2PpZ7YD0IQLkC
bZRC429HpmOchP2F0WhdBQ4JEy23b0AxWowN08p5iBFVtLiFE+rVvABnmdANsuKV/CoLAbdFsEBQ
FejWVymvst3nDhngVQqiNIVCeGmrwobKw5CUPVt0NUL7pT4uJDSP6xCP+y/Sfom+EjSqOwXXGMJT
VMihwo9VthjCJrmzY88w4mTMeEXeoF3xymxnPn27zQNvqia3DHjkf73KMIvScN3tCIzCwIM4w7R9
MfE07GODbVtXF/i8ebBChIzvUwLiwQa6rF37s1VWLN/ipoGkf5ARDTASuqwzyYDmGX95rPEMM3cr
WSgMlKx2WSemfgAKHujH+TMbrPCjjRKZ+pOaiGeLMl3VMT9qyLCbgMA3k0Mf+cUB+gAkPK6cZg+n
wyur5WtzNNNr05Jo2aTKiGQWeazVnmdq/cqkCAWstHqZptXBgIYvI7l3qbCT/Ikf12DeGpk4g1Pa
zl244oQKVjMJhM0dWxLZk7QIL5CtVr4UGIpIVNuox90G8JhQ/IvTxAnBrS2ZMVB5yuPitkMLgb2P
DC3nuLI984f7N/Mxr/R9h3JuUj5j0wNvUFHfApmcT6/xnpQ4L0ODox598u1vOViEvkE82XF4o++C
R2i2JS1dG80PM5wUyJcPbd+cp0YfkerOPFcSeEYqPaLF6hrQY5wkC6r8SPq9B19/fTtMJq03T3nO
HlTJ2fmqZsruBjSYwCsIc7/3C1BZ1p+sM09cPm78eeExuuJXevxhOkv8lt2CCPDiR54HnvwmwdF3
Tpa6wmtm+HFq8B7ffgHofxnBrsqFGyjaP5uWRf0SEox56eIZjPQSMaRJxlswDjRjX/exZuhj3ziN
BFDI4m7PQtCxjRsZLfrXjQQZwOczdtGg1Y80oSQB0yKurv8O2khgM4NMbKiRSqUsj1DetWygD31V
Ufz5/yrtXWVAPUUggyP33oiklSE33tci1JE5FzbJjlJaOqq41zzrEPnFnliks7s6iKUU4ZBFylT2
CDRNfB3Nc3rImgYjLTEHnuVEbXC+b50ySk08jF2M4DzsNLluBJ+V+hh9Zc1+UwzBh04fKRIWnmNO
9DDsngFEetvObhhNt7ecJZMffZ7L5PGdw7DQw5T5dEembhjWFqTsPiKqVl7weERo8T1cGApx/OTz
0LCgSeoz1DvaHCMIUPzFj37BV4muZBiGuJcwNu3TML861Ja7x53vgoSBQaiDd0b2SAUmjfdu8jaB
i6BVgS5MKahgF8R6V6jFZUS4IKeesB2iBMO0zwOf79+t0SpGVMYgQf+FSX7XcK5M1fY2YWDQgs7L
VvEoIQ/ecvluxl1NsIhPqCcjehCg/lqzMsYYjqaKygHyeK9uCPEcgyCTNSN1HMFG1LuQ8GdTQux/
OF9WBiI8Rfk6DdaWtX5QIRr27Cwy6Xrmbq1O1V+GnKBzrnHQ8M2O9Dahqwg1qhKU7zB3etP4HZGK
XtdCMkcYO08DsXbUymiwyF/kKnYC92I5MEtbO/i27s22/0CDXvHc1sk2uiOpbjkHDW7XMkPqaiUH
SnZeyUfHc5wlk+wQ1wunbpecpNA4YUl2scR+b+0y22vx5ox3TBs3b6pSPrWaaFWS/j+urjPKuTWF
mpGxWItSCXu+RqMXKG8rVq9EnJP9DdRzB6CfMiisrqnd4kAlD/8z/Q2gNCSvbxe8b6uOC8KOKeTZ
mbvSP9WW7YDmw2v/gDSLQBoBzJMUMtYTtX+uuM0fughnUTxl55fOSy528iLdlfmZF1E2Ub5weMPC
ZILuuInG/E1CAlJy5wGQZzYoNX9XJftTi5IP2bszc64SpYSP2pGrd4vec6ph6hMIsWsMfRIgD+DO
oH7I2fZnYJrEmDUJSBJ7Pr0iZP0wsmIBGLIIfYNoOslfi5mI5gbeOrNI0nPfDHP1FASfcErm0MCq
UbLxhaWzCi4i4+V5RxZZv6bDEV5TJhQuGDOEp68WfnCfx6vN+lWjJNnkZaWKN4Hz2/Ne35niqoie
E2cOdmvV6mm+1Nm5wQ5K4O9UAiz1X3KBx0ZRlV2QHDD0WeK71jhU4UuiH1tDsNOXZUCfnS8tM/Q1
6f1pGC/QswQk0GjwLpDJOjQAN7NVkdv+SLz4Ls1z7dpIi4qkfX2V+Ep9e7BIb+lvSIbVLz69hURE
vUsDhxMmVNxoVsRuYQxikeekmDCHgct3qLnzFv+bPXYQmAW/lMfEDbm+JxKEbOhfP7ueZRoTRDm3
tm8z8+HCVJe1Ad+EV8HM8cXNoMHbn9QFpFUXJASwljLT2BV/eQTj67xspLg02OYp0FHqBBhsw/vk
ozykN+fxsumCWLo5tRsSky4R/XpoEY/79pOQ90OrVZGNECdbQw+LA1OkGA/lS/WOd1Vesb6Mme02
O9fdkLu2CkUfNFfzN9CmaMGjFv4XtwVEK7jk4Sboyen06vSY1PsumJB3TPxr8oM8UvvAPKqlSzbh
WRN35eNCdI5tcAU/gAs4rL8hhqZ69G6WolyiRuYti7amaDnQNYCIhtEn732BPrOPOvzZn8ssFWY3
NyTo6JiNybN2rw6cOLbgdPi256ulUKVxFXB2GvIUsWxaagBy1SgYraF4p+nEqZ2Dg7k0hK8Nl8/n
WmCD9BWr2yMZBPDYJtjMjiYk1Uv0LCdSqrCD/Ax1daaWKUvOvQ4uwU6bdc2bnRd8WcozooRnjLt0
Z2nbB0RjtIO07wRyMKlKjigijoeRZBEYAxO4vGQTQsJyn8LdU8VpgpoCBJpGmZhjeYI2VYVFZVEw
RW+cf138erwWgnjV53LE8atWBbYiyNPQ6B4yA0VIasJcue2GYl18O6l1BKIGASqpUuEdR06Oy+Hb
79O4heyZOqiM9LvmpuobUcpvQU3+edN+eEYQ1YPlTN+IaHx94SrrQeU0ThlzY8c7jBN+gi028ca/
qS/RQYRo9xwyQDuRgoUbJ9V82IVUD88+fnQMR8aWvNTtkeKKIOZw1N51pHD2SJ68aWNbCuIc3bpf
82MZr87RTXbhS867p2nlaHsNYfkywE1hRc7alfdypXtRv561V4pVqNj+Ye9nLIMMWBmvXCTrIDBH
UXKAhfarXh71vh0mdYUJ/lW7HMkshOvorKrZYmyahKbV2xe4C/5C9MveIWRhOSKDJw/zKMeeNQ3x
O6Re5DbQ3gkIC33tgu8NXyL3yhlcZ+INEMT4D2vgsNu0OGBzjaofZzyHvbay9IKTP24o8fH7vk3R
cD/XbyC9meqYHGQpDvgan/hAq5gs8834SBzNVGHwlnZtFQTLRlV/rGBi8MZu2sTSjOkks5dJugGU
n4z4Dqn4gdDTfxEzxInlBccsgtNnBgispfx8mz31sCH3mSnVxkVbWMmF0ko34aMBcc+wjpSW0rtt
0gWDawgO5OYTDhOfAMSHqBIHAls+NJ2NKNjNXcqt4JJDFQcNDZpcQjUZfXgu0JXlt37ave2M1+hu
8YDNDYhlmJy/K805fQeDNiRQTkkoPKmiiuTr8CrOmuovVByrbFlGOZKOwNa2n0QprccTPUimSU+z
8FQSJ91catZqAosz4YK587YQ3ZN4gKqHb6KmfvDFlA1WhS1gx06j9Mgwr6kfriRgO+ximYmB4yTr
uNNT8+7ioBHkp21xmI8qkpd0VE+xlOm9r+xShhB9vNxXm001n1wX0tTv+Am9Q5bGIhu7NfurO6lU
rVPeQQLQlaaRh7VQSGyizMBJ8F80v6PpZ6MQBxfflJpGQ9mI5O4Qb6n7Ac4q6OoU3BJfucsaYnCw
WxRtGgkV+7OZIlQsqv1iGbz6LPt5fj7HYLHIs0QllQtvvCttEM6Gz6hRselJZ8wgNq8iv9qf2qjY
HK/C/A9M3Ipih3dmv6AKuSldPCCpJfSezpAJpW/i7KrTkgJdAQSKQcam1PsYIU0gpfGzFdM3Yirx
4EgxhuGLl5jp/lX5CUED/TsTw8JbKFwL8/s//5P+v2ekZb/g0P45onBrP/bOUCC+IhrN0qFRd0+0
dSxZCC63pmt6c/l4abPe0nhq2Pp133Ltmr592giIXV68s9TjKwKdZ5ubPH6iDAcDHVxEJZDSObkz
li4uu96rOFFEwfCGb34BfXQgsDLnav9SmB0cqjYGMHomxe5wYO6VZymGvXxwOiCbK4eBXmy8cXqr
/vGTMPh9WbApJ3TTMxJE5Hpmtv48LrG0owpA60FQMj1PFGEFkxlx+3Hd7vzghb7DyeCmDZNqTw/9
c0eP6zqD/SIWwmhCbn3fSTLDLNq2Xlge3GScwBDc/wNHP9X/S7qrbbhu4cbgG6yNqGR4SoYvm6+1
Rw/hV1dFe3yhm3MD9+BLLgOt+2Jthn8W5eZAXK0V8s8DhShMk4jK1oxhI0YSZLLSPFtRTMhl7qIJ
JYnFs+NDukfJQGArGwEIeUcavmqmvEJpblvLJYdsnDuPNlgWQlfp4R4aExsjdubfMVLsNkOSIBwU
0hQ0nJJXn+LAE0v4cmFZZus6QzPyj03I2pxX/fLV8vjLlMJaVowAtPJusbaQhxKn/4CTanRvAacB
/PbqVE+Cc0QDNGn9hJhuSIR7poIoWpWeuGBgYizrVA9qkZm7lBLIncd0BPz9p/GgTMQ/887rTuSw
IgINa2SO8PMebh/kj3qkrFVukw50PpgvWHHgyjB6jEqM6a+YlNXe2xCZVWBavCAbLXNi1oBFdEoT
BWTJddZKhj6CKieGsqpcgeDv3mgEYmZXGzNsO35sv+D/TUKtpryfXxgjZERWNLPU9d4QfmvoSyI8
RBEFiS/71sv5yGUHqbFD5e2CzP20XIM4mXHbfotVvkBSS/Zj7oikJISBYBUiw6bQ+Zgx1mrkLESN
InkOaNcfhrSvP5Dp/UvG02XPX7FNzkXb9dwRvNsGX1/AHAOPP77SncQsCau0Y9QmAYigMFppTvqa
2no7JaxLpkAe8+hdBLxLfm7uaLLWz6sk8mkiWNDsWgF1DDOoJLXcRX/2vA9N2gewZZFcPszWzktM
Sks9WmoQV0Y8f1Y3TZkIzOolZMMsXpATgbwTCOGhz4CxAYIu6k4lQxhaCTi+bqDAbuWaZbnK8rG/
TYsz0Xq/E5nVZdQG+9i+iP5E2+1+86fxwfSMp+JpogIMqmlfPQxTJcTrKGUT6iKbwVm/uBAId+rd
O+vPJCHlpeMzltuGWP9V+OqZDP71kkwuppzuAFhr+Z214m7mQvL2x5NbPwqSK3yGbKjq388CPnLh
l91QIqDVpkV/fohYAHXkshIM4lz2GXfqe5ElerfaRTN2mYmmvIYOA7BbU99lGWS42rT7pBGCeGjb
kcqRkuwrn41RzkttJJB4sPlT7QM5F6oyu3IHBAvYB7EeuTUASz0CpXByC28BTfn6D3iIbSOO469V
XcA8fTtizG5APHh8HNfrPMQ75MxKi/FaCj9vU+LHXe8JkPX4Tp8XqB4KHCXkELGOXrOYflCCt6MT
hIv9affO3MFkUxeK2CGuPTgPiN08iyn6lV6LRsBCpRC45ghkaBtraQxpnWxfN0/GJUHLNWay5Q/K
WdR/uHnfFtVtMhMK3AIbZUJE1cqvmqOQSQJyqIjID0O8cn9dn8Y9kX3s284oZcZx+89y6nDjm3Vk
WvPpoiDKtM5VhOGOlum3AG0Wr3DztX8oGtgVfaTudH1sfEJl1Ygi6s5HfSvFxS5XYhh5kRfgn/CH
ZZ7H+hwQibfj35tKP2QFa58rNKLlWJP1hbG5hcCBg8vo9st5OenGpl7fgXEi/yHQbY0BWlL6KyqT
3Vg1r8OiP+N+luq643FmO8lNslZDON/80geZb268ghlcT74R2WM7+Qr7Q+Ft4ADCq8dlomSse4/p
9si5AdmYRZ+GEPJSOZkPcRyZab56Jflt/oeNNZXnRM+iHsKNI6jOawQ4MYGk9hdsX0B9vHFmcU4c
zmkznyA0JGKhwWNHUgAVrX8VmZ9Pb1nAV529Ko9Dv/g0kO+dtKAycR+ADBhlbREJSkGFBR2OszKF
0epAF8ccUj49uP1IRZILseU8ep/0F+a85dMxrz016txQ1uhgFarU+h4cZ4oxV8b/xuCi0GB8RGVQ
r2SyBmDeLylIV/0iupwZqWbEC9bDWB2Ra+TEDNMy1MmNojWAy+Ofmg5Lhw4RyBbbV9y3gTSRzW4z
nDytrS9S+wUJxL8s41nVbfQnzLLBfztBEHw8zb6YPwUmfA+ngoR6oq7qKTayDt9+EWf1pJ/+1n3V
L4FjMHIj5NR9nVCghQ42EErIcoNozJxKj1wPPCYdEKxvaZKamd0myig9XizJ16bynPPbLjnG4LQ0
+eTK0XKrVWSiaAicCBmOuQiPjT/i99EIuOHwEZgSHRCJ9tKsA3ucMFk0GKoCBafvzlH/rMnTL6Nj
NeFwsGpuQ6lhdENW+4XEU/1Gzdyt28JHanAweMw3BriAfuQ7m3FkcjKDhm0Lfojglpx0V9UDFzRU
6rckGOR7JUjMnBp89gD5XFYpoweEFjKxM+FgzZ02di/ckq+SxGKkhQgVMAryM0kZaaHUqCVASUKt
1F9JEqH+ux/Jlg1hknbZ1FHVVzZCnSteuYNiWucUciLL4NSNk/adr0q/8EEr/6xUl4xaQjQ9gKHz
+3/qPfNRQsO7rfO1CErqxplL27Uup01tfJIsCPwpp029sGRPvmXa+TG7rxOq54wNNgNKYjlK5/bb
421pH2Rvyg5P1u8NkkUX1oxIrSVWsJ8FO7mVDrk/M5rjpUfK9lS4UIfo7MIJ8d3yVoXNZgH8SN9/
4KBYOtChLetcR1cBhXDlDTY0LdXc2Yg6QLFpY4vW69Fit3Kyfh5rAkXT/RR3oZg2uvXF9xuA0ctz
5CuB4VhV0Ys5dvGrnqgIoKbRgKw3Fzx81ZAivSBN1oZZ7sE9/ORSUaQGMu4acmIszYp1pC47mF5E
lOQ6QWf9/BzZ9uxSVK9VD56EjKQ7FdVjSoe1ToIm51FRw0nRxuyMy4n7e593JIBB+Ltj+fjG01h0
/l9QX4iB+05PZR2VSzjU5QDDXjH2IgV3mdzxs8U7GHemIfjnqcqEolPA2XckKf59DOW5vXTgKE9D
501E4Baa7CGBKrGwl24KxeHGoFpuWG1bKA9NU3DjKHWRy2S0Ir2fREx4mAxTkkDrUVwpDa8dxXqO
Huor50KlVgeHqnuiOWu8L15NMIAfTa+HewrR5Zv170AoZ9yY9SUfZDrh91DkhazUBWmlSjk23cky
ZAn6mKVBhqQA2yQIFmqp3ETGP9cGeW3ARnShsbynXkUc3kraa81tbsQxl0TsnZrwqAQwRFju1Aj5
sA8kq74t0poIS2zv1//ucXhvm50xPwcexJ5nOVHH8HCygJdTDPu9to3d89ugDLzdVGZNDhoH/zLK
xEqhzMIxpKiHsH4fbFQEWfHLcA5vglFjSLngsD4N76e/bfNVyZRu2z5lwuXTc1TQ7hgvi6BnECcc
drNP1LtGMkjsaZ8xPSsn5Vw7d9ps5lEyGzSm0MikQEMKJE7kJqMos9xHZS/g3drEJV0CD6icwCR/
rIg1Oyf2m+9M4IwSCQralitRzd+O6twuYJII096Umuooes9WIv9KL9Qk4xBlRa3KqU9OoTLMAlWk
cPwMGKEutltslBl0Dol+RiE0/y528q2KwWiZeuNfr6u5wtpJ+Xnjb0TT1NMt3eUxzmBGl/1LuV/w
AVOzS+zuLmh4iohz9+HrltRc4AgZZUXvSPujqkQFHX9bXWN7kcOu6M2iVPvSolMM8Cummxwz+LMT
NiRyeWHF/JiMYhlaUt4tJfKFeH4ZQkUj499PEkPWnntPts7niGEvyI7cQPKRIkaGW1Mr5CpyS4FD
z2yqPNtzsoT7pM+4wfu9LY2KG9f5Qq+Yt4y6OdWm+1vkhzOfBGFr58abXpO1Vfkunkx7rcKtc7bs
fxGeARVsmeaCcyK+6vahxp/GKmJYhvWjdketQJQhrcLEDn+JGallVFx2/UQHmdtk2AZtoZc5rPa7
lmnjQCsHKW/vZQRy+WKACAQheRKepmDCPsH68GhW6OvO3lJhCM59nSitHBS/lZsJopaAVSi//7Ol
TgCMLvlfrdVOwhPZgu2nmYsZtrTpyFZhSKlG9Uw+eI8lVCTWOoBnzUM6M+TW0qZ3N+Y65b/p0bCs
cJ8d1koume1lHXeT5M7Rhvb9Ci5/hsTHtG9rCsYv/3CqjFpVarbqDt1ML2ib2tWZv3nbYvsY35nJ
f2AsEUEX+tcPgNuakwNzytn3P+mgFUHtXv+3medzK4DAynhCxttlDvm520Wxd7GcsFzx+wpMYixj
lPh3oxQHOSo8ElE8Viem593rD/NRJ9eZduEyyDe/blQMjF2Bvwsejdb11DkjuE4hx8oo4sb2Wbx0
nVGs47BitwOKG8Ic6blSlbuGWdNp+ckeIAuVb3Qd/w0A9OKpn2uOeA8kKhdzJnElAks7EZZCXjx2
zLkgvJBC5cJZNFqAa670XUbb0K1hnSRgqKoaOXTttVp3+Uvra+btFfCnp+L7fvHFl2t5NXlldlpc
RI7mBX/FHa0WQVMCl+aGar1rz7x/G3+8znEgIZfqfVAehBR+fNm5mjVXRR3+QtPnSF756KQbzVyY
OchE8xE5E/0wEoHdWaUFsYM+x5Nol+UuMEwnzpZ+rj6fUlS2YFV2+072GvAbQCTjN2L8fjKtxrbC
zBi8U2E60oCm+fs/ugYSvU8Ghknuuj1kkEguOSf7AwufYSFMElfB6X57MSLxU6TsvpIoMsahSyXq
ULqnZiA5ZG5uMBpGmor41bWLm7UMgop49jb/mEaELMJsrArGr1YwfgcTwDLfPnXMDic8AaAgLugV
JjTi/pgDT3pFbBVdUA6usmytrmG1riJItzV7VBJi+qej2QU6NyBtVIQJWPfsYc8ooO6UJbpnIdi4
47RX2nhm3iz8PrY7ZDBRNqcLVKIUPumrbE4+AykkLlh2rgVS1aUinP/PcRqd3q+clRaAeEHVwoHb
+NtCPCaVPmdLp/LuoDGnIo01UA+SxmzG8ad2NkdoLLtZrh8GZ++PpCi1fSlU5wz3kKmqHl88KLpM
DqxHGcCc84f4qRYshPRL9iVAlezUS2FRFAT12Jn0ylNUuUaRlRicet2ja8Ds7v6HeMSY4hT9UCmr
qMwgXMfd7HRllYfRy8GnMd9LFC+sZ5fCXvHQkRRflpMrhn5sSWT1ytHxp5Og7DpHBMxCNQZjPjLc
B0dmi/En8bal4pUgVuHfilHAFGtZ530B8qYyzXwhBNce9uwg8H+B0ShKtg9/Gp0m/e3sHHl7f+1u
Sk6tsmCXpuOcYBvOBN/aHv3BFj5/Azn09XGJAZDDgNHQxxB4NtD1RYpVRSAhqAi/5DA2JscJnvBj
XH2ivw27OA/mijmPtEeL50wmcJ61kfYCwZCqPIIBlO/51LN3J0Gy8OyXuYOKB2NRbkwDJdHXMMXu
p+y5Z9+iSSooCZUP17QiDaJx6EcukksaXSglCnstAkyxNSuuB75AVUeMJ/Y/3aKcNBDD/RkUQLZo
n+N2SYdmJqvv9GKdxR0Eg16DmLNaKkAZrvrJQeQYce+BNktvKSWDG+U/HeWmtrmWvosUbQZRPo1N
iaQZO5ELZrQM7FcSF6ByXoWWFTw4dAeHcgSqDwE5Siyg/z3mw1hVX74EZNl49umLihj9c1yElgGH
XmXvmfIK53URZL1cYu8etISmQZt/kSt82hEOELJaiSPLca1FNvaC88s43or7c5eOBYXoDknfBw9A
+H/YqHwW5lekz9RTxzUTLzYXT/b4Pvl3hsJFOUoGWVKWOi2Nf15jn8fPOd3k+/0zGhPYCYvKDcpl
OcKiU/SpALWAoPC6xbJ6chPKQspdzmcLhlhqOsTZw/S7DDi4yY0vVqIIt453XtFxLl4A4D/C6fh+
G8OfKh9shlOtAexFHYVVZRBkuEpCnxzbNCnUjGvNLcBuyA6wXX9sArvgJrYuwA/2PidY0PjAA+QU
3CEjsM+nfHQNovQy3L/Iiauwd9oA7pNWPrWOuWigJ643xFWKGKOMuzAD3uDX4c3cTXZ9oe/c0kbj
dndQh4PrA89/4OVA9EEmFn27lZcxCy9QAWZrhsoFuYo7f3uYH77zymqSsHVeEiBqwViWc9WUKpw7
ebZcZfv7cib7f32w6DDH/wrAEFEKLdMUT+Q5s+fbJOB3IvTS5rEDZHn4Dx8tXk4xjFW2OYEkCKKs
7pD/ih8w+JGVs3uTByq0cbzZEGRJF2z2cydQqZSmB4uCroABVHVr37a6bR9/1v846jTi1xBzf1RY
WifR6X5bNc09tIXobfE3SuGfK6gtDrecNuQcrsIblswQdiSpNIzjJ/DCnrW0+Mvni3ZLsAUAKGbL
MVKNFIkHLOreM7EqvukCfLDU2Y9G4MVcgjixgHM8h0swQGqHi1K+PeUmqk7eI197UdTQVuNNKwTW
C8D6onwSe3OAScTZWCe872rT9kCera4bRStDfuTRa+1dx9X5D2lHONSvd5PQhiKoaFhakCTWfFmJ
9VjDSc4g4NZR6MYAsO0zQ/9jNvMpQbvNKtH7mHhHvxJ31NZNTq4C8RdI6w+QVQj5B+5JUlo7wzWi
4iLimhA4ua5QBH0sJ4k8uV96AJbHGav1KR4dmgbHhT1lIGsk1C+UoMF3Gm719V/a5zssgH1eX1Pg
Yz1yMugZVwPyj9ev+5B0XkmAxl+Baijl5LbVNvpUbzC0w9ZbpiP8TsI571Fe+pcuWm7YcAlQ4tkw
a0UmhdkE52xkk+DOIhGUpbE5jW/1zFMT+wwZOJQULkehxBjZP8AWQydV5awDKjH35FuN9u+X2nSZ
BclLj/Ac2oT8a29q18SQqGezutRvgWTG/Qw0ZA6+XaQGLjAlM6vubhBpU+jN3ztokTA4yAvm0TKL
daDnCLTJEYAdCwlyaMU9bX/Q5g/7xaOlJ00kYKkdY/2B0lvjf6rabfLyruCV6p8EOAmQaaZ20ww4
GcDCLNIlyj3CvJ0GCMmlBZbhDVraTJ95U6OdHJl4dSqs6USE1AHnT09oYjoMlagY3F41YIkGrOJu
EuTKnH3TxDfoU+YbjBTmlBAaUJNXJXYsnkHaQAdeeMkDty//qsayadzpV81+tg4lnkpm0VzRwUzg
21c1zjLPiCRPbW1yhLNYt3xGHSDRqXGlSrL2Xhi97P1yrHNk5L/pi7vHWhHWPwu3aCNguyDwGnPh
zZh0yQwMqumq3FLt8l+Lz39muIHRAyO9q9B0TKSovWUwF719Cv2TiCfWX/ILB3cycqlEw0D6lgq5
GNTh99DZFCdgGga7ybPAVmIub8hDDNMg0F4xkxJqY0PfkgGBoyhvEnxTBrmOxyrSCnRpym3GTK/0
Ai+aRMaFjsqJ0jLgDHYRxnQyvl9dgVuU86j2mYBSwTErrcHxEL7uqn/x9gzNsArzicvWjnmbt3k6
itDPRveDyGW3l2al/Cv6Lh0+ZkoCpRo1KzxKnKzRENg0GZ9B6Gj7Xdhk6mrHDO+O2fC1VMXmxi/g
juWzpSdFzAhcWqER0aLIZly+SzQ8dL6D3rMkDa726KAkDIX25tjP1tH5taXI+yydVCEWtde95KVV
+TAmiGfFQg5KCT/eB/ZUoqj4qmDn2PE01KxZ5wa8sX6duuDOW2tZWaFZzPWaimxyXg1Bosb3n4v3
mQFgcCV4Z9dTeJwbOsowU7Tf9wrbPJGji5qRjoHOpYxqXtuuAUrSpBvSngczwo5hPH15zSPwvnjl
gyDH3GTSvpjQK07DqZE/EQTSmJnt5YiNod01dtPQPO/UBbn5MqSWvL82Qi7ZjiEMKx3aPbYNSl6y
KKv6ff5crb/HCnPsS0XKrbS1lGCfnWlGTuWPhwTszshnMY+RonIZ+owdVTcJeagpeutFzzVK7r0P
A/s47KhgKzFbrW/8zPke6qVSWOjJ7Qu8Axv5yT9/WluwjViYfrZbzGiZHBneEsc1MdrFlJcxKlLk
f8OlcxcoKXFdcrhLdBwkIlpMd4rmPQEJrXOYktddzmpawfVGGl+T+N22FQxssbriXiOAwnMNnB7M
9xGWwTYOSZ72nrjwOu1qUNOLMTkAlahAdOQn2+dkaBTfC4516rcxtrhlJHpQrXXi1/5kdUeUQKjL
AUPltQRLe8spJaguIYCP0n93CQa7Sa9+2ydxYRkL3roXKddpk/SR7hU5E1xU6XKuwWQdbmgiF1Xs
CCyC17O3mmTXXn+7xGK7YA2tIidUroFNoeHRO3ZfaMXlXPqKkZ4CRIJIoSySJh2a6KGi8AN5Fae3
kNk3iSiQ/s1XioOoicKP7hgQNdyFGJUnjmz+DQ6Dr1cUEmqxrVObrRhDh28hZCffh/A+zIkZzR6e
x5rgMnm9mtaq3YAYxLd3xNEwGBeAC6JYaXnB5gaKAay8HwED3hBCFujgNimen4k2xmJAxvCBpQMf
dhdd3bSkp4GIqc0h5j6bC1g4swBFSJkXuSY63WT8evaoL5k7ljDrg+56j+P6uo8fqj7bf9kV63MF
Riwi2pPoOXSlIQLCjXdrEWFJ3bfDvcZUKacHJxtpyHF+oQDBG+ZbaLGcD1jfsE/PdWSz7DMUXXLH
2EFIg/5r8V01aq3G50incOQnDkyalpg1/n2DDC/IzMNyZvMbVJ/IlNUY2ehUxcx6ROeSpRu7R0dR
tAxnWf7St+YpRXJZytQA2+stc/3+2XJORmi7+ufMoj2ga26ED9qnzi1S8/cp7qlYlvM4b3RsOxDb
5ZK2RaXwu+Mp+jUQL6XweQA7UD5LMHm2BZXnGCvWtP08fyLvHUqK97cjUj6LMdn9bJuZbUGriZf7
x9yl3VD1Y0ybCcOfVwBDxmkCAtvYrE8zM+0EV4/yH0f/P5h6MMvGUt/b3qtQwoz+083qVkqvMpQ7
jBVHkuCgxF1YbqwtUoORnXunMujunXjYkuiBTRdtwXXSsLtK/7PlrmqvLixeI7Ykjwr0fbEk85mA
Df9L/+FiwXiaITAuHwKCjIAZrDcZy6En2Ik1GP/qPHP0+AKEFrFXAZ24rSU0Kz6fjcAXQG7/sWyR
F6tfypcmzvnzmuYlJLWZKruUUAAjAEhL8EOnaGc8wcejP1mMtD4THqpSE8N/d/Z6DE052vHbrE0S
BY1ef8OQjMIdZUEZqaAWgZ8aov3k/Hzzar6hfbElvEEFiE2/P33oGyjkd5SIvolefArgQfRt6gjb
3m1s2QfmIVszNUFr1oBm8QFv7Yhj3lGoxdTrbKLZxFJA6/xFZo/qTdnA1+TU9rgZi+T/sHHDHzR2
bj6IDZ1Rbv4awATjEBFXagqYmq1o3vK4o2byMiulggdXJ28ntT/s4cgKSCct8+X0vudGJakdc6sq
LIrVWloV/58y0vNjCSidQa158NsQq3Ft5oswg6RYem6ZJl1Uk3aUMFLuX11CwaLpnyg8JaCAF/Xe
6eztC0TdCUMYTnsxEqPPitEUrnNn2kQojKq5av/7EQUfLFKV+Rsm6+pZjyos8fg+sW69Jmzg/Unk
bKtm6mVHMrj89sBtOeKwcVyFAxlSekvxvrWVVpUXdqX6rfnCXxaUMVHz920JKvaMCP6G81DkkaG+
NReLUh6QJgAPnYSeBycjbdhHg7ZSSqpueuKkdje7WCM3guLYId536a+mML4AMvYwAIQ9UD8pW0pZ
+UZReuW4Zpuh8K1OB47VvYQWkEEoJX5ApR2H49Lqsvb0BMiBa8bmjoPI7fZVAtAz8xcr2dxM+f70
DM2hSdsC6KouKPeMqaR1Gwq4N0iYzzZQ1zH2Cd+Q18cmANSI4Wy7Ysb6K1AJoLPjieclFI3PKHsz
FplKfz5Pv2taaiswmHixOQufsBaGbHRMotFQFJeeH4IC2Qm1n3Sei66UXPe9JU80ksyx3e1D694t
NUPmuDvZncuOvFvgUf0Raws3eOVd+H87dTW5bnFVA6F3gGSklcW9ae/LFn263s5Ei1R/n0SqYMzI
v8xRLRcNq3AFm5vVQK2iTZJHFLYYbeZUK5I3LfA8npKAa9OdpPMzdEiLgD64vyGDF+gg48+l3JUv
dSSx/As1KBSVxBRSZXghQVKePgwoAyOkISdr5BjV86sp6EyV+SfhrWcx/q7hvZFm0RS/Bl87TPeK
GOxIkRlld/RkqaK+qULpoICz3eUr2JxSPCa2ZS34MsidoGUUKMTvCfwPjvB1kKx67CuhssE6Vnj3
jOKbSgOrktSKrU3ZyDKNsrUMBHu/aM9qI6dE5NkE6+fPhYXhWb4Rkm61dcCWKs3ZNBfZRU1eHb6T
aWzQunApvcRMjso96yKsxmxY5IVzdo69LhmdYZUuhrbOK9LFTq8xGk+g+CwW8EfoirNhrgB3/5AZ
SOSlkT0PfGIaYLcMxlWN/8LdT4aUx9tE0uQCBix0OuJrCPWaEe53/DVg5Guw0IsaDpGb3JpUZmf7
dRpy0ZebHnJ1JwIB9oyNkhzE3ISB6Q93X8AnOOQPO+yDcJRfESyzdyk9xsf5G9wqJ8LkpOF8hg/i
/g335Qz+4gKiASaIAIlWFObWTkNxsyH3f4KWyF8ycFJSghCdwkxKOgZHHGUlJh421ofpxSNDML+X
kXUFCKLDgLLT4Ww7xJPpsu643MowCw2D+fbOC3JPDo3SWsv38WBnJOJeoXAcEM5fkH4K/J/aZCK7
0tONSAuILjOl0qpKgDohtpx47YwnZc8W1Aq88H5GoEv0hWrlOcUdiknT/Qr1utiycDWxF37wvHOg
hUhSE6NZWwjMsTURgG+65x2Q+1kfYearoHhN2coUT5Z9lWklwiDPJDLkXP1Kr7FrKA2PytBEHiGr
VfkUs91ArYg+xkucMDuHksLBHlKEiOvfEuh/kaGumBSsLMeVZQScTUVDcGsmC57sA+xDt/duFo7Q
iyxM2JXDGq5Slbo5EwxPWqZvnHYhciYGwPaLUT2aKFUrgORCVSQ/b7SHbTMk/YZ5oHujZSANRl/7
43ezXYHA0XKpVSex+zfouR5S88vmNgoT+TPpI2So4FKPnRANUv5tnc4gUTjwsBt8q7ASihS8V4Kx
4trF7Ut/SJO7rYbVbNI2GRH3hsqNMmScFKa6MXHijTIV3M/4qhbTx/+mYMeCOJjwaOZjs14ebNJE
zVLJ6AltpnBidXLrbJqm8IV3SKHwsml355uCVPFjQVyeo19o14whf3aoQyfmiChFcZTQ1CAh5IHB
i4eDDsXc6AZZVqqXuoOtrGNfv9MWDaf4Y3Zn3BXbV+oB31EhbetpcmfdT7mxGaMw2MafFMWDEi9Q
SDO0xXZeKn+AeCEbH18rO2SObbB2r5VFjS5jOruA7aaBxy80+rZUa1NYj0z0kQWH4TOAhGCNrHZn
dkxsybdL4XTMPyQdWGF7KLE+fZ1jmE8o+A5NMw3WeXsavaXt4M834soC+zyQv+H0wO59O5i7bIij
hsZzKLC4Olm5/OMHzg+negT8HTzVJeAn4sJcurr2e9hFZFsf1e9nzUnCqBXd0fWz/OUdvk6PdTEt
7zKH9lUSZ8qANSHPhVk9JEjP/0LWM4sYRrc/SMF0Ee4wJ0FN/xVxrJHYnGscdVCUW1dt52MqPBed
KH1bBM58cDXpULIllW7WXsFICvLLWKsJmmGbQPgxDpCAbMTxCARif2gK4izahx0Tgiqsw4IvyNwv
Vtpue4xY5TZslPkz8oDLdoEmiFhK595LXWNBHI4xlpIK8YnjL15J1yHkNa7wEu0CAQrmwO2/gG1o
NKinvIe8zqDP8FeVXrlTCp23wn64LeFS74OFwoHSFwRmt3QV0omC1x/ldXb2AKSNzzFh48HVvih2
kWgKo+80+YeEVIxtlGNJdzlPxwIcb8EaL3IeO1VIdXlAyFOY5JVT9zxgOiMi6WhSCCXlxqKzm6Bf
aoGIlt0XYOHKI2hQlrL/CyctF+JuNuP9GCp+O3dKlMDNhv1P+8nIjWz8sVKwd4VEGqnOtLSDw6fT
zVPv6QQZj0R9UTHZ6ZrmyF4NBYVZOzerAp5Tifp1aJMld7LdiVa3S1uVK3JrkV3A2wzFvu1MbBxI
S5velBXotx/1xksDE7gb+z8mgtvEiXeY3CWNTdkRUK9j5oQXNsoXdP1dkJi6GiNfnrSuwGIxoWyv
MVixfq5/rHvrpBH8kehjALzB1gSSJTI9ZdYEXJ5g5TeWOFHwRKYKXXreeLBfO8FrDmvakxOOMYNh
QAONAhcbCr0cIRuXcoSQHXEfkNXClTLmvibTQidyfr2Jk1JXiMwTEhFOkDI9lEKIGokEMs1PwboU
W7M3wjfN3gG+AKvbZnKSqGXKobt+q/75NeHjQZtBpoS9HorB3/bFD1nNPJ+N+lMot8VG+mmB9FZH
P/FcJunUwDLugHhqnawmezEzO5O6cvi/isZhLpAAfYRYU2irYIX4zOjFDfG1dWv1W03nll3x/zSR
ZsZc53DI3CQK+fkBo/GU+CU0qYmTWmcIzeojUO/RA0tkppn+YoW6m9zzY4P1QUuRb3ka44g6/9c7
1caXBxpiTfTjXYTuVX7IFfK6XhiDKiYOhlCt5eoaV2kgB+5ZqjJLOL9yY1Gv334+cKmKTnkMseMm
0ubKJP7Luptxzk54l0Yq/xLSqurYVZ/o5ceXSEvKWrQBZfsk0jbvqBbV+X7/CIQjBVyitNzvgVUI
QYDSxT+NHc4El/6T4sXBKQMvQzNtuzBA3RzzUfqRUyrMS16EERx5vdrG+3ql3c53VVwjiVnvyyu3
zVmOYtbqKeEGR5EfeETUJf0eF/4hmqIfdkqgJtBWlDcQnTcnr4UggKIYZ9MgbmkELqAMWwv0iqOJ
CNL5mGyYKqdqg+bHdIHiyyxMhcmD8vVla8amjrxDqSdQrOAKt+1eD2953MIpz2srL9KFPeMYjkwN
Bw5MLobST/OENGA9AF3PvFn7bAe2CW0GwsaqqsBSgCFGGvTki+SPBVxuIT4/Hr2DmrE6vqEa2/zJ
5ekI+MLKl7Qm6raTDen+d4u0Hoa6UfdqDrxHyIdwu7n12A38lRZH04JJFe4Km/86J4i/TlXUBH+m
gvDD3D+CQGT8AWgWeghxPaggNtIBER+o2Xi+QcEtuylfo/I02E8B0A3tvh5/BmLshoAZgtRjY4Er
W4/9XsyO8Oiw8Xpe5N00s78mVr89SsPrpUIcMVSBB2TviMizrmov7vzbs7Vdlc0JfFaTSUz7TTER
nMfbcZQik73t9oULBxZmyCii4JqeM9zhdnhccvhm3cK7iStxUo1e0n9o1GhJNbhfzqU2KyUHqjJI
9VkE7G543/hGYlsxzVXemGnzfrsmZL9JwRWqugBLWPw8V+Dbz+OHN+9dOtso+b2tnoOUMvW6o3Qb
zp7c3X6ztbvIhRxTm8LH2JekW2ZMOBKK6KdtM1UB7H1blQKIWz2X3f7ioKJAsOeQ1YxnwpoEjYmg
sidQygPkN8zhEaVQyvjftnGkQ54ySYkaoYU8yrLs5hkMVC6bhUiDb5W4MFPnaayf3uwZw/eAGuiP
KHij1nchQ/i55dI0RyZdGTMCFkR/Dg5f37YK/e3r/qvVhkOuPn+UQxUvjtPvv9nbkhJF4W8V+McM
HHBHZZNQfmp7IbKL1pT32aEiM9lp58lP5PFHQAvr51XNEzm2JcuSyewDtrvRf3JKYirXqYRqJyrx
+aE=
`protect end_protected
