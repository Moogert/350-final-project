-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OKFJPXoPhYVRQiwlKY1VxvWGAiGuos8lJTexq/rdRZl6/WrWu8Cw3isF8l3BuA2WWp3OuRBHsSIU
Iw+micKTV9oxqExm1lX9Sjc5gQqGsVcNyngOCib0lmgu3lEUTueXN6PEdbAjrHMGgotnNeOCAhxq
bDSslTK2CK33OYfQG/c0N8eUqxMWmpXc8wVIyN8x7Lya6rTTn/92fIAcfUZliOvDhH/rrWqhDDo5
J+NYG/5vlKE26Ho9RBVoaktMcWfaraKU0/Lx3sN84QXOsMJPJmiNxW2GDvuTThd1pS+/R6bwE1S/
iZkImzI+h0+JaHYj+Mvq/RxuDqgeWw4yy1Cx7Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
C6Um+XlgFhUVmoJ7Hp/tq23Cs2epOPR5u8VX9ZemwG9JLWdmhac116zBxbYfgfIeyPGUYYZkTn5H
FKciDSZQqP+Kuy+IREuxJ/ujzKggwoRwNbdW6z1cxW6XcXUTGRpBsjf159y6MMFE+jQQotiBqP01
NkJkS3U+onl4+NcebNuM3plxUDojDNS5zy9a12sUnlcw12uigJaR3LiwG7vf/+Ev/deJpwZ6U2ur
8QEkzqHCCja3PBuROjJhu1VptU0zqkz0Gx8cSj83GwN5u4UOochIZK3+IV4B8Ea9k3r9AA0dC5VH
jzsxyCfhjgWVSmfEPMi58frXdtmnLYSSBeM/XYEXVhr0uu+q/5gqPmBa6j8eq8YmUqvhFScgVm5+
CpFeweWx1lra6Lp6r1fmc6GnNE4GEhYUiyxyvhizXih+hB3tqcYw0UKCJx64lkTVElYu+bj9X5A0
yELOXMYKou3Hr858UVGkKEhO7+VXRGF4u7ds99jZJ6ij0baZivUzxnNXm8qNbedCHvhpXexUhcbF
kwY6kxld1FrXktGv4RXgi3foV0g03GR/uqT9z3KnxoQD9th/kUOFpKUp52v0ZFioe2bFbt6NuSn+
ZOAWyZ22PuS8iXxihFkUO5LKeVDDBEprIU3TL6luJ6lUcveAfSSQ27ozbSCQ6nZ2C22o0nEsUA4G
V1vqBG1AYaS/idHC/SnFHv37+Z9ZO5CzkKsM3VMWH050LV7ba1Sq3h83C6/ybNxk3YeBZwKEyFmn
+Kfrak3zJ8msyyfiPcwHInKB4ctDgC/RAAaWD1vl6FL7+OjIwlwm8zxUVMuUCbwpd3JDFGJWpr93
dPMlGRVbrXXjfWTRkvfxGTijak0nADJNYmMT+erLLFJydSS8AZhiqX3dzJOLz+peDvDURn52yP/E
TRB4TOoCWL5+IkRVGMnJmh2pcHvNZaR5ykwyYF7V2/ZiCSjz3xZhxgfFjtbWZZIqzvtYTiK/fifp
Mq1wC43z/czwL0dgqqsatlfwnqJ0MGhnuOyB0lTAkyptzRz6rEBdUSuIxYc2v25aUI4DSoaA1R9/
Z0anZ8KKLkknHqzyQsxCDPqFfmeApF2DUmdQ+GqfcgGi03U5A4d59MtB+pH9WcE9nf0JbG8DoDMR
0VSpOkt8WPPAyKvNHL5s5fwQBYfE22G0T2FOzDNKEXIyPUhBvT886LKBjnBQ3XNqAL3jlodEjicD
lo5RDgrO17PO3CE2yuiqmNIT+Xy6M234Ge1Ud6xk92rSECmoC8iXV02bdZ7Vy9ceevX79Lyv+HxG
ShDBGB/AGYqUczfMVWj5oYl2wgFSJ7P99uy3nvl7tO3HuxyLDLOzZgwpTyPmZODa9h4hUqWwB9eX
M0ivJPZ5Ori9qp3DfnuPJKqDUQydfOYGxF1h4fkQMbNbltjKOEEqNCopWhOocDv/Ed+RVSRfDTgt
6Az2fXndMZO2nlEySCIh4IiKGiDThJTuPwe3GescommtCVVkHviuNj2u06AIzT13jxCtqG9w2eM/
QtVaTVxf+PmXd0aLKf1ZHCo46HEgWxT9rVQjMj1TAApCrqKvMuFK7QugET68DVp1Sv2hxXAw/jU5
xsKkxj2CkTe82JUPMnqdkTlBgApsN2m9pwNQMgNsnBZ53I95rVGO9y/diWLA0v/P8kC2gRgh/Ykq
DP/ZjMkFSkSNk/IvQ/hTFQGsB7btrLjx+h3VBoYpT2XC/6cRzEXwyTHR9nVfBPvH63K+HRU+H+4Z
eUak86Z02b0ZoO0nRsbY7gA83RCqWX6EY/PEmFJede9OAQ+F/FRuqnQIXlPlB8c06e01MjSUmFlw
fkFiO/2QQQHDltC9EOszWyTGpUaW3PrCL0ttAGEy2M4kC7hVbMvJh6CE12JFuNudGVDH6DPX64lz
l6Wj/ZC7OP0zm4CPLl7KNxdh5z/eovrQXH4fJgRnikcu7Y0TbpwczBiovG1lM0Via6t4sW2kd3uO
9iOnwKnRTUwoecldOkV/By84/7I+Bd0XWUJATGlHwdkU3tRz+fE9fahwGUsMT94wQU6pF30Llbu9
/X3uhvtKkn1DrWuP+/5tahm+03RuYVa3IIzn2thPk3nBd0QgMC/XsFD7gIjsg22VcnJ1ub16et79
9an0BjIEKOPaEANiDD9VylQijM3/wZ6L//yQxhvlAHpaoiMuCZ2pHy7jm90DhzrPiKgOrVd6WrEY
/LkTvXMs6bmu8DIiCYPiFa8XfPNNJh4KtrLDVVhiJm5TaiD0/t/a5raIVJ+gWAwq9rPPrVOx4fAd
Q59IgNytHvyv/h1kUMxpWF7F+VwbF3IyJywHNYTXbpCll8QwKymNHcafRCzhvjnMVdtXuSpl3voj
Hlszr62f/rW9LT0nOXv8t9ZnEZ3CQLVMijlmsz9bz8NV0U59z5ElEPE8V3ED1GfHylwPJ/pF2+VZ
O0r12PDm/Vak0GKx3YvofNx1rA9erWaJrOC2v5C0vlZt3xG0fLzeQWNev5knYUaxe+h3uEwH0LO/
nHwbanLeyoOUNid1TJgZrBKEmq20iMdzPTiSzbH+L9Tve3Lb5DFSnGn8y5CcEwxnPyxNYiOMrT6g
X33806eENJSwffVmgJW4FVmr0yAsZzdSROn5AmzFm7lPYikvlgNmms7kv7mVvFuIWb1Lr803ZnuB
UhEPtJ0aCs0IwuS+Vxgvst5wt+iBcm2uyzovXCy22slGP5rkC6XPhzzCog7k3SNqTc4N8yvtgm59
9ggatc66Tk6aC2ypD13lZUOnmDWlFq2YJa4KfQBV3ADxzQx+J5+QVXlLpPP+U7pSqcEU/hhiC0fa
fDyjoIjrujPuhKGDxhPwnG4zYRYL06WJ9Df/k0F7UxMYGlrfzZiqdGJyfirOSeIjXc7klf524Yrp
8yv9AyikryCV7clkOtZH6EvGz0jsRJGg50q73KMRslHvGBEp+P7KePClTVL8sCdE9D3fAs22Ud9p
SPWlWCz8CKbJVshgziFO5oQgF4lfDQOLOkJ6RIUYkq1UDmK6/vm8+gJ2wUVOD4KgUDDhNwCfmVYz
XM6lnJM7KTJPzrnXgj3AJV1dtAjEywfncES2nug7EzzuBddqJOpBt6iKCsCiBhNmiRChhBuJSaR1
NGDNgmVsYgXoN2VwKqRoLQPWcFvUpLFwOESAnY6fE+gGZHYinmYxmsB/zK9A3pCCEvaEgPlgIaqe
f/AeMC1ix3gmB+NjPxG0tKCsmPrKV0GZt7OWFIAxJwsMjGkQRQoqczpdUSi9eh8s3Spuwbu+RLsR
OIrCbXk73jun5F3Wlb8b+r7dX2z9yyHScXiBMf+gbjnAvTC3iKNqVrKsezfOKSbbRldpLuI6dM5v
4ObVPNw8BYcVUWo8t17ZnFkdQotOK45ssz3duzJq2aeHD+wMdeLGfr0ZoQIfHpL9wLhrPolLukLF
oqrUetj4T5lhth96o+v1uKXTHRiRQ0CDVldzIc0jD2rivE7fI0QqBw8tCmNeuO/FixzCeuYvk0Ub
QDBR/VuVhh4kRQ+qcTluEYHzWcUVjLT/PCTKh7Xb4NjUiCaxyLta4J1EVnWrSG9VnXOGDx6dI/xz
bAUJvBPPjlpRyhSe6wXlVSieY3k4H9qPOKAXP8bEIEudPc+42Nn+eWe4VXVjjxqWdEQgm4zrn6+5
4mRcx0tMXn8i3FtnlE4/5BWQjoIzsGfRGwRt/8QcYZfzZa1bKUuR435N7hCEuam/d3TX5440R0e1
Gvp2hqDhO7tBl0fLxa+FnCHvZ/TNI5ObDyphXsw97DWhn9eK+gHeVK+0UrC2tN2vUAPb3H5SAQsk
DoqewgnFYPq5iIyvhhdnLy3qoPu0tn6ZTtCiQoodoVR+QfrQQHFChMxBfTamW1IruueCsOQdIB+y
W1lpbBQWhi9cj8/gNB5HntBrTkUaZo3YmUjbuIsgwe2egrYGGrsI/siVcUqDLD1cIBHhOK0iXFka
yPywfzHjSBz3moebgcFnww37wLInH8dLHIdpv1v+b7Pp5PmJtSCeZtmqU23TeFYR2eDXha7Tx86o
kQK8jBJvCPybobUN9chjKWgRcoYniuN/KJ406S006CNx4M7LYaSJsRRwYzDQ/5c6jXdflgizNj+o
6DQqZhPJWAPm0uiZWgRId1IWYWu9/PzcBOJzxCcfBmpa0OMzyvN+LkvvZ2GcutOw8zl7E6pBrO3s
z1W7jJPLN5rxlSb5yhPzSfHqXm2DnYxsOp5EC7nayUJxMOFeAxqwJIicSZDFyQky8voWbTtTPvJH
QEbFCibAEVeiN2NX62ziqUW9YjyjeXayL/QbhRcjyyAqWfu1PeBRosvEzPjjIY2k5o2KyAgya5Ip
sgsebug9YrcCpcFCVPuSfmS56sLzHpfoENUrq+K1kQv4dBOPd0DEOWFxfYEbhUpFRA823X9LXedF
23x3eT4FbEZBb03zhdzFR0VJDmjxAZ/Wk+u+jY0e/6OQJAFYZLVQJq/1EGmUT2FsgAnPn/q6sGCY
mptvcfxV6yy4LNJyK3loF/j+MHfN7M+ofSx0FsqW11C8di8dXGNvKmDdtdB8c3I7UQ2claVuAjfT
EVD1Un27wRDL/kd4ANZ99IcmKiYhoV4cCUSTwjs4R7fyQ8AML5kOsTUXzW/cGp5EdZqiUPf3jnuo
bWx2q04FVaTk+DW0iSyKeGusaHPOdfoOIE2T9fjeXl4pLh6nh/OlEna1+FuFLn0yb7vRTeXipx14
YpwrtxQOMF1WVYEXtZhW+XCotbvGxgS8mm572kiyzikjHBHwjJ9W1mdu7Gx+hT/k0jUNjVcqG5t6
YuKXaRY8o1l4G6HOkjxrM1ako6SUuX5D3ppcoLhxK1/G/EQ3enQR9c31yGt4FrvTkrqQJP3SdRpP
C9L7tqGp80EcgIE/bd6h8a0XEC1V2hLICJdpPVVKDAVKHi+ChpuXlfPiX/9hKESZMLaXT22s9Dn2
ieUu8N1ooX+OFezHMFmi1oB+SvAEvapi05QynBPu5v7XDXNiMWvjiV5HALgZyOC4K2C76yoHDc7n
3G60KIoQwyhh7JSf50tBBN7WVQTPttKjQzG0l8FWgZNsKmYmRCKND8zqHtJZj1yVVj4hEUYCrkeG
4Rhi7Me74QNJOutaUiaDx1SjNTDp/AeNY5go8N2O0UDubKDJsqgatLgVDk1Qklk10WXXqw9WN+r7
H99t3Cd0oTTuCUoL1PMQI3z1LRxaFLxavznIijy62ISwOLVWzI0WJ8mFNlv+sUJivFLERO2fRhzA
BzPU3VMk+8IRHLKPfCKQ4G9qAwHCUAuFCwig7eTaDV4BP4XmZg+tiYmWHLBdSqs9PfekSbMOogV6
PggmNqDBmqQWjdZ86m17rPn826MJYprVWdi6KlBN4Rms5Fu/Xly2R0W5ezNS4Txf0akTxc9yPkSp
SVlE+VMz9ut4oJkHHKP/5xUf6/ZHLylwgQHymXnv22Yqu/uuTJ//LxJS9gBdbxqE66WxO4rqj/No
diUrQj2wHYAhuLLpZ6daD76Ij8/OF46suZWNnNoUz8hNFMEV6wrY39yyHgKcmplDl8e9ioXqSI1D
2m6b18HX/CfeZCsbSrRJafqyYfzHUi8FKU3r+FbCpJmLC4M3wGRgivdpQu2LlmWwJnGUtv4bOHji
8nLdNWDYrvJUbgVaHDFWwp+XJJ80nilIOGxw6LZCLdqwSyhe4z0cV04dKqx8PFjqTevmyeMeWfO2
6V+c9Q7/MziJcfKnF/ruUu6Ir9nZi9gdG8yRehUzj4QNt4mK+Slyw2xCTvMM65m910KJKgvQZL0X
k8sLoq5IYLIyNrPF1w8X+f6qIMzkvEbfI1SQ3mbrtqRg3H1tcKFXNvpOCi8utp8ZdW4NSuuSXN0G
Rc/aTz2wTimcU7Jyqbxv3xvYXcEbT7DloJjaVmCnv90S8qWL+V2LXPv3jD1lEDz0G7S+CbpLebud
FW1ftFzr/+JSMCmDlURs9zyAqMPgYngvtNdGYp9C8drsUmquv5plE9ZWVhcdpvLdC1OWbRJMe1IX
DoRQ5YrQ3vDBJk8sg/IHTxa5BBl4I4FWmNqv/7ivuybpeQSb4mFnR5vFpMJbW29U8ktUzu2HO6So
rn4hPmZusYluffiZG/r1tXc97A9L29QYm7NiHAoOdFw5Lt7dttZWINCiPKmNyTlE2hhxbjJ9MIi+
DQEGQZmissxMsrgfupyNrfLNFwtLh7os1eR/LVBLz42Vg8BneK2I0IvPXO9o5OhgzGeZiZK1BLmf
e8mk1P1P2NSpSYPQRx7uPugkzl5RbhJhW80oQcTjqOycNnvgOhnSc2VE218J5IoiV5khhi1GEhLp
JWLK84B3oLw9Oefjud6av0zycc4OKMHQWHnOOmDRWvfZCn4hhOgZp0cp828QVjUcqvdSn4UbmhE9
4x8P1Ru0ARqJZGvW3KFqC30AK1fehDsTVY9oo5QH9KSfskoQ0MODAR5l2C6D4JymNxQVPo+AU3XS
9MJd9V0GL5e4raAhqssV81sTZVeZBhw26LWKl3+OhyY7MJcPQFR0IHcg9YAsqKREfHI7sEBkKVpC
M+AkT1iWKNGhQWtcHcXzunFw3dm8QVYnQWl7P1KqmStWg7sCHG+UK0hbKQxteroAznHXoD1dx0y6
S7nzXq9JODt/QKlxo8p2oKTRYoWvSBh/0IDgzvmXFzmP9NwStpNq2wUR5Os8aZChkqefuefPDcFZ
N5tr69QtPNev72NWlBQV2qE7oR+2Ldu+RkPw1SfiW85PqSvpJovwcj/IlLFGn0dysSKgaHXocRBg
vxNYthNzM8l+tuep0axdBYL0hs2Fd6sfTzocz1sSfBfu25MdlWAQLtOxtJg8HArmbzALDB67/4Fz
Hu0bk2jBagK04x8x/lu0h04n08y2HeZKOYa8OU4eoBmhM329+mKbPUbr+oz2boOqzMewOke42pBV
oupjKtkkA0U/GRM/9Xzo18D9XabhCMlQZnlSn20A/DoCXW45+vREmdRBta6rjYb3Xn0gCNg+XFT0
OB/qx9VhQ/P1hALd+AvhmdzVfkUkpVva4KcM0uD+n8vuFABiF7T5ibFMzFjC1zwVjBew6Z2t1Zzz
8o+7WdboCJGBTmeH3GEX6e8lF7bF2lHIUj00cZCKHV21rhOEKk2xTW4U5ojxXf5rImlCJiRyBqdz
5E2kjvfRTPMqu1/A+JyeH/t5l+YH26U64D+Ln/1LD1fxAnu/gwyXj6yag61W7dy5A4wL+O0ARCpM
kGPnmCGx3LAPn8mAq7oxfzmy48KY7BCxQ+8jjG3EaUapdZpnYyOpOxqpmv0xjgvBpDpe4y5ibbZZ
cpziOemMRgxFP/CXC66k7LbUzT1aEkVFaF5+asw2LdjZ2NHskpNGFk9ioDY8IyZa4WwDweKdyNT1
fsRlUDZ5p1CNKFDc3VgSsfmbvoqjRpEFJqiuFnfPIOultlwsdRSzONH3CXnEv/NyXNxrmLfbCWvn
xZgAb1q1S7Ix85khJl3n8+Ua1R/WgXA+gGh0EGEyVrYIVaoIKUYOIybc/kzEIs99te84E+ga3lfe
kRcO5eQYdYCpRkUyLEdNKeJ+Ier7cMeBcvcdezsZVTejLTO7cLOzirW37e4JMofH6Wyi2LPTjH9l
w8kYBSDbbWDe7S/FThzmD51Vn2dBiHR0AcraYh57wN4iE45upb00kktJhIO2vILJkVmKPejTueKM
cGrHM7xF9ujnfXdjz2S3hV9Fnj3Fi6XFyBDKm6FypS3pFD75rYZremIoOhmibQ24dwgXhRimG1bw
9o+kbUzK3EYFYT3O1oEwUyHuF80AWIJs8NAELnNEVnncMjoDchR3w9ApxsTi6zH3DRTL+eTrvbQG
iM3Eh4NlYV6c7uAoS1OWZTo+ZsVwDRQmJE+xXJ5M5D04s7W4SKAvIoqIpuy8Nn8XZQxZIOxArVxV
POfJlUHiGWaUB+VPr9V2XWRPUpO7E8EnK9t40APJA+e6v7y9R+G6LcW36/2/o+PL+3AsQqYIJf1s
9qWJhTlAu+qeQiTZ7/ZD5Cv/Ar76jzmwB9uQoG/ie0osXHhMPIgjUo3OCaUUl0+ge+X52fpCBvkA
u9UgXIXDD3vlvCkwhCLwooz+tr0I5dMBdR2uFMTPvi3PGbLkgij2J802hTGEkQbKKOt7LgEtZvsO
wvpjTRQveg0uFmgaxItxPgIIoZsWlgjAsYXw5QPP0BNmp0bQzZvOvjZA06qPrEpxcHEJawGs05zq
Aa1P8bGJzlOZoovebh/fhLK53qNVCsCoCvig8aXHOGTdwUj4t+UhwMbjusgzYK1EIjWTu0z/nWG9
Xn1CsN8UoXpwAjZL3bkMJRs6D2Bl1mEAI/AbTa9zAcB0b09HaXdoZTnZbUT3Nrc0VpUexcnFf/Og
LSXcfB9Zju2N9yJVuL+RGHeElbypAKnUiEqGgtj0fzGwpPkXYd7lGonCYbzwZFZvhey2P6R3X8OW
wIXdqcYpcoiBYk49vQeT6urrziPPfMJug9HH/gdNwfIX13uhS3gAP1dUSM2mXa27K7MNKIEZUJW/
9lx7q0gyvSlYM2ICcusjnUdvl/Be0I2s7ef0hcwgvK5hFJp/STZqi8Xq+QqV5KKcptXnpAjuQSRD
gfUZCnTKshK/s7pYMm0uMUerT8rroO5Xha6UtE+m26RUilnGJhQfsfaoHbpbUXiGeI/2kg21VThQ
35BUP28aTD9NfUjFmn5OMA24iHGe7kQKg/Q0O9PBEOHPqLgY9whESF3ioTSfRZk6K0Wmk8vNKRku
d6oKo0wMuuK8s8bU8h3AvCkIjqkkI9RvyZ80LtQtc6qPCZ2zWEDIch+4xPhXCq4v3jAVRdds4cxg
vzVO5sPHefJserlZzwTj5lOH+jnqgI1l7uGa6dBQAEwWzB1JnVbO68IS/rEIPmmlMI2GsaBTsJMD
jE7/ZkEalrJ+hSFl8aAFTN8txTBKeJzu0WYHprB58Ke/mZZXzslDpuUk83CBlOz9KtaThBvC69Mh
YsQ1EnOI5VZYEYYRfiY7lDC0GqS6IkIGGW/tgMaoDELxq8eRpfLJUqb8ciNPrAQ1iQ9xBYu05rEo
zuZx0XJuQiNhRNkEm2w8pXt03DkWwu3QFJsmknxHYTiP5tgjgmyAFqCH1Nkyqj2zYKUK08XIf0SA
6fSokCc7mbyF6iexERrHumft6/XzI1ptf8B9mZSxb9qrMmC+reB2ltRvG7HN2fXxiij1aqw3JuCr
YaWHwx31nsttTHhJDpTbZorKsIYC1aOayzSAkFMYR/rKGo2rIkizm5/hRhOvR6R9DS3yxAiXuop3
Lu9iNhQHVE0LPxRV9AJUTsTefEzTfsDhY8nyyvFVOzJQWhFKFmmRdUARXlEacbNIn+UB1NArhGBS
W7edKX3NQ3W4unzIB4oB3/iqBIcg9jg5EzP8R4mjwldzxZNPQVqndmDBOf1Kl9bUkukA2Xbm+1nv
v8W/akz+XbZL96XCljbzvbKm0im+rtD4vPaAGHujXVHw36mhVANQ9OWS01J33so83CMtDqZzOq5v
ICtGLyNzbvQG2qN9QLjRKMfZlx/76Y9QjNXj9wLIm7uUeGEfZi6MEe98nmkY09FGw4VdqAS3JLwy
4YZKkSAJSs+VcXXn50DpuJYkTvhD9rMxQjr6A/JLlHzD/HV9gHJ8TtRwiZMdlYvab20FOan+ofbf
E5u3N0J02VZ/3L3QZF5g6Td0/OdRK3/vvKc3cQdvGIf+pl6QUMUUVLg/a35JmC1/6Ys7Ogr6nFo5
6rfZuZpKLJtRClSS632d6JLnPsGS1jYuvIo0H9gikUK8WhsyZu5RVP4P4GNHB856QGKpJmm/p6m1
MeJqbcXPNqF0S9YsfM/nfV8lZFVgdx4i5ilTtCH2vBrGM0djQaOdLNkBgo1YMLVBD8j6pe3W1IV9
LC/rSeL2p8/OSVcNv/8lC9y1nECYDR7my6+960rWT0zUsY+MD5VjBvDopenCf16iUmxRFPJ05bT0
jiYfFPyOg24+3eRLunpZ/6q2nrDscnPOjsRd/ETaRERWVR6ltnabupKm2aKI2hclKGqPfUo6HAYU
IlrpgRrGWn9xvKud6boMgs8cC/euXq8kFRM1E58JSqREg68OuTSOCHu8a6Rrlh/Vc+SHVOiAOFfV
4UgvNDeMr4JNhtfKxeCE721CqG4nVEYMsALOFjseHXBYftS/oEVVfUlaSw+Jx2IMDGB20iwYvDW2
WqACK3q0BH4vz4fFnMk8vWK9LNJEG6ZioGUeEK/qBpHvQ+CmbSDuReoJglkys+OHc73NPem5ZbUT
UuBLM3Twb7M/gizmw4hIYyFpKF7f15mNnei8awwP1nllCSiRcRq/vct3AIG0BhaeuOj/abw27CTQ
sDFQOTtWno7Hq97zn8OMupjqCUZ1RYuRKFjtq+bLQs19KodvcbZAT8bNnw71Dbh+DASH0zs/VRES
6Rlux0iKbBYJvFzRFzR8hsJ3qAkWY5nARTmI6cz89DUAVjKgRZ55NBvkuqED0CUfaBI7ZR1yJxbe
4OvcdNgGwY1US48ByGobotKsAzgovqbuTVCb7M2cxdfDqai6v6qVq1B3sa4CW/dYajMD8awcKjwQ
TPUgiKsAZo7GTxP2PC5GIx2qJ9BWu8QpNPCSFszHstWTMq4eTHwCHENrdKfZiI3o8JMMnZI8lN38
4izFxyo8XNPOF53Ab0/2xmwesAbV+nUQcxCixAoYSKCM4lZCAosGWctEytsqPsz5aSrjooftaXGp
fucjazvL9yr591sY75/BQsTYwmqQQOZYlFkhG6FdIfa+TplpJ7c117Awl8sZen8QhTljQRa9TLDd
PdYIEDidhjWJy8DaFdbqtZDIsIKeVSbNvF74G9jF8euESQu9SErCZIhN7wwExzNWflh6czBBLFNc
/piRLkFooOzvoEi5fSySifOAvPtUbZcWYV5XAuPo7BEh48qMc5FrqYRUHf8fg8k6umbRrx9D2KJX
y9VhmfCAdvjz9xBE4cZSi13ymb/RggAeDpnblrLT59pG6jlT3k+ELWvYi6AEZzFSe/UtYVw/mHOb
NVpD6RGHJsOQQCnAnDnzIsF2nHC35aN4vfMDjMWYR7g099x7Y21zsbU23aRY7HYb3hSiz0YsPXEM
oC9bWEzGE3h0faV698jGxGDLbTZnQS7BLH1sL/iQk51MurcriHn+YKx4r14ZTtWABy6oVT627U2A
udoU8Ms85ll+Dk5zPA9Z4gTb6uvuGFEpcVDcaBFcBtEs2Rgp574dLVr/8juu03cwyVNmglOtQyS/
mmYPOf450MIwCCfZdMYpoNfGr7qoxYR9yAFBm/cBu74LAsHvRUB/ht5H8Wh7DAHQ1PJBGbiihzJB
iUTbu4U5mtOc5OptGKvQ09ybnzIL9a7PxH8YSsHeIeHNqjaJbE8G14aAGp6QMUgvEwqMNdxFOikL
BsqsFlx0bwwmKMnwrciJfWqDHEaLoD1LGOF77d3+QhEquy+bpjlq2RHCaIMWabnVOFL097Ln3yWW
Fbm0pn6aH4/PDT/EYQRJTrJHV8WcezgM3bJKI8XXOdoND6+hLsnC7IGaXrN2o46e99GKtoUTdiaB
YD+YyW0JMFasdKi0bR/xM1GeMTTpLZOJvyjgzbJdD35AFALjPKou7pc1jyZUKIc8ILOdoSCS9AkN
f1ZVcfNXl5Y885AZ9NkLRepJ0lLorqlnV0wA92lmMBLiJjIUIrgw6qHxhQ1LS5Gk8z/V1Jsys9KN
+1jE/ikSviV7SF45q5XWIVvflJLx6XpPXEYKPIYVKwe3NITuLDtjzEQfocmMbMqRbzyFtd9iaKO0
qSPjwNU+wwCefLgLSGOXmtd8eOZoau1OQ4kp2kzbpT7dGQidO/dhwh7hkSS18LChz6Y6pwcZne9p
ZjXQ85083PLysj9HFRELUeFNQvdaKMbE90OmMbT0jFZsMC+Qr/kVgr3iAtX+i1VN51ECGcFOr64z
NVV12H9E2y0c4gTpsuyYqmAjGMzJAGhrskrchzxca8QS2QfPkwTaoNMt+ae5eyQl+t8CQ5T5W38X
5U391Ad4u20RmEdD7536k4DgO7ciA2xDcHsmMR9TVAHOQCVzsBfbssiGMvc/TnX/r23Wvy5st7L5
U/pigLvOqW0mEH5z380DKPQO6k0XWkImrhwScV59tJraTdTMo9+z6+Vm2qXhHgTEyKKSmHWZ4R2m
zoNks6s1aEKF+7fPFfmrWJEvDtncfUaOKkW0Wuy3yZpN++Im9+zetPvwOilTIYLrVEmPO7Z/urbs
dBCdloAdzh95vEumkt+5Q5x9XC347eXODQtcFfE0jpAVu1g7rzzkOxWtUxTHvEN06nd5XJxR8RTY
xJTXNx2vIn2QXm+55xzXmALixdd4r8OvJ9coBP/DV3VfNvm53DsUwRrSCA9h1b+jUDaQ+aWSdF/b
3VKBaJ4cEgYG16RADuosXgX7b1LPLqiYE8gEVEbTtdL+LeYZwbVSSFwYWqzWjp1PVjv/iZt1bjLM
OKNysZGDxin7fOQXsuUPpRf3ZvbtYszSjH1ZsS9F8pw3kB1WXvPAWNiSIjz6DsRHbPqsR4GEv5lp
NZH6olkCkKGBOUysegE/G4TXDjyNurNhMMIw9c1++19X0IbaYQ5KUJbtoPKfiIzhlwIKtwS3McfI
k7sRizaKFS6WNzLBYSFjpDjk1mBFV/SBiZv3Yf/DQIsIwgWfG5cqenFJugqAt1xCgByC9uzLq8Za
1YCqlVC0k2y1EpSyqkmq9fU8u55KiOljC0CM7GNyB96Ri4EO6mSsGVSP7nWIfvgQ3GV7eHOQ6EnW
JrU4qAESJqgKo4F0PW5nGBLV6tP7mo7R5xkFSAPnmB6hJXkgLbtOlZnARFRAUyjevYygtwemdpiY
Hr842gUHxNfPCGCht+rASl9jg9z94LjIgCR92vs0WL/xedQByJU0WrhWwJ5LKr0yWekZ95i9M3Gx
BPz4ARa6DdH5d+2FDlnbuHZAGX0GC7AH0wV0Ts+DVewveBEidQV8844fuLt3RQyxLDY93RBv8Ah4
kECdMZc1XT2Kw7kcD6uG2PcP4n4c8lKZp5kWjE2nN6DGFatQaoQqZK4cSR02iVFQGPa37p+HyEix
+yeXsU0jdW18VmSN9uVupi9YKewY4r1ojzyVl9kuTa/PPoKBpK6zZB7ARn3DId+yc2ZJvrEC5eR6
8vL2gEIGfG8P3pk+LmCyG5GP8KhjE0TRdGpXUc3ubYBvFvCDbKMBhpfO0m3NY1UZ4wou60pajgZc
evkZ964FEiDxScdH/e6BKwRNJ6Njg0UwodkQEPJKwMmRGaax/BCTfIp8RqAxuoJ+ba3chj+UTzyE
xExMEeved61hZXwzfS+ebSrZntXxkPrVPYdPwPeBM+vTgA80rMJfE71NQzZM1KzxrJopJORVa3C3
kxazcWv4IsAbYNSLi49bNohHfmIi9wusOMPjdEHRIZRrhdeRxHc6K0iXzKtzaBWLr7dfvilN2pM8
pSK04wx6HSuEChW10cnO72td3E1VkzLhMMOAL1wBJJfMxLENHYa2hbdmSbqn+Br/zVOWM7VJI7uR
FstySUNMv5NEFJbxIJxTEdUf4tH6zEDo8JwflAVikCc+w1SfHSEwf/yLmEdeERGfPAxgAnib7ZA4
H4fjvzWAJvQ5nO+oMZlxXtjP3O6kix9OTrgxZ0NwF+cXrWjj4o5kt7LJFJidgrmKdkI6XjE/k8zN
vsMAPuqRooIoDEug+GAbuR6Bh6rCrEwdiWIz1rcnZr7Bn/xeDipjLD5ggGhlSFsCC3EalXfx1Q1K
PNcyJVzR/arur0GYyLZG42oxgqYTpTqCG0iLvEXdxhKC0sU+2lkVTFLw+UfikDkjSbGO+CejjLj1
8tNFV8vfc8TtDNkVJBVQ3Ir62sCF8qgXdt95tDYVPZH0lEDyorEoSVK/zYk736+oCgbsgtDu5hyg
DFD10FlWwvRXer7QP/lNKk0SP9FhFSXsMGKCxEvuRpnNRRr+hHXc5ZNz0UUMbzbpnJUpA5Qaq6+/
9zS27DXgW0BeMRJUVda7U6CnA7hrtbTJfKqLJ4/l3gYDuFPy2pfzBU/Zq3cFSgBkhkSyWowOTmiQ
ngSFnpQ/pS8X7DuIQemFG9mkY5S4oy21/A5C145Z45tDOzASklGX965ugzF9mzSZZDeCKWijljnA
l0ZQoXjDY+lKJqvEb4CToj/mI7rN2ZVejN8ptdM3Bf3u2eSV2ZsTh4Kyf8Gv4EXVMlpfuFLmV9/3
/L1RK981cV7ucoIZqzHh9xhElXx/v9O+jtxyX9keJjU1HoxGesZyTJbkNvHLg9JC38J7wWJIIgLc
hQWkBf0nMxPmKjHHzK1Hs2dw/1acSwflQtV+LKn39pE3nrFQEb8APfptHscRjVKSroOGWKHUvI+k
S1e8M+0fwK9kZHowOmAAvqRR2ZhAWSRiTpmlHpNfX/8rdoVCYvOGRbcu8gpqFhrM3ffWpv4g35yk
K8BfPdHpB0FowHs+WcdfQDkb63BgbZ2FckYCQt9WYpkPjdVttbxLwkSWpiO25Q+0tBku41cdUIzE
BJsrHYFLqjtG/R9TfUg0jTQUiwynQKIBn37vbU+kmzNwGrVNSysJQcW9JafgEW6/FrUmRFMWbac4
w9pniyQbhllyYN2U6IRPeUYi51x5CZjST4I6E4mfJKh2iMNMv5eQ8Tvh34l3CS3yrPtsKEnDOg0J
je5eiANovVXwNKZXsw0iw5jKbTDS132ehdTPryhemgWfj3cx935stded9NF5HsDfNd2J1EYeQWbO
S6PEw2HcJAdXYRc0yZKZxEVol8xERrWBCyBExT6a7vSwsXAQOHeoJhZs7FHKS3UZTy7+QBFEHcMu
jtO488wrIfjY45TfG4pT1V3Yqo/+KhGbBd6f+2MQOR1pOZi1erMZ4DoNCMTJWVCdxeI7aMN7qP7R
od0lEtjUcpFbsbJ4UowNZLVxf4PFdKLb+NC2Vra3ofvfPEs6rtMSZX1ErOYzlUnchvsSDo3pvyag
wygSCouoinFgp6/ElukDCf3e2Ezm5I92mdomP/bRrbrZ1QTfohV8+J4h8kM5wEwam/zwPd0VQabW
j6g4nTkzoAfIafvQ2IH46V20sE+5bxH/VoySmac0x6obWlC07aUk5+NCWe6W92bxmc1ZUmaITePs
BgJb41wIvbqB90HCb/IKp1G9iT5z3GouMh88hjElqyf2YIuCmPcZjzRsgPJQvhBe1CWq8vRT58Pu
kxnLalC62uushVtMNpjLCBoxoJ11W5NTdOEuBR9ict0M90BIJ3+ZLfxZMv0tJkBAixtyg4Xq9YSa
UQp/1H/8sTjHNf6r3p230/o6N5S9WUG5TagormtuyPqsO8l0oVXQrqBZRA4j1rA6YyX0WRSJ0qf2
hy98W0tTyMMj4dL/5enZTsy1FrQ11AOTJoK9L27/kPedleL9f+RM0XAgySbN4lkeO7DRnb0BuFkR
a9Ui5EU29z7QqANYQ+deyzFscfH9kbcWc8+8Y8gJBZYBvgsEi/DdQ62j8FLI4xZyEjMz3dbrUeDQ
RlRfApvaNIgAY+U4b/KUJHqaRDtMvQwi9NCuRsmU5LZzsejfXbmZnOJnRUUn/msUyw6RaHh+joci
WMB66pwhAoDsMbKsWlto4PxhFqRzEav9ZzyOS9kSen9+tJJWJUbRFqTcxcFpvckdDQ0GOPXtnVs3
aO2PJyrSb2pyUUgzJGr1uqAshmvAq96efGeApmJPgyCSwF+UzUTxZf1ZE5Yl9m9uZIddPbiWQMX3
kjFSo9gF9VPjtncFhbHF/V9F9rM5ps+1yuMJXRF3UCvCqTwEmQrzE7xD0LI4TJ+quBP7FwDWxIov
GvLG2AWI8091IygU7XFyA/FqU1hVtEmu6vP2pAm/yrUOs66w/CojTarH4W2o8ZpafuVNYGJFQNv/
cVFy3hHHpSsVZbItnE3Mi2byqz26KahlFMcabsSC8uoCGiRIwd3aSy7+Mz9EeOGM4LvsWcIkELhH
4reGwDRXEr38Y5ewedwo+NiEg2pDl2XkIAuaL+H1UXjwnrTG0zeNwxdlBu+e3g+ckR/uDBw3WCEa
1RGvEqa10ysQ4HYi/T5j1lU6RErtafsJjt3OlFWU7BMdQiBRqZoTbHTTO8/aI3WZMwK9GcSEWdn1
YXcCPZkVHhtOKxpO7JaB2xoK019YDOPTEVmY4dX3OHf2Qn77eRg2/P32UFKUqqhqOQBslc7GDuRb
tRMiZuxzp56BdTzyLHxgGDxMcyitrvMz714MXbJsLZUOSt8LMX+DydpekIF1+N7dZzS4qCahw5t0
shWiFnV/FswaqBs4Yv7GbP9HZf5FAzmwzrrLgeyGBn2Q7ouDsCyoRYKxKre5uO1hroETqmNRrlAv
94SvWNUio+ynrG1oMNRYSLAOa9OleOrDtI73vzscOeMZpWrfdOOFh38YfXpMlQu/htaT6d3vh4YE
EzvOx29zg5Y6e3NwHJJBcdy5lRMbayk/NjWcPHoMRCFO/bYNuo88BTccuWm/aPi2Dsfaas83nX85
eBvP5XgzPuVNHbMc8GilSrf/2Uk5zuLD2nr4WQ8tUyhsfq4rcIgTwYYj2u2VX68gSOwEb1ADEGyc
qD/qIouO1uDBdtEQ+Mmdxumaaj8wovW4O6bZHirfuVAu/rmuEtsf2bmoA566M7Avo4hKKvi7hS80
mbtBlMQB16vq5c4vt5/aXOVOh30Cdyb8vF9O8QUft+JzPCbebVcXVNAbg09pIX8RHj8ghv5hLjY5
Bref0XsTNxwjCqax5MnySeD17tKvsfYeGvaOEGTg0duk/OZ/dR4ogZtTImXb2IyCMWF0oXicXUn9
8Jx0VCacy63vts3/j5gxJyvWCsHlXNuYKvoxVaF48anxCT9J7v6MdfwE9zgSZpTt+RQQLSI538er
0L6Snen4uvET9+We/6gCfJnG7EJNIKkRo0SBkZyQxZrrtMk9aj1MkwWF73J8wgAqVuNOKcoYDIrV
zfq3qxkNBz6DMAEEi9UY3ndLvHJRuyOPARerZdCaGCbBw0Gp2M3VS98rIOVa1gB20d+0eo+GkkOS
nBD3TSP10kTmKcZDfWABIy3nI81aLQqA/b3xIvjponQ9wbmM9yyvF6GrJroVhqsVX2KLs2MM5CE9
OWruGFwEksz7eS0MXOqNa3xW5uPTzzHOHdtjL1XfxsWl/UOnFDZXElqtSBaf+HoUezF0dT/3n8dT
ebMfHh/6Uh4PGybh4iwwCyBlS6UZbAAzSLyWWHnhupuArNIDhQAwY9OtkIk94UhuiJhWd+Rl15po
gjDmR5trJVX9XB1X93KfZi04ThLUYYSmB1DgXTxVY3cOlMazWDEdW6GWzPMTERUqks4MaAuMUdx5
y/wszQsmUvv8vj90fPWRVr9vaAUfezxSrsbbg6cytY+SnAWtvYdsPpoQ0jataMm1c3MCiNHwG3Rp
0zwNBimZgMjODq2kIX2x5KjGp1wFCFT/U5qe5qTiDEKz/4muLp4OofRKALyC5kEL0kiwFghOjM86
gBRr8Ipw89Wm+VAU2isJLjXbBAZRkC1A5o/PZzPGySj61SnrKDN03DF9MoxYjEpnv1usKaw88byx
PZdL3DDjcd9nUcAqg7+1oU3Ff8OZbGM/LnZnTiGaaHAQN30ADFQ5y4G7oMvrkvGmsjHZbrLSXZMx
NACNCvQ417DMzEadgApWWsoJh5EFygA0jFppi5SRSwvhCwBHcyuc7a1RJp5jMb8a/NMKZtixgiy9
6r7R+Uh5VDijlKlPe57HQX9IXwJgPDqtK4BzqYC83Y0LybmgnoTLpO3tTvoFHK3Um5btS07kEgn5
8+Imlg3bEepQET3Eu854zTVj38SZLmwlieSw/AprpmcK/F1U0ERAWBqLoIDUerOVVMs8tWbXMl4R
TgpWC4yWn3nTCDSisB8X9nnJXpWizJ9OKf0W8D1SHj5wjYSh4vZDADbs2oR/+ZSReuBabwkL86wV
iFBIuhkNqWAd6enqv1SsCvT/kZTJ2/ovImhWqgoe1yhHQnKEZKK6gaSfYmPM9Ftvavm1wDtUNWee
Cctu0RxUBIO8XBeT+DDwP6a49Daw2q83q17McNzWnub5Osetb0f0XMjZmPqCDRgwi093l5ONi9ej
fJaH8Ay/cwl31ifOcj7Iman8a9gdlBf8kYI8l2ZvIoOf04MquyGJKLvdVpWCyG59QJBLXfPhwAsJ
f0/74A7rlEli5IVy+/kvRqFcUysAT2ONhKF/YJeK7LIhxz7yfkpdDgT+X9wvdIEiZneSprUpMG34
S6rGG0hFcFnEssd2N6ccjwn+BOXOAosMidEpemtJjvLaw8QMuq9LvabGo6uvhwNbp+aqX5GE88pc
DCvrWT4sCk3m1icZYfHRhl/j93pjOiUlHa5+3ptjCCN4f0Eigo5mA9dIpbjDydBB7sKGTcQGQ7OR
/EsgjaW5Px3n1tzKIxO13OzWU4dmRTUpHCKUVbnsvcYZyNPPF7a5JocQQpofX86im95dj4cqbMXJ
WdgJngW7gJRXSwRHTWDMYU7rnl43VWfNXZd6TBoyrGfYz0rzDHw+b0+UcXsUPQiJC7lLk18M40vC
OOBvbOiujzOPOnRodF0vA0S8IVpKSUMzc6ouwQoN266X6I8TGEXVMJxg8Hyx8mUnHdbTZ0CEfCdM
D8lrk1LA4pE6eiU+gfV+k+6QusU/Kt1sJVeW+4D6fXuEjfNkb/7WrpQAAAjtzYJR9IruDVQvBKf1
h0iDbKEKhGwjo/KTho9aKR4Zq6Og4ubD9KYHXNGKUTDiNIjZ5OXR/FbWlMQr6iLKtK8+NDsZoz8Q
Af7Sz7rUYF7Z2V4AGdGJmdqKTt63gj45XG3RAnaT9FGLw5RtQDcyQjkcHZWg706dkymxFcVSEgAh
i2ZwlYlfKFvOPdYdseDPfdZ+/TNi9ThYXnmHAQ1ib5X/qJxXBL+AV07WLIC3WFdFIOD8JiVTpPxf
FaHuc+D0kfsmLvjkO5l1fLM//d5ZLtN7PQy0ihEB26165YSjZ80Hr7/RLCuAc3YEGuixSdSVJVGg
8ck0aoQM/H4YQDuKwi7vmMUMtUwG9NTdE8HfGjdwuCbJLNoET0tQYwgNsOpxg/0l5JkOd3pPGwms
flTMWYwECc9Cmf2ZagiMibeke4qTx8TvtizGuJNWX+wirE38m3C+eJkWbOVVuG+oln7+MNpXYlTc
gy6JyljIMxXObH6S2ifq2vN18o3DyIW8NCYXZv9qUD6L2IfhwHVuyx2RC6rxTBl4YuqNuugFqzx8
AInMgILhYVurEzvTfz0L5y+vfEhomAjrWIdUmmsM6UXrbIIwMiWOcHWi0R4hM0ImdSnoGEQP9hp+
/wMdSSCdbiXcmbK9XYpGqSAgCN6e2NL0DVwhPSe59oGREajkZNQntMBvc+GVWFai+Ez0pOTKLnkO
cxdsLxd4rlFZ1USQR08yPESIyiEiaOZIYJ64b4Lzo2LcUW0+GEjLt94cCH8VeViQTMpcJi9NN8Et
fMc9eH4CHTVyeoWFxMdPnoQDhzqjCKPXJA2gELqs5INb1yilN8qQ7p6onWGavsw00qmk863okR+u
luTveSyeaUAVLuZ+83Rekw9huNAHpkaZlo3BWSEEVhDBEiLYFilol06RJZwDvMNxL3ZCDMp1Vjvn
zPTsi5/0j1BkEmfiqLLdCyn2MtJEioSfC2qcuE62swhZVI0K12r1jWLLURH8nZUnG+VG8x/cPYli
yb3Lr9Kcc4QQKOMz9vQwkGhzRVOx6CD4nQl0hOD5++oPchsEqMGoe5kAYNSefs8OZxewhBfuNmyn
Ze0sJMrGNAtaA73v4HJUusZEIZFDqN83InFg90pwgMDtZtmBx4USmhGVNkcRwYt93XyeNSweUqKV
ebSmlnF2dk1OrqULc3CiQ05Lica8lb6oy87wEDUGncAKPIfi0Puki6rtypLN/GvFDGuRDepHQMP9
b1y3s75e0aDF9nx0e1FARHuc68AN4SnDquqgHMRVGKDwwLpDdX/HUBL59scQTHiciK+4XywWeYTx
RQAF01NUB1LOqphgWOsMgQGYenkXFOjtwK0i1CmJy2IVEo+AsimxV97WtUBh1+YZaKUs5YsvQ3Wg
XvOOegzJVWj4TKSLBQLsre4YAQ1/KBxNjQTPyHbkjKZFSYsQ96MT+TpC2u2Q1s0qsfT3u9pe1/Mo
rhqVltjwVyoqF0/eFIIYP44FWvcwA74HZYu13zmIdskNzpZYrO4DrYXO9DSuLyWPQkdR74VK4FgX
5o4Yg1Bp1tuqkxHG5MEOFxHua3pu0Pl2H6ObfW6OqPBnBEDX747lgPCJeFDIhUDTZFBf/RkS7CpV
p7K9dZ3lMXFNUmJKcWO+/IjcZLEuo1bnRa2ZeZ7/GSVcGZoVTFBxsMyrP5FeuQTqy7Qpy9bqq8wn
rGs+NRjRL1CVaq6drkSVq73pL1ztnh5OAmVnv6wNEc1Qo6rPXcJbikMQUuxPT0Sophsc3M+yrCp9
P/QewG+EcdZHxBtAXvvnlk3i1ObZiQpBrhvqQ4Vacdul+S0scHtoR0y9OcZsQnbo0xhG53uLTQke
HZkghzZqj+ijCLMjqUHuA8VJwqPGi9cOD1VhpY/Fl2u7toDof4ZFR+ED+kEbRtAordOJBx59WqzV
J+5CqdnXJG05/27c1yZAmOp3KQniCJkb7YmPT/EAdNIaXzRhHFZ0h4a3Mzc6c9Jql8FPcNl9pXoX
aHe+/bq1AR7SCcFJ2W1dkZ5s7faCYd5TSfFc+0rwtok629909RoBVx/MUEvysDGd00Dow1zsrsaN
20uTdg2CPDkn9kaowfBjgcW+3PtqLUlrBzyFCANKhk69BJg4F56yf8V3LySjvBQg7Cl/Gr+np4Lt
f+M8hLFXvSaau/2Oi115H0EF7X5tY9sxQAWSqbe1ErFE2VuoCMKhXH/8Ae74KkNlAIoCGu+SD0NV
Py/DyX5vcSLRa91773eCIrEAQVaHozOFHovdW2chQnKWU6WZrvXUHsbE507owKHkU6xFsFTlvBjg
xnpet5fkgFdn2EhA1OxunfIkcMEl8plZEWdqG/3lpjyhPGGy0Vov3uGkt1/TqmWNW5ZmoZ5Z9TD4
nDNa7gX9UJXQzsOrz1siBC3NKnRIYLrvS7icD8zGjzRkynM3mbkZ3ZEOtIg6+vGTnd/Hz7NMJlGx
bQrzjTDe11HO7VS6qbHm81pDOPXTpTTIKsrjMxCtqDnjZPGbzNYjpljOfbaKZMr66Pjx+ViINC5d
LZ8ZcnRslNdwWcUXAinT80P7JLKWeneytJJVEZWmk2qqnRKQDHEDvwSWSYSlorj1DTN9/0MJSypJ
56yNqKl5LiljYz+WTJt5KpvRg+YgizMFG44sfFRLUk2P23n3P6UIZPsMavG52HhID6S4Yjd7YxxA
L9sgIsmnVuKK+yMAMgs0O1QG5wWJQgI/gw6bF8VBuhr7DkdmotPTPQ5AkLVxvrgBcV8NNPPWlmvC
z6N32F7G+oQOwSTVMOAd7a9xr389JphAbwWBDqUKA3IaJIyu6GpWXUuDOLmwVq6aagNINeFTinpM
6KVeO7TkUjV2W3NLdPnDQVIfD3yjzr8T/D3uMUn4zRWVfrHgFXt0dRq+aeCF7rFV1WnUwDxyTTb0
9AgS+w967qFZkkwYenvzKbyRT464Qzn+lVcPKzJzMMXl7lvNy2N6IGUyFoAiRiWU+O0Ii9G3FKLw
/aJz5Z4pPNdIbdwm2bDkavIQjow/vTVRZui57Jnn2aWudizeOgE6bYC00UV/qmYp3anFTUNv4Nt1
cFaxJXElb+SW3OvclNUporS9GPQAddHYPcTj0fA5T/T08joEE5x3ELlbB+gm9mnO9D0vVSMrue5b
EuQJ9z58uHAE4dMZNJeUuRfF3WD8vr0y47ji29hJzsw41SEmd0t1VuPwXKGSUDpljNHfBuIjB1K0
/9MhXiLybAYniKxPF51keCyMwjXUoRTRQIvdI2cqMfg41cl6aF4QYOBPU0SkwWqQ59eNu8yphJ3L
fuNYqhHI+uBqak38yMWRDh/yzgR0uLZ2oESmLGdV+Kbv35xSwwzzDhrLI9sAjaNFKIXgEa+E8JI/
DjtVI3+ZMqIFYFmg6Ge77b5G30HcPN3lTEhIinGE74YYV5cJYMVKio/bT+c6V7EdC0ym5YLbV+sG
xnVHm8SlZ5/+6RxpWyU5PA5DxhLtX6xI8FfUR3VNw80icX+zvxg/5ZFFALJ4thDvRrAnRaj25Gku
9tQsiNSfxbbv1JlcC/LvwyKLVy0Vuuo7lLttD+ASBgvg94X0oJkTFQNlLv7x+LMQSyzcgTEH1FAq
3CQGpPI47jJKTlz67RK4krMVH9SKeaxBDc+/qx6OrEz/7Of/GVztGA+A/uVtOXmGSF1ZQHfRh16r
T/CByOKjlXDa2PXgnG0USImEAie46qytsCvIRh7uQgyPdMrtyS7oT9Iv4D8rjTH8bwq6z6bdTZLI
+Bu4CRpmjdLQ/JvBjMGV62+xfKxhcDXDL8D3S7/zwvN73g6Nuj7DbsvR5jH1zdnQQa3LiyyzpWe7
BOIjTce/gDHJRhwdOI9hupGUjl3TXQW8P3UCHSbLyL61KQC/w3PUNHKsxQn5bt4XckRTViLriMkC
S3y68GquvgaLlJ9ugapD/mnPHRQvp782LJSEHt0hL4y7A7vVajTT4cBtpQSWueEzTsuLKrK5VVcx
KYcv/bLMW1eHfGaauwWVzcSagupxpsj7M54o85Z9ZpkQp8gEJeP5D+Y9nSUJxmAX1J+L0vIhKxgd
2z6qxp1qig3HcMMxFDXoiagGUr6wFXmuz50bi4ODB56lrxmTzJdeMbJrQ2vwT5ru/cvOoc7MFGhX
bYBYBT4gTRM4Qff5kj4Ya6N5K39lT/bSAVCoOz1iveoHu2FTLe8Ehduv5leFqGEyb/25sju5Jk0x
+SYFboFT82Dx2nJmhXdjZ/XWH7VLK/lE00o2fNTUDcvtOMmKuENjvaKKdnovtvRk2JyaOF0xWyIB
CW15kAU5WM7MG7aIcKS6o3IdH7qQJtsHk7su9OYcRY5HOZOCZmbI1vkYNhajuvRHPDo6wll0e5bH
sD+MYVif1BM8rzwJYItWKPKu/8yoWMA2k+M6Z7D1idRCN0o3lCZe5WuNXItKbV7+X8HfF5cNoGuL
xBj3SDGyhlc2/WLa0ShE5gKGeIqBg1PSFLtzwm9neqoO01rGZm1av/Vw67/ua/tAcrikBKBANQTP
4zcRhLu1jPCzyYva4+I79gYBTQ0s0p4AXywd1UgwXuFd++zt/O5nlfZUk1RDk7XgJrkBQS1qtTOJ
8G6Rp3XSNaYNbWC4cVX/5Fp9+iODSP0QjrwYdKtlVq+nvKjhTrBcMyNRhljaZA65PdblvkQyM8yF
2nb1XQ85Lcm+9EBi9QihxeEhYgvSCMDAbngJ32pZ9jHzSG4aJzuY+PH+orq4S2dKEKoVxi+RK3dY
NZkmnHcQ3nn8nrW2jfEi15Sawoui873MiWHu3YybBFxjD3s5GDdRXQyC03t8jbhIvVRu/Rw02Wn2
NRWGyc72/J7p6tj35L6THsUmbk9TNo1imEIRfETAsiokRhefbsAYst8u3052bJUSWjsV3yw3IAz7
n/X53PMegejcpFlfV8JPEea0LHP2BRnx37nMSxn2URv0AZbxCOpQs7nPpXBn/6NmU/cY6vzz4LGI
Ru/iH2nIYIuWxsWHdW9kaR3YBKyqBNiAKyJb3dL6JguVmYE8/FGDSbfeCkW2B0+5ekvcgya2Zyux
fmdXfcmFRLOF9TSAaq1Qb7I1e66J8ei7sEJR0RO5Oxa+NRdU/mzjxZqpaNG8aq1YkZRfk/XKoHIm
tEU03BDuwao8b7yTP+/ZyXVxVSOzw+l5iImkjAHU15An08IJYWVZr8p6x+3IUqnOq/GWJNr8EJcf
5pj4XOzwCRtXyUN/KD0MP33jSkyxaN+Y3zKI/AwTYJbsBndqXWzda9kJfNpfXnVnyPIeM3XkhQXa
skx8Ri4BpvS9jfMPAwTNcvIXPs7sijyCQAhkrKiwznLoy9eVhAnnvfPsGkCn69crVPpkjBB284Wx
EWBAsB2xPiXJBMdEb6MF31knqVwFVtu5HPTlCLhyCb/EJVgUXqePTrfwN2JwtvqVIL1gZ+rMtsY+
nxy0B4fsCpx0cUi9djPeUx5V9zETtzv0EbYUy3RiwAyIYLSDe395vUzmdAcEz2uEJiGGMMCOw5pY
NM85jN9njexNNnSczJ/0Km/J5Jy3VmHFlOUBhTzBpKaxbWv4z0wxz2Pt4GoJa3VS3pqgzJtwzKJp
wmkzzBSlKoc/dC8PXUnUTuwtjVR2NwIlV5PBDVJ8HqZLykeck9Vu0SK2fd356RMRd1KUasw/S03Q
UqRuFdL8EiXdqPO7POEdgNlLpHwXxOSvizqiW5ILQzkBtp/mc13cGpMbXEOB8/iUJAXND4g0ncoE
i1agIknXV+f6NURXJUs3XttiGcY6GKMRFNrtSbSriVKCIoeroFyo8Xu1hD6wvmsspUEcbc8ea9n9
446MbC8YwkReePZXCSVVNFVbDKapjhWAJ41D3bE+ofnq0J81I8jsRWhfBGkSB4qgOMeW/CBGSfHv
7HhxcksOalfaC4yjoOkZxaDR1zzXXQ8v/ckjRnk9Bf2+jErqq/BVwSQzEZIZGSaq3F1DHtw4Wggw
MREKWtw0/71eej2B/Oyj9uuh5DqqmB0ad0eG71AJFuu1IQMQhIBzw/girrFGYJ9g4PtFcn+FFZzR
eMedidgbFnSmwpXdBddBFa39RM38adJZBEr61hihy5R0AqTdhBdd7mLoMYsbZIB8oup0WbarwH+G
MuvQgb/vP3h3rai4RGfklIFcb/msFM64wbqOfRxcbQl/W77sjLnyD8+KEz4VDIk6uKbm5IUeX4Wm
pYHD8ioD0qnjprEE4cB5lgKR/3MjmGXqgMiCqoJT1iY+PCJtHrr4jdc1yQXfzF8w/xVDARYpIYDG
YtCkK2N+6dIOKSb4zG+FIqGpzLRh3tOe94Nq8/hDbY22OfJ8Aejf+A5gnll4O+ViXCSkDFn5xa/h
661jviS+t8wp3/pEW+tnimq7tGHZHqpP50x9DNkvK0IazFEP6kKeBMYwG45tu8qQ7gTkPx6pgCyI
8uRHTG3oyXysRRBn/EMaJ2GhVLPxxVxh5OJycgyTtuOs/P0WURGBYypbhs3TdL87dhsrAccW8oh1
0fCd50qGNHzfpjHtSdMIHeoc/0aWWlZHNxV4M91NZazjZapEQx932T1iWYjIxmlXVSFkT7pH2dpo
gXIb1eSrcqBrJjeKnjAEanQk7CSQcV9o/U5aJHsTLXbOz9M5YcEdGBBCMJI+LOKOoE4nxI6LSxxC
DoXnV0eeuFUTZOwAOpDA6Kbc8vRA/GrSYbqwTaVvAiiH0l2SrS86QEDspsvDQFaHG4y4FCy0tKal
Nu9EE03PHSnV0fK6l4ofU+435aR7SRlay3GwJgHAmClQV821HPNBa+K8DzoDZ4+Stid9kFlC2c5q
FRXMcVXf1sA4mlRtVpd77cw6s6I9f7RZtMi+hmpW/JaDcUMTziUxrfMO6nIhMj297x773F4KXFjO
hEMMra7LR89TXzYXcp4fH44mGribIrG9P9LEk/eW5/pu9E3JG1ygLvhtYdasTNhKA0FFHFGmf6le
zlFI6dg5I2MJI5VOWdJ+esER/TuYfgvaRfztwlVsvMaBxkj1YLvOIPukU1TVzUFbf5zFP15UN3yC
/xjvKm7M3k7j7eCh/WEbtO9xRO0fydGk6S17/pOQkeYRKc0dyjHCXGPX0NnmOFQU5KISFRzrh1rz
uciZIP8JK2vM7Fp2mJQ7K61Z9sxU5IIqlMDdmBXBs1cVfxuqp2KSWxoKFondcFCB79a1yBDPzEdg
uyhEA5yLdkZYNBwDLXiFfUBLeAaKdFeTxtsSIRN2yFkcoefWKCe8m1dWKgfv+g7vGp/q047DCCM3
aiMvxKx+d6okiKkNIVZe9/F2TJGExHt4cf+NfMAiMW14XyXUHEmdMR9cLTPSOof4NdVVFEe3iX+x
pgPJPN0NZ49tGhjaGuG4Q1L5wDTZLm9oULzii9Xdbude490VAza0jHVhfIZDqhRpUXm3NoYNy5qf
zfZgs7JHfFqzC5p6L+XXnMdPVVZudvUrR1wGnoYqPs8WgQ7Tv/wIiAvc20XvAE7rVKaBoTIfMV3M
NL5EFYgdrTaCjS1nTJNIPP6O1S8oj/LicTJOgUQs8oz74jcvuiV7QB/pWoKtnRpAn1E//i2/sU21
Lr6vdnGulvpuYI/t+XSCtd9U4W+WNzfsd2Oo/9oCCYVNIHHfxx2G9vatSfwIYDRqG+QQ+l4VYC8V
KDPn5vDdm641a+BAWcr9W1EC8r2bCqkNyTUg+gVDidpDVGdhf9/rai4exgURort//VF29WLt+TiC
c5fXMM3HVrGDOTh9KKJ4QJ7ehJeMH8OezMWiL43ZXBPtv/ciVYuCdE1FDTV0NNduqWXIA8m4auYb
8wrAvnBt/wNGiD5yAsW06DucND3lsHJD+JZ7p3GYmWYH5pg/lc0PrV/cSMgdXhLfDWWP8YdsZxYc
9e/+q2kCLjE3iPX8Ogb4gI5g6x8PwUipPJJS3oD1fA4qFcmq+g231/0efBiabVJrEzmNdEow/gqc
lSwRlSMih2lchLTNLfJCyanOS6o7gdibKu3II/b19B9+2++FKNKy3iSMC5yoTL8D2PYxgow8TLlI
q4kA7WQfy6cecKkkf+nWXIm70teWaANYWZ0jMpLXYts4RusicDwdOEPZeGg9nQiAVyzEvTe54pi3
h7+TFwbx+V6gOWoQxh3m9kt4kjDvqndEev0MJQ6bdnm4O/TgJuofOGGWY3YT+vJu2uyWyvxtXyQ0
8UThe8Pq5D1FB/SOsCKjRXgc3Yo2wu7PgIrm7WYofqICzRpes+9vKMjkes4QevcBnr6+5pYJ+DI+
kcBRQXkwmbQ2/NCgubdi4bVNUhiipFSCSyqNFNiEkvp39ksGSq9Xl/hLFk5d1bm/ZRdNZf+3JL6E
ekYDWRUg2e3p/2r+g3agmNm8bBjIaQL310B+dXfN4S5IIGqO5qqZt8VKuI2MsvtA3/gL6cKv8Qaf
jtLWI6AsVob5EcVLqZGgLQxQ4yLKodOTTPbtu5g2guBMM7/J4mDAlnIFGODUbACDcbck+icRlP4/
t63MquLzI8pc+8COVt7dCSOF9bQKCFO9lIyhKrnooaRKbyXntXzrKv1Q4pEN8CXhc68+lu5GuIkC
bb/jOCoZcwytSXIBxt+02JAVcFMFrULNCH+91YM62HeaSFzpiFdY8cKS7cWVn13GTPXjS/B73G3g
p2fKVbWfOuW4qqmOGojdXQpmnFVCRh1MigWH360ZTP5pOsNtEq5HMk19aYYXEBcPfkQWh2FXCvr4
D957Oznw24B5t/hOH+6rdHvnuvRSMfsyu3mKu6md/ZEXi9EhSJSdYL4KkjNelWWOr8vu3siQRHTX
I9Kjz99GyCDkStSJfx42a3MZJOEx2GuR8d8hSnrlngxTjYpsqjbQbDXVvO1mc5kuG33t9XGbMgKV
Tc9HqkFrPVhmwOlnGrHPBi6bi3wn7vDRmJLT7U3Z2Nb7SN4vkLB+8Ux1uChiHZyGCErDGaZPfNW+
gQn83UX41j7Y4q61Py0xj1egVGbAjRW7qY4UrnW3KspiBmxZRPlI1CvW4uKfYn7KEQWum/2EGzfw
/2sNFHn1xAhfbwI3qitfGloahP1PcOqS9X4DKuNeaMVP0mWDUi2P5kE7u8pCnflkNWm8us1pDVPN
gsNLhqZCQV6p9ZGk4UCDlqOLWuzqF3tjvqCyG8zNju8tPXxBSogYzz/o250aUlZsFwx5rWeeQ4cc
0KMWYStxx6gc2j+fyGNuviaepWWeFvif+EjWdxGw4LAHIXLStBdSYI+LjKJRXFvcWfXSUi3rGj1+
fml/prILtNhIk0A8UtrsW97T6ST3NuyNbuM6TA3MxhBIpICOaSQT9wywpWYXLEwltdVwGbrtCoC3
AuOgzanWHe/YAVHRqhNd7ao+yDtdmRSH1YSoAF3Rt8AMo65uwq6+wqmb5Pn/7ln9CLCQMmdAnW9w
jYCWF6f8dsJnNqIe892rubcpW6QKgK2vdh7d0VyrLuFM7lermsR3550UM/qwajWc2e6qvZ4kzywt
aajxspL5QvraJvuDxMFX2rIGKKMIRP66HKfkJ/PeTiJzVIus0d1bGUUm+wozwbr3Lsikv+k8IR/X
f+cY3hmlN5MEZgP1+lec5lhfeuQtBTo5I4mOu2Cr9H5at6V1dbKi9JdaRs3d5VEyKQF5CDeSnGbY
/6RDIwqzUSfW1LOP3vvsTBdJ/hi6RAHmAjQohW7+z43KpeVr/zId0d9jNXkvjwL5sYb4P94p+E+y
xOUufU8SOuiRCN+I9Wy4pSaEyAsWW2XOAjC48vPQPC4utpZl4Oa5sqZrMbH+9CFXorsOisYTQav1
P610lQnX9yqZib9N3NG9+zhTZgx3Q/7ESsrZj1GpKCp4kOV0WJx/TD/jEIESRFJC0H5drQBO/qEp
82PS4kxY6IvnlMhbWxGhsUBpt+e46Z1PfsrSx++lu7xAiXZixA2CJGkO/VmvgGE5aB/PmeaZ2hLg
ah/rvhw4aPl7+e/0JovHdx+zfmkzmHJmR3kZJV+Vdoge/FChMN/kDHMqFCDJIgh+LTtGeeEpo/Uj
vZr7vUzLlMRMbdQdgcDHdxZrl085dDBt5nGHrXvXsyjwxXiH2io1tJZ8R2YHc4Yhe/gTws31tioo
tXbtlHJ9K99RS6k08syZDkbpk4Lb19d/FO2CUkD6BYKwsp0aKjdESzIjKS1i5uzBi2CMfv8hbaST
QipbPsIdR0Pdtu5LxsROT+HvCj0Pr2Cx4rTiu7uepL4T+a1WbHUFzUjGMtYImJJtn9oBpnSxNqd+
bxWlowrkWljbmJzG/vTa8eLB9KZKGXdqnS/Y9DrNgPL57t7jj0sNqRBn9SBrcJLHsR8hE8VzM2Wg
ricWq6SEyQUX7U2d84a38Ja3kGcakNsUIy9WCnddYa9SNu2wrWZad9Kb4UR09Gvc6ALtn0JK+npG
jcSfsLtP7RWBp3s6+mr62CgtvXzULjIMUAshJcAkqr2f+AmLcFnB/21kZSs4WAvg4UrPtY6YtFJX
f/HHfBAJCi2VCWUYW0y55iVvNjG3Ctn7RpXF4nOO9CcyL8U8Nuh5zTxXvUiOb6cuOsxb39JRf4RM
UzVkcOLoMrgpxB/BRWVr5S3mNRwG+omr2Sg2vIwaLTq1+Pz1NrprByk+D1+/QnTd615erxLGhVrh
TfYtHwrdnftax2MwhN5W6MHf0Q/skQi9PxeRHe+0SPhYW6z7tYI4GwLAeaf9LUcg6qS6ZIEJEEtw
jwYPDbJjaWEHrkA1AbUgmKBhaOlQv0l55RNvWo/zyUiznzEC2ZMvlkkFS7kzvUssUgqRpQFkDVaw
P6bTKYqCegTLyQDNP93/JE8FdtKS8R7KNj5QU02dmULwalb/y3t52AU5+OOwGVz7WIgQQsHIbCqc
n/vzEKJ/wYSMotROpvPGqUjHv4uW1zLQad8DhDHluRVi5NccJw1egWcwEtOr19cqVP2uVuQL1vN0
k01jzD1feH485BGcdTVg8hg7IqKiZl2IAYy1I15WQgrn69x4UX/CLG4lfMLUsFdmAbeNsBUlifk+
R8YLEkTyd7ZdCocBJUSb1EvwwvIHHFmadqfbArlo9dH2tjTpGgiG94crPc49xHVH6V6cZI0V0bc9
PXG3X5WHwIheuJmSZkR42sluyu7EQGaodY22n0jkjV9tlIDRq6Egej78chx5+Dg+WI2y9W9BQDXw
YiNyH0dqr89ppzIPpAuY4rkuhEDSNkpm8TOyDY8IUbMDrPBSKzhd3UmbCMrtg4yge4+pbbkoxNwW
Akico+GFDHXc6N8Y8NVVoH1JCSYiIOZPj1F1skeeUQzHc93hSamGQLg+XqfbmfH+5XGP5clmn7W1
jKr4mM5B13gZPvFt90GwjgwbwGUc2jLj2I+4ia078u5ALW6XBcsav4ENff2fSJjYv5nCPHQ6vXnu
19May+sYqlecW0m4TWvdc8Or4iMKlXjvWfxaKdARrNN9oKJbbf5q+pjBdnDh3QOsA4eHGAmydTSK
rrr+dVScKGTsK7Rl7/AwXPFgj0erMdkeW4nZ6U22CMmZlrLEihd3/U+GmmJ0XtX1I8JOD++S87jS
kThSfTXSISWPg4hr4pBAIYkyhTia2QMVk6IN8vDfsfuiF+USuRp/pQ9XxKVoFgvhlzn4MMUpuN1U
FUyU1yBHUAydQujUuvjgVLHYgpo1JEvGYJatiAvLqxVBskMJCS4FzQwiNYyb6fpb6Ql5XDpC0Xfi
DGN5JLf/qB3RUafYGYLmlOIV5jk0+gXEPRhEv7lJjA8XuIdV+luLn3l6heABnrAo8dT9OdwpckdF
C7ywpct0e0KUN2xgt9L0Ko0PNbJY2r+0A5GDOekKo3USBcrNDGbMNIc09cNGXlQ4eJBUxNW8zD4+
3Mb6gi0Nx0m5YprmI5rDGNmm38oxOH4KtB1fLeY2xENxut/1tEcY1VmOVEhT6KIPXdS1dCPopPeZ
vRgFVNVWj/CeiutAe58A3dRc0hj+/ZC0HB+PVCU5GQZHhokmLdMgcvCRVIGUo0GeHeCm3wUuDGkM
M/0enAiIgFLrywiqO/AVPfAoL8asMAMMpwS4PiXz9FyXP9A8irOI/gMih+dqsbaAp7n5HV9NhwA8
Ag9a8DBPOYt94uGpQo+0wI4+iWCd4knJPAHQq05dpIe66e5/Juldlpif4ZXwk/Ohi2RYgXxoytjN
lMLaUNprlOdJQLTuPxuFFk8Mi3DjMCBnblrQtIAzmqCvvqqclwSveRhv33UtpAAVlIv5p6mZRGbM
LtEducu0rkAxP+YXrild6d4AGL3B4MF0WHtC4dqR/K9el10SNZnhqBtL1cn50ibZvN1A76avdw1f
EuCHOqqcZ70zFtI85ZJEWGfWNU79zfxsJtGSuWP5tM9cVnZEH9lMKkr70UbYBXrvkU2eGYWvtYj2
8GB3nDg5UXy3sVZQGIp58/vRxy1+FMSdMdbHhCpIyja9Y4cyDeqcb9Kv/yVNWH79QC/DU7fpgIzR
eKeVwjdVyS9t7BYSEQO33JQb3WozxQPa7+4MiEzDsS6ewsFRA4Ohg0XaWLNOpVY2jrAQkusucosH
89XLeK64Mux37LI5cAe5ZJki9BtC3kHyt63QcnCVY7NY4W6PvvSOsb6ajGgTJhAsMIgMS6rVn5Yt
afbLeAuN0w9RjFbdpdsUvaQUzMiywpJ5zlacmHj68Aqhys0VYfDkpMMhtWDV7i9yO4rrXa5AyTXr
U1VJ8wRO5UzjmD96eFL5ghph9XHSZ520UW9rVQMGOvadddDrm98Vmt2lg1kElcDWERW2kkonL2mP
zC1/hW3bU4Zzwqlo/kPog2HosKvT03I8/iRUz+B5heXrSCj756degYfreQH3/x2HrFT80Ywf3cPm
nRLq7+JikC7X9kZJjClggUlkFjBCc/nw9g/iSqKPR/qyfdfkQ+j9shr5PrIaVcsdx4hAv3QCoBmx
XZjsl4ETPfFKwaRDkPZdHKw13rBrt3eQ717oteS3TgA+oWhXuL7akASoG7zs+Wws5I9BLolI+DuQ
VNMKlowwzrU82zOBQ8dCAVp0zIpOWUP+RzsN96KbGLnHZJJkplJPE+Gj1F7EOvj+FCx3bACDsJkM
G8d8+dtK2WTdMVpI0DMcAN/wcPejaLdvQYwsC0leyGT7dUOv9UrlUVIUUJzL3NSX5f2KGFFvCsvU
/M/8rOTyQzo5YdAFi4Cc7jlGb6kxzzCJqYaAVEr9NwCpwYZjkCBWTKpnVhiVt/oCHqgtUj++hGsx
4kyXwi2kM2IGhkj/gTQokLIJNGwxHSO7iU5M+UZMBrmztcRVZVXQ7b6DmgqxW7JfIsdD/cXmf2NE
rjfv+lFCGBusQEqT44R53ddmSlPtnGcCf0Fvu5E3yWhv7onNQ60prwHOGfUONdHyuHvyijvtD9xB
U+6cc/jrdKbjpsaCNBsW+24rKdi7g6GBAQgIR4DKN0rBDokujK6nvFY9+QYtMEO9X8G1hCbrtoYc
XX1FsKvOsRwS5tuimcPAuTwozhVZ5eWZ/PdiSMqmQ2E9VkgapoqGTMUmqhLuxoIAyzaBUz13NKuf
DPTkk1lfPFUxfKhA8VCv+lBiaS+ycoL7kRR8lBMwKAi0FF6J09Bjyy2SijjC7IpvskMyZD+7iSdF
YfsL6ggiH9cYIhevF/dJ6Xcu1xGvPfxcUvMdvElCkyOmpMXtn4nLJB2UoobQ9YHeL3abG+izXO/M
Rzwo/iJFAC/aqI8TWeO3qDmkeLQhLY0ghL+PvInXosXY8vaqlpJ5/2uH6c2/SrHT5g39GUtbb6vc
BqPPT5jij9vfe7QyDPkToBjEfUPnHDFW2G2KfzHzF5tVQoZLjNwkxidH3zHxE2zRIc/M7VUeB9Gv
GCDSex88LVre0GAwC7LUCRzqqCRUhfx4Zyo1527wrtUJzN35+4ko8aZDBDbiup865o86MGCpIvsB
mgFX6sql9Bt6a+Y4g3K7m3DfMqcOZgP+eaPXp6g/hBvGP1zpHDgMW+GI/w4fBFYHu7LVArmGTKR+
1slImI5X5gE6+Ii7+HMgrcrS6UdUIfvyxhe3e71HfqYganvcWQ+YQrky1hmXSDNp5FsXvt2Dleh6
/M2dJ7XHUJZGrB6yOkpUpVqKBRSPzrr5zI2DKC9xi08JPKYY0CyiWu1wneX+XoLgS2OinYRDaCf4
EMInFzzjI5KAz6WHg4fJwSpYuwLlXYVcUprYuWugkvi0HIvPxgRaBZv7AauKafgRB5EPlEw8sYr/
gDmBdnLxPCMQJb3BdI2GIyPN9BiciY1lY0qNxVT9dSatoOnNcJcK/xf9vc8HZcav7ZlPZuJyKG50
ute1Gb4T48DnvZpxfHUAkoeuu6HfxVtkCPdCMAbeFQ61l9lbo4e7j879s02Hio1NX2QKUlBuniIQ
2RQqETXpBURqg8TrNptvmdJySBG2xbx+JMhETXyNGveCxmHZ+AwZVXM+0s+EF9S2j7XTZuJw7aGS
LoSYtgDA1nBi6dvX+lKc7Cwh4K8R9xouKGQRxUdqn9f8AMWpcv5dw74j3tDmPcFyMVDXzr5DZ93P
mWicqbNhTCT8tQZjKkIHcXdOXVIF7A9+QUevJCPcrJeQGls9ywH7d9ktG2Xst4D1qZE6EAt8HPWB
kbtfQ9uVuzWhOVfmc4zxAyglENXRCAsdeWfle+r9PLhu0yMnRhN6SoOCDeeq9TYFX4uvoM1fq+KU
49KcpiIfWzXSkscDc2M6s/QmkU0oQetlkZ4PVezLElL0xyAKCY6YgiLInadVLy/cJGIohHDuHDZP
/aKMgZOEUK1/PgamfGcNksoN8mbOn4UssAji5XaRD4OFLk71x1o/AodQ49ugYY3k+9noA50KgCZl
67MYY244rD8uNrCzyabYcdSSGc2vEk8D2LV+b6xCE2b1B9amqATEHPOcaJhnmjeTCOri61NzyZNN
Zl0EuiTNiISeOAau0wEhSRs8QTbZmg93w7oCABiQMsSHlp4iECK6J0MVgQQqdeO3i/8/983VPFFK
hO1JpbdTx+hjQZxzvORG40QLmNpZRloSTFHvRYsXhjSWuHvAbTYgnlaA3HonQcP6cLdbyclBpqzV
JXs2eJSuylbBD3iqaTw6dHtfYn5hRLatXKODEBYhSGwqTvfiyXm7rS1aoxJIIi2pi62bPRjrd2Qz
/cFKC3S4davV2ypTGDg8J0OcNh9cJYPrWZeq0Vr7d56Dwab9Jf0HU6fz8FDYzRAl/j26oqt3xGLQ
ZaJn9mneyWOtp08gd77UlebaX7TCf82R7p1noNCP3pGXh5ZPHeh8zpiDx1TlhNBa3klqLM0a5Xbz
WboQolR8H0kvrUlomzhRpcdcdVJ3xtzi5mj2lCUavFfiSysFIlugKOqDIRFpoZMEY+P01pHr/7xu
3CKO4xvQwFmrCu5aQXCctiHc7WCikXDkJ/lKVvvUe0k80zNSzUWl0dBM/TzJmpfED96Q8IFfs5+F
GnYmPO+mYCBpFg80r+uPrYqvOXXxK9RJ9ShW1M/lwlXMWQVb0y1ARVSTBHt1x7UcqN8mipfe1MVg
4n4w2Dkh6rMKTZ6MoA+aHnfqOIqzHj5D3DEBGspyE1UFd7YncDUHk104FhF/i0Suws6k5sNW0dnT
3//zR2z7hCdA9au/Dbftx2ifbIKU7XNhPtLbHV+P1bgci9YCPd20ix+OoS98Yi1L0bPx1ipSZcGb
LA35/VXVsmTsDctGe01XO1J99VILRwytmeCF+NsNYQnPEkWvvfdeyr1tskIIbqLXPAcDA8I5DRyf
8vA/eNFdEAc3AKfuLEEQb+6Ek9h49MIl4UOqNLQcGnGsxzXs7Gg3W2XcUIj39TZ/9IWTo9Al33CE
+oLX4ikSCZQ2uBxM1dcjdKSoPFMA+mxAI4KIw/ORdiHzTT7n2zuCac24Oxk9MTnuHQBjgKuIMait
rCy/iDnDunE1b4+cFtYdf8hjmj54wjoYHzZ8ItzF7VCIdNniU5eCiquCEPdILjREBYiY1ObKYrdL
cx7mMvxJk2YQh74c23YG0thCU8GODUtPLx+IUQKuIJLZ85N0wZ0AFUMXZ6ispuc7ddfXFLC8f3YN
wXH6n4gXYrV6wUmQ4xihN6GPXWLeuP/4aCLwY9X1WgsGNXbP2COJRQkE8sjKCoE/+8+wD0LaMFoO
NQ+A5a1J+XIsHt7t7JyPRMcuBJeNNCoqbLk+gU8AcNm7yl2BE44XRjImKN+Yrn/VvZUuJsZuq/vi
7k92BJfTxPBVkGLaG72+N51978hua2lYbRUZsKM9ntY9NE6MYUIohkyNR8+D4VukiWUxUFLXIgDp
CcptI3sg6b48O2Rs1uP/IwQagfdC+lV3lrNvF1ID26892HXAGPx1qjUMJfXQwmaj0mIibhjfifmV
YX1o6blQ5TbIupuVIoQEBnhJLJubCV+5ZnPXrZcW6oxSM42VKyzLVwKm5+kl2Cezh6c/V9juh2x4
WuzqJMhC5pRpia3NWAMUxuEtKx9otFGXbNDVcXQJOz96t6bRJ1zCs0AmHANTenKVTRMqi4dSO1or
sv1gA7yPFRuDwSadqwlQes2i148EyANRFsDSpjIYYK4yhJMOhBFCHwH0SC7kJtpzj38Uacvl4U2F
BMmz97yM12gSFode+SWiCdPa/pW+5uR2KrA0A3saKVL7wsq7eZ4oX7pB5IfuEBf40H0JjafhBLcm
/BcNfn7wQVTG3+YtSGed0vZ8+d+1oMSCLbxXG8uLiEuwRqkRl2y1zLKQH98mpH7Rca6jZ5SP24ps
lWrbuM089AapZ3UlsgrT3qAQqQ1aD3+PxUUcg0iUmMsDArVritKSquIJt2jY7j9NvWPHUV1xp0De
A7I3+K8vCcclhdLU8k3awTHUO42qiIZnzUMGxDZUUEmQ4hQMYnnhCvkvJLqEP+le0ZpWS+EOrqXn
pwdzGco7cN0pa4XZt2PqTTNWeM/pSNpIpDprlW+XV7adnZb6LeAPHBPk6wGTv59EH0YS6J5eKtiQ
ap2I663SY+QyF4qsmnpNAJjeq8wxdfqKPl6TDjI18EpvSMJGYzbQmCVVHhn97PAS8CrdhctmWuFw
Iztmhtq1W9OEnR4GVbUAokvVEVCq4VCY3RZJ6piPJBYH9HS2iofvRqn65V5ANn6VMEOQjV6TdFIS
iMr4NEvlMSL7xAXOF9DUOWrR0U5XqL3d0AVvDh8fGOgzU7qqT+M2kQPNNSlOJytOK0jwUxT7EmXY
Sei402ZcNceGYLOsB9/IYf0kjCQ+Z4dEoew7/VR/BxLVApCXyjNkHbnEUXg+se9kqZvM1Bs/UCuH
spGM0i6YTCB/MlE3A4pE2CoH8Gluku4kA7phhPoUFzOmH795plC6WP1kRhRYdYTcAoM6MFlnrCnT
CcJAM4+ld7UFB7ZdvO0FeOMW00XfhlhCoM4EMvh8BMzuEVFX9VsacbROtiRpUBUeeXiPf0vKZl6h
FGLcDXddZmBJbJN4NerZb5WNEdxRONHma9tu92wFpTYKGlyXsOGpYXi1QSvIcO8qzPNnegA9oNdb
RAt2xFYqdkcijQKgZs0ww19TcKn8hgY9nNbrVJRlfyCfaFQkcfc2T6rtrQ4KAGHMwH1jg6aYZJRO
TgTP/e82BEuqOgXYKDdJeWb7HNgNovh7Uqpaz9Yp7XdyKO/v8Vel7s8ipq2wTe02+Ai7R06gmSlb
Aj745qXu3W+FMHd0LgDzumtZbzQSsZj+Pi5TFqjyAIES3ktxMXPoU9QIHF2RXUOmc+1gAjRMmpU+
u3PaV/qH3K82qojcxApN+JXWs1C7nM27HebP6JVjQyZkkNfRtVvFemY3p52tyHb+LicA9467YcWq
3fIkX1ypvoL1Zqvewowitq4UKTONK3hD77d8u32h2goF5dbgOFT9xEpG8/zyxM/88Q3g17MbgMh1
GbjH9KMAmJCNLj7bWn0tkVMeIfxGWehP3XDgL2jzagbkvbgaae2w6KBimtMOyJqX67XZKe3MkYRP
fQ1gmmeoboTo2I7qvLzC+PDEmdRyD1t+QEmVPcvpEaQGNj9XjFaJlS0tl9a5hcoFFTgBl31UYlT5
dIJQMCiAyJ35m1SCmy+SRJE+94jhzhl8SauUnf5pwPQcSmguWPEUL3mQ5rEgO3UjaC1G2eQ8JHt3
GAO3W8NtCEYJXvpPzi4gPBBoLZEVYHTshlZBo/kQDfCT0FGNDSEq9BUlDp4k7dzS4I22z3Vw/14w
uF0VN17xSYHBk0aFELnxCW6rKkWzuUNI4qQu72jqzpEwADVXG3etoUHlDMuzMKL4S40QFuygYs8l
wHXU/cnNZSg8q1G6saYsyhgTxDKyuu6uDGT951VIBWUttO3EJSZvqrIw8JHGJ4D4G7JthXW5Nr3x
sEJP555Ce2c8NW8jek6UNzfaWQCQkdYCdiC9TxRR+xAeCcy5T2gp2mRaxr+mK5YsnYcNrNJf6LhU
3Kqr16vGyHW3n6GIAchnLvYiRq+coVRKPEqUk2HrNoenUTmCLqFxrAxBNcep+zBvd3+f0RR+4Ckz
i0ZjNZ9uPsb2dlnJ0bo9qy52bRQ1bOwIIuxyLvn1VPaq7G6yADQEo51dIGIhb1meYIu4Vmt6/IfS
9fVsOQvSffvwVz///i3sHVmX62sxIk0PNgajFixb6/B/GO4Zx00EgWTBe/BmGeEULh9c9MZHYtSf
R/gTAcDGCBwYBU/tBxWwiOm/o3wiXGxS2MqHEPaHmCJ1+TwqrV8ca8Ywy4+k4OhjDpO1xokXDx9n
oF/WTs/cv/4q6Qm1aZ6i+Xcz7DliLWg5cjX+fbwcYFI+pUaVkLJQX+IOaFAythER5z40MfdiYK54
tlZe6JAbTNTNv3neUkkwGqb73HyT0jHFIffTipaSy70UEyxQCZNXpfR9GA+InwSTdg+6EqMO3tGd
wPshgC4bBrC61fi/OijNMXW4AOPYvBfZ4yPDPbIbkncmva/g+o5yJ+v9HnhAUM/F6n5gIyIn4BGO
cUVbmFPQd8KJyxUzxoXJ9RM/09iq7hdZ80ZfDF6ELQIqQWY4amHr6ws78oEnl5D5JRtEytRY4DdV
j8K5l36l1H6N9XHwc6Wp9Jl136DG7vYiFVAwt67hYE0TshJliYJ49ruegGgFZILwhLm01qjaqpVk
WUQTjBE1pMu8ALt10S+KkPbecRKN4B3VzRUuyEJ1W4uBayDwZhaCwEW5EKxEwzBnX6KnlV9iALFX
DF9P3D1IqEGuID0Pl1Hj/TchiABelXm7Qtslo12DWVKzZPo6u9LvRtmGviqEHTQ3kqkkcObl9ee1
r2jD/iALoCEwQ3wA5bA1GcmaHNZo3pAGkRCF2vF58hgZQ8l9yE1SbE0OGlDQrpA8f9TEq3w6n22l
SV8M/uv41PafsNyoYMhR6WowL+YyTD3bMZqn9v5jKVoEUUL77chAjqATEtoP7FPascQhN/9QfpOM
L6JNImyBUrqBW0JXekKOvO+Y8xlG9pRQsYE4N2tsY8OyBsq3DsRroFyAhlBFeTmB8Iw7o3TWovNB
SQ7n66uozbojTmLXkM6jmk77xOyId3S8DdzvjeCqmD19mqLSIzhdfh/G2eNt0AHq7mokFO7+mZp6
LE9aYWdiVoHUb0gFQ80M7C6UzHIekxgdtOZCFBYUT7tVrxYYICI7IfKTIS67RCb7RDHz0hlK1BhJ
VRSrWbqDg/Elv76x1Y8YawkGAuZx4oxv3cLlFusfsfdLzhrcAPIyxDRA/qv9TZ+dlcEIZV/l41Uf
v35c2jqEPRbl3SFORrKs4+ABPjrhpbm9eNhRYOBaQ68wSwcj8nuCMmIVDVKdl9GckIegRgXUZ+aX
QpE2Y91Y3EbF/U4J6SIKhaBBN+Ls+Gg2x/Te8fEkIOGll9No19nes7WULR/3OvncwcbFEnPP2aPW
tPjuXFcBaHC5hxgN9AjtVHO7HDWwEejsEk8Ikk1wJJBY5ACc7PHFqWDF7l9QqFUOdIjK7SaQrVuW
dgCAM120OYftCPVuonmauoFTCZaIdTVKSeXYRxwKn4+SSdI5BPLccaS12Gbq5b715JMbEp+/3rGo
6XdzE3NbOhA2e16K9josAnIhOWdzit51yfeItXd0xhhkNqAXUOjRqYvpVzW6F1kJKduAx9x3c4qF
2hGf110kWsDKE/+4OfQqVjJapiOo9HhAt6pnWIMpYZU7BzkE5wdKcaJmolEW3M/ELw3opTymuaQW
RPevoHPscfvIuj/v/UCQpur9kc73IjwY5eHKsgD+opRDkegrIR6GBtnBhOmITXxQ2/a/UtQwmzxK
68u2+Rq+SB1j6za5zB83QB3TiqltZafvZ66xKZJVnXdMhfDD7VubBpM+uIRjcEmooQLvTSrwDB7O
SLllGg/3fSOXTCCBGa6I9bQSDmloGOMDOr/m8mJgT4qYC91yqnPQSE5DqDfQ351j+sYWrznJSTaj
L11nwrVmanN2a7MgSA0AqzM2NeZ+GqFCnU5CA96almfjqsGxwbVsLEytWhzxlRUHiLHek5vPeNDM
sXNVTYnHYpZsLHBYwqS7Uv0uDSWKzzYXhWavBKrT3blz9a5jX47JT3wb08AjxVJfsGQQgz/VVRtQ
sS8WHvr0frGhjFYHHfEiCMDZx0OVX0UncOwdbQWRzeVXbAcpyyJf1Cn/k3BbOPsu73fHAhavu/IF
7Kjja4W9XBlUJP5q4vt71BTpiNPU++eR+4/E3F6Ax4bwTcOaqvuySPI+CfbzLtWdFM1Z4mR6hllb
2tn3FMb3wwXkjNtxX5Pl6IyLM+I3vZtxO7nnZ0kIJUqS98twbwXWCHAZS8qEC5nZBcG5BmE99khJ
DLumh8eAGnNQmtNlEMtnH1zB5RgRUQw1cQAKPKaao0/FGpxRae6vlQ50WPRT/AmroxxjvxC2iFXo
j4PTFXHHr+LCTmMheHgAam6PprSmNQXa4FFS00T41t2fCW/DjZPV7ADtLaKV7BiKPACxZbapB/ru
1L6QLekf4WKyVKVYee56z76sJieUClT+OaB8zx6Me4FAwAzQIq6sjP3LFb6IEpoG2sU6CXb5nGx1
sZpTUJnob+gSZ36nnnax1ayVhQ1V/kKISJQTL5HZKC+ifH6EWtrek8R2ezSVJLa7bykciTebSVhD
m/3tqONukhdiEbvKnkeh76HjiNga5+aL6vBsqOBIqG6g2qpDfK4LAdq2e8Pq5KBkAYQD8Ed5P6bZ
F4CFhu3JLe7BPw2AUY2f8h/DjifSmPSAL6n1tMsubMXEu7h6tL0kV/bOSMsPVoWdnyMNYqkdD2im
sK4AU60b4TdK/VrKgTSAxi4dYcbDyZiQEUKKsUOjxfhidgO8j1gtkRjsJCsn2JkWYlDyuU9QdeKe
x89CgaOTC0H2/xnKzssXK76ezLpgW6pm31PB698nKkQD3g4B2IWlPpVON4XQh2gksZwFqoQlLkh3
SeuRcbcrkcqKTg8H6nBtlkw19Tt9upHdQ4QYa+z922URXh0qur2fX7k3JzTc4VozReQGyPvHq8ij
9gAa/L2rIXOU0vC0F0PGjNdHKDCzxZ7nLOA/aeCUMJjIp9MBAhFeUMmnYoBK45BbUZmz6vCs0ogt
T7KZ3TmSBPPaB6/xIw3HPruBek2LaCdCHAtt5ViqNB02h9vuPQMJ+UIV9HxENHL+gG4QDcxRjHD0
za+7CUU1+mPhfZNYckK0uH2/+3DgFOgfU4Pd14OwmWYVtUFrdmnFNUkMkvfcIc+68qjxoA5GFC0L
HHrVrNXIR1oy1CgW5C2EEuCQZXGiygO++aMXk5DatsYgw+bn/0W26uuhNmzGaQGSnhf82FhWtYgC
jFsNXi+CiJa7BoZ99b4OJ9qaf1BaVKDsGfiRXA0rbNWxTggA2HW2pwGDklPb4KU2EnMHERzOENOb
h2yqZt8J8njB2OLg5Xc048Uv6DFypGnj46nNMeYj682Gw8Fxcky45mu+YY+BDRDfcOpotaLW91x4
qUbeRQLaVpoG9gyaKHdvkQdnZkfr0vLAcwA46/GTTgo7WJ+4iQzsUo4KtFVcz9dpyklvWpjj5DqR
vYnA2anUilFow7yREXKI/kAWFlGKa5RnN6E/6fpMx31J24mBfnm2ZWoUK41BznzQj5tzyqaUL8Qy
cEM6tzCJRA5DsGkuHh7zFSpPQ1uoJ0L9jQ9IzlXf3Bbaw8zdrB5CYWQHAbRSkxEyaLaQ8+hs3EhI
3j81F7Oqek9TjAXwlSlGLR5kKoIQjOQG+lvjMwzQyAqbrz06dAVP2U90tAw+HKrrz6fxHWyXNRLt
xc6pBGQErKlzHspZk3kGZ5D8BJ5IcpMjJ6e+kLBLItcSxOdII8+HWuBhgoV2BbkbM1vE01edCiDx
oX+ZdtthPSFYilBLZ/QHuAe9jib5cdllJKaMiwkfyfrNenh6o29ip1mteZ6dKBm0NHjkletTKrj3
lHTU50m2AVU9ggj6Cr4hbCHMXicbnIKTgwJ+vIoMEdEZ4YlXoYyBw+sF+nhM1iS2dAZlngd1oo3u
KoPMLYMY/arRyGhVd3l+oBRwhLpqpoeM0xIrO3MJ4cdTQvA3RqtocWczzc51PLGPB0mamdlv0Fe0
lAYxTtYOchm/e2cnt6R0ntoUfKXM3ru/cYpq14x2MruKOmW01//uwura59LTTXE3vk1HTKxtfubk
AiyxrgYDpb06ra6prxKG3VBz3LilerQi4KS+fN15bLt6SpqGGKvXMy9sM77YpSGHYvQHmMtNG3yn
T94rEcICUfNNG+dMwp/IRF7fxoUvYbxX3rvM42vRH8oWVg2WglAMsuV31MMZmowVhrxJm8jAsLXs
rQV23yKXe7K0v0UrmSWP3Matw0usPu6CF5tu/T2pjjn2a7BpBEBAUGpHrXKJr5RZjYOVkMmlVvdK
aLBM5y6GYiFPAqwUk4/YomQPww8KzXjxo+IuGsRcvTtQbbCekFAOxA1VB3aH1Icf4hXRj4GNMyb4
sHaD5J0GtYDr+Dj2gOAFfbppk3hUMKeZUKXFL4WNURB3PiH0k7bdTIwHfsOWdkH0XfoUiD8gvvUJ
Pe1k6DTYfr+kYQG9z/V4d/jUKIzReoGRDJjZ+w20JWL9/hkNCKWjOw9jMuIRoAghq9p5/JJuj336
1S+5iysp9tyChfPAmLtppcEXZ7BXS4MDXWVsWXr6RlclhkUuzBQcLX3IxwlXr5kB7x6pPVDldG4h
wU7l9pZYq2PA+CpUzljjDmNkOYuVuV3OTl5oirq4X/yeWliZDYaGp1mCiUUYgaOSKM4NZGT3Jm/H
RZcTjQyRegst3/qZ/wmrssh/SI8jH9sD6oyBAns1GJSLm6s9vTo6o1SwmC/vP63my6kRrXhtpK3R
/pDB53FgxMKQ1WlupAsCd7sBAk8q45RbNqEjrN1FsmQbPilwf/FN5hJ3hKwubpw1se5pGf7hOf7t
Dl75b/jGRGlyiBrhx8taOmDfpny9sGcCP0defG83xciLxmVzWyP08gNBsrUm05QKg92pssdd+Je0
4Kb33700xRcPyOYt9Pbzim923vHrmi1GUOidJjrsMRMbeSAnzJI2HsM6nQ6KQMiGZqo4wEHYlkdT
lenKAKC0SDJfC97crJWvu5mCcyvKRH5M41FNoVNLqeJ8SctTAzhsiAKjmgiCFMzqJ5osWzAe+5++
dUqtqkFP7RfBcvREAB7r6CcmADVicR6jRwqhCkStiRCn3n6w5k3zaBptf4Y5ojggj22xpWn73ebV
mwys5Ttj6VNlCcLmI7pfDgKO4pAHHMy7gLj6rUOS0JdHER1D41ONVbVsSezhZdHl+1to1g2qurFN
Bv5HQpZPlKKCUZDGw087CfBiwF1JJUlZSHe6n3jXEJ+3DqBKtxn+FchtU2HWldEYgRAyQf888maA
FmysAwgVI23hJYQQfSi74bCmAhiR3jhM6q0of4/Mjbx5oPwDji7Zp56NZ1E0aBrCOdlc/34OQzAq
bobSA7Il48BkOn3Ur3c/w8d8XvR6B6j9hrIBfvn+4qgBK/UsBqFy8/fbXLTJGPjtY9z7GpWL0IZr
r12y2x99IjNyGgY/WiLInKriAPYF0xM/t8VLrKbyaVne9CRnlXAVoz/142SX+Sos65Sc9AuxC0UP
i4tGXGv2TrKJbZIa1otg0OGs2BiPrejxPDPNqu/ixOq/tXyl08pN42Q0GYhQFpqGuRg8+e3h5Jj6
AOI69ZEGnm7tlc4KFOKZGt1U5KefDT8mlX+sIgrLRpe342qgdqWEI5FGi9a3WAG4H09eYb8LAsCr
6aMq3Ce3I5L05F1Ec8MPiXWJzlNiDsAybSd1Iq5j2BIsTf3oYJUNe42dPZu1LxEqBtP9rC3NDU20
RROS/Lxzrsv/80vzZMlzVsIvRUYDiEqQBqA1a62G4Jxv2UY0YA8AjWS4CProop/lQQFDna/oBqsW
Mpb6awyFehI8oT7Pk6NdMF4VhXyDtarlj3IdeZcBgebPjRF0k4vPSe7qWKBdTuNn1t2eHdmsWX41
uAODlITUZ2KuJg8prx1UM6NBYtYN7xIsYaj/l9TACzyuAio4YpNHOo4/KSq0eTzGiC1YoFUw2tyA
FVTMg62nY2hM1uSXdJdfzuLrSawchmKxIoNV0Z1Ykafe+y9+GmjG0NFymBD7Eid++8bhSuGqNou7
GJzVn+uu1pVCfJrFbA2C4PC9RTxwHqwesqOTcaw5TD7jM2fYk+OMF4xK7vRFypasFNjU/CUSpYmz
q/2i4SfZTUA5GX6ga/y5zeBrco0kbIPTq1l6Q/8aRgQdNdGopeCR6231XIAttzyY6RxziR4YkuAO
G56Og3z4BrTyLMg5uhXNlsjewKuigjQ55+peQqHBa3V6n+/zEkWskZQGP5VmhXahkivQO3fM9iL1
g+I1fvg3YPHtCPokFB+YPGwt50UZw2Yt6nZZYimSSM77uxTukxPpEmm5r7Iy6nCji9pXCnjjPJ3Y
5N8ypW4zmBSNHUDpXmk31/eexOaTpMsZYwGDGbY5zC8hlu/JWFvYDJysUfXLFKJp2HAFzphy30gp
hz9rKvyOXa/KVKuikExNvZl/z7PJXPGD5xRAzkCFmeh1TRz3ZfEGSlknzmYu0NiYpETYARSuvWcb
8HWP7UDbBqKLUtn3zkdXkztrIbuTohNq80ZwqbMa9CWmeuKyMSQ7p/E/5UNaMFYoQAKb58/8eWWD
BUruzrfIdr+Rvu3LOAGLFaBa1lMHwLfl878scW5cbn5wFOPaNShhPG3gtcaijDDQ6rC92TtHG8Fx
Vf4AJrYzZrHjgEPbLF/w2/2uMglEl+x9No7s34EyyGX6AJqfxxGw6ENL0r2PPOfKSvv51Ly1hQjS
rH/RCYlQEYevdfp6hRoAseRvYYkXcGSFb9BQUWTmez126v9j6+0j3QNk7jmx8vzlXfBHR0uxd+TA
Hz3tiwq8NXu4V+pbjZ7QDHmPI+EfTxMIpXFd88ouPQ1WyDehRC1G+1Wxu+VNlBD8XD5zJplZFaiv
ZBGpjs9LIDIx9XyT3rlEczTOqHkvapfznjLAQdP1bXfAO/R9bZtJ8t3wlvCJ12f2S8sPo8XRP0fG
rkJbVYDwxNdKVP06JQ3IK2eo/jPTHr9RemSr8D3m4iKdiPxp6V3j3qEQJ34hPkS0d1qQjrA6H599
P/mZYelV6roKDCz1yegR8zGWX2SEGwbXodFDOM8wpDc1PbFyK5mhkBkdM1hl4UqcTfAgxNcVOICt
5ykoaxUi3uT4s4VkPF4UcLQfUVDtnz79Mm/csA0Zzsv5zNRk/Yk0OR4wizxHO37ulopHHj+RfmXo
fbKYWhYC52hnE236m9uZJrsnD+AYTzGAx+Z+l80ChDLzBccdhUO212RC097pj2WiI1RFlILKUAh2
A/zcXLBdD2Xb8H2psArt+cC9KNNJ+iFKCOW/p8IvpRqQenL4pULi8FFfvkz1XZzvotk3oZ5ybrvq
7GnCKJhIFwM1KKjMXvh0UYv4ttRpdks5HBAUPgFkazqBqbjvXPZ3dxP6Uq0dGZYlGoUZ2+DWxNTQ
gFvwL6+QcWW8vz5VKNjzZwvmTRwR4OM0FD/J3sfpTQ0pJhrw3CYAAhkFv0AQ4aojAcaT2TNPFiEd
50tbTYgRV01/uKiwkJXa3ch5HlhD0RyGVCnxv7odJh4UecU+Gw9txphpkfiaZcudB3cGBoz1qyUy
7KSh1ZQkHrJo2vQY2PrIhIu9XLuCK9aYupBVQvsWLhZfZ3OWr4lcMfHFmYeuLUh+GXo5TKso+qUT
FG63kPsbTB2yNqVZZC3GpX90JZzAHXB1qke5XiHAq3tiwlrePADVaf5qjyzoGEK6Flf2S0xbe3Mz
839rzsB5SAdZDMjeiKZdK/RAw1WEjNRBM2mcErPjQ24m598/H+RIqzyVNxwpwEE9IU+EVF+GsRJY
ZwGcFIen/WgsQ2d4XXt21FwTsX1m+XxWI7C0AJ+CxP32WOQmZSIM9NtKMZZTTyRL1n5u4Ey+V7ST
ezFtY4Agpn/2gib4dfxKj/JN+2AfdV1Mua4YnRzjYEMdBlOVUj95EfK5Ennm61U0SHxxNu1pF1Za
yZoIgOreZszgZgk6+cKNpujYuVBCEEV3gKvH0Q4H3eXfcpJqb0eF2+gx1RIsgLstDIiDdd0kHyny
ErjK5cRsGSlTVN50HDVh0jzoMqTQ5fdzBk7WMKT2CWhXl5gHKpPvEg+XFuCGtEta94RLNLkq6MAg
p5y0IN7KJLudvFwbEnrmn6ae3QM58CGcfCJ5iDj+lVVL/HBrFqayauYuA1GX7aTUqaG00g4XA2q0
R1PCZxR2rVzF6AZW6A3wsyeJJCrjE79ovVYGpqN3FEX2OHkqZVWsdwiFaUI7EzdeHbELojx688q6
Ke73KBxtHz7F2qSR5VKxRHxrt1ejczU5kMB00Lh1AS7W0G7aj+7BbWpar1NO03pQONE53lKBUuUr
4OaPGU7VSeyBtnBmSOaxcsxBEHVfPC9zwV2kWkK6RwTdBH9Sh36epo7oKLvrgxLGpv4/UrZUM61e
8gv7McSGB94hDWrrim8g3OrNJ0bW721UNEMstKhygAn0hqzQbm74Te0sQDnIasi+U0Prz8UFJycZ
W2o6tWxMRnFzUr6jmRRDnd7cKVs1Pees9QCCQjBy4O9LaWZBmcsyfHl75CjkNzkOCJVP3LgqLn0t
5Subx9MizFeSq2BEF3h4UaItH1HDc2X6NoIX9KHd/dtXqujm9wpzjYXhVvhSipJvvRqLd3ioy8oe
HUZ7Ca1cYsgXgNEin187z2mPZ1UU3mLQ/EpHnDbkMYB60PemTGD9BJTSYuimhU+j3JtOymDWpGa4
oQm8Sv++hIsYPaRcoqL+caZ/V7Kmm7MMHBEMeAdTSJAS0lO5NnaUVv+FzgCVQSSOvCoZsoT9NhcL
hvtYCHdbJIVcguQ2NuesxgqOXcLOcCzv2rKtpNh7/BfXZIYN09Px0EIUz06czZf4PIqZAV9mFqzk
QL/KxIhaotcq0Rxnt0PsVWYUEF94z2nbNJTJscLS3NRDmHm3rY9F1iYQXhUeFqDH5mlpQkV7rt1Z
TX3veDgaoZGyX4d7ZMpSdEGgztoThi3zBdl7AbHn4pptF7AKgg6bx8CnKt7Xc5u8V3udChTlkTUU
chNU//7O13sTqo1qOc6hfeecv5NYzKiP0eOs6V8rfykeq5PURzAQjYbORMO29jOOG2w71lRA4DLN
bhqMGGtTgjPzuO/LQtA2e+XCAH+QXKMWq9RAgP1n0R7q2BCAqj9sYMNkJ1+/DMr/ogVQcDItSuRD
g/xO45ak7rKuTe2//Y6HAJBHT7RE0ZUtiHXXlcwpRtDHyyh1HJPzr0X4IXk/Fm+R0XkHOID6n+dr
vGBiUsOqF85m8dbdPYGDpZ/Gn439P5CIjQSueU7iSPb2m6nAGBwAX/GA3VSGRiv24Lh6tdDzWhBR
OTSvr/E6tkoJDPtM9zLPtEJQH1bUvmfO/WsbI1S7vIYaS4KwuZtJvad+IXBqzy5j/effMWfzNgLv
HDIzO7vRKWz08nFR+uBl3OWJ51oIoQ3dXMLmDNcBZc4Z1EEWUiiJGCFeOGDrYX3iVSlwdHyUu/mB
DzoG4D7bBxqVVYorB38xsYzmZoCHpk3YnLLrqJn+piDyr07aw/OdnSupQsdhP5I5OQ6fzjscJxrC
2uaYl2dG1bxnapsVVaO93HkR4xVoHcoQmyoBicgmk7YwBtuwBIp6pPC6f4yy4aqeHb3wfUojmm2/
BDsVuByZ5j8q5H7L8taO5sfRqBqDBe/qyq7Xq682CILmoTpehJ1m5uV/ouFv/OBUv9/x0A7lqLRA
urkO8UCW4fd1fyqua7NXKFm4XWCUHNHTNTN4fnQTXXOG6WW/fLcX2+UxMOL/cbJO3EQHKK4/x02k
VI6WOcGcGaPgyPq5c70oFPZUqSipVJlhiyDELepF4KZBSwFxZdEARbk6zI4zK3nTukUwvPspMlLX
3wHB49KOBarkERd6x2hrlOc+5IdmqeKo8mv3fOENcn0kSzjhR+Lrsk6xAitjhtDeQPPA/Nisdx2s
FuD0B7YXjQZnb95aLvJ9pROh0VVe5Hu+vJLlyFGeRnXHY4t5/f8A5Iibh+5vOrQygzpw8vXvRUBz
Vp2ZsAWll44anlFcCdp84cAaWV/idI+JqtW1kUhCvujjuqCh/MZpklT0jVhVMgD99MgXTzXE9fE2
kGFPdCB7CshpLMPp7bldBCpCKSTEWJui6W9qXEVA9RHMXtDyFWkQWXDpInNKl+2LN3ka4QJcYHQC
yO4LSbj8YwFRQks8+yRrhMxOuo1kvtqzwVKDR4EBdHd8UKOKhdtbrNg1z17CE1dWjtJN/rzDR7l8
aiNsAHBwCTaTk3kZPg9sony4aL3KsSPVf7pp2h8iY31y13VbcTO9FTd0M4q5YsDPZtZbHnefQO+L
92F5CKh9zNRybPjeMDQjuUOiSz8Ha7hbZfQ0cJbWkPZ+28YU544fzWghoeUxNC+vIChRKi9oVeJc
v49qCOfnbivlSfXI6dPKnjUynfBOT+zDhcegaQ5AtLoE097T+gcCQ8tdESTsr5tOs+7bXEvTjQd8
s2FtDibrVcAB7n4nONEST2ZdHzB2hSgGVb6+XyegtiFW4IC0xeqHnGkrG1qOjxZc8qwlGJ4Wrj7b
dilJ7tI8E6s45eapWZ88wDmCB+l+zi2SbNbpFrqeaxovEQPGGsjYe2z4nt2WuCyEKlUxZZdjP6xl
A6mcHlw5lorLJJdRxS7/kkPCq/lo6dqXKzwWikbOi9naQU1Su9g5nBwIeHDnvLk+Q+Iv6ihu/eAB
3W+nxkZDAxkanCXQJgBl4erqIwNNXxlZy3T+K9lyFHr9+TkaDCYiDEHBNrVH81J2pQMnzMpthxPx
X8TQ8VIe9ICYW5zJACurOE/SOi2q9yJpijQ2DQawUJe+BixmtYTuWwpZ8fMye3X3ZGYdKJ5/fNUD
PpP+BFfkTlGjJGIiSbeTFqczJFKwbt+ahCyVqd0apFYKj4gRVvkgmUcoUD72DvbsMap2pWTR0tP/
ZyJakkwauvgeMSCIubyNGnkPcLC+/kM87Ek3bS2cV7sh44dW9poh2c+TJETbifRVLiL/QPXzi0gh
9WxY+NPbrpNXXnoobbtuiuZHZzfJcPBMK+ES4Q2UqGm3xHgZ95dL0Kx1me+QCJlpjhEjI+YZ5NPG
AmqNI4Ptddsq7IqfzOxTskCcBck+kx7zC7D+iKCbPVmMrM+wBVWxzLCPm55PJrWd8KMl7qVJ3PYS
O2mfQdnc8oR5WWxN5dMqUXbGoZk3pVrO9LsAxr1C2br/8sbUlVol2g4RRGVlu87YVWUf7Hkinsc+
88hmxOJl64Y6fiquwTkcLJgUWL6hHmghY4HnDk62gTk7iihqYtDxqHlv+2GyFmiU3PaznW9T3ePp
Ogn5QB+nrDRzzw924e2nW0ITmOVudRql1Y5VWfXQUwtG7j6mrP74+P1rMIapi1EhDIGnOhtUishv
90Y/jwoyUY3hugnzrUgTxBScQJYQ8ke57pcnsTiDk9eUcO+fyrwY5r7zcJJZZtg+D2yWKOIXj+Ql
DK5+wYZxGBlunuG4YNIscb97GQNlF7DNhLiF7gKsSBqNonHPurv3a1Q7afkXrjVcsz08n2blf9lM
ogEHTcaX98y94a/CATaOToQWNu376G3UdnaQ47hU2JoeKQPaXS5joa5VQWLNY10g3JVRm+5LB9o5
gMZmd9QoKEsRS1BHKiKGvGK6hbnR5lQGk20qxf2+D49q6I0mxpVYD6RB/OO2lCq6XgArt+1JqjiM
4nEb9adcXOztFWKyZ7gHL/yix9/chiFR+av4g2EQvUwhWESwTAYQtGQgMS6DxXTFalhytxl30jFM
6W39uusZVw37zZU3wbD1RS7TJfaB6wCVnONuAhU1P00aVm+EIt2S8tS5MjlBFwOR1l0viI4xUZgq
jT9MmVxRwNbOaMVpc3B7XWGU+oDD0bM5z3HX0sqD+WAmhEzzMqXU7ekMDKHI0RPfR3WFclQIUpfv
Yc4MTjg7PPzYdxu12qy058M+7BNADe602qiH4SepYTAeKeb1fAjL5cI4cWOU7Nw2EPl1lPSAmJu4
M/tWRcRna/bmLoAuT7wNL42CDRSBuG+35MVza1tD5bbUtNnJ7LndJc6sHt/7/H80syFFV7uAF3t+
LisHP/DHmmMvXATUxpKW+VutRTU+jag8l1PkZArJ1woiZRZcf3x2xQY9Zf6PAF4bfqKhgfy5Tgsc
JMGkGUfpZFP9C+IS/TIT4pkPUmx6jp8W/56h7DHQVfFFPVt/0cpf4x82Z2r3d5s9AOU/Ting0GbV
rbNVUU4BzD9SX4ZBdiju13mj7rUcbIqilv+SAQd0lZJQI0uMBbIVFbfIFZpB3LkEnxMEoIScl9cr
bukyJkJ51LtWVNAQpM4FbgSzsNrvfZyQR4dsLk9iJAzmeYaL3O+ebnv8IK8KOLvr+rVkHj/WfxJm
5etffCPvwSl8pRAGMVEhWDoULP7BWkPTTH8m8mVSpuYysIbJpQ/T/FMBRNsBfWIuYS+5Qy5e4dQG
/1EN8Ly4biMW7KhuQjoWeP+3I+bW2D783TyxZQcyFmYC6TLRACwzAAIqVoiW6rE+f4i4giQGvbiV
88mM0ouhZ/G33AUkrPMq6VtSJbLJfEwiADxF52/2by+5mfhOZyasu0tfz6nxsD1ZVcbBr4fXIFaR
Q+2HN+sgHii/sPmk1GXPGkROyL/WBlrReaOBPb75GzOwUmGd9gV1aG8gvMlXEbfKs3HvvLcIypgZ
9FFJYD04+es3OFLG8VuOhE985Q6+Z484VF6GUki7TQ/USG+ALNDOpi+cgkVk/SSLEJJ2p/As8T6X
Gt6vEQcFuw117xOyRvO7S65PkgHgZ6KpR+ner7Qaqr60o0QKEgvTERMmoPRJQfG7LUr9uaMX9HsE
QDEq/WgkO5/+0oiXId2674G9fD7zZWAdaReL24nU9tpDC1oYMFVCBAWPCi0i3wGB/HQJFfY30WBe
LM6ohwGkBVvh0rsBgUoZrF07++Rb4UA01Qs/oLqUNklpRk+tbh3gzsmAS5J5RzAN1uRnQKNUu0/+
XQR4IihGYC3a319FsNGcldlpunBXxLirzTTMb/wBBBrtjJmLNlTf4z2WQbimLpJ2Dqc3aXiPG421
IHuKfIiQLBP0wPAMHPZ3Srk4KdZUUT/hMc0Eg9mdx9+TH+CkBVA+1htXzL8yJFRrJTMXf53ZfOxQ
QHohmfjMT6+H/lLDg5n6EoT72vcEKSpY+PZXm1qwzGjRdiaqcDZD9HT2I6MdDut7TfSbWbh9Tsx4
oz1A2f8T7gcwo9s4H7KzOxVqtZWRwMmJEWPt21VyLNsaQaHdBTj4PCwa4on0rFl6CvCtLCZvuF93
rrziZdwK8YQA5CyA44h7C20a1CEkWIVdeJ1akqX07lcRtV8mOeb6oC+VvMhMn1MS4EJISwZ7EnOo
XWBxZqo5IN3zNxKFSVN5XNWctJ+buU2kbKpwfMO0rHRsAc4bQXnEAkuqljH8uSu4EvSdw1obJGaV
+dX1TuNZG7Nv5TDNb0ac5Ef9Q++jI+zlOl4CfxQFZuKAHoPkadgxzARMaqIs/JDeGDLy9fAJCDXN
4KmLOf4SuQTaeFf5KNbXfLnL1DOIJn3zfbi8dg87ZrdUMii76MzjgNnqpdb2BnkLNEvg2Z/kDzy1
RaOLdlUKHEB+kO7IOrN6Dgafp/rh8we9q5Hige7BZgah1Ka897YWEd3OybaNAHalJ9tAm9MQ+F/u
B8wCO9s6yKBqEoS/QM1tmxByHJ80ButaosBxhLBgRgB/eQs5kcwGP+JW9/3jCAnJWPoqMNkzymjt
ma4E1hzXOtfI1G4xW3/CG4YHHrcaIXJkQqO19bIfs4YaYu63BJh1e2kJXdXvm3hntydJf93T62mT
91+ob1+znRFBNMJSvjwx3QA0asHDHBLzXTergMvXdV8mOvxx243V60XtjMuxgwTunXZDTUaTYeT2
jXegHGYq6jimS3N4hY50umqyVrwNrKwXj5zFfEreLV8BmUFESSvnH7LJOCsQ75Iz5bAwTZHYF5cC
Q+IZntP7uokyKef3wPnShSlsbAFWBxsW0gdrCFcMnFbo2NbmOlqNq5rvS3KdiwT244F/8vTjx1uy
YIdCui1ls/CEeNrRCXRlxLf8xm+nHM1Zv2k2GO7TznILZlmx6Jpe6gIeAt301bApa3HXTWrKs/DQ
qbZ5rqxraQQ3RK6pvOy2AyaDkllkPnhZgj1cE6xSzw4HVJkLT4kcy/m5zKUlROTMNeM1hB2+OkZV
yJcKSN39NolQlsvn3IMP3JzRUCt6CXiETMJQ4VXZfcsGHhgX7030kMeTiwANpOgmWecwttxZCj8w
QHH9WIBadbHXsCddmxfA5urd+VUD10kPv19SIcMqQn4lW9Sk8Q+AgRXyVkzZpi4TviQR97eYQiNc
N3zOWS2bwtqTUTYIGOwcR1uCigGd6RdmHnvHg0Hs5H+fd4JAdEI4dEl7qdRPC2gqGsF0iYiERwL2
QfsK03oQFKvxy4DDo7XZkuEY/MapT6RSuP9vJfp7A1mLOie82NufW3obhtncPnUYCIzZpv/PvFMa
IWzEzArClmqGJY7tYJoL0vcXw1wX2U4h1sXjz7mnpNOEq4iyfqxy5L+rHqdyIXFPyXt3fQsyEx3W
g25J21n+awqm9ExlZM8BakvcMA3Ts8VoOMSnwiMV+LNVYkQv6hhzvj3/JXdNuuDvmyfJYj72tBsh
iuE08meuegPzVCdnY2HYPVQlKs1JEebm36fVQIkH+wyVyVKQwDKf0bPDXx7nJq6Ot8B9GsFnyzul
d6xcOeUpJoGqsW4jcRnKG4Igc2h8Vj/ow89TRoGoNxB/pzYOHO3EV6EFEXxwDLYniQKhkTYKP1fH
xai21YcuOPsDh1zwas5GRvZwSo9rSk13Zl1D1M1+ITaU+GMZAUJkdsf1akEkh7vYhPQ+ULts6F5O
uv5/MkCrwWjPQCdoNhIByxWzWVlT+SULx1+imOM0Q5rlikuCndsiU4C+Cma1Efpa0AsZ4DlSltw6
GXWkc7YAWbi6acl6z9Z0T0Er1EGFh8gVnldlAOAuBfHwao3NaJN1SX8Q1Sz/BmRJYCVDcZjpWoU4
BeMe5ZcaUz9tv1qbQjlHto0JiuzbCmL6NASNbNczp0qf2OkluLY/iJwY/F0ckr+cDDTPP41rprf5
dqxDUIWgcg5dvIwcBCA1vFz4arSbAO/4gQuydULTFH6+W7h+qk6ZFg1qSD7W+bPtcFBQqwkx4KtK
IHADOwmX64OVhv4vZJEKIZxpgVgaxS+kKe8NRLgNnYSpvGluHZQXll4w1kd+yfoPq8SYqWSEoXQN
k7KNjdcD7u5t/+Oh7F7PzNKdpi/HNhQFssXtZ3qZaSfd5q1QBC60itrBBzWFuulSMJYkgw2+99Ek
2jz4fwLs7IU4NeLJ8oE/iWQ0KYVexi1PMXN1I6zOo+MWEWv7SNEgip1sBxlsLjbOyniEHikDuEz9
YaINU/AwZgo8AlcgqEd/Kd2cA27BQo0koJOrkYFCN9eCVZ6EC5GMswG2fO8siLIfSSg7ybCk1DpD
cyqdC7Qoy8HAqVbuHpL3IG1eL79HrC5fwv47cZaSuG/ZSy1vHK7tND91DGMo9kZ67KUIxMT0J4AB
Y+DTf5guVy5wW4AJ74zxhwm3UHOhMiKC5xeVCizppdtfgvHeN8MgNx5gqFgPVGywWI4g9TtjpsAT
BvTVDRKo11eoBfJ/eCVk37tvOlFKRo7PNflu/D6aWi9gRTgFnb+OFh7O4jj84fKFfMDNRu9zEOBV
hjvXvKUeiFfeBqxDD8PLrrlz8Euv1BmIq7rimIE8r0VP0fWAC8y0r3mWWqp/zx/lI3FLk5ORLZ4e
xD4glkYST6dNbaxHi72OdDvILLhNW1jtyLrWXjzVrfsFn/DkhCUE5IyNHJzATg5lVxlPua46yO92
Z6L/r/JVeBh3ZxakV93GRLKD7yf3sHngWbgXDjla9ynblpKoYJak6ph0UmkXkhWuU0KLRriC0idX
8Eo3cn6RTm79fOHj5G0BVMp6nzuxq3eG/vExuLQUqj4uCDxuB7FaoEMtzd6dnTpaNZUKcPuUh6eT
p7lbkOIK88MgxOSFUkTmYq9qpW7aex279W+iTmKaGXkxA0dAvsH6dil0I2neUbdSdUlANLQm9JDG
TjTaW2KBS6vD2YLRJr66sKH9XfgFvU4pZIoQZUtNrmrJFwwfLUuCVp4BmnFV85Dm6LNxTuRD6sX5
mCYqBsRj/Htcr4EyubGGkoKSLhuK/nNUdgQE1Kn3kfxv/N0iQ3gXx11pO2M9G21Vjwr9L7dYBu2l
GBbFs2VOSu1SEYoDxWwhNrIFVs31oW6HjFID2WpmAwk1jKqDAmTjEaMhPjMTGeIvtMo8bJVjsmM6
7dwVFEfEPg5ex0STRQuySW0h9Ox0dV2qg17StqbfCMHay6fLlEYqEFltuoSi5NZnadxLfVb2an9M
oZ4jHUi+x8X2g8SSWbY368XAJwiPjkdfryWHmr2FG7ie5aUcldHqcnxoEesq2w6OjdxZ+Bdx+9sh
rT87qm+62uE2vwfx0hta1KWQmXHpc6SD2WMge4ZVqQ6veLySS9ck/Tw6qvRjZm9koF+b5pNunC/b
5lxKOcLf+Q2gQIZDXgDAaPYjAqKckqCzVkV8dH5g9rBIxHKUqxVeYEpBz1Af3YH5pncb5Ni/wfwJ
zm3BF6o5OkiNDg06bP4e2Lum8IRzbDm2e6PWYkyLtFD5OUk3KyVwEY9Av4osnRA5xN8cgNLWtdO1
+Vffu4LBLtzz2TbMm09kqO/0To/L2DZMnFbKTGqORhFglvxvrsXPtR4RvWgAP+IFvZzHt3nXUikf
C7yrnP3bmqTOmpieSe8kcV25JHmTMbl83tpJusJc+ZnwfpjpA6Ilb3eFiovW3OmyaSGz0ylAV1zt
S/IktXq4uhkYiuu8Gl6neFA4vVu+7gA0UDcXtQA6+sDLFOgViRBTIlZ+KTXLmX6w5vnt+mUoZM1X
zXWe8COBT5mkTPFtoDRQ3WzELrCiOHW0KVhwMvyytDdngfwh4aaKi4RokNnLw9mX2k2J0ptVGvBv
tQhza5xk7HUtfZWxZxPU64rVBs3xu2nLUZFO3gAPd8tD3xMCGLG6JHMk7dx4ivMxP/O/xJCHnbOD
0prI3B25xCTPQPAopkvWdB+PyrWqSktZUB6E56Op5NkyhmPCsPKX4JzixPcGx+QAT7bwPFVcPQmS
qjpHrEeG5uFij/RyrXKZgslQIG/hnFhqp9evLZLYdxbx6IHRiW47871ohUD3tRPraSOjhA/0UeEx
mdM0DGMhJRHBDEKOtDrQioo2Q/6wHo4dtlWd3X++rpUnRqqqYOxp/c3ycXn/+ovzmhhCaL7/T3EH
stb78fpBlo+nPI4Th/wEMxvOI0SS0H7hMHY2yqeObLCEzVQ5wI56q/XOS43ArBlsrvZ9TTvwWd8k
c6SjcqkipSQHpBh2bO2pj/LKgYIr5T+s5b2Bnr0KaguZ5eoDWOcx6fSZT2tczo0Q9dXJQAdRbX7F
x9QhyH4nTlhh010Pd6IwAxXER8po+NOKcBbpTY8SNi+aMy4BmeroHmBNbz48tRFZUZ+1J1U+d+O9
v5e4D+263GfENIqx8ks71Kyacm5L+55Ly4GYaHiZMBnjBkRybAxctG5kvI3sSOxKhTL+WJLGWDSA
Hju63822QwEhMisax9KFobvdyTtUZD6rsUoaQs10K2FB6BmrqnvyNHdXP494PUSwfBS5HgZO3OLN
zxKC+Ag6ynzosS+J9Ity+oqkx0/gz+FUI5cCnXTUcNFP/2qQiP3zxaYW9N/d4RKtP2S7fVyJjUWI
tL+xJi0UYJgYnOJf9MiFeSnQJjtIz6+XTxcvzMml2nMJutpN0IHaXJCRusUAnJBjMUIXXy4A9GNh
0umkShCb5E0zJxTYgYbrQhLT1frPd1h4M4GuHkI3k781JpV7crZzZQIeb8BZopheSAXAq+2TSSv7
qWLZKVWC58RFyM6HShLZdRQ++z2znsf7RGVj0cqxNH0Vd6OYOvce92duTtkcYj4i20d6liPprbDE
nrSBF5kWn/Uca2hLzrd5pBzg+gpR6AbZTUOvBzp5IrCTPSwJ1iX0kc+saTvohcVzhuIbpWn9Wwzj
o5OWLyl45mgbRA0bD94fcV2pr0wpWFHlhwzKPhNbSc7waDuMJse2T5FtZa175OQUYVxodKH6ttKZ
U5uvGnfmHAAqK9h6hJY4ss2+NhOGvRMR97nLNAdFq8QhybZ+72EuFRwqICchyoskeNkVdbirGYiZ
IWk/KdVED9m/EKaxaihC2xLl/VgMXrpNmDMwN/dM5m6XlZdw6XiLt3e1CenU4gM+U/CMxEFp4mrY
X00PZiOmTiqE+8KcJCdZQsrnMkeUXVXsRgJuFi6m6C13qp1T5blvn9tvlu85EU5dW/WEnlKBcMY8
30ybWNSQfbsDy0hyss/V753h76JqxbwPtDIP44tH5aXYfs/RBecxZ1J4fcEotvDCyiCQEYcPxxWI
qwtz1ffIbAvMkymG9DV/dITrYNq0hRm4FYbplM3+01OLV497yJMAyc33ITFZ8hUh4tfOFS2mpzow
cU7TBkaBnAiD9ba0WTrI1wnbcwwYVYC7rg8OKJOv/9Qp5wjMU4uHVxzFmvxrOcYSF0w3l/q4n57C
sbSZVYgz8boTTlSB+t4mYhzMPIRqQFUTiuAQy9Dvej4m4rqrwOGD+EKNxChgtsiBbHQH5+S9zCaH
SwECzfwp6mn2hH85e/GrPI8EzyHABZdAidNnsUMtiuoc7eeoLgNa+VX3uom7NdZ/HRog21dT6PjM
WWOPMfLr9UHeKmVNOVvpRj45mChRiBl4xPsHkqoLu9k0RFFrMc7cjgvAcfvI/dO8EYejz1wUOg4c
eXExASMVypoWE9QCwQzfnXHyKHr0rVScf3sQ8VyhxUtfVXoBKVsywW0Y//bTgK80l/RTEUtAzTme
Hl9b83uMVVYk9cDZcBUS8cCGVpanoR7GMTQFFRgNeJTbuapDa+WIorMnKvXye4+zXboIQlSJx/Re
AudqBmGX5w8598kqi3H8pjFaNOo7qFEhEf72Km0o9F1Bqk/RuREDUxPYrkn7ErgEmqfJMw58bgo4
wNxm6kYNn0YLKhI3TZKMeMFMemWxfeDAONUUrPvnp/bMQ/NcOxg+A6Ee0VsotI03da8UC0O4N6wP
JSVgdODSDGNjQsgjSYvoCPeFhwM5Chl6y0Fl0eXvAqcbTSKQH4kSdZu+gZ5K0aGgdtdUIK+OyVQN
Ge/tz4OzPPkiwwRRHA5brHG7YE+x2L4stdGh8Pk1fbgkSTludPRdUpgJSSXvk09/xdupANtqAjXz
Yrqb0kplYgck1KHMQBv9yhZAKap2zHfEopDKKLtL70BWz8DbCOWI8svqOxdLxHdDX60iTlPm1kRS
RX5cXqcpkZBAPECNjz8j2a5Sbu0DjKJcjnrwuj+c0f3LvlHJdB3zSrzwX4bM3JbJRDNKIVb8G/8Z
ZSdVCsEq1Pqhd+2XHPelcoI1g5Wf05lIeIjXYYXqr0znyoL/ES39OsEGRNUmuaVtktaUsYMWykng
jeznLmqWQfP8yz0qKo4L9QnF8u7F6BmRSsQObeiaaoo1WBYvA3X+aK2e3TKcOUxlHdQbCCqMtNl7
QW1O7FG/hqXB6eTMPFf5Cbp+LIyKDJ7rE7+3UFz8eAfrmVxyVBt2YJrh0NQlbM8LcGikv9VdiQmy
nAp2yC62HW1b4SNcRvsmhi9zCIOaVxPNXrqKpmTISP+RxFoWzVabf8ZDetMTh0dBYKod39cNq5rL
6L7sqK5BVTvP1As/fE0W1YER5FRqAI0m7myvHB+8+dDytPak5u7Tu+RuZ+gun4XjS5lS1uePLhtp
warCBKMPCZN//RTY2UleDIznomp9l4vmZgLcX1LBc5qzpTZxap+EC5XMI3cNHoQqGE2N5GsX2mrW
z0GhgoL1u4pLvf8lPFlZr0drp4pCFjnMQ7pGaF21wbGOopr434O0Xci6e1Jr89QNa+ZCKc6Pu6fa
CW0MfIQm3EhMAmYkS0TrFcsRD6gXs+Raiazhcp66C/qaeOn+7UJnnfnBcWs4gOtw1qcFQN3QxX61
9XhM5o9AI4F4bWne9r/f25zmWBxbX90ubeHCpnt8t/yJWa8a1D/Rd6aTXsUq38x6NTTP0a42tfLz
Udgu9RNwk3Ps8aQPpjl2Q49kEKCiOY//ezdvaU6pYicMV84l7yZzOmctGNh95ekSKDXD04O0F5SH
Mo7aPXCnEPedsQQ+KIw9QMgj9/YWDz9KXSQaVhTRfA+52fhutl6Xb01qcUO40C/1+/Fyjeleo/g6
v1srB2xjIrTmDazIP6osEHBrcb9azJlePboBKk/j43ZHs9P64m2vRn09bYuIgoBL01cADD41BfWq
55lTrDQzsF9kXM7vGppI3thjAqEG+ed8kXVIhyyPbJPBspO2ktkpfOySgxB9jlktBhBr3ykaRiB/
jz5UjKknjf86tpESdCMa8Qy4Y+OrKnEZ9aroVN4z7Q8F8iQcHF2vwjT+Bl/fV69PgdqEhCNg+zz5
afIkdrnIEng2Rny+WLsiAEWIK/bI+gCqFwPxuzc/RiLx+dL7EeIWfq2CLXLpw+2pCzlHDooX5dwx
r/aN19raPNU3JToJan1vOgzxefDgnM+ZgWpSh9xTA/W2j/pUkgUsdTBs8Sfkcs58z0NYGu67emWC
P3Jpv75ootrqMjrhCq1lzUqixkYvA+oVY2nu8IQwhihhTbI4zv2nTb1gML7aUzAyhDv4Cy1IhtMp
98I0f/x6V7DxgNxE6OSqvnMloBwoAIDzeWvStQyJCKCFn7NYNFymDTjs9pNIyJXUiqztVCEGwR+o
cpFrxYSgUPA/XUxG7Q/CHzKkZ8n1gqm46tBj+fIwGp8MqJLs1RjBJFIywE0C+dGn5t7Kw/9VPiHf
VlB4qW9gRQvBJJdUnqbhHl/YBhZ6YVEIG1Y+uUOxd10aBN8niL1jAxlizXL2rjBbOX721aJlONnU
W04WurQOc6blXG5qawL7ZJy69KY09n9Cc7P3Amu/XeZLosQzWj8ojn0UqYC+HXar3arqOjIZut22
FvqfevWP6X1SXcdsvS3S//yFHZZFwzPgxwBYlwwUTPIm3w03OhVa3fqEoqJzyTcYjbhFomrEKGeM
RFwBMqn/+KWxyFByrd6ga4HUa+W6qe0dqZPq0OI55ODnWx4yeaIBNRabRIXHGqS9OT2ehVlTmdI6
cMBOpC7GNbvewp5Km4n68qQUnjACgW7Ks6dyHZ4ohA0clct5jhdY9Kd7Nifx6PtHtfI3neqQFjyf
9wnGudSoY4++9GDBagybDX5AGMhJQv6GmS5KiEdqwuoer/Z+oHL1JnGe25CIxOrqS7WhAdv0juJR
NFLoWuXh9hvM2HRIB2QtGOxrazGQPwiyzkk7AdG8L8I8lmFSTMKt+QpKbm1RzCqUc6YvQB0vlr6e
78Xay/wpy/G+xH6eIupB+UymQC6jh+gryi7whNm9ce/de9NDQcqrnORAMHSpogD7xOrNzJRHRNa5
EIzUaR0g0HYK5rY4lXp+I/sKy1asn7w+eWkeMkGALd3rNyQ/isnd08COBLQFsqFXJF5ESOjQseN6
og3fIRWJTr7kf6HFGWKMxYPw12anx38pfK8Ht5rzaKKscr5lctaW1ADXpueUn+YS0gHSHuZM2STL
MqpbNg7w+3X9Pl8W+RIRKkXoerYbVYnRJ+aD1Qi9bzA31yrPRD8tfLE3EdTfqxZs+vacSZySnHMS
yxewdudD25GgqantKwZ/Dcctp3jfLAVNJQySCktF7AEvgDtkzBR/DI1kjajH1Eo5HdimuJhg70va
XemZM7gPE8+rTSFRtyx/PYq437rxlAQLFaBDycFt2AUotpDCs03/RzpNdDY4xyC7DJVX3p0hVHw1
ogaKU2wVGWPwBDaQwKPeAdaRsnC7ipAtTEC2Z9gJ09zZTr8o8TOmEtu9jzJV/y2e1vAuecdPEMTW
sk4yNLjG76YwZ10gpiKWkjdhKWQNtDDYRI5Juxx+TpwOTnVuxQnVVVG8V3ssE6BYPS/qmOkCen9e
CSEz9xbtHpo9xfVFNeWoXUrULEQRBoUthBG0kUk3d8+OqBedUzfKHD1fAy6Bv2aLUPpKuFrPZ6ru
Eq0vTeRjMNR5w4nhzRnYtI6LfkS0O0T2vDTsprtGUS91fNLuFGiUojhfDlfP3c+rMREGGYHBTKgq
YjogRGCc63iSPMcTKk2DqVf7etXEz7iYJIRfyCoQV0xX1x0iEu4mgNu4IE28DbEciC/pw0MC7l9L
cesgnvJNQEoNLv1L/OV3dxx761l2uDZoVMzPMbu2Xcaep9OwbzyGNVnSd0KgkUg5ZimxNIagXrOw
kFboARqjjWS4H0mQLMZrGWPRJevOuvK784WCVLHE1wY6HFo1Rioyh5o69W8+ISUS03ASWMiEkjZs
MEKcdFhxJJw6EfNFybzMfXbwt5EUSOntNB+E0uofoSEwbwcu/BvBcZXq+cOaDg6lmuzEE5WI0x7Y
sjzOxkT3Qzds1GPxNMuY6IEkRZOLkxUiyQMiz41FM1XuQP7peBZ+5rBYUhNO5xybEgjgpcWb9xNL
whs+pwFUjLdqdXe2Ja9fm/dAamm8wLPFjazKQoxhWeEO+BGjHSGoZ+ERpOeyRypSfATcjqyeTENm
YtuHFrXT1h7Nq3pyuIe9NNF7B37eem6lQzcA1CPJDmuMOJKl+PrO086vvAGd6Bz00XpFhdBjLdiE
p3Gk4zm7MHObpuMwV7GOZYK7geMuouWLG4OvumkhT6FTauYnG5+CucBifv3XPj4ciQTenmFjanyW
FAlwE340nmGGqFziW7b/GkO4g73ym7OWvTsDkKzebTAjAw75sqKeCfPVN6w+ZRI6vkN1iuQtcV3J
RayMHVP6DwwpHKlE8QcLRdnGaXgUmgZoXbzkLX+eU5TPm+VUnKcTXiEUYpnh4kV9pObax1nzkyFv
DtLki7OVBFWpnnVPgW9DTdvQBHe3Z80KPbVjMHdRX01vF/Z6hLwKJ/r0rFZO7oGx4bsiCqr8Stg2
NW/QxWxxxPEeym+U/8SrsUompuQaU/vwoeYskIx8S+7Oae4n4YYr3ynioDNM0l14lG32j2FIWYI1
IXralGaEe6FN7ix6ZXn0dDykvZz6vvrjmVhO0ilY0snajh6w6IU/NvKIFCTLs6+VuNv9P7M3/6aj
3IVCQearR+QCaaiSQOJaJQLkwTSj4DcC/Ny2KBrKd4wIVImk5crZKwRPuOoDx6369NmHEDxmcLN+
vV3bhorTJNCLEne5yk70+S1gLoULrVQFo6DH2SjlYeOOt9zi/AEvaS6ude6okQgxpY78/DZ5Wbhe
u2jBkJ6+aMMPT7QAVguXUmVkll0SpfDmmFSavxtCWlcs53NCjCSwHkob/Aq9j3c06G1Mz+tuwQN4
2tX5XkJ6/4IyswTaMTmwdb6q6mVbNngCjVPnbob5rlKEDMdxfTxVlDSiUVWzFSNn71uLkfYj2tSr
ny82PZhVYk5IGt5M5xyruVLo6g0osOGvdsjxUzBgcWwtqHGRE7LRURi7M8Va1hUB9ZMvXw54Rj2g
FooOYbDeUk0VhWwVRIaWU9D+0CRkZpJhB8mDHtfYLrE11VxPXNVaebKUc4x93++GGUHuFbe4Mpy3
8Ev3JgFoSq6Vx9d1jmW/HnYqLp8Marh7hvrvvwntIIVtPJpxc0PM/jM3kEK9bSXhH8fJuUg8dOr/
7EBiwJrW0luRXAfwCCk/xsjGdWOXu2ftLprdoxngGBwxnQXTIzIwka43FHW64INN/g7CC9UfNzu3
Q+woUvbEX8yjiBkgrXxxJ7otNaKodY4cFAdaIjOHXG6mWDv7EFRkkh4Qe4gsI7FXyB13H0tcGDOf
pVc+1FdyeHQuVu+bmhIF/n2jGezcB8Tt6DN6ZIWs6u6qoL7jcOQHBpoYebGpHOqIljF/rfFr4T8J
MRXU0oA28kiZLG4Y4/kwxqx767CsWXthm/V/2YTt85tadX8S6oFFVmGIo9xTi4wYiSyalzYCJjUZ
8+SFtZ90bT8j0PS0DYBIcBcdcEKFuuoveBALI8uzhV+mzuwAeeNOf51dE3sT0Jhkg3/DwzMg+07u
KjqcR0IADqGfGmvmVa/40tVecDMpMLagV//rqpEVZp3S6QLADgPjLufChi3kgD6YNJkV/Yi3Y2jQ
XazwYdfIR/bBNijIFe6oynqTHoLigvjgntO8Gj+XahAX4W2gnMPS0OUp14anTSYsZRtRJonxRa4t
PrnP/DpBrIbPj856ngWcEcds8OJG4jzmT24BsLX+X6xJcBbV9EvdxvyhjVy6WQdTNrWoARpRApCJ
yixXQ0VmAg+tBKgKwSNbQZC7rCRYNGe0JXBbrW4KwOsSkt1R3G9Vr9t+COzIYB/+oQ8UeRWG1RtI
fObg1KmckC9WphJ7FXNz46bKRrIFY2nTZD9i/1+XkUQtsVh9N4hEMqWL8WDPhNyzB2CruZNFU9OL
I3Oh8rAh0/a1yxpwn8KF0cqHyNyGM9eWr7Rw+h3aOTxmhRqkUdL3uywxVXUSJT2SgJPkIhY09v8X
ltUS/e9f5XgleIcRYamKhY5pxpXyAlDLdK2rWJBvR974Qb5vuLu0AJPln450LIY+5iirNnTMyPCO
GESswKJRaHhn/zwdPBiK/qnq6o3CdSLOfp/oEsL2YDLjKuB2iCRLz08kKOgqu14eoO6V0Vm6t+tn
BGAudbc3F0q4fgSSlb8GaX+LDGxSlIMXAQNGe3XyVlxkfXm7YatnYGPiC6984bQCegzWZORUfG77
yHLi+pQi9mxlEaDuA+GLCZFIQZ8+LDJlVJs3HWLWURJ28+6qK/stW1eaIdEN0mUFjraWMTOwGlbr
2qgtnVhB2XPSHBC26dvaaBVcfhlu1V0dqyNobaQxFqvaOnPUF/thIsctIYhO/XgWX01AqUre7YAg
5sPZT3hPjUwHlelVu5TlVhM/5a1n4hJQZEyiZLcntw4w7dM5wv8KNpy0WVMCKTODZTGDotsKtIXY
7Goj4uTyaqbuD+ljjpimPJsx+zaUjlIzIlZBlC84WL3TKOMpvJBNJ71dd7bOw9BRQxU29xS4fjav
u2OPkpGGuerXllepoYFShIRybx4qoZPd3IxyGbWo/x/Rk4dBOVWxLeBXcIheEF674DNjPM8BqjO7
SmhLRmutd8O72LJ+bA4pOyoBtAjpI7Dwr62LxfQmJaVyFPj++fL+IJk7cLE+FIBfdL33eGHoXeOc
KCKSFDTuxXHDHHA2VKAMbpuVzKKruvpto37opvMG9yERmXp9Uy3fN5+oi3uOkMyA9nIzjmW7olbR
Z/ECwuO2B60ceTlcz39m5fFpXMergeQZFYIAnmtL4GzDcm7g0NYzlW/XT8cOq05nEKlhGymmvvul
pVOHPqTYRse05zC/i1k/fdB2yGL0/u5VvA7B3QdjeqEz3iCF7Q/szW+So3QWBKU8ZvcK3p+BUXzM
CEhnnzKXQSKsItRLVUnonqsxOpyntwpPKe73aGDBTvx0nEnc8pL9Q3qY/rfKkYgxs8Q3sa7PEH5t
2BzJvolfqX7lXtQXEQyClKE84hzH6DzBwfqF4xJIFex+FSK4s2y1BbfDLFwBbmDpeB0WPi7gMjVX
SkOcljwNfzIxzgbhw4jOT6YNUceU9oT5Z/XPfsnEqoIlobkRsWSGIEzN7zyEnAJ7ShX8kFBBgj7Y
wAKr/q/6wCX6/5CMuduPpPG4YRuj7x6PY77dAPBwmc5u86qo0sBnxEMeyQyypPBs2QnctsqGb1Sn
HI3ndW3FgEABbAe/03DY2MCpUuTR/MtbyImJkGB+dWYJYM9x924t5jM0AbPCrhG5XiIZMBqscVO9
TRZ09y0oAQyWKm2Ym2JT+66/imNSz/AhWQQu1cX+uG0jjHCSlTsO8XU/YwIp+yfNnAGWnWtABr+9
BoX1ktvRhzjyNAApA8sZMPeap/5dKYXX9j40bl68N4rFJoCOAFv0Xus1NAnIhNEJAIlHx0T5jux6
DniAEHEbLskxyMFffjYZUewmA2KT06NLGA16W8xnv0wEtAr5Lpg2BmqpKNatZHFEcAAg8+3wHC4J
hk9PZ98200+gqzUrmBysbNyxYLT0Y7gXmYaABmxTXcRoyA3JHv3wyiOnG1goctiBePWODpsP8cKW
MNg7VWzpHNaLkiNsgkH8AAEMs3eYhXd6OpbCbCzs+TY6hNUM1sorblLKF0uRYUg/zbFpBqVTmZCu
zJaDSARmPjlA/xXw84xNnWguyCBqQIDlHpQDWMbuvKcZwrfrAwiG0kgf9PHvcWPPd7tcyLWuOd7z
BWBJ5FHNuwVHnLDGpnSz9hNtx3rg25ZdWEtKw3rZ79aW7Y77u7KLjHvpwh5upSusnlN+zszBcgQl
gBv/B2tXDaTc69c5pHTMhZIATzxLPDWZeCL957M4+2AlgLvIUCyJ4OdQRqZZXTm0pFhAK8m1/9Y7
9jFmVRK348HwB5OO45rpoE2dTmwdgDKLNN9qZ8LRL2iHS5xALDXCjW6Wd1lmBVWjuzyJ/nYdCNl4
59zCi9N1pdQvWKiBWA0u7dxZo15mfQcyMBIKFvBaLUk17g7P9z5HgBJpqr0Y9AZKMY4Dc8/qr0Oq
Qrl65sjMlBynHLskdzAlwqBAuuirIu3QpKt47T26QQqMEpzvsRkao7QRP0LioTa/XQEB6yHgSYc3
mM/ovNMLJADmjgx5N8OYJAU2uSEKfNMMpHp9aRr9s+ChS4jxQ7z9wNMfiqtsqVir0UXS4ESMt7q2
JvW+/fQqsM5aSnk1O2fNeNtsK0LgxcO8vtI7Rb8LlJTgQVdxUMLtPAks2GdjOgXdAnXxsq9RWTo4
0uREaxMvI5satUrSXmAAOowAr93MAFNuns1NnP4uRxhyX0TddHQIPmE+ZAJSX0gFG+1huNlyBMpL
XoFbJFBNXBptkRkLanj9HjkySqUgCDGSn532xQC0nkxS74bHkjFfEVPQRGn+wwVrlUix3/7JHnhT
Ykp3R1NpvGr4DbyJJ5Pf0ue87ki9v3UD4DQBysqYdlNJqC+oKQN1DnC0n/MXU1fj1YhoaTT6SXK2
pFQkh5JjqQm9cvop5Eg/AEC6Bsmrfj8Ux2RVbDZYj0HEEMgTJUEjrPmCEwbI50lw7UyUTrj1niGB
zcnD3B+rFABNuwEk/Vk8/ojecPGXNyYNcsJ+TaD4DYohMWnkYR9HNDZYqIUu0LiB4LzoM9oLd4ZP
OEWT/6EBcmGbmzy4Ftc/6LcoezLbbW9x7BDcSgrloHTWAlTEveat8ax4piCuNlpZ0Q/cZDoa5626
w1OpHB4A5Q7b/SUbV9FMqUBm0t1o0sXxqOgQdq3kxaVR/41RrF/Wy59idpiQJ3FRNgOmtidqG9tb
xa0o+SIlKTzxjtQr4VhGt2wQj48yF2vavpMsXZYQlWg2iX6KPKOivhXY5TRBKpK6RtSZPExCCWOH
qwTl2UX7w/DBetQKNUhKZX8JpJvHzsEt0wAKQ8EQUjJGHFOu26Lv7Rjy6nWx8O5DVm6MwVr78Oib
qnbYE74XP854K3hOKC9Uy7uf14xc8WhGgep2AJQM7ixrsMrtmIR++g1Q3mdTirhJTIMDcuFjxFNh
bwB9ydqx7nCn9JVRdVtpRI9tWugEP9x5Hr4MgCU+Z4rng7/z9oYDiY3ru6/NPqvo0GSzQCZE0QK+
vUzsWUHL3Lz5sFq9bKpqXvE9F4lj1AmDqrK5NCXtUKzuLMwh7UJg900f/5jt6WrnhmN3A3SxEJyc
5PLEnUuOg8oDDi1CYXiCgJzQ98SN0Qsyb6CjiREsUffQHtbLz0nMLKS5AImbALYqF8KfpJaieJ1L
3tTdWR9qZNTA/RzXQMh6d0FIPIHHgc2cYHY1KqhBLEndemcoiof7BKTyVuHNZWfIzd4EzPIw/st2
c7yb4NxHXqiDdEz8iC7+pL5GNeUQMODS3SpYSjOOt98gWKYMPa0dtIENRnctBY5rJZK2FjUHDKKQ
Fy7kFvYdPZVsTuHmMK1pMKuNi3LIrGqwI0xKGquY3VemiRkPL8m4sjrCRHPd1TfQ7SoXoupu+ni9
kMaehFbnqHvBPIrf++Rv8DMEhsNM3IISclkLBJ/7/JFzlGFSRKrWfonnZNjUw8sPKcVttqGgZHMD
4i+IB/t+Ow3mdkODmzJOEU0S6XsdNXK+TwYVBq6MxSFEZE+UJIgcbHDwAGC+ikId5mNh/3CMk7/p
QhJ7wLbnVdQkhOYfDie9txYZix/PmnxbYueWGUd6N3DEXnTQnt7LDQMR2pL8+B4VTnJf3+MOE2Bx
zH/OIy+XzysKzdMtxvF52cy3XN+SSLqlg5iL2eP2Jn6htFKQxzGvmk8UJimTW/8nhCDKhAO1BtPH
Uwhj//MutLMw+WkD73l+5vvFJcvbYE1n3FAGgR2PDfMQJkb/rg0f8EL8TDY67KWgKjbEOQLT6lq7
A1NK5SDb+QmuDBN6ORNdgqJ2puMPI8pTsZOTDBX2zgiuOfDtvYqaTfUjAWeGs/f3QNt59/tOy8uN
FB71emThz8p1M5eJOTlDqZp5j5NFWW7H8Puqmi+YkgoEUzAx64MR+lC8IxFbhTIW/9MNJi/NjgB5
5dkSp3m82a2mFOKvlSuhZwRNM9hb0GuWnzbK8tA0wu+5/YTNFAkF01jkcDLN4Xul6qmOk+oKrP4l
iWC6HENsozbPs+MccGlCWnLwcbj3Idkem2VmWnH1xoo6w59ktQX3nroi3J58zAx6Dw2jh8d0AxtI
IkK0FZ7jW1nyBjTwl+ftQhlh8170KvVSh5OGGaz/C3neC2cDVWgu/ZFiq14zYpn7krAV4SIAMxv/
+u45VJFjhvmjV0m1GYrJ8A1Utvxk+VOB6//yakfbEZuBpKSQefu8aobaYIcs9/aSyQQOtx7YFFnw
mi17JqQLWfbhcRYzU3MoD7yYPKVW+VcsztgAXMcPiq5c9wsF9qzWPSAsTaMtHmT7Jv+GTtF83A06
WbYDwLfBreXIz0S3tuJecIf9qH1SbM9k2vJIsBssvURZ+jgWUE7cQACUl+jaw1+HExjzkm1hjg0U
LtYE6DK9PhfiKPAbmOHM7IafsCZp/zJuzji+ELjfXdG+yTVCzrIGWoJOF+GFneWJKpLOlE0bKOx0
9CXGLTxfO6D/uPEMmNgH2kAiVNS4G2y5ZWXAZUNFj+pwVcS3fVZB2LhJe8LO1nAJ1u0f+qhhHbxP
b4j40dWenSVKRsSh1OtRowuYN9ZU2/N+Rixd47sJX1KPHKVPg5Zae9MsAhaAAQwkUsg7Bpa0g+ZO
k9/iMQ84aRUqGDwVuzzyb6cnCrVwSbr49Jvu2POo99jvQ/34X2y5YkHjWmVP5DNV3CFsqFIJalUP
J5P7COIhQawFbgujpmVWAgIKFLcEjN4pcyUsZbrZHyoWVUQfbmUE7fDNbJ2QMpuPbTKwqO6M6zej
rEGT3qojfHyx9Oe2cQ5MhK8IUOhWhi6nWKc0pq+gZFe05fy0VO1UPV+UvPoQITEZ5FnGxQQTILzb
tnoRxkE3VaWaXOTdgAATpTLeaO5GF9V/Rht5015ST40LA+rMtGtYUYwiC6JqWmGOzVdtHvrYtufm
MSxhgMypW/o/Vl70qgU/ffw+qaZ/bYZD4aqfoPnNA33OgpOl54lmreC/Yyq29057uv3/zpzIBpwR
n9VxwIUF29V4wphuotOGPj0HFgvl5CECcHBYGu1905P9p5o3kSeEAM86tl8Ny2+bJM45PHSGKTIE
bE1gP7UzD0eIivucwf2QMFrg3s4a4BtTXkqOPzyI1ePpDpzMtY/jbvsjw+kf7AR4phNnpZo2H5h6
6RcDDx27UmqEunNgeLB8DeiU6+jKzWaepPRlcQUVymzNKfhP52j19syI+rfhbReD7eOWctreRvzu
UrIN/rNPKOwhdBQzPS4hG4ndwc+CUJ1tXj4CXExWWWdH7HoUgxLqnL7KpIeEyHSkjNpn6VE44UM2
HcDrd6xPMl7v3UkP+C60iY0EdRfJn5qVWRkAFRbWFTNWATg3U2aplj5fZZHOoiTaKHgqM8SnbSab
Zs5FwbagWSORdBriKLWYTRo7n5uidh0pMwZf5U4xlRGRo/BV2WmxQNnl6ZBWQDdjWCxwJfKBrrt6
c9GhN55rk96pjVKT1+OMQK+oj2Fg+sMtalQ79U5KkFBH0w25bGFX7hPuJHeEeadiAVXMYYIIznoY
9eajFpFT3GTvNA6eUBithXAhiaqcaFMRqqFjbdlui7TZJLDtA13pZ4s5tacJUGOIvxkFS4HEXqss
wGaY+msy6/F4jl5GFwZGO4FSyNQkp+SEZOnl8UlEAd31Pz6EhffBLdBmSt2ZBtydA5cDHsG1wXm/
QUvUPS9mvMQc3LsRawPuXrZSNRoLN+fcq70yIQylLTZcfG6vxTHWVbimdnewOLaL+2fPFgI18wxq
16l9/Z2I60oVS3g1+AyTq+IA3z/BFf408XYKGxnc+j03bkIolZrmk5nsO34sjD0TSYjKFeBUpheA
/HLyjpmBU0cUOwLYqvGQESe7SvOd2cA7xjdyBfRkJM2LTJ68nyWn+X7VvRL+616PXMK6ErfuHS+n
YqulODjVrc3gnDR63z+1Hj62YxophenQUSyn+IY3juY/GO1uHrwuiU1Qvcw+hTjqSPOe1SXxZZH+
d/l2hk3dIjCQTKZbJp29zuC6+SeMnpfRTmaFuUqiQ67pdtnfMlzcmwgUfUzDOUJn3QgVBjR6GBst
/QnH2vN7TkpNnZueOYUU2ymXUE6zZj/IcFJTjm8Lu0YUnBp5/s5KQLdzRIUZsUFCOZs5Hx4eW4cO
WcP/m27YCfY80/3/eLFfdBxSqfHdUEW391Q0GWmsC0tIt0F0DPeGGQXLyBkv6Ra255bReAg15CZ9
FjWxpd0kIk9WtfvRN5sPlg05HM5Y2zvLGACgh0zCsAhJc8y+APW1FxsR0vkeHb7XGj1U3AUoQbda
fs3a/ARwkASbP4S8onJdcse0tIJqnCEjmUsNEkZHF8reRp7jLD2cmn36SpME2GJ9n3YtEW1+JMsD
PdyOZvF1PiKnnU7o9S2aTRXyjTFpNJ1jydCGrB93tddK1VtNFdLavyw/5lIBWsRa/g0XB+1Hm2jt
nhsaRXTD9uQ9oquNGIRXJS4H/yN7uewGFOC5dQFYz1jfxcU19mK7dtgLGn/4SKXIvTBOWL8ekNkX
AmErYc7X00Q5SEq/1On83nqegbu7WpUXAEOYpqCebVjahhN1RAcMpYwiTrGbWCJplnduqerqY6NZ
kZfwAIMj7pNV1RAZtjs42xOgM52B9p9OoH9QEOtaiyxQSXgfHxCiSjQOWHMEL0/dqeRayY4V1Kcl
urMbw3NmD1XBtlZO0G2tpsPj6fPTPlgym3AOPz65fyaE1Y4Po1waJh8sKgaYBzsLTztgWeigem7Q
hgMyeC/otgDlh0SX/L5EyRyoDWwv1ZNAw4XCd/WzEIQ77A/TxDfH80Xz6zkSBzTunwXFteePrTij
r25Tw1BbGQm1hGL0rqYeV6FWCqY6jG1xu8YWLZVyXCSgb4bp1CYASyfphUFvndwMpSmjo3OzDmx5
9a664bnDqSNg0A17Us8f6O1hUydCSgBDEDMESnww3JYCNuyIxAKHMdgdfSizN9fqiBRNQuDWg1iA
NjjQhnzj1SGb0sGWcOOn308rs25yhUlm19h9QaMes8dDVJDJRgLorganddhO47BsfLVT83P7FK3h
9G12l4Bv/wD97MLHZho3Uo0xvSf4Qqd5PIpac6pmLWvfVj8ZXN7D3QAlOZgasSFU0vlBsVeMCFhw
bPPGJFKe9zNibPgTNIWMEv6SdRWZZirxIvI87fN4B4VtQ0X3ihwS+Yv8nZfKZOCiQcG92qG+oflr
WMx29OXfPuc0qT3ZRx3fE7Ynq3c1dAjKSTYbgdHNW7PPM/5UC/xFDONYyLa9kBVAk+uUy/gGKV3K
w8+zMzhJqXNCJiWifUodUZzQhkV535zMAvwnj9I/U7oit42nWmJMkKJg7kNGlLRq+Rso5FtbSHPh
+e64d5UIbWnibHwXmwmSfXQtlcB5gvpies3a5Y12ftVu7kPPn8uzILi/crdWzfXwiP0esQhuKE0i
35959BDCx9yzXyJDkOFkPfwXg8exGqr4yCqDTzygeFgPcyt+AGVC3InZYCt8MYlcb3EIEgJJ4tA2
DKy5ip4Sad6e8UVJGd9KukbO39YNYFEFd8ZI5q3JN6p7NtHg7CJeAjYwFVroab7I2t4S6W4c3Nkb
9StbRYfkuT/ldFo3ELaNQhkx9HA10avirpXK+JnXm7ebi/Dztjn2jQgcXtIaEBv7tdLK/rzgyTZx
Zb+nHWdvNKKrP+9tNp1aX5iULxBq9byRSuOmlBXSDLu+QZXfJM0iIAKBUUDCAl+7G2Ff3Yl898Ur
tahCyIqEwHijuwXeBNQTTyGuY7L9WwTWLW2Lv92Yx1YFqKrmHUhrbxFiuKxMkhyDlIegFzmEOXG7
ORbU7ibSRaFcEFECTgcWjjPcqw9Lk3u/m8Ih6TsnSlU8vws/yC6cxWK2krX+aARjKVM1wxsYnzQl
RT0YYLGVwHnGV/oi0+9VGetpf1Q6o83KWoDYW7uxUQk3kmwOg+DJli75XreJG0UhDL/1dBMVXXvd
MKv09XV7VLP89zhymuCcjUjHX0yxsIpL+Jb9K7FhQwaek9g8Mb/NqDWujMHgLdRJN7KJ2c7j2Wty
GrOYwYt/PQbt7m7miL129gbQIpu7dwaBNpKrNtR0HDGClTUXCYpJIZXDA+wm4xx2m0SSykKuHyVc
4Z1tS+bz+2CK9uRaaJfL/mwbRm7aIjN6z8rGQsqdq5G6ooAhBkaATwZA6hWn2hkjcxgL9+1LnQ/e
0ycUvshb4YbJTJ/CveCKzw2m3A7A7c9grTBIqYvf+M+B7STDEdUUE3qbjq03lqUcdY5cCuBCC/EO
J2ADlnMbMHetq+YBHZypjZyj+pXJi2B5o7H1JWaeUGl9wYOc/2sd01BKtK5v27WesZWuSLHelmhL
f6Hd1WHq3CqgONGBL3y8OB/fibW7zbioGKGwB+OzihBIqGfPSxZOteDQJetSRCVYTpPm87uicYen
NRqwzT/vbzutgMautQbDEq3cS4/cFU0C0tzGaDsQ62CfPK/sD8XoREx3WNCsgoNZAWvh3+rvLfpU
wMmEjPrcb8nC5tlWlOxrMOCcmf2vEz7XwZ/OF0EL+nhW6oismK4S0gq0x3/L707TeWagY69WH4a+
sGWUotlLfHWuV01T0mTXalK+nvnsfZDXXzgBm491QT7qqMkjyXkfX6QnScRqgDnUEmYBcanABh2I
HG2LIMDWAY4L4MmHbs5spkR9dvn4EPsH53ahfG/qq2EatFvG9Qa+2cXIz6D0svSYq3RB0G5DPjcR
nFlPWrJvgOvLlnz7RaA0M8sayk5HUjs/HqMapHL6jQ0dp33SIIjJtEOTqicmZyuLVjkG0z7DH8G3
B+vFGI7P0nMjQF/xt6DB3bz5sd0ARW9RLIWYlv9esLv3DXUNDkFsNmm3G63z363CZdZvMHKF8pzU
V/oJQFdVNvmZcv8Ub8n1DnNwwycbQjaUUBxO2BfJ/6r7TARt4KGBBz/485e7W/p4aB7/ePtWXFZ/
SYoFZ/4X8e4qJTx0Jyph7G+6zFpQItsiWNT/VIxb862c8GjgB8Wf++6nzd0/w1XJqkIPLwQ2Nqaa
+uVdIraH6ad3687dyCD8U0EjLbamINIoiW+F510pSj7pO9mhLY8YZV/Q2N5XaIEJruIOLIwQk+Re
2SLRNXvij8vkWBuRCfLwLBs+Uu0xbztFtTUK7e5TharFXiQ7VoBBPnt1d+wr5rT5Pzh/EpYVUSsu
/dJW6U6M+mFupJmJDkVsbC92+EdVtvnm43Kc1AXlryu1aGaJNjuujthwHVrwCKdaDxIkr9yu5ncA
y2vxBgh2vY+RhwFrwA/sioI5twDx77mpVr5Vhe7SN4/UFoRDdrGlNAtUhP1fVkRcQmwMkrD9GSst
wY3PYkQJnIy1VErY2EazwiYim4kewyawsTrt7Pk/NRrHZ5/KosqfQF730BRJXDtS5yrCYzlWy/nI
oYEP3YPGlSYTeknEN0PnDkOZMTuQOWWOpLufIuc9yAzhlM3wQPo7SWovmVCdDgLZjxt+BBekD3E1
7hZkBimcJJYdlJZMB/9VRkPVhc5uXpVgHDAJqYculc4N1aya2fNiRzEZW9Rhk5zYs0Rnw60Az7cf
3bTBYBXstKq+Rt6SnL2ApqvgJEz98CwC/BauHBZZgROlBqofWmpKQ/UDIxiqExbFMF9FzP8WT8dX
e53ztad2XwubQY9bTuPnN73z9CP6Zfg4znsbkETn8zv1E8pBOlcWrOqkxaXodOS0TNF5b8fXjsTd
QEohpu1yRy74N7cmZuaZO7qwRf05vi3Z8qzPlQIEiPNO9/fDz88H7WcjerhPdDCvKvyxTtajLgzD
UOmmSAXfSNtcW5j45uPVp3gbUOwJnzxtRX4+8LqD1VHy3R1xbosePLN033nQtDTiH+icLwulTy60
mfZ01smqsNPwvjkUWlc7LxzaYOyzFjaWSvXbb//76dizDdlReW1gAabMdusBRrguy0JAi21/SvVy
Ug6ZyLtq2Uk3VWIEuxtEXx2vLaApSEqu+J6mRjBlNvvs7cY+xMpkCuvn0lvqG/4D1kyTvv/0aMT7
Kun6mFPYXtQKFA01PnbOvvhqXm2S5UfcDVlubNfooptEZFd84pxwolSvgvjOrKTBKtW57n5C5eab
57HTna/TDpzskGXlCCsXhHdpR9SRu7/P+CDQqwsMH0S6+WJ0wnN/7QEhfXnT7UN+aXiUlZv/YIqP
PeCEUYbdb+Rz1bzhSprvXHebrms+4o3iF6nqHE6cyTfI7CJW7lvmurTbMpC1I3ZMbE+pNC7dZQH3
LczAickvIVGIyxlDJNJC2iK5um8193TM206zhKmC6g1YIt+VP7VwaV+huUUIlhty/2jkJ73iRdpE
/pWwv6CQROtP7GaS8bRaFmfEsJdGHQv02d36NCHj3u2bSdjJwmA2mWL4pquYmX8wK7xOUfHrtyPJ
z2FJqqxHMVoY1+K5/oVJz4TbT2TfAvMCuR5Htz3TtFuJdGF0r1gfJKbW4y5Iw3DA+5wu2vn/anR8
at8+y5uCM8N5jHKMwhgYREFn4tVtANsxHS/0daYaDfCr8p6e9pfMAt7CmNP9HXTpnfQ5jCZRn79F
Vwiz+YVI7uQIRkXafUosCdDdVXkAAZV+ASVUB6xw/ZNpK/nJLVmx3I+PtUmIf+EHA6X/YXvf5Jni
j7Vsx/2l6ax1eH5ZhnvlcY+kBpRJM0wXVAQtVX/bu4RqVrZtK6gDbT7YDBoXAEffxSVMVvNoKXaj
gXskmus9EbqKT/NojLYFNtALjLNJkI7fsewdH80Xc5DnKZss3AMqflAh6VlNfhVo/WStycpnBDt5
GpGe0drhnKPrPaAlT234G/OGt8UVy5gtMqLhQS4uqxxh42S8F9V6GLlaUNLlJecEaNGgEvykEBhQ
xbJKhTJ/2GcmmEozYTMmWMwWNxzRjn1VdMkSf6Oalc6lRRLCWgNzkKDwranT6bYx5LQzOsJ5jwqp
UQrNqcxAbOgu9RfQTEK1aBUHXRlz/Ir4z3uwxbuhLI2VjvorH+XW/TocxlS15JaGThsLB/PtXLad
s4tKgGH7wJUGng9iDr55DN4aSQHwWwcJW+9hFB8yFmhqWORJqoC7ke1/da/BeFMfSt02N9aw5dOf
1Jyv6eEYUT2HSc9n+2fxnJUze5FmKvA/8U0VUxzbHbZcc6dg3ukvbNz02judzBFLewYa9+l8zSau
h651Q/VfIGzslZ/s7WEXEyRxJzzexNmQzjmrS4SaWSCefkQXts+wu8VAAKtjlYlsSb455tbk9fTB
KytLFfLZERwNyYXggeI80teesL/ETTvrodcpqUxC063qa/8l8juBzqtD783escuBGW8ETlT/aFTZ
iVV3EDuS3mjyNUbOFNNHArMnHKcVfVIO18k2IwfKASn/hg+zl2uh/5JWgtPi2fKVgLpJxTIkDE7N
PinaqW4aZKplGyr2C7e08tk0ZxCS4srR8i3cHjlWpZFneazYHYJrlf5bJhZ4Tf7+hXvA2w/JNCwJ
Xd0sFfiq/2x82D71YklRI4HuvGUA6Yax3vGFJXy7ktJXmZDxsQTDtzUcKrO1Vm44+A9+/vXNPQgd
9Le/VXmtxmpkTXtzhYv78X+g4ALy8noR7qoxCW7cZk8HnBRjVNPE2YLaid2iitumoDRerixpGyrR
T8nxekRbrJKkvdm9CvDV2TDcTNitlztCyWu2ri7R7Icjc+Wq3kfzMDiiz8cx8cwQ5IL9KquV0Ih3
NtOuhuqF1TKJwNC6c6+9Cf3BVR+bO+nhTt2zEJyr9+Bzex/1L2H2FmSlqrgbF5aiIM5/B+sn4Uup
giLgFXB/g7qW1ZKf6UeDtTUq0U0jMPxd1M5JXmtAySms2nU5JI08qn8V9inDM4Sk+C2mXpP80Mp9
kwP2lvxRp5eNYqHPDrKuc8/0uhphFyBdx1wVx/qhDuaTnaFF7ssBCg4gLwZVY3aFHUW7tk/WuZIk
OUMLP4ly/ii396dEmgECdwfEQlLkbEuQMZk4lRQ7lCV0yPSdcbYvfsLPrthMBRUJ8lL8Cu0BACfq
mRN0iGgmoKoTwnVtAj44zwTUEpOhJ5Eb95YasLObsCIcNdrkLMRDi1Odlj4C5FYkEnBjJiWYt/hH
1xGh85Tj1QslpggfHkbfBPY7AcnLaCiyhHTPW4FBVA3+QxjeYMcoOeI+I1V2qeXKcn7stuOAy/6/
ePB2QATUUZxZBD3YMLxkGpfWBe9WtuujaYMVKH5Z+CMnmBB5gYo5Tilauhv/l82GXSVjY+VyUy+D
M94sqjGKznAYzYwzGNk1YMyt15L6V+zcut+CYEWxNRdCyP82qcZ46Cyc4TbPk7SR/XV1r3ZwM50U
tPCLPXL0e29DrlqPcP/kGR9FKmEvhtKMmQ19cVZMm9AVx01ivPyRiKDpJuIiWaWL2NdDGKF+XQJI
LsP1lanTaIfy+j9XwEQUhVT0a8MeD4daG0CJHXk/39HkK/kV/CgEpwM1eDQX/zcJx9tgffF+nQob
tyLUTbkjPNjI6IQvD3JO/15BSh+pkH4/4imPmSQCuienqsy6knF4dzA2JFihqcSmeTD/1DgsHOhz
U8gpuS1ksmjH+gqNanmG/gkk+UFdJpDlvzKealGjLCWWK+73XGMydOWDqld0YX+2KbRKx31leO1W
ZfCAg/+3z6G12rUbrZAplyPF899jumObDps/moJ+odSaWGIG2R7ulzyOT922wmkFDUYnjlwI6sk9
ZdvViHV0q+fuMdxVnBDDdbetl+9p1lSWQPnqGe34ArUmnXFFnMECL3powP8F7uTtgZqLwDwBefZ7
THmiPJ08Gfuly94ZGXDUwlG7xZSx8TWT3XigM1xfOpvIMBy+cSFk9J+ud+v30AN9AVVdsx7UlAw4
BWFcyAWlUAkIpBeThDewZ2GjlqduB+KYtsINjl3Bb6PHdkvVSfio3Owimk140+97jQIoUISaQyJK
Msr9eu7HDB3tN8ZzMd4r4ERX3yKRpajaFUeg0xq0xJg2i/8gpWkxy4GuIgWVnmH/QptuLa5OyGDk
JyinaQTPfCOc4j2IGasbvs+sn/p1Yj2Zng7otur4g3pyyjfr3qj0kWh44un0CA1u90OyyGbnkpNp
dBIc0B06lQ527nRdHVSH+ErvyLz9lo/o7srT9nEC+UJ3M7duNx4xDFaxxGbjtEq6ANu/Qxhf5Zy5
eee6ZougMKvsQR+ZgL3Jo6enh4H3wVNoJAo/IRmV5WSoBmKGJ0DsufViKJlhK2mBymXxa22ndlJU
BaZR9BUWgsMOBy6we3JZgmWBKYaw8/Rkajs9TY49pCD42Dut9X2+QdumP4ArhmL76rI77Q8YccY9
x1pkaDIUOn9fN/8bmdk61PHd46qxNy9DtnwSKhWaQfbSn+5m2f7vfeIAaFRRRCVKnMKJW1RPDU6e
Jokt1QvCLFzfTh2pm11J259vJEOKYTJGin+XpDWAo8iQbEivCnJvAOdQA13SXIgvIy3cdD1fJ+At
GYI8PfT2LUAeg6AWMJJbUCsrDB3ZDsPuZZyykAOBtBcVMAeNnaP/wJJbKoP7pGTP11Md6gBliWp8
akcmafLd3+zl/+0DCOl/h9wiMKE9WJ/Fzu7kc8OcisYdvtCj4EqVTSq+cfIFKF2u3jQR01MDAf61
w9M+kTrdZ3d+UfWbtCrUe4l8BhrD0X0tSQygRUfYfvoz7DB1P7q7wocPweC+NcMLO0ep9L0ACixu
jUR2UKQZwSlQ5ze3mMyUh9VV/1fnVSm037zqnu8mTsxf2a4b3NLF07RQbkGokz9LuOFVhJL9vBdJ
hdnHW+QeTeuP3YbYunAsbTkX7Ml6mGKko6zx4PiYRhFY0l13pNIhiEihCpkAObV252TKHr2CaqaI
KNPOplVrSOzsprVcZ5swjtdCLl2B1ybEp2h0EvD+DwY/3GNFtWSEsR3Tq5dpx8tUqHXa0AxtA6ga
0LjwNxr7xTh1cRfiiSe3sOeY8TCRXgQuDjvpjq+XT+H2G2+3BYgL0yntl1d70khMAeMHUGU4YPXm
4ovfUVqLbtR4tL529NMYHmtcxxoosL2ityQ0QkgwtciVKnA3OOPAEtCJDiRzH4tgP2JRzzP1s0Y7
q6o/e/TxrRMoxPfxCGeuC4qAuJtvPF5v/vQHr2Z8aVCviMT8N3RFVKkKXwVPjvXPq8GW9r0Stogo
Bh7Yjc0toA197C5rZlxvcNyF28HL1X9i2WmYFPhf21Lk+6mhgl0wBvFxguzh8UlsKnfel4wXx3ho
rqqFlQhSrtMjcm/tfApVebPyR4WZG5BnPfFb5/CqKqVfizD6fwkfFhWlKH95bgnRGbY/eqEI9QdN
ka7paxEsvdMZmBg//qmuhmYQj51vK7JP9jmEgVtrKMBmlEA3Q93vOP8Ci2MrsOY1t5b2Q9nkXamG
8UoDAENXcTKlmn8Eqdzv8jS/B6mzwUG3mlsw1dP/aPuMO6z3tidJBIoBUSdlb0meodJVwLgtqXwg
qQkd/8bkcakbKaP2bWgLK3yQ8XWoUuJZjsTYdnrn9/ZQ6mNSCT7zvDn+DUusZ7IN/jd806yoXuOy
NepEVOrGCdPk2SwMzbFUPPBaUgYjBYoeM182hOLyLMZbp1UOII37NEg9h+p5DX1iCAWajZ+bmBPW
VO3dxjDOGEQKbA/u+FJlhw7MfYzhK8G9aEbhI6nUXWiPHTigDEhPfXHWj0s1257jNnDKtdHAxZXe
F3fJQ/iyZkibnTkRAp0KrQor5Xb5/KE7Pm6UNTbVI5Di7JO2S02eHW6Dyym36fP2/D2YK/6IM2Aj
DvKNI0Id1OPMPFxtPQ+/jUwLw679PpOVHEOxNb0doR3/VTvi2xEoGjyjY7cAwCyX8sFDCNI8b2N4
MpWXlKMDCKBeA9WT49ZNcllM+LTGkVZwQskHenuu53UnJ1wFm0A+ucozhPhp4+6/End1whtgbKY2
xySQ0R9bKurHgPIUVvStfL6r8GVR6Sh7sKDHHe02NQkfwwFYMlRYCpEox04K6izSBhb88p0M2g+0
76Pw6MnwlfzzRdzwh/2obe5Lty0di2IdDazuTeQmJxf9OwsY/SGYj22u/90+T1HAAtF1Q+X1hKIo
F2zc+BE76SDTuXKLqgC1UTchgNQJfActjpAp4ghxpPc1egEMYbNuwWbZQzt7SXlFPiJmTdrdKrk2
GfCwc1aRFS6FBbqitcBe3/El1b+jwb03Ax1kFfSisLw6elEYV5chn27om1r3uCZU7a+46jO/d3cO
x7Rbmogg6CmLhaRiFOjFASBhXK5M4xqhSLuMLcxRlwmddJzeeE4htxiHviEOZEXE5qS16u9znz4F
m+MCJIxxqIBslWpbxuywcFYs5fXuasu8CBwATthDMOBhDp2aKWu64Haif5gBRAhILm2/FzR08IzY
NoWFfnxBwMhKF0s/MZqea0IVx/XxMhhqc/p7OGFznjh3eVg9qrv5zHnnRx+v51yJBqAA+FXUCosr
2M7K8XCkj9x10fE9hTPLEtQE9OIPS5y6FaPFoCPa89zhHGaoI2DkZ66FlBZ4ZflKccT2fAwTu/on
jSrbI2/hEQasyw+RRkE47A8kS/x/NO/9xY9u8BP03jkzVUs9wjf93EVQmvay0u+OZjTUu8PLjYnw
eUVB5dP7qJaVs7V6F1+B0tbMQFhXWktW2wWYgr8DEzCTmeiJLxZNRkvtWN5kFxyVlddE35QMh2DZ
lE8p+aY8OjUTgSJdDv/0gpVNsBeOJocBdVzqnrQ/xjwBp30wjb36hZJfTPOiqrLktmkd39gOJIdH
ApBZNC4WaQjKDQFLmhdMze1UV/G9fGKfOsyXooN3H65S05b6JWLB57VA9M6kt6h+zkEMd3nK0j35
jSLrx9DahCOoce54YkkxtF7rW0feHOiOgg93As91f41DSlJw1ITrOApBvpLs3cpRVW+QcLKC3fzv
vOZert6A3DRzksgZ8O1jnDZJUBVj6x+mcfiyg0ntUXprchd/WTJNd/r7kjl8i3aoaVsYrb56gN34
6CHunGe8A2JGrNsSzSbgja/mMVrehy1ByUraWfSCvhTUZPcwmgfjZXctBFZvOBXXxUCPmxt+rkRJ
+MPc5JxxkL+hXA6gzvbIdIVE7ubFwtOcBJlMMd5u0QAYYOVDGTwVh5xPxBX5dt5AcxZFzhciYscb
rMGAIJQxmxd1kmFrs+u0YuiNNTZJ/8nUO8Ne94dIw2PTsW4hsna0OtWTzRmCVSjbgwwn5TFqlAXD
H41wVU7VQGdOC6JObDGdW7AYOp9AAc9ofuMhs0uN6AN4bsm/ARfFm677Gm2jIjcb4zGRSkTeu69/
e+sjV9PCTt/dDqvbUoZQm/QkZGfAeeA009Q1ZZA6v5S6RxmqbbF7t4XgHo5GZfZrJvp9B6nCfrI5
TEn3CrLc9sA8edA+xED5xiSlr8q5dJNhqFeSfct+DwHTCpLCzoLiSJ1sftWrFBw9eyD5Qh1HOafR
rdDp9wtBl1xDfojsBF9K1Z+VMewmC5bOGQtf/+stARgJ6PwjooadQx4tXnu3PjiODjywlUsqkgMB
FjPn+IahIuzpOyIO8I1KmowOIQuUmNEFeur1xMoTM52H/fcMZZNfxMHcEuQ8nGTMRBKgSOty8hA/
CkO4Mva6jQP1n/qn8DUYpVnxZadjvMNw+U4PftXIjlelBnKzOkGGPAU6d2VdiawikenGDzuvLLkk
KlPXwrWbXZUAanhmHcqRz5HdcxW1UOYVsZGUoWALz2EJAPlzpz5v2t+hcsdCLHCE5WugivMSOyvf
AN6JzSnl/OGHQwFy99/G/WeWqyqOoBnPR+uXYVnoT3VkH5p3xSzFmXKs6c+iEs4xriHU06FPL5zw
vf6mulaMpobZp/CQf/Aue+sz+Ynh8tsj/PJcuPpLRV6dYrTt3O8ECT0VI2jrXj3Pp5uE8EczTUnJ
x4mhNOOxbJ3OjHlAu7RC9Epo6Gd+HBVTTbxoVl35oUH5j384Q4WGh2hKxZXyQ6E6hkFo3MYHajul
lSAiYjhA61UbOl9bzBxNYOAcIeKFqPTGBEdJE7V4gGGyPIY2XdecNBkNAama6KYhO0dc2jzF/GX0
xX4RhVxSiFWq+K0JTLnBGaP5uaxU1QFHzoe9PJ5qbz9Ezwp14q3zQsnvVtG4EkK6N2QayNdAzj7f
YNEUpEDirQTHfYPxF6W5NOjzPbdpstORdedRgfEAhfjt5w3H0tu5hAb0MVaaFoI7te1QPm2Trzz2
gdLs/XOcPUuSOQvcz/oTZuOVrX5LQfde0NKqb5d4JMQpi+/vV9Pw28L2+BIzVueGi6MRbIsdI97w
/j4zTzmGXzjNYk4/ofd93vfD5p42/x+4X7Tb5quUfNakH2FFA0HHGK/hrX2tpPcb30ipiuM5rQV4
ZwxE3lwIOgPtsMzU5HmCPoF+8y/5gHDBI4nWYOm7zbMjbJImL2FQv+9LEbhJfG6GWbaZgmpxkMxJ
1Ov/sIzks1grDWxBF4sq7Odw+7vheQ3Kcx1LZQ1Q/YLMFYGd0dJNVJJWJqZbTxT6RYEi2ZxYTqGb
jp162FxCOREZckbQAHArL8qy+SFFaV0eUhz5r7dSC31PI7cy2OEhRmefuEEm7+TkuRo+cq7KlRlT
csEpPwc/KytLMYrWHGIgTpB/ZxaHwm3T5/CyaxTRCPFbiGvRStHPd0HR8uHUytH1+QUBQwSVWOn6
X7dsRhudmoLdg/4kO0Z/96QiOUcG+HUB+rfT396ChSaiNY5O4+Fn+JVwaTinApbjuO07HNj/+xtP
UYsOnjjCIQ4iRSmwZbyUlg36Q4/vNGPjEPiczyzRfckFCyAjH/mxoZnpn4VBSqFpHVBjTyPjnWXe
2X3t8t+ewr42Kw6IHPiVF5hcYme5UbP4aVejGddNJx57r6zSXhQj6ElVEihZ2Koiugjk/3YTlkJJ
Y7eFfGig0+IJUyDcEd1cIzdSMRyx5eXx17AP4CPqHn6bpQotPx/DHrfNtRIkh7P27Z2kVTP+cMks
NoaaMh6bI2P4i0mUXFec/4NpM+c+7X8emq4xynJoQUoHVh1iJCtfrOLDyFKLkU5Cy4Ob6MbyO2NM
WKW+BHKOJ30v/AzyL0ilylvqxY9xh2GN/TDlm3OvxhR4u3B+9tOQ9zP3Bh/KvGk1FPuB1mhGjjxX
4nbHzabi4HtgpWDSPhv2SoiGj4/obH36C+5HfDrwcjdg5jM5eG5pmCdmapQP2+HB5gQIdNaN+7nE
lb2DyIbPm3bI9VIzjVxSqsiCvxtlUBso6Ug5EPAiBb7lqaV/f7lZ6XPgIeFoDzmd5L02lidnF+HZ
I3DFKthakJMNnY5xHO/2BGzriQFaqZScfF/GosM33YXmltBA1zCa41kKOffH4qda9agJ0LCQfPXX
K9TUjyjAJXPuSDoH/xQFMkIB7gmnSH6lDwouljGbrrDLNivAM4WP7toy4KxQGwV8k/ezlY7N2vKZ
2IGycU/tziY5wrsHlsS7WUOcRC5pD6zCZx3fGskbS15kJIv5TL4iSbP4cpHaw0+XFJnO383jbXb/
qtsqr/dDMvd7/4ouhNgAVsZ2j6FFfc0As8VxyXViZ2JoRejHAULeEWFZTXnyIaSbAqoPvlljEL4m
v3G/qWjr7LyNTyo7yN3FDvVL4Ybi4OthmDjwqqTfr9IMYXnGVN/EdbvDz72a/H15BVgZvYfEaU0r
WSoiPoGNJA92FjV9fIDbkuqZhcgc18lar8EwcfDvztEYpJpj4oUUnbRu4Ul0NbtEq3El+HWZisTL
/90v5z6DDiMWipOYNBCi2D+dBzLyDTKZKaN8T7sDcbO4tKyoJgozrX5TJk82KxD03y64FNTdcVXp
/hYEIoCGtgoXLwjbk79wjrp/5372OC1ls5DadlsC4vwLGZWHHFu7sOrVKmxy4itP8mrL2ILdhptk
B17scrt3eh5HKBp11RZRqsaEK3nkfh6HiZjEn9e/kItjYryIQBq8e7UQBuFiCKJL8hlQEOWjvN41
Aud2mkas2s9zf0crPSuzao6thbIs0NS+JbTrXILNGN+KOLj0sE2nSqUOH0eRcGxTtkrOr257VmOY
Viim8dsZI4KtEFyZOLuB0bIDOvqpXRMxTEW+l3DSarm2ZlgpoTdwwqpryyFFMcFzwKfWxk86wW9W
pjn/MUP/ZXFnPHjhpa3/muaLu9HDP4AZhdRySRRR1Pm0kbpuYtyg544xbcBhUUtQHwxP9989piuM
YTxF3593pywjpBB4IHxcwZ8wfT/IDWpkrhs3qsjJPt8B/Y+NRaGNoUgh4EvVDOyDiU7Tr1fstknL
by4bZNAyrGshOAz+m8VIXVMojpHhfwGdKjjrImDm/b8xWnQrd4LjqLRIavxSCeD3XmkiKVc9Gdtv
HZzElnaPNXUwQ6x1IVqDJZsG1ZC0Ucu8DZdwnlzprEcTftOKp6x+jFaG2YhlD+2eSsbPQ8RNp0/9
Obsw5KIsJ14MGsPeyr1AlZ21187pN0P3/+2deTKAeNa41Q1syv1kVSCs0RcBteHZkYNMBHzjaBVt
0+2OowkLc2dsM4R0Z/L8Bsta6wSocjTbZRvtOYPSyHfU7euLrOSrfFHgMkuiL8eJ/4d+Z9W3tBGm
XuNuLx3jbFvgy93HV4zaoy9y/UE1XuLlOq8MMG3ju54aao854+4YjAwbDeARQlProgziwvjZtJ6D
Cd11uzgBrKUf3FoKsj3fuzVjDCwtsYv0Vzje20XdDIHqKUAIbtzprjJZ3Zbyo31Moi08sSphpBly
WbCXEeequQiNPPTh5T6hLPG09klC4kj+bJYJJPpH+dltVfy+CnkXg/s4+5naOizlDIgn7D4sYbQm
AaJJJpwW+foiJiLshfptmUg9TSrb7iK+qTbonXueQjySW5ev+2JA9x3c5/bEraN+2QQe1UCXkm3Z
AckaYlQ7a97SuXQEPaX8g3LSjPZRIvwg9TlOIJj0BdjGEvLBiVz9/XxHrH/rjwx02hpcjjyFFcZ0
8L8cjjsnPP4L7TwrZmVX3+urUp+AehQpNUF1oPnv/JaLlo8jsMyxkt2TZg8kg5Po86Wn80Cql7Vz
MBos0Otk8BIMzD0W43ZzPaxAp0mZsoMgspAJiwotzxKh10RMGUdpMIVs4YduCnEdugMKL3n3QLYN
LtF0qHCyWstTDv6AwnEo+mtI/F8MdYTkWNokSCisV9IFgxqjsOCdM7bIse6CIoXpmaOrSSkVuewG
zjYdsAQqDjxI6oCD0DtrTZxIVQbETyL/j1YTcAqRxHNCUcNmoqcKiTG2ftLfezvwxRp8BXIgaqMD
vg1bLfBowK414uMTKvsOcNIhyU6gDW3XHzs1F9Jixc4uGWBrr1aUnQ+kNy+1up4BZONjEbCwX67I
noLjmBQS6+iAWYs308eWB6TAzOcDoRgQlzu2QivMIYaVaIL6mZjuo8AEvFXXytI3MF0bwq92vhC8
8F5WRGv4J3n7tj/y/SxMVmge09DMAcbMx89F88DdqiDUjR+krFO7T7WbvXh/j8rPeEO09huS17yC
9DikfTEQ7m/mZ3WhEeoIDOk7y70Vc68LbJzdS/q2WukfajbT3MhZQvFcMUp3lUb4pyF+y6TAO5+j
8eQ8MO/vT0tL4csxTsmXnZKcy/PnrVl4VpeNDEfHBuRk613bwJXVpFDBnIJveEOjSCCLRwVFNEyq
J2SsC2NMBxNclgGzZe3HyBMBloi3YS+uWcRIzUx5XgQDRvqJ/SyFMOXAIbhYDTrWf6X5ZZfiHDns
4muInkJbnqjUlV+PuMHgUn2We3LFMQIB+1Uca7wSi3D1RBh3MDTexb8hkycx/wbfgPa1oFjegeeo
xfQcjwUPZrD6hkEVzEjFCJ4NjhQz7ZByKb49O0on+ClKE8XnrZheiNTrnj+j3pVcY0sGkW9+ghfT
zuwtVtS9cnymWkNmSbbKAEneTsMuZ2c6TJk3hFG70C4QNJvtdcxuNMVgmL4lQbxd7drqhq/6iN/h
N9P7apXlwMHckKyth3nGLjPyHaIeUKHN46DkwzIz5eC6vgg6GCxDG//bQ8aowDzaDkCDL15zHVJQ
3BVMjxS+krve2qrt6IOJheH4+0xQ7mfr45MNMs7vwsfiVa4Z7ehP/J+Y834QgLx89TY02Ipj3j5K
jK8uSrOcg+2NUscapsQgprSz1izYW5XKf1bW7IUg0kyo/VNBJEFji2yqx+SHZTjsV7wMNNk84ody
h4e4b4gyqjvKR2anQYq6usKdVOCTY1dENG6KqsSCJMJeQ37wYYubodx0kA5Jav+NyQc+JYHACtaT
7tFGyz4Yoc6FgqgWerxcWKIwNQjFCw0IR+q8yrUMkHv5VzlYTaOMnh2d9HaroABDHXXqnN/HjeqW
TE77yclHY0FiX9vkn2jARjzPLOjCDNiZUjpQeCOz4JEZWgHrytaTJt08Ai/g2Ynqfc+man3uaiMX
n7db1nYXB5d7XnEjOWINcqf/MWAWhki+XSZC9o0Qef8WIeg+45EI51xCZN0+bamgWv2JM+0OkHV8
VUTp0t/Eh6Uzp+evoR+bjcSSQigJvFxxRF6YfgCYdUyFYhnxm/0hwrSmv31ZThi1+ClrA+WfI3tN
5Bx9+ZTREePN4f0fv1vQvPeBTS9rJibTwnC9ZjeiDZlYUZTQGFj3pXPCDz8kNE6uxD+yMFUOQd6l
cUXLCB4iIy2yyDhdDO/n1fSS3qFnHzLbpiZF1R2tGV7OpjeD1N8aY8RLFQW/92RhJ3YV//MprukI
YC5d8B5qxXZG2yb6SwUX17aqiCjimas8i/w3KuHg9ixYaLVQNzTL4fAlQMPgaQcP1j4lWsicn6gh
YiX8V/CxNs1XABWMrO3ctO0sBePBW9KNpnN4EYEi5WQx4qbLl+ACv8RClu4FW3SrlrKMZMtLGuMa
ymyTzonP8+nJMImY5e0oWGacjyTk2/WMAIBUZYoRX/CL+STquCEYZfv9K+AuS04CPsLGcaqa9Qyi
lZjNHltp8U3eWM+X+ByiZWI/oleY31zmebW96wnu5lacnqBI4pvz5EVlZj1ypnFswrMBQFCXivby
I6NHJ2tUECdk0xGOs3Zxyx9cwfRX+tpoDfl+3Dca/LYIY5cu4PLE0oVg50nSLdrUbZvBd3NSGfF9
TM0Vn1y/ERqVGvP2dCag/VzOZ7LVvKX+oLjie2W0Zdk/h86wLC0zm9eJyp0OSUF1K3j3T9gwzVSL
Vt/qryLc4hsP1AW4YbzfIS+JAnukUjcS0+HM+UB/w8KgLGleHC34UmXb/23FEPTN69Wn3HISzTWE
YjpGOCMBcYgfX8FFQV83O1FiA4p+uqGXeMu+SieulzWKFZW3kIbvt33fjsyU3VEgMZ1T7fMOCXOR
6VUwSLhTFDNCJ2Tfhtb4a6nik5cypfdp9LFbl9zB1ILDuSNEKGCX7GIazT1W85G29+mFkp/cy9L4
p9tUOePHJyrSEWK799mc+MUnpsLI05fNO45oiosec+d0OPEs5IZv+zghO+5n79ZMRh8YEixM2zbS
sXGqF/hxQQrL0hbyAXduLmgfA+kSxlWVvgcj1eS2tgRFaDVHIs+kf4Dvf1oq8J6P+YxYagx3CxZM
IpuAY7oVZqbYHpGahCQKG4A9pfZXTKZ15I4cMxHU+1dI6PEieDXPW/erzRLvS8spyQs+yUIxkEbs
pABRshfrPJj3QPA1GGwgJrqvtF66fx2WJskDatM3SyBZuJl9jsNMJer+fYnSRQ9txBdYRrJ00t1m
6DJXD3ADLxwU2BhlhEiF2k3nTzG56JuH2LV20SEBXy/JuOv64gcqdndf6bOEJ7K5ASZceE18G6DM
Jk0AUs8YghhaAlUU1AYALF5UFQdPeJ6cSKyP6hPya9n5fk8KWxuzSU9NwISSnAq3PYWP07AFEhNz
BZ2Wto5Nio+/+l23RD5iZ4aF44zV4K89WqLVvw28UdFDVsminEGcZzKCaGnWpN77FmufoN8sKWfQ
ZemzANDEU7s4pvuVgAGlN5xGDp94X/wK9Js5fBYmV4Htmr+GtNQOkFa3sy5/KzWmVs439l/VAVNl
oKNgC7AajF5imMwWVJCqk0MF932ngScTVJ5axdgerLQGxZc7mTCqxPk6LGXunJGJV/V+pN2vl4BZ
mXembXdBD1u/36aeJt7jECX67JHFdIQ8rwI0K3Fb8S188zonmAo2t8XkeMzDJlJXtkBs0QVQ+6A1
s7GuOPiCOZdWu+6Pqzir9tg7bd9nFgliceFdpZnDgJzUfHQIgdoysoK1riaNsdXqI1MCJJWdory2
T0eWIy1ItdbpdEii8yeo9nokJiYaxF3s6kQvDwtPE4n3HaaQnGoq42O8LnEisGK5xLJTMzanfU9n
02uvcw9sPLXTrabUN3GEhPiB67UeaULx0JoBbmpB4ib67HYi+HDsaY+x3/w5J9Yj0BeEQWz1vGkW
0tLOKnPjCI9uXnHg2BKQZKfzo2fqkH6EQqmnFIfKNTVSS3bHSzMbvzux77KBKV3JSQMop09s2hX9
cLBCZvzHH+MsmOPKCqci9fI4qjVUpyAvNfe9Cm/U1lZyDh2BAJCq/bHKf5qI50kqau5Mvkt87mp8
h4Ej+vUB0jQ+pin8o+u5OfoQglooeyDyT2cvK2tHRJefw8/cFH2RC4k4q5FXhlPycmSigV4ty7hQ
0gEQxRTrHPpF+MhrQW7Zu3bXHuIb+CocVHSP3sredc6mX3OKpWQ1QeUiTU/rR1SeHm37vrx9k1MG
3rTHIgfFmBYM2PDeyEp6rZnuJNDw6Gc/7XpfrlwusvpNZRf5oMq33LZqAGhdwtp6rmxp1GrfDdx7
wjkLBIIWVv3XZGG6GU32snmRkmKbruJ/fWdUUt1EN40yYAbyO+g2neneho84fb/wvsV2KcXSd5hS
i064rEmtUrAZMkBl2zUucTyILyO+OPVvdCiPhcjlVNZSgBI3CDRfhlc695ytm7GXsvoBhSt0jQ6w
+1Ekrb7izW4R+air7E+lfFFy9PT1STqE08mh4FVNpyCcOrS7Jmmq90+TUEzPDxP2P+aduXNW0HiR
niOzEWj0wgWn8wuYwJV4D9fWQVVtvDn6fwkqyLw90YZPUvyuQHi04m8rpCg9SRz+uOygKl4X7gAB
XqacRDQce3YrREi2l6btnLTSXQa8bB1VyKj6kaovE9X4qSGjOfxW5IUD+Z5WReQfmGEn7vF8+R+F
D62AZUuR0WiLjt4QODnUUAh4MDwxCMS1iAC1gmo1nkETQNZ8L9mmHq8Wpl2UYQfy1lu4CYCUwYUd
wuNPtBXiZ6xKfrtXD4gGzOa7vaW3K4aV1WCY/QmlelgvboiuZSlmVY89dgMxlEbrh6ONdPa+7klo
gIbZv5rQJyGiLFJTovX+0MSwkWl9Dkwpc6CudT/1vuTRHVcmI41C1YSr+YdT2jvJ4o/hkG0DYv6T
lAkUEJYn14QAzYGBJ9OnDjei3N3Xa6R0zgKkLB42760TBx1n+sbr+7riX3eLM+8lwZlAEKv9l7B6
lC1e8I7OZBZdRZU60vYIap9s3GarKTJat16M3MsxluVXNrh3G+o16Gq57It79cOv0DdgAXq6cy8g
DDUyxORYPO1tw7NuHGWazXQcqqsUM1WOsQaFMF3LXlmpQ3triRrGQFt9moAILmZF6DdQ+r+pAzmq
lkLGVSYnGD3QWzre3v23p99lV0Xx2bPiaqk1DlHs7Olb0VzeFmboUyPdq9FezEUK2b7l1XGwiLPn
M1r3WvlLVLrUYh8l5uGRglLmfHIQvxVyWn2x3E+Gqi6r6YftRCg3BBpC01d+i1InLwxa9QBucOMx
kReU6xwFsCS+BQchsKKLrcqd7kFn65Ptyx8ozxXZle1ZawsJy/U+97fHG6WTFRAhuRVilATM7G08
eYmhOLMAG6Xzbe92JU1H8gwSa1umxOpJy65uaObt9OeTtokR3aZga9Bxf6cMC2DtZNe1wQL1qjvG
dQpCG7C3dGMTIlTZOPZXJLa+NekRjt60NIL9B9bqMYDnfNFsdw7/+dk2QcvSMuh+YSIohLeHCEOF
UzHZMJsQsup+WXVtmCMZI57LivUTOIAQkqFeqFO60Vsg2v99/TlPhtvVAIrCcatx1WsUd4+BFD0H
tSRefwXqZb22FCtMMZCrxLM9YFF7lQDqnbmlb54sqYpJoYkF4PEwiePvIbF4MW5qj+dSBDXch6vY
Ah/XlDTVSkIElrY8CbABm0oKqc37Xmei0doArbI27ZZmyH7RzyUOTc/2COc5/ErEZtkh5/n7n36U
JNyWczhsZGOvWwlSLltTC1TU80tgqJgtDwTKuDMxf02RpqzyWGCf6sWhd3NTIK5PVblWFJcPB7j1
AsbOmi8mMl7L0QqfOLxNoFhqxHrvoU58nHL+HmqVlecrtfyI22EPRqCN7EBfEFhaDPKFwYGH2XBb
H3dBjr4m5fSSoYkfVKFLm5M/BXKmGmTAEdhtARJT43ym+4VT+Di3u9M/NIGPUKSiZGsuKh0p64E7
1fY8gxjHHKOvFt+zyb9fIYbKm04DVNb//raFefVdbSYNFnCBcnXirThl/sXFJ1OywW8+/4c7T0o9
aQ1wq2OFEqg1hcrRDmT4x57F+/n9IpVZq8sFrU1O8pzrh18gnTepvlOhNGq8+cyYSBTGVN9m9bMZ
U6g0BWQ/lud/GpGavOpKvcB15R2NH4Lhj/igQLdP7/Tnyi8haP0VwRopDiDUb32HqPoQKDAHyhaC
t2IbfBSBkht0o7yFnMLjCpNKrmVgNMEEuqmMvD/IiEg8tYszmaNUOOqmrrnLryn60V/rpu5kEbvo
gIu8LDFJ8KERYWdfbOvSnqxLRg3Kq1LmAxSKHja+JO2b8P5vP3YQMjQxczXjPD8HRoCVwy0hqQK/
zATgzs+JnS5djwH0Q5BHxUcFlcNSa5iuINaeWVBAUHsRzWwK/nWHGQm8nA40jmIYiMeS5wwNfkVb
NjVp6HKVZzwWisS6rXBvvFzSY0DDY2pYaZnCn8o7dbwzZSyoEB5ZBL4q4NyrcX4N6AWz6RQ6ttwa
vmRIKi1FUzje8TzVFVIrfyGkx9TeY3BkHMBXrcawESGbaKZhyqh1YoxFW+By2f/heht355hkVvzT
sTE+yJa2DBxwXliRO6t7s2GFf8upCTzvUKtGYjSFilK7XtKMdf02S/ui6kfJyWSiqD3jd6To6tyJ
T1z5dQOGtQluYA8RkcyNxVQ4sufM0b9cQkTm4i5czK/mw165k2iBcewJMii0vUto0wrUcg9x2T+V
70cQprHvNATy7HRYp34cpUOwQ/szMxACIxg+zwkSjWkPyqIO7+XMAVeRbLiGzAUVmorR/Cry/FWx
r5HmDUDpImqk3MCdph90rqTVzMrGaBFoEh6VRRm4zi+PbbAI9OgC9xAL1pdJedzBgQoDIBcdFHhq
TiHatHlhueUV/F/8np5HN1XyTNfSV/sitbZX1qfJJHbL8hNXaUHl43p2/bwM+Lf4Gxf9Umtcq+ri
gVb427OXPAax30nsy8ZXX6oIdbBx/EemNFe65REejOMJkUBJ35upqbW4QRaR3EyNResNgsBeIDdm
OOfXAUBPjBxqDbxIFpROKXLg/LwzfUJYQu2HmCnVBxj6xG21XXcagXSUj0eNbYR2i82F3tYNqs+I
VJ2gXxXFwbELSAI6MDXzF8m5jvfEHM64CHvHNr8EgJWMMFajYu9uC875DYDKhLJDZzAn/y2Y0hUC
q1eQM9RVEu4uF9WLGmf84r6INeTkYOP7ao1WQ1GiUfpyBlIo3CmKu2UbqnbH3SLcaJ7sIqiBQz62
o0sOag+egwEf7j6/FXIUVcfwsuXDR/1ZyV4qEoxaeUu0TjO7IjzBJzIO2ntjoC7yhohFGlYuZTaA
d6Jx+9adPN3KKYMGdS9Jn9B0PZUZm92crJcwuSAwUntxaVgHXJP8WWwsaor5QUK+d529ISiYANiH
9cDeSoqwDpVLwUHq+PNTzJn0sy4MXSS/+EsDUJNCkUu7jYjTSRkA33YmQD+A6iAeZIhUEc72PZfV
CAR0hugjg3KiKAS/NsPPdIAxOEVnzJSyB8AKU3KmkH3/Tg8JG9uBTfNlPyQyUSvu2YwYSDJq6LBt
mOfl0sXiPWieWky0ozN/w4un9+WYgoTKYjpp+6xfUv+RIG8PauE8kuZTff1J9ooZHp/D/UIs3ikC
s4XSLZm5j5wdOkDUZ6sIL3nj3SSfnUOvmldqCoD018qoTBN8ZBahw86yUUhnvj+SG0GxZOhL7Pn3
2pP9mswx9yd5FduChhNfW/N81ylwLHpnl+GTACbptlBoC4pfUGDQH3tIBBOXIFZRq8ewmKWEk6qs
B1w8m/E46FulUOuX+SGyM17xGFYr5+5aLQ68e7nwTsOd7QqdhRUK3m4BrnMmwRU6nAR074OxLEFf
ppQluX70lM91dLy7yBa06DGLRkuMrZroNVnTc/n1zippfDTWwI57Cq9pp81CYYlx4G6T8yhz5zfV
ufhCVM7CciJ7UdMiSARl/oY6DzMvxrgAopyAIXJ7O5motRvtlrSSSirQLQ7HfHjdmOoT6vlqfIe3
nICsa9TnybOSLVFJFjriaiOT+Lr2U2RsaQANnGmvEFF49RiuVjDw9y7/Aa12z+AlOJvMilGxxslJ
NoXxoPc33lG4ELBGxnZcVWkk9Zj3qCUWTwUEqIgMvDMnEqsAkiQeqORxzX95IstCyfBYdR2TuxtU
BXlHBqF/cIwNeWrJQQsvPSqj4LM46H4DQPyUmNpNrQ/OVqroyPywG6vWUbDIKS/im2PFWLzLsxlp
+cuvSBIhhf2F9KX+cqb2As06h82boj9RAfWav27pBuqu1fDbAEMc0oj3Fl8fCsxGHQE3S20fI2Cs
PpKS5MiX3zCS3Jgc1YJR7ekbg1yOTPgCBEjqW+rT3VdpZAwPr5AMHRgdt21ZolL4hY1a1GfI1GvB
I662DF84TW4WrD5PF9o3TFTim+y0DiMxU07Xwy8pAlYijiaJJb1+cBkzwYt42d9N/F6VxPLo2JK1
pWPwhmniQlIcssw6M96FhwCVglhTnJkrYWRJXoyYuXytbk/PTlbgYaDZe6AWJg/dxSGf7GCfRQ5C
2njDTaW8jhXFNdPCVQd+9lRVaE1xtmESRQ7gsUg7ddqm43bYmUulrWS0Rv+OF0PtxTncjipKRaM1
ZyWD+tv3SFPWQxXDGhBcYKh2576/W4KDyrvP0pwG/1CkQmez43HqLoIKqYB+KLryuDtegbag/V9O
NxLfkJjDo0ayDQVbOhrBc5adWqpbwi49j+sQsnGmjVFMHs8qDnwqc/NQ4+2zF4T3FX2af1Eu/3/C
udFtQiciibhDhfCa4fXbf3/+SpHEFEFJGeshlf28F6AdWx79vPWgjihFXbHgjgBSe+4ApgMpLgWG
con62rbEIAEoBPmzEJG89WbTvzCNd/hKYL3c/nyXGe52QE068XecBzf8J0q3rrcmJpVAASXea9c7
di5uCuXZ+FkzmIYFvqBaJAvKr1SMldzFLFC7/02Ig22G7N5elk3unai7NDrSSv/qw4r7mmXIpklo
Qz3WzJR8oy4fWlt38BszDTvQ7991g+mt6Gdk2E8O/K4UgpFAzG+vEL2ZZ30n2IYxVU8tMdsbxraN
GN5d3i2bMGncxhMBtEzy74Jy+SYaJnXlfsipH+g5rmFeza+ZhG7BFkLk0Uq8WOh5qTHhhJvdFoFc
RZBau/b22dloeZkFhXKijAjVVdlWia/dU5neEFrOPzoZMZINd6mCWloSf2ZJoFmMPRNO5oKamkbs
heSqH3yTY1TilMrJccwjKrvdxXUWyrOu8VdbVXccintgsGIX3cKhurKh54YtLp0XetvG+D7pLpN+
7dJl5gMr0gD6UXZ7k2wRYGUGtUFIVtAFTdBLntQg92nIMG1kTRzj5i/TqDlCym/Bk62QhkwR9tUj
OPyHPNxgAyBnYKLnsTDl71JFBhryPIF/BtqLMkZW40Wj0/XSUMQANLMM1waLgiK3VFG/jyBPgyM1
HsuSuDm+K2kXLgxK9Saar+R45kt0b8ezMnOMOnO2gDJFNBo/0rwJKspyIdMlTG1pqrZ0VlLP9qHo
YkrNoHZt7E9HWnSJ+M/a8T5EEn7lZQkYGBFuX0hsXBbXAFAIoeD4oqn303K2dW69zJ2HcEGszRxT
GeG251nuk+wxXzvBoDOp4Oi/VnM9vKbZY03zwdFkkoTOgFVyZfnxaVTYzv+ye17l6rwbOlYrl0f/
pQCV5ysp6y7ltDRs84mYq3w6IkcM6UPocr3dQCDh/s+I6PU8J0er8V0DBuezW5tP9/CNE6qzJjN/
PHrYbVJJ7MLFrqUmZq6E6wyVSTF+enIkPIkJgFohJHs1hvypkzfMttVrePVlZQfZPlFzV83K4RT4
CqGslDMd/XdC/d6sQymEPzUkoAiEJs1hPhGkXtqubp8pz5EYOleY5ZnAuqi8gBQ8IqKivBtPZ+dW
b7Ycd8eqpv/QfQY3uu+Kc58K1bBOxcybiAGD9FRqvQHopuWdke200qBXKzg+ZDtnLfbJbjNJvEsG
o0d/5I8DDx9rnNths0keJtU/aqteZBQLgCDNNxi5SGTrbHEYf3K3kKqkwwgtzwbCZnVZ2Gon4Iev
z2K69a6nykN/26OdbUiYSVidn79NDIcj3+M65nLtaKQFAfrXOkqDfdgnwnnCBagaBhEJKhmme3Oy
FVYwfUaO9k+/mkLGa13dxkUMIRAKx6QHnVJYaQ+6KEXn9Hy2qtsu0NkCk48Qk34CscAphf9Dr9Xy
w6s5D5qS8G2MF1Bq3CjPGB1zaW0Dome/ybTC/45m0dLXsNEJ/Z42yjh/a8Rg05qytvBJjCIWawLw
fCaP3+mHpITevuV8xZcS93zaPIft06U7cIZGKDBnABYT8aBscnpha6eXkoJ3iovpr3GjBrczBaei
8v/vCCs1LY8gg0C4d9mxPRI/Ge/lsPDM3u/1wpOlWGnTGtu/Ze3ukVK/11/Jjm/PQ7WbH6h3EVQK
A0GGMifxFy4j5TeA/mxh8fV9GLQu7V8awS8oAk0GARf7x59MFJCPbBft7sOQrk79xURn6XgDTpgP
x/oShgXXGcpPyIMkwp7yL6otj+3AF53PuzqZwCaJFXTvp167zYb7NIUi2GpUBnEojqXmbS7k4Lq4
oI+h4C6UQsC+QKlWvNRV9TNTv1UtFM+mRMxGjuSU3Nf8oeLs00bCAJ8cJ9KFh3YfoN7a9gmRPOXQ
EyqRRe6LAWjAxQzo+opJHuyTR8EDDFNm2I2KtlTjvVRNGGwIO1ThIsGHQHPCuc7UvPHGGYC+jfeO
XWJMRGF2pQ14dTNEXz1DV7CIG4Xf/DoijXOGxHU2MMSY9YgGzJCNbggBffMxyAoaZaWcVCfWRMQd
l+tJtny3C4LfynjDyDEfwlgvoNf0HmjQzETzhpaFAkLbw+Vh/jOWMKDyckI5h+HPbKkzyU9/slQm
QiqgjenbKG21rz1AgOxZ2To4oWDw0UXXmwlhn41aNbZc2zCDnbUZixSCZMfoSBhI14g5Jc7RLwnc
9p/FND+xflN3c+reCREIL0FI6cxOz1RxBSA8rOV8tOiyq7pfDK7vYdgv4IkxO1N9X8yj10Q/DUcT
9lnoL8BvCmA1MWS+qWibnX9NGvHxAz1LkfMbvr0472GFmqkKeAQSi2L8FbRQU3r140IX3xGAQtB/
VthbLzjhLtjnScbci1/g6yGxI01Mf7+ZYs7BUi/MHUOymzSNsfHSmL6TumVmeLjayFdAssJr//UO
x8/OYITDmXiRyZ2+nPBZv8/M0q4k+3CahZFoYGK8nu/y6dgoFH7j6G/l2gBWz2h0RpjNEzARxFaM
aTutu/Dgd0xxKeOHD3kkkL2WMK5spvhkcYZ2Tp+ZVX51ytZvarqsHjbrPqAtHOcPmRieTqFxEo/a
sga/e5V3I7JbXGfVHy5HbMpcSmJXVnQq3Wv97SWk1UES56CdZp5w4G3AsB9HBpLH5hMrFFXiO8vA
BrqSgiZmTh1QeBPcw/L5VEJoi2mXN9SLLfLmJrcD1vwYKRgTFh9JDtRsiZNtk8e3mCefZmVCcs8w
wHzsfckHESOBjHxmnU9LZ6jaPdrHHvH4EJlmJlL5XHivnM1Gh3HsIrNV1OO+KhKU0IUq4Df7h01k
15Pzr3kw2Ed5HqjtgX8nOINDQvDdMOPQmyv3Pd9//FEhKo56ZsDujSzNSVh3bSpueg7EV9ETVLqf
iR5AspgeflC+FQyV4a6q54VRdegx7G4oVECbylP1sDEy8C3eQtxCcWe2i2Y3MYnicY2AyPeTY625
q53WCve5KbixgGq2G9uqTV3f0kYw7/wJ+KrPQwwAcbHsSIcATPmRPeNFZJVn4xB0MZSUGbOnxKtR
PJzZQvNjj/fA1/ph6unroVqzJ07/Iv/CiWY2zZjJIawRaA0GJquIPsXvWHoB/862o78+nujCjy23
BC/7kuaeki9GPjz9d3/Pr/eSeTTziEZE91E8CgXnS1fm6I6v0mL4Vb12YklZp92TzGjvILxaYSA/
7/UH4phdZbsExFbI8M1C92X3+BaACO+EOLopHxQvPtGo6ub9jL+GDURo++IVq+bP/rm9OzIt9Fc2
XbJiscB7Qyzz/SePO/tlDrYQCFDZC6XUl82aC+raXTh/8JbNMs+V098zi5EPGhsKw4Z2UOF20mHP
/2H5NUo5c54+DBAmiBkKgvdl1MpntHO2S5QUwFvKqd0IlojB7g13BqdphTbdSzS21i9cBl91cDoa
UaaKJLnHA/CFOZ9iiPXywfREdtaCrsvwHAAnFCYetYFOqHSK67ZNiRePQZXynZXUkO2pznHg3iot
0jqgI00AIUTAp3fW7D4j+NRmhccvfofrbk0EsSlir/2N5DgjJOuJPSY5eHldGQ5HR942z3LfUjfB
B36BeNQYUh7GAJ0pRJ/uww7ZJAtnos/wLIJJfKETZ7HGq1W241RMMz6hz62uGkkk7R0lEN2h3nG0
bceBJJdUGobtzJjXbVPPAdc8oIA+64Yg5qhncFBG/pqmyFuFvDr1ePCL/KL/aXc8VS64GuYUS0eX
qFyxox4BFF0h8qk2dfa+Yyypv+X3N2YK6OsgF2du9dsDEarGDv+j1OYDaBNjlWtR5temMtZehVjS
kQYfTRUmbHK91EvUg7qhppvc+IXyXclYdzjlE9Odf/icEq5aVYu43xFnlpNh9OLpk6Tko9vHj0ht
N5oB/AnQKfxBBb+yypgCWohTdgf4DlmghGGSc7AtL9dJipiPjDWrXubtqaFsbqM4HgphgO5gfa2z
2ci05z0/MnlqrKHVYY6uoAS+qiUx8m4/5gJ2aRu8BzgkH3tMO+CAgwRuAttlJ613FCw159gHCVIF
gC8TPCDVopO80aPhjgoefrbTdHdRI+6SwOx1sGV5hxnkO68SPjre/WVGhRobzVAjBd8rURN/V0MT
AnXgjrlIG9gX0qBoO8cykp5IH0KJPbe8kyICRRTQeywIPmVEiMxReqn8dG2r4Wlb39Qm4PIWZ7ZK
P/H850tq34KhIfJLolhdNQN6+xZhJQ4iAQQABrNiaX/q0y/mjZT9gweLmtPpxyEVD5s3lTUxuUfs
FlR4zZqj9DZrWnFQJ4hr8yvfPUS76gH9MagPs0wST3IW3lkEptd0Z8YkMP7FvSySuJwah5EX9ej9
CccdvTHCo0bCjtsn7FtvPFO47TxHvJyagTC0SWPdUfIUq/Dnrp+356o1/IQNW/T7yp87GUHCQDfy
kMqeTBpbYJTFFRohh07A3uDTKE15Je7TFD25ME/gyOJDnyAic+X+EKYKE1ayU9JH76D7S0oXIRSQ
ibIKJQjsOXV+3X2nOh4Rm6Be6LdY6vz6bUu4/SOBhqVSjfa1raxdtXAZHXroFSpXz5Ma3yeejNu4
xXzBG/7zQ5xfeOWeiWnzaOT+NzGYTrqeNNDrXF66V5V4HfQYiY5NY5kqTvO+fAscidFk5sNwq3s5
4eS/CdsmzXIE77Xd1yG+etBWupQCGvRSqdCDlz1m4P3/w9CPwARJGfgbM6U991os1NZlwSlgdspk
DjmKVsGXwUfF5+eFgpG81Ed6GsDt2nZYiisXA3YqFgSoANRTKQ9BV8RwygXfC8jsoLDRBYFRYV+C
gFXx4qCu0kSWGzZW8r7ffU+PT9RXVa421Ldo25Cwu0bBfTV6L9p4IS2B733/srLsNBYM9BGOk8jt
avo6yMQ9eVhIE0KjceytjUYTvzqmHYrhzc3bfUVUT1c6RbWsvGypYGYUGh9Hx7DA5GQbeqHcMKtT
+TbomMjyuuyL1xpE87R5jcfZ5QypNe6YTttuNPJTMBIDwV3wmDFVjIdNQYVtUQupN2+KVKhihTfC
7RuUa1iN13+yydjqRMaTPQl/aePvoYS5nSHJzi1c2xYXmD8I0mO7jgeWf5WOWAjF3KKIWMOMbXuJ
ClfSNEQaXlWer7BgGLpDlkgVGNCzUuS5nKvn7/loiTfrZH9YnNc6nCyTui4RUJz2aHkEon4z13Wj
eawFCfnD+jaV2wCEZ916TBArJNhN6mEJRSB2zt5faUCE9KIFAwAXaSSC7/3nRiC9QLl1fmG4HfgK
aCuiQ1b/eGIUEikwCZX9NU2bDp5KIjYMP1XVAuipjl/FfBStcwm6kP1kHzL9i0ihAW0fW8tGrL7N
9gNj2xOWIEvfSi6m44U9OwOhr90bGPXQx/9KuFdcOgbMgpkXl1eO1SPkcNQFdheaj0yoNB8fNnbu
24wh5dzOhJ1LXs4ZWm0uQGFp5yP5VprT0orgOQLlZAx6ViyHqFpBhJN+UDvW16P9U7nW0YZZLN2u
kMFy+6XTQ52QlNe8+JR6nkXy1ymOTUZOVH42Px8AfZdn+zBTw6fttTX8EYypMJRgdd+ZFk5TJyq9
MGx/gVUvE4lY8+QVbT881nz/961gwS7IOveRNTdU61yIPo5vRQqWaKiwr0PuJWmZJio9kk46SnmW
jY3LGPm4Wa7FssIveZD0qU1Vupl5J6gmNS4TXgP+oIoEGbq9s3KnQp/dxOIwY/4DTdU0tL+kgtl5
IebetGMxqu0SvLeq36MJzbe69MEova1xI0PHXG9vp3/8tA5lzKKDxaucPoJz0RMguEdK/kAUYxBT
pes9BeTDOJjFVu7u+F4RPPTrkD3xaOSKg0A7vrAXS/WYNnshB/eVNmkLROHsWHFFOZyuKtcAQd+o
1emvkFMfiCvaM40hIUFH7RMvhlcfN4HFlTUa1CDGp/ySJM2kAQdQMcnxGAeG5psEfBtMKXeXWnRg
aJgk8jlOzK6wAbccyeoC2o7mekO/Zew4/yNGwzydYirNc21STcbt1Sl/csJiJR4Jv96ek/I/Zgu9
/F7noW1TGIasawtCz44F9Y/adCZACtg6Bkp/ZD2FKML65IrvZo7TafUvnQooMvFG82nkpFh8lP35
ehrs8ZvlQULL3Zb/gC1SGnIce31R+h/3U0N0QiGsQTozI44xY7lCzjNdOjoQY1vr56dPHyQ1SRKb
2iMJJn20emrtmU0/hDV+mGLS8gXSbkVc+NJLD3KWXK6eEK6Avn8rbrPlJquHQKIocYo9ezNf0KUG
KtAFVMIVBlVwbRrRQCqdO7bBYS9fQD8+Hi+5JWW1Zrsi6qedBO6gdmhJTJU85Otwjvs996YmNDAm
I3A+FRhAVyje5m5JR6eQ6GPOxV3emE9jacssLAUgCknEBkD7gwaJKCBk8tQ6Qh+nys98NUKZE6f7
XvnVnnAL4T5ltVDf2yK7/2NRXqKbdT0F24Zh+hSX6UGAs4ZwmIeHhr8J5+fFlNv79dQvU+2Ulid1
gB/2YUwDGLWy631MpaNJ8tu5uO4nfc7lcVsj+0ibGpIxTlGIheJXn+LQBofuzYaYL/oVznttW4sX
H6pF40orHUNsPVV3TlR56bEk+22GksR+0Tvv7kWv9Y3c/5TiLTulgQzx/x2/N7jbLyWkj34Pq4dj
Xu0Jv0bNEdYP2XqBFW1SqRsnwKwtbLj+Lq+6VZvSNAVNS83DJBofdBUiiI+36nRwaXsvaBF28fQ2
+nwIpnpGZiY0/8k2rRgAWiVp7tLAvjuUGtGaadmVd227BFthFlwPNVsdzZxNhDOfTwoQFrdaL39a
LaES+yU6XsG0s5NQRN9UJNzChq224NCYPPeatGmWVsg2ucC6NSs3o3H/dq4J4RwBXAY7CRHeATKg
qloe9gTd1Zxl1Q9QG2LwVkQAMeGrd6byoZF9Uu3HsnUxkDmWACrwUDy3eK5uxx1hWHqbY/U7y1in
PXWfzi1VxcHYdgkxlAqZ+qSuDNxX4VmGivWxdeU6AasyR7TGzGVKoi+DYsOaLNjOnXmIWPa6CsK5
HLdH9D4a0dJakQK8/r2eO617sIENaMyrfDoiEjKUtxvt5X1ZXieNu6WKzQZBJqP69Om+Q0sLo0QS
fHGaARxOezMa2eCWddDu8KsVQ8emzlH7iCdYKtmI/r29wyz3U0K1zw0iWtrYRjq0HDXM3jzDUIgz
Q8QoQjO0wDD8UbMpJrHOO8G4gE9h2I7NBZ3XQk24Tr+y6pMu7pDY6O0PQi5b8/RdVFr0fhZYcRFh
t+834ex38qBLt4kwnj8xlDUuQ2cZbB2NQ21uqSd975EvAYG8FOzjmp8Xj6XAkVKYAwCMLyhlT+lc
43Psu90moj678zkUsiL3ZAUe2P17nds7rH9jmZjWoFB7aIglCzRMO5E1Dzhf9zAzMgk6LCwTjUKM
SfWGT2LAtPFuMNlERdQWcJsJWS2r78ch1sDz5C3FGVqDoQHXi/wmRKLIzVz7Vg7V9JviTagHq+qa
n8lenO0kKAOZI6zGUa17Dj9xoHhe5kyYhtfN5PmKgca/1F17xrmd/xsdTen/N7nOMlqHDTn0jC7/
8js/UPt+Hx+XyCs+m8uw4lU7CdEh8iUrrjt6926fNH3n8G+Gq6hMTngcbEhS751n1t/X5B2Co4W3
xQCTmcmifnb/8oqxqEGxU2DGMywwxa2BRMmgTHZyI0pxubXdgysnna1zZiX+6/Ks+4z4+93b36XN
c8HA4/kBzsQR11wdnnpiA1k4F9yrJvbzVvNpYyMQ93632WYdbcLLyoDlihmmfzLXTMnyGDqXvSHT
U1hOfjwxNMTWA2T7YtnzVKCoGjsa+CKsFJ0cur/4Ceokb4ofbqJ+GKQmBy7RXmn90i1G0OH58ech
i4Wtr3UXN+k7B6zQvhk6wP5tArXn+mMKkoTXyssWzjeYQXcS32YnEBeEN7xyGKWHKUGrI1s/s/xl
dtXPl3MfMZvunej/FuKvsf7ryqjlwxLfI0YKd0uFXML7myy4UBaZT+3PN44lrVto4OIVmlSh/Old
DpFAdsgnAcbpaXNZH8SHSrxPOcOuK1GI9jfOr/YRriOBaeAw/KwPWix78p3Ir9sS8IqI71yEKPU6
Saed77CBFG0N6/0IvSIvpQezpummd1lCsaauszBmC8e+IimQFSSUfky4CcNwCwiqfYuKIBp46hYn
+dTYGZ5kmBtLv0UV6jY2Ynp6uW69NMKiesxOWxsWX/1sBae7bUnCJyKDLCVHbRZu09RvHfU4wEyF
ExGj59zClQDsXvYw9fwS5nDKE2XYXi8sPQ5wop4dweSfrvpjxDTLOgAP6RJOanTBf4DuWTiloFVH
bR+rpfYbwvz8Jhl3OUUV6lkBCVT2qpm4lPJnFKmb3TItRUJbEVqQnoyovQ/2JAGEvx0HWahi6mn7
LtUi7cX2TLNPhgpUl6Zgrh1LioNN5qpmZgaVJfBImlmdZPZDOTORXCb9ReKuMYxVs+dXi+3xL1QX
SGpe/hymKTsXBJ8UqZc4Chy0DwNH2jVeY/KbYdNh3y3l2YVbr6zDQnKBvTEcIiqYlldTkrSigXh8
RWpMdntkBFm61PChO4AEN9urp6nVgsHrzMWoE9BIb08OrYGQDZ7pImtnbJhV/3wIdhaw4K1tqQl2
CwSSvWZh/gWB3BG1doZyKelh2ZdZQm/5D4PhzUhLEU5BVwpfe8e0CL5lzzcMrZSji1iTcax6QBL8
i9Wd+SnhCeHIG+D1Tk7cSldEHPMeSUo63F5XhgLXInJSraYpb54rXzDNRiYJaVUNdx8oGcmfg2wi
krpRv0evVysiQK4gkRFxDfUglNGd9JGwyIyub9kaN39sPfvGgs6/fTk/xtiMVQ8xYQRICbWSrlzm
zH1y9Jd5olyb7fExrf0p8VnrG8ocKx9q6mLlv1RwCq6th+xIjbJN2882keXu6k+pAL3GUc6qH8BK
Wq4nKHvQyuVuzSdimWXGLgGs9oeHxyi3ig27jPP5QPyBncQOwjnzcHw4jPenSphwx8DOBcH8YUGc
k3IY9CiuOXir9i1XouSo79sesko9Iscqo9F8huQKZ/b/uJ2YFFDEYYUmIH16q2x/+lIULTINIvyt
RNUyGrNprtPzHrizZ4aZNvsAqQ6cGyNIxJBF8rGXbI27DiT2ioGtBCXAeA3RUATRI/eo8VEqXSGR
vSZ0ZcNkdO2xQeVFvqfmy1JrCogw+S9H25eUeloEVsL5FArMPCj8NkFynM11D9ZmWUceVrCb2o/1
L3y0i0/oaeWCOtFjFzGSeOSp7RuxBy1I2X+Ah7p0LJ2P+3aBOWlJMbMbhFEIl9/CyPfYWEVMYaXi
GfjW0wG2/h9+ZdUvoadyXPnm3Vic8NOE/ncV1ytkEj6HGpWj5JZSkxK2a2iRKlQbI4MkstGJGVOa
KjnNAyMke/A0GC8Nh+B9pdgd8Bk0IV/OgZP75rJa+fAoy1bF4euDbqlSs4bMjyxWuN62JKWZT3SB
x2kJGJJC9q18zfZM10O30zs8eSVy5mVEAl2xYX7Tu42yXIr/hq9GPimuXq8bc4fWz3UdI9zzz3D+
qBvZV6yeb0K2qCg9ebAb1x6bNKIXCMpK1wbUMXa64nJKTbdt0aDqDjRe3W6sQAukf1qXo7iEYzkx
WgVErqMz6T+aWx/gOxSRrMlaG3vdYJb5LMK3EZ2Znw7rwhMK6SdWkcU1T5G7o2sgxpU7r0yzfJMU
JEndYkL09Fq1RvH1SkkpSZcniU2/PiMx+z/S8Rmym1LV2wDg9i85EZ6C7L/SI9d8PUSrhgSvo209
1IJkDjNOnqPw7hTxrZA2e+XVVweRnN0abM6elmG+02JaZlbVc6kluSPKgcOzUU2LCc+gbCjDN+Wu
v1Ylc3cRPCfMvYmU/1WUeZ0jvSjDvyaAvsdj+4WpOenYfpjfBf+JU8FlKrvTqSJoeRO81RAAuEQI
RL7tDN6PpydfSfniIaF3lcAmNKRnF6WsLpRlcQlE+S8etOfaNsWo7BuwnRKRvBskegHtvgMoUQTr
OTl+i7CwyiaPlJ6knEd1nT/AKxU2ee5hqHTzyjrzV7bjy9gWNAYoapb6B5a6wNrVLL1SfABNIMuS
XtZ0VQKEeoAcIF/N8fFith9Yp7T1v7x/9w70UWSbnqF0GbI4aV73HzhOEI0mdNzH5UOTFZfTvdST
+GRkVJoiCY1HNbJ0ltvDEThMa3jP51mUOznI8cxAC8OlBGvUX+sS7aEDcp5NQr5W5hCK0eifzz7S
r5gYLq5pHcKq50O460gwHjMrOpCq7MymZz7Ql7aeJ0uQdX10i5JhEREz3svffsjgCLQpaxGblIXP
7iFPwgv7fPJIhFNM2t41iflm2gu9Hzo1d38PR0sZAOGmRYrrFsS5jmgTu4X939grhXoaZjWhbFOo
pcEOIrfOSJDnWMDda3pVtfWp6XX/Jm/9XO0oPw5lAgkkUKSy1roHG6UeHWfeow+wWzIY7TSFWZKM
E/0r6UOYnkBU3wEWJUjquIt7kI+EfCnUC8B6hdmSziqawUdsR/J0oXYtgJg4ifNxQ/vRDXKvb1GT
NAuX3ff4U7z2KbfYUXf+01G7XvfbCF7byi4LxfF+UuE6J1evAO1c5HPqDbtikm82gUqqf7JPPIzj
R3jFxSTBIiSh34lXKE/qqmGCa9/6f63pcccOdwiEhNTVp5Jphrgw7iOY03WgAYPoCOJtlFw6H0HR
ppWgqIhx/kY6lQ0Xf2u+SryTZbP0/gDb/BD0+4/vK9Civ9UUV7QkO3IKdCR1llXbUvw6u9rlCIKZ
7jxtGxhZes92JvyfmTHXDcCcmu06rSrkGS+EfLL/aOXFLqLdJ4oqbP1IITXziEVN0UOUpIXxhUJJ
SH0Fz2PcA5C78KZNwUPQpN5/7v6v3ALSP/ppIRTpdrAWANrQogVECoF9uIcF3AclZR5bvinH20/X
zGJ0oi+NwGOVpKELQ2teubZEDk4aoXwn4FlHmlV4In4N06BsywaTfTZrDU4Ow/9DBHnnrC15Rrmd
uicSxt42IJkZpzh/Sshiri6SCmY7MOE+Po3ec4kxJ+ihCcbwemTUcq+1f42z7LylWWUwh3aQh0dV
wExhrNTPNO0ieQkfaAD25pouGBM9j4gtan/IIL+mUODw8fnJMxVcNmLbF0ZD4NxRC+HPBgNVuZS3
4yvyblbFUAakGj/Df3Au69NmmaOlL6wqk9Iod7ZrAF4gJuOxKLBtPxo1iKZFCbt0WVmZ5kGNlf8a
hgqrscgbUWtUX9Va6bj4Yt8aPUyQHgbkMwyH6TfN9xdGWyvOYeic/2F3IdezkOfJIFfoBF3a7rdl
e/yBFMTNNotaOAWoQQxKB8xB7GYlMknzxr+AOLgbMTwmqTgDbWrvejpNgMVxwExbTyASIfMLetNT
u/oPPhgZXqpOTOcWMx4UfuNRxNlBEbCdF0+pOh7W4kL9P4eAKnyKgX49xJpGlkjwY8aEoG3zU5Um
j/MCBSXDh+riWELD3BzRE4v5zK8PeXimEIzAIn4wjB0EfUDQEiXQm2QrURCevHGdF324CX6yQwgb
BH1bUggAh/54qbncWKOiD2zqJyBv5OHD8q0I1SwYAuGaltjKj8UrDZrZIy2GBmqOTjRiettkLFHr
Cpa9BKJLShYMhu8UH+ByPshd7kZUI93XucasOq1u29OkF0cTiSI7enmiz2VBRKliXrR4YF+QKn4f
nDF66tmgsGmOUE1MSYJuvNDZKGkfZ01dtA5Qh8Bd77fu0qCLCLOEmNrDpaqhxAQDGGIaRU2QP01D
YRBOsUU3HJ58GvqkDd2eMuAqY+G0RuxKFCUmVFK7k2qL+4GHPVJBO3GX/jyginSLV3E980FVc4NQ
RuJCJy7lYjELrQxCcUKeegoE66VGZsmyqP0gaqaS3jpa5PshdZebwnVGksLiYTWdFg6QvMI9mxfH
jNyUcFKZ/VvQo93mDVzcpcloQ8Tbzm/Ef4eZS5TK7L83xiY5vxH5tL9c4nCNofYLUmUvQQFmyVW3
CcfB2ZVbT7hEOqrpgugLcwaChqplf2mzly1tKlwBnN4ylbOczQreKcTpmrS6EKmOCOXhDJw9fBjJ
wB3kPVkqtvODDNm1CBz4tMgnkebY0E/th6F6Bgo5wmiclF2bZ3ZUm7w2o1nsOY9QD6m8LuCZQnZm
MB/fljUFfg/93I4oUWa7RDHXLDlB4waqcrGmUwfYWIMxP7la/yW8H5QYf6hbckDQ1N+pFxWcMIJS
ITtqujK0iCw5yIYhgnlcSqM6uZjO8cbjqaYj7cxlg7Sz6CxSwFVRpYfIa/CwqCJqx2S1jn5jTKkO
hADImJirdZDQrqJolnRvdb78gKsOCdFcK3Z2r78N/6Bv3IP+iwW2V69zzW6sCKvFjZplE4YcTS2D
HATBV0gzl0jGDs+774LDMbzEllW4GkzUJkSo61gcVxccLQcl4qlncdTRdvPu3WAvhtq75PJr0tlf
WcnnqcuXSF1JYwuaS2RDpfm4JomGDF4EXmD60kaGVHPwE/bkXACMWoHTzBiRMCghE2ARXARXR0SQ
nh3dZ5TmAVLm10KSYPu+jQU5g/eHwBphkkgGCHYwNMHwrs06jSwox3OaVlMSt3kk+4huhVELZpMt
JIh+rtAvqkSdpO+UGbqwhMmV9w7Y5n7wK3+/dH9ZXb2NGEP13WXgxFMf1iJjcylrX+bFPWftrLDh
FrcIw3QsA9pkDq+qoYsWie8hOBa9mpFxU4NdhyZn2UDWWFEhNhxLVcj1ujpAxNVVa13IhoO5mKkG
pz3X81aaPpx7m08JB4uN+reaYaRLSUn13QeWKg2u1O123fquxqUKaZiy37Ff9m0oEuWlqZJBCdX2
h63okxRAO1AL50T7HKE+DsTC5Ai26dh7+FL2ZFvm+ma91zjNrnyYWZTioKrCbWzYrTr91HSkJ+4u
bkBRbRkpMmLbMHt5o93/BujLTL+VG9QYSGLGOrlMUF9oowjmKqS8HsfOjuPHKVbD4LoXLXk20adg
YvP7DlMobnB1jl6UMls8kGJ7Di9bSrxQfKCVab0cJeeZ7mn0T6RZVg1t7yd9fKcuefDgkbPAWZiG
66f88/EPsVMzO23SLLIVl0p/P3cKe8Sz7J7XW0bZzqf0HGyQdlmy7y1tR9w2MWJyDLunKrLaB0kE
bEJcLE7/stkPnpWQDoPOfD0ghbZqyQeEhkvmqRx4dhTJKtbJ+59rElVCZ6UhSaoyNjD10fDGqyly
4wOEHRvoBFB95M6ueWxHfgSF2kake/zDlvG/UfUgzmQYwPp+Bv0FhoKCA/RWzs19g6e6YrllcvIf
xFMbp0EQB2IB/gTnRVdkeg9ZLjXIwiWE8mO0KxD08W6n1gaHZuaVc9tOhNYtxeuAvMagOMg8agI+
pGIrEtUe5FGFr4SDGkgUl8ba/us0KW0zg8dp+oDh7808+HuVxL1xzCVoqzBt1JRPWFs0SA3xXGcb
DSmAP+T6JWvVESLloZG3CzIYzSM/fxTVZSkBbgrc/gkv8womsz/jh5aHc7jIrgQu207r9s1slDFQ
ormcACmXiBdcIGa57X6E1a7D7puSb6s/lUgmXL9KhhaD31nNgcaT7EAEDPREOtII9UbjZhGspOP/
5sayhT9RvCXOxW33A+ICbBWcgTNy8WZUGs/PzkdG4HCYpOqQP+MJUfQ3qL3lK4usGYhdQFwWrZtl
b9cQo/YGCUWskoAJTrBTWDBD8nq6x9jEM0iVeeaGo9v28ftrUK4Nq6aoglZNM5jEOP+L3nOa2aEg
EG6ew7UWuDadEZvvJwYHpe6IVI3sEHugFzB4fH30QwpOl6BncuHKLx1rXaAOU1mqB2eMH0vhLt19
pwTLQvrYtk8ilgbRjJQ4nFeB4y7S1Hdp3cWV0huT7BultdCVx7b8GXqv4qrZQ43uAoVGrP/ymyoT
eobQYtzoM+V/1MuH9oGX0iyLarpyy4aZvL2jVAlzj20yaxgF8dCm7pLjVnKhR0y7p50zLtan+dyg
eXMrVLdsI5DO9JAOl5p+2zTcEm/BCh5yPDY0D+8/8Mwbq4Sh5LCVFPPKscuLdjcEmH/wquzN9Hgg
05/7ckw2CpgtUhKieHnPOCwa3ewglH7ESLGsa+UJEscXOYz33eK2QS20lCK5SFz9mAUYma54Eejl
PVxQ1oYsPQGYqxLUUwAsMA7vfcqzTnzIHDn4DX/33gqle8Bve93N2vmdA3JTPa3vCL761ZF4NAI9
wzOSTViVd/P/zmH233H5RnnsKOTQN4QDPGwZSfI7da974oGTfVbbidXTJHl/DKrw/H8NWFja5trB
WpcuXQEiVISNJmWsNPOymeSXoGR7Jtv06wzJLL019gnJ5uUZSfWmyh1UZIFQ9XWTFFo6Y1VMjkBe
YMU+1wfWD+o4qoCAaq6E7cWzWDGh/Ldwz5CUwz40nrseIuBF0d71c8ZPS+5gGuSWQzT/r/j8scwx
RYWNUt+72YeA0R7frxjgjrSxsfzbuwJuElxk337sgjOIvI8KjuHqSIoifwhFwdq4Rhd2uu2IITbt
ndy+aWL5WNHZzqW/MxG/1csI4LLG2nPi1mwShA/hApfkzhJ/JujufTukRp+T+rX2+L91NxuC8C7P
MIeEB2mjw8GrCVFG2oF4RAUs5vi9bW6iB3VTvnGylXMqTuzY6luX9EjR2Tl112d5w6ggYEfjQIFc
m0mUbEI3Thsi3xeQGo2RgTZmo/keDHv9DlfciSXSrvtPBk8w0RnzikAdP2DdsPNI1qDE0rfesybT
6f9d2b8V88G47lUC38mYkyum/9crv2C4HerdK9hrLj+GOrPqmgh756Z+hiGBQvz3fTfq9Y37zjoO
awj+qyc1r4bE8ttuOAgtIfBykMLCDqsRFC5DXi48mzYOsrE64jyDcO8PQghNaJQbx2vlzo9aSatN
7FCcfGI0S5ffzprZOBZ1uO558Elu3AM2sJzDQfkJLHzpEwOrGP8pkgofjyYJ3GNIQJ5MeuDdEjLG
+mWyWnAXZcTfX8xCjT5GyiqeAmy0NUgiRXIu9hL/QEOEmDMR++HPrAs9g/pUAYQjfwe0PC5gW3mf
GRJqt1xl5KcwZ7Y9RLohDimr9Njy5De7ug7Ig616ZgF70ZcwtitiTeJN9ulgLOB4akqZ5+tJ08Rn
PQWHOPMr++7MHc7nDr75FC1tpiHAe9qSCU/DCTE5frY/mvpVOReTddzjHKnvRyiTZ8GPwhP6aofL
gSxySwghVe99uYat/r+1m+V7gPplo/GpSYyWBsa4Ob+dANf78rAMNqy7AyYI9m9ZGYg9lYOuDfbL
iCxKet1ux/vdJ/GToq9S+V94G8MeZWn+futbs4U5CODDj8J3psAOVp7+VEKV4EQBFnyNZLSAh/5p
UMHqGkYsjvj/cUwE1hVK2SRyfRbDF5La8pXBUYQgwN9Aleqg675vB3DMOfQ0Auk9RpRp7IkX5E8h
/hCo8wVw/C2Y6sW1qi1edSqEbD87T4Z97At9k6B6QY7Kp5uzyscRKAck878NJEzXUc/gpcSz28+Y
jk2g5B0TLaZMNi2hL6csOwOT4cIE0dB34nfhOj1mEG8orSww8ZbpOM7mZTgoaf7maC0V6hhWOclR
txSJCEE8MDKd8KT6SFrVyF9rFtyAeTFRQO/IUR7ZKy2EgxW1DQ3V4NLImm0Gcq7dKefEzX+L3X+a
RkxR7iCXMLmYWjTretTem3wfVLAcSNka01MGI/B/Z5l0fgfaVubSw+y2utEdCNTDiSnHBJni4Wca
b+ZVn3al34ebenKqoalGXuof76GQQmtESXt0gRq/1IXtgaPKMzsn9lZMaB6oPhdNahOZhSglQdiy
v/WKVfsWT2ugWwLWHI4eAkSmII4GtnsIsIo62ZmCyauW4r3csGhqnfwJf8pTcftoySqCK3dG8PEm
XVieD1T6qruwac4QWb2Vq3HX5fRuYmm14DSI+e+omTi6BohNNjB/5ygkYNqSBUEcz33K/Pmu4dYK
j97IuubsfKmWFcZIF8zMPRf9ckdQtVp4kM0AmKrSyYns/i4ohhNMUtLWTjIHVaHqb1FM3FbwLmpq
v+U2f+uq+XKoE1SQzbVUY3K1FdupEDg3BVia4A2VbHSS5N4xpeZhiPyKV75yVgmuFledjB/h2tFi
LAqM8Il8VPxpFK7Y/Sr0H1OFPv8VM4Sl7XQk4pTfl+FFbTxTs3RuQdJcxVQL2s13i9sgp/FYASbi
FSf2DbvputRChNhXxfPlt2bveJLoorz/Z+bnH9EIYZdATYVSAcUd5kJ3zkrNPDW+lXqzRFI6eMQE
vH6jkNmKFLglkepHFEMnKnitUTKrGYrpR0mBz4Y0Nv/SkowpBR7V4+dckAIEUxnBT+Vu6dkM4mUt
BPG62F8uDRx3w0/h34jbCNRBuf5BPM+vg7HTvSrbuJ1jFQlA53JiiiabnVh7hMBZkbrXbUPz9LnN
Eu/OA+ujm7eQF3Ynrkpj7SUARwQcXwfAJj1wpo5gsfbOFLu/Vf5WtRY/lwmfXewZk1XOEpOWN3WX
A3Q71MfRE2cRx1i+uLaNHkzj5lke9Fdy9V0hnUv4u7+Czql4M5vPRoZcM+DbN6RlmAkqfvpHdhjR
dOk3XgCCbbKjr8uwSvCHpD/ISARVs5QJe2kuZNoZq18NfwkX8m7v99Q+eOFGfKaiWeNeQHbyPMp1
TOj3n9bF03akbc2KYAyFhquzKHRjQ0ntOO35saSkVKxwiJxthg2xkIFn8scIrAs/eHMHCA7Vfiv+
UsQ4/aDdUkipSx6L3pUjXEdsMmzwdqsKD48a4YvBzd3QURbWRpaLb18Ndpr2qtoNWQVNuw9exNA1
wFJ+BudJOYBZmIf2g3MHWvC2fLZJiQ0IqCk/5wWz+8lUW9b+sDOdaGFxn8B01jg0ReReCbZIlrdy
jT7xD0r8+XfrAKW+CXYRoGav8l1468wHuc2keLafRAQv6gIKJEFmk4k1C80jdXhb2WABc5z0q+KE
cz8KQHtjPbZeD8usXPjspEnjLU4tQoQkyY1saB2AgjI5yFsFAoQinQTegkMJ3g6c1XIlObzdAUjC
e/nWJbbisSdMwjUXtrrYejEIgT9roCMwjIOldGq9E1DzGgYCkJiLmCtE5NsrHcCoL5Y8F0+GRP9a
IPvPmw/bTQv2Os14aqXhK1SOkkT+oZRxa5aXMmh3+50DoKSTcy0ZsaimMBRjLLLucIFvz1g312ep
5Ka5/gU46k5hOSZp7yLL71VTv1pLSL9jRgn1dPohqQ1Wxch8K8u0lXIVvZZeLaMTXNX55O1oX7iz
WQMcrPFYEH6NFuurcieBcprfRdb+8NbxI5fUJDu9yJXzSniKeP3OOLa9KNp7tVV5UyAERpPfmNra
AYd+UFkzn/TuVoNh8a49g+tV18FtSPA6tJDJgnXY9vZTOBPOes3W3dJMEUc+jkG8y+yyHEPSoSrz
bozPINOLcPOHBT23Z+O24jHwJPRehJL12CIYwvcY/W6271qMjIpcK2M34rWcFQDXYeIe7F1NyN55
xBWxZcipmkz3dvLc2+/Q0ZaME7SQ+Q9BromIp526gyBW5pqLqIWkRQrGXNK/uavGK7eoMRr59xXk
gU2A+VTrNaeOdsHlHeNQTDYccHiDDcfXHhptRrCRYUXfh8ox7CIvmDbtPpBlWKCfYBKjIwL4YNDO
tJV4j4AuYAeQsLi3RMsa7s2pe+W60av+mwAD+nr2OkWNZaYhbnRNi0000ANjwCkFB+srlGr7fdKB
VKDbPiNjhwBVp/zz5IUePEgCzycym9MgG4Xt/DYiIjtjMuyBm16g7uE4JCtWIoF13ZhWR0hOMT+k
0/fZuPMQoudoSOqUFO5GV2gH9Sqdaqlk+J5mpaWSihtkvllEWAzJ+vORh7/Fw2IHEM1nZhyGrlfD
m9s/TAwPSf2O3oHjoBCNltvkUzaNV4r9WahY6Vx2mGzCbxvZS2xLHI5E2ikad34B9ccR0UtYundu
E8uKYxp02Ru5Aaae1BBPgkJqzOdLYSlQq/fEE1V2gG00yj95h60PklqlkBZ0H4Lf99D/9+7dMImQ
zynsL1JIdu4rRqZdm5/xcATd3b5Ou7bNF8dmuxuh076tnPzYZElpbYtSaIpSXL2hYdZ/DO51ppYF
uaWQToK1Bv4gObPogGPeLeipvtO9QdqizCl4RjCXn6anHlVVUpvE4aec/LnrBXAmLEQ37Eclarlj
BlzlyZnQLaAnfKu+LA/P/N2aQA5jKf3BoDhXz0KCB/ljHIfur5Hh4TLs7P7PwCIxx/kljTsssNpx
2Pa0WNJnZ71QXbXVGSvyauTe1cJOWZybXYiP4MEexWXWf/Xg8dTN8imEW/QIzhU8AZ/7dO4GN1+q
p0iw1jbCh5kJvQK4FJ98mmR5sAkpcrFHRcDiu7Twdh/1bQfD2lfq+l1a+bR8Baoit2Y4BooLk+T4
jGlUYNZb/T3CoPAPgRYAiZJ05aqpsscWaCmNefGX1a4XmA1C3e3yJVaPPPW/F3obX+acUhHKEOXc
NkZjBzJIfbA9cjsskSRW7xrkPpSKLfsgPeRFzERPBCBi9lz6r6f6Fsmx/meFEeBYsMZcvT1yHnfm
a4cxWWt8wj1e2PS1pIufdo0e3PQj3BtcAhILLpgMYe5SMWaYb3WzfzZB6bo7J05/jG5cszMY4YIZ
55lLDRmVTmYMHw9R8j8jkgMrw4eGLeZ8yk3D3fb/CNI5kwdBM1v2uUo/1AHcEZWL6wXcEOEqvxjp
n8+Eg7qHHa/ukPijDA5vCz5nJu7L6K1hmtic1B+wOj2In4PGJWZt0al7NGDlRCYSjl1nhZrXS8cu
aeTmpgPREP7m+NgnTuT3rtWJu+HDu7hi/W79jrIoJfLF4Gl459SatiM1sq7aaG6ou9JPtCESJFU7
KHvkhFeTTUu63UMx9GiefjuaobMMaI2jpkiM+B+6e3Xqc793t6f+XibPhc06bZiOoleVEeQ5OVB+
Yla4M8KpbnmYooYO5B7KgacLEVfoRpq2kkwePrxCNbk9ELRPhBkZ+ZtgNNg/RTKVkXbdT/GgEs9l
265kevHgeX8OUrq7G5yT9uL/0TKmuC2kwk0xEZm0BLHO8rW9S1EcSvI6EIEQM3LfgLfRMjX7cdkO
6yLKjctHJB3hMjiudu50ypkQ9/cQrxLql7pSnla/rdjcGPfec4ftQH1z88s5qAbk+yASla9aOedX
OPF6wF8wWsmKMGxTh+lynB3cz/MFXVyTAO/E22yGCZno8JYjeCXCN4GIYfrpNwIuCm8lgDEEjCsn
ZS1ziIzj0Zig0dxu0QKtgRoHPw9+m+hohlluq3mS+pj9c06EdHnVkU9XfustOo8eF1DyVm4TpfD4
tf+VAjcEvD49qkaLeBIf0RpiuDitV37NamiFHmoHjbsRTfVTr4HUld8+FN1a5P0uFfBSUTYnMfnz
MXgJgus+8LzPk7OLtSSEoFBX+WI/XsyJoE8gHLusreas6mq2XtLJKEfxJLl+kaywhbfNITQyWpC6
TztE9EYodBergTblBwNySobSEofSPpORbLEDmdZGLoIrU/BZBP3hZXpFrRtildG32n2ENOl3exyz
j6JSb/o6nxfXha8DSKpRICWpbTvWAhE6Cjp79KPX97Be/0FkTyn6yDeYOiPNyoIeyIQYBL23IN8c
5t8y0ijUMKcI9wMT8xCT9c7qbhO5tpLQqeJoqE3sf1Yx3WwUxdULwXF5qI0guzKlnPkkAKByOorB
TI0f0cWTNcusDn+NM06pJheNmmeehI3Gk5LB1+Nwo9kwfzouubejjS3EA6dAJmnNAjCuehbT0DER
41OevjDI0X3RecEJF2KcjTXWwbBrgMQzh3LJwzJy+A1OlUMa6F4l7tuLkn2U99uPYdplRwGwbvRl
x7TGL+PRlgC7+e0ITPO9ATvs+lZ9U4p+ubUte75mPgZMnDfULOTYODtERNPvDNAHbedkzqfAEeTZ
xnHHKAh7GhE6guZJA2aOsjh95pt7sE4XHaNXnhhbzmj7VwtHr2mOgdjmbcvt8HbbIZdZCP9HdmMz
1TE5gUaxJF83aUCmFcXuPibJzUDZ+rrbW4RiKZNNGtg363dAd76Znggb4U7Y0FR3padqZ+o/z3wa
gDLhlxxd+hRZh1to/Dxbh6NtYGkMZxhh58v9Ql7192wcKhEVjjgE1ensHEY6DnK0yuhDfGyWtdoL
aMt2p/zvlXlvH57ifaK8MjJaNkPQSYbLTeBIG3+wwkplZ9+YD36Zz5Hv8ZMN33cKSYEVMSEcoOkO
FCBRP4E1YAAZ8to1diMdCqXm0HCM7jdtcEaMxvuOfrvRSdQSLT7hMmDqF/52HSlF8eHZctnbL0Tf
j11Pym9xe7GemgTTmaJqgmWuH4KreVcJg9/i6mqLbb3Lk90Gy5P/kCGBYGM4FKKwcCrbz7hfbao/
LtRbmVhKyA3QZ6Sia7bloadVZzUWiCEpyq4eysAT1y+D04JJaQa9KrSfU/HZO9E6ycCic5kAAPwo
9zTLqNAwRye9GIAeIGslesOTNKcwqAeQptyTGm5sbyyqxv90tQpQqS9AdpNrsL7lQZMFcZWtbMhu
d1KwSqHkABPp/hi91C20BtaOkE+tmlEiqOelTgpgLQ3dAxFgpMIhQS+XvKX1eohZIjfdJi2Owxhw
YVCo427rTk7uHf2Ht9duov76QnWp11jbBkU3aOUk1bTKulihP6YM/JndB4/4mHbufxAJTWlszF5P
vQT8v4PnjGu+ZrEyHxA8Hx8l2rvwluB67r98JncYFQ81pmHEzkmxcK1vYF9ByI/HoSMpSscuOiub
w7OPZZsMHFRg+Y90ikUB7lrm5JsG77R0LGwPTXjwtdizkkrp6/AEv2AGx66SnfsclS7Bwq9si2fX
DHQZsfmc8Rth4d4Klrao+C1FWv5hl5fbkWayt8HbXeIp9KNa5USgbWt3CdygtwlM63Ad7RN5iZ+x
+q+RpeIjZuOfBRPKvjuibGwBMLkCANsraxn+TSauNuyBsjLViweN0LI6VU7aWS71nHli/UvOmQNc
QdqhCSyBYt9h/nYbpgPm9M7A3EKlEo36qV2rMPgg1mFKTB22nUnGYm+xDW4WPYy5I+kPfZIxSeJN
LvOQH0ENSSzDiS4c1kSzH7y33GTKYhx0c0i1zrtujhWhSaY9Yxb8pdFbeTfsRA6vS+oP0Ct9lNvl
ElNhCziBBuxLmuiNqpXbgkCzZpe4h3WqK2yBzzZDZOEgCYDhS8s6HJGp8MHpUo3sI2+Ds2d33RKx
5Y3OB/pkQDAbQuutzyNl776kGybADllJ5UyzpgJfmkmK5tQ+hDbJmdcKoWJft4Nf0BMekLkGc/lt
pf2wtTcWNbqwKUsI80BRRVZLk578IGcp3Nu5ZpGGfMDx28t5B6br8vG5nUL1jLEpco7zOQ+gZTV2
WKeA3LKT+oXiyNA/mUWhdJaCESit6M+GlAIRflRmjPL1SoYghJUsjajRP81fj/kd0N4VNkbrsY5C
8cIWVjC6XXQq5sRtOiYm0/fG/1z9K1EUwKVRfTLx1+LZdR+wmmk5gwM3+wLN/YuyZGoB2bxtrBwL
Gs7hM3QEwtO3DwEj45xwXLnjfRn46cklKIhaceW738epCI6cBwL9C6f0PJaWTjVkUqNCsABQHOVn
oDNRvT15twQi2waElAM2/WUGIpRMz3eFurCxUyRJEyFLAGcCe8dok3FtPA8oQvvVOOIoTU+jWWM3
tzzw0YtmnziDvxulCT2FSyzPeZWt9+7yzGSgK5TvIY1GM/CANAlOkVLiz4fk/ODI25ZvLlGSxjTR
b2OHiFPQ9bTlBEXdOHQ382402WumPJlWYonjTSTRjoGIAU3Uux0ngRcQb3ku9RwDHQ+7hVb/GL56
+kS9GyWZNcYM0FfP7U4lvwOwZHo3COPQ3v9hlrh1ZBJqoSTOfEwrz1TS/h4/Mr+1frpoEoaMU8/2
BDgfG+UjeoYkeyD4XVWADeb2MU77dOyjth3mOQWgnCJOi765T0/Ikb5di3kE+TRiDr7QT1Wwtw91
6n8i6GDrBFsiSxjNBVgpwJat+VKa6otNw1fgE+lTc3dKlonwZMdXsc/35SuNqte0iBxS1PBaIRb+
GepUQj+ZWUBSTtzYPOKIH6Yx9Y5BAFdMeB+oxRb84/XxWuUd96hS0BCNGjWpn5G6E8ZPTF1QiXXS
pztHW+VhKnKOVgE8QIQf+HNIfMESSbkalqR7hzSiXZdFmqg8inrGEaG8/r2qd0phGRnXAOwFYGiO
190X1IdXlZ929urK46jHucrjhlvzbEW4tM5yVhcZz95dhtbQ1Cj0Ryxb9nKuwl/Giu78TsFJDd4m
iR8EJXVEFoQ+Lbl/d+2gB02QtVe0BnzjAGnUnj8XU4IL4joD4kyd9uOtCPH/on7r6cI111WS8KCS
3COkQbshxi4JeVefPdU3IUdo1LdNCLtx1CpoQJcHaf8VWWJwINGJlTbIqIB0eu65vT/VSabf2IiQ
O3aYwj1j6K1vDai9IsvKWpQxehthLIZtG9ClBTA7HphtelboF18IIzsKya7TTelWK8JxMzo2icNq
v/4/qYEn2mR0IA+4Ru/8jTGmqXawHeuE3ylWoVydk0g7VGA87ieffqIWSPeC5enbtGDt6xSYHM4O
Y9PDynAEBLhDlUZq5cKSC3m8liG9n6vbz7GlsFKYavdNi6KW/lsUl9biF5+PfU9AxEfUN5UrhHoV
G4YE6tzvH0eNfqnff6XruNtMtliufW9GlzGmUBxt9YxoBrl0rST/pOEzYB7yzbGmVH4OMN1oXf0V
xg29V+WEUPLY5dh2kGpRvYxKyfuPbg4ukYpU77+rZCXF6I6HaCEEn9b3RONQKiWyuw0Q+3jpFL8W
FW6HimF240RdCiD/UaQ4CjjL0GEYIWWgU6YSOKRpXurNSYGgBrK5xhscYPoRXM71D4SniVw7GpNc
0FHD0kFeV7/LWDmFaXFmWaySDwKBd+/yuGJxXWZb0QJKknzfPHRjJ/5+i2SrGfGrJoW+9vPeaTaj
tjZniJXhuG+Vp6dk02O9P2KA7LoYfIL4NQSVsVU9nUwJmpLI6V3KVj/dT6VdoHZZEXqt4rZyfmH4
hP4C2tyU64NfxmOsoxWNkUDDWRogfVA/6WjppXHT8rmO8bfxlu4FgTNeyiHfbNnssdPG4Olgp2O/
oIyCYi1hALBf9TxcoRlZLV9UoPWUtIT+/v1g1pL9dU5hZvNZJRbvyZjyxUBtQSlWJ7YkkS9TS8pP
wl2jAWp9BOetA9hwScX7lxD+ccGG7Dhh9LqBOwv1/pwGUWMtlqe7+9sbDidlSV0uH83Kk6vsVzp4
iASdZgibqIOZecwuORzWp8vZVIm0VqXosmE4nRWip2zXHmb0Ddy6SabNvv3tp3Wo0R7ur4wOn8/3
miT8KiOB0qbFCeGfczXy/0hiRk1pJW5vS+Ew9x6dHxlyJ5kAbSB2d5PdVhKr9Ywc4weVN54lvhwM
Qa2DfKiQQlzQu8KLy2ATEqfOyhXIA+7zlutxKSF09hsRdmsjItKssndBR1ZBW6lf2kGp1dvPD/on
V9Kzp86pPd19qwCCjQIUQlSTQ7fqsJaioM3U5Z6HY6c3jiiHEhUF626fYmJmQBb7mgCNB+sWme6J
yjRr4E7J8OySJ5U0Uwj0bzUAf8pg2+m3o0jGt0YbGRR0zjd5FO9cj4FxnvNnfKfUUbkttjRtcr5g
TB6oHum9MperRsJ1waeMR4XI1JMEoPId/yHMtQ8I8nGYhwyg6OQcY6wzNEN5VF9eiYMBug0chclZ
IZscvJb6PTLASfHxg6QRzfgrfD/E/gCRfMVkEasVpUQ9B+QdE/5mJbWAjoISPfTcNxHeAWKUhnFs
VyQ42J/gyRpV4tQKJv5Pv8CNv3dSvdg68gKGLOnsipnFZDWCy/rpVqehx3bGK8Mi3uWdgYjGpZpy
gUAbwdax1BU0lSe6xNXP0kVqWLIIQp+psPjQw0m2ZMhEc2yZawkWo9wuJQurcv0d6iVIVBGg8NOX
49gL//3iJ+g952dr9YYqucowQiNn5Aaag2dIfn4ufNQO8cgwJsW95omfEW/To0Bysl82wUCkWr2X
o4PN6rKOQ5C8nqL0uS6x3tQf8pk1eRx7rWk73Y1Zj1IwjPn3XYziAH+uIKspDJH3pACy/RnBMKSs
Ivme1994LHagiM9xGN2z6TujdAenzhOljY36MpMOCOrElt8+78+Vbbt0WIPVpxU+ag0EJ067V5hN
LShXVs0Z9zcgYVRStvBk/pTBlPmIaEUaBz4Uy9NQ+KImpkeSlEgqI5UQq/OUhBBdQGN5K53Z8NrG
gD/hC5MA3W6SP/rp4GWSsxVerBFAKmOtls6JGB+Fb8NwNwOb3oWRIU+VHKtOazF/mqYK9YhvnPd8
LkCHMh0py6VYvddXx/rEWZkqVxYfL0HLexLo5Ydo1rziw9X4dQ/AeqAe0+VqjDkt3LvMATqu2kHB
CXozJR7ADl8XqtxaCsNFCbDhDGQMnGccyWyyQNBoxL2ou9hUbpdMFxD/ztqpMNtdp62wwRY4E7DR
KO6lCXjEPid3bNLFybeQUYdG/wP7PN5k8hhNXaUCIwvx/xLCZWm4U45WjcURiRWs4QVjq3ec05A7
LocW7Imj7LxMlF5ksR89kquEbXqew0NQoRq+aSGI/D3PXJ+Plmh6idw+OwYgzqqHCoFIyIWnYB3T
e0ptPQTmQmu1YWGDk9qFR8QqYaw6AlRm/dIBpr3Rcxdq1Kn6SHUUROYOdztlvqOzRqpAS2NbVYRa
HWjNRzz6s9yMzINgav34z61AIQ68CtM6RQOy2mMayiQpSixyG1VbKsmTmCKi5fBPyXCOWmUb1LYF
W1VuOX3qTEA2UowtUblit03ewj72+jSFiw8iqpUtiPabjvKU04OcaWoQwLJH/it5vWU6dissxg6y
Rx8VZV/vOLSdtTFdyq5Q8JbP+gZ6kPwOCysQEFbiVPqo/KpViScBhpCkfclnonX4ZnLDGXhrf4wG
pBpbdeCQH1RrTB21+QIfyj/jJb2pFew1wNaO3nSTXJQtmOGQilleXdN0JQvfb798rWUpc0S1COg2
HIAZklqV9Z7HYrlLoFJK7vmiF/dZm1gmaH4/g+lXqXEER5jjQ7CsMMXzMWHCUBvxOJCbJl53e50u
rEyiYZPpRvxiYz0X8FCt+975iOeywvk13dSxh+68fGb3HIDZuQzK4wHMOVBp0BQCa4OcyDxLx3uo
KDxd2A7QFK+5wu039YiAS0ifFht+drWeaImE7cvqx4VeLcAi8sgKGrXypWptaLwsj9mnlHnS/mBE
ioi32+I6ZnWtap+4CeuHgbzf+E0BCZMV8CJeo6RJvrki2FGAyYDZSxc6ic6AVoQaV5fwFfLey/Fe
XFWyL0Y+0oWnDKO3mESr/U+VRcnjmkLVMA5GaAr2yxp4hzcJuyH0u1+qz0jiAHvxqsmUOFf2NzJC
Fe6QZ24UYoC/x+dSIMQNcLeG5hGMPTeB7FhNUS35/UrczEeAxf9qzF/ueVlBwLwSFJXRMkqtZXNC
aLorqHcgg0SzQXougmjgHXb0+77JalfJJKASqAWyc9Cyw/41dqKK40TK72In5gIbEEKCk1Z6yuel
qpd7oWnw51vu7X5mZ7zY1mrvTuVeMZI69AP3em3I5ZnIOxBYXOAsA2U20sIbxXxTIWFJT4yek6nQ
EAqhDjqcBSpWO5FV4NZYVLf0xLxKzmza4/koZ4KK67A+fCiPSpx/GmmvXgf6/XeacYld5vKtBKLf
xaQDVGBmCoS3/hUlhRFVwJjrds8YNDtgBsBd/Prs8fAXji5ha4q0/IZxo0TsRX1k15GwQVQ1uSuc
n4ResJ6bxSnQEj9cpmwm5tkkj5VaAS/yLF/BsFngeogfYUccU2tQwkyA3sofsk+PHcIV94t4rpvU
2mJESVqbL98pqKRMW3yLOuMBGTSoWi2n6UOMxCouwbJg6aNtEvPva5Eov6QdDgbJ0c+xSSJB8oji
nhLLh0hVz4KLsQ3hqABxutMjJrTr32zUYWEQvRnoOZITCJxArJ4eJDD4p6qKFkhZMWaXhIgeu88b
bJth9yDX6MAwFiiY3wZFniV32r8NRiLzroZxKzgSyN2cj2RrbP18YrGj6bHUxMX/YBaZ9a0+q7b1
5bzGuTvZhjGRFgggExYSftZJVQsJxzqQW5rydOovsI6muMQVwM0H+z7XpMX+qgmNDWYM47jPtaa4
zuqvvlwqxYyiiC8qR3Fs5fOZS0gpu61/GZThkO03V2Qyt2F7gAF15F/SaB/Qqo7uXeBp8hJ524B6
PVem9QniM16PMYtJG3++zym5e/qxZ73zefIjD8Y0q1yyqM9umbRKDAcX32P/vbNwWFRC6wXwo1uN
nCaF04ToHh9d0WKvv04iUC/r3ACsZvJ3yPC51P8ip2bbmCnD8fa2k12bPNHnH7US28UKad770JBQ
BEHCDDBhJ6raJrsVLxcyFlZR+x1B/3w6XJt6ax9v4wOPP0aPPS1uxBko6Rs7diW17ZkvSDO6ROI2
CJ+tYkkSRwZlTsno0qiycWjRV65/G+GW3JJVfItYydtSZXtK5i911EoF33yizV/jmY5yH8JyjtKX
zHIW319nvT1cn3TiH5lHukAHUiTlwXsq7yZWQd/YoxWKz7ghZSb1zrOTXh/laVd1Io/72jTJGaMA
Q/RYSekkRepVDgQRy5eYhNHjWPlh4zLVgJgK7k/2TDWveCZRkXaHU3gv2w4IqMPZsvefWtOpuv7D
W+6no2adLy3QpuWgDQ9QUEjU+ogmKyd2a3YhpsIBMOYe83sRMQDfOmu3NnNSsDwouJ6lh+rdvWr/
c93Enls2a+dEnoNe/axKGzgpAS0I5OBZAK85wWn91f4+2bTizRxrkKZvRod/xiN/Ai6VNAkH+eLc
8AF9H96Q2vkbnqaWigp1nbMswbzVGyVoK1t2ZZasIhhG/jp8syOZthHor78QejPohatTQd5JvdYM
AGD26KzJIfjzV8We7uNgRoJcrzFR4zjkVoV8pqCrmA4F1MTVngyWH99wHqG3xqDcTVgxN6909BB5
byMy48peB0wQcx71cxFXQpCmSREyq8+eGS3TO0IFHOBe9XBtbVCWK5OFEulWE6iNIEPTqZ/6z4C5
Xvdzb/sT2kJniZ9CAhhcTMu4aJhf7CnufHpJIRacs4jFsEfr+IyMI8xjgQQQgwUOqXx+TMvqsRJo
Fy3zsO7CC09nkbuiDzqHhaarGucYaYzt+v+jAS20kUiLeqfbAEMqmxOcH3YjcjIOc7S4JsvkrqLg
FCKM8KkpzR8a9VH2Ekr3MV/cNsq4FFprkVrX2KzYpRd7RMaYT9kzcmg/vRPsApWBIrN9TzFPukq7
pD9NTvyFE7zMO8R4FC8fZ7TF/XoWiTbGKE9OgZ39iwMMw6Dt+9OTmxCwrCHQRd8Bmhvcsu+zOUB/
UJ+1QiBklxUpzRZSVxNNQsm/cna1jN5+ZSkuEMtvsjc2XUYJ12/SsBZS/ZiK+xfRAoICKBXY8ZLC
rh13pBOtfovMZc4JiEQnfqR9C0NY9Mv5MKF6V1k20HFbVQuGfLxHziL7L6SypTP1pwZDjfzGt6+v
d+CNOAwJzKd2G0iDapo8b+g+K3hqrtEC2ovIWScXxZLpPEGGud/epru12ObejOT3XvyX+WAsxJZI
Kci3Zfdoq99cmeIzSMamQ568ZCP0rKddU47rywCZmiBMFz+4/GyibzwQGIEH3LQ8750wS49k/6TI
1WvhuYPWgC4+LE/+MZRsXpdxJFmUX0SDGaBcgoau5tnq4QetUvyF0JFZyvaqb5V7i5tblBAB4Ror
E/uxwXYOpT0u7vxS0tgzBzlXfug9gBUHmCqbKrq+jvkVyND1RnWFjgyljWSPHmkUpavm6mE5ptOz
Nvs45c3cnuli+v7GcJB2n21irX1daob3KjYQwSoOD/nnuJ7G1vKxJXeup+BQR5lRz0UnS4JithJG
NftlvhZNvUuqkj2H0AJ5d8LDm2Ix3kyOlmyv8hMMSIW1Afk8mSzdcpOUGmhf+fScUMp1551acuVP
fzbeIkBfCYrBS2qF+dlZhn3mlv7xUdRfb7fhZZp4fPZKRdV4Tu/SIUToDc0c4OU0XQGTHxTPLOXu
gimzxBM/5SSAtmp1CUAEVe9nuUqz3Prf7/NM5625Kz1/hnBBdruz01VRppIo7VaEOHDgwqTynuvM
mkT6jbxwGpvpUs5CSa76bxcoGVMXIfh9xa0xTNPRzjKYaaKSrG4gNjMZ1oPlbsBacdIyFzaPehao
fd5n/RgidmrSHijrRzH8G+GlOWrfADF8DpdsPoyiNXllJeWITaVkyf8JOYdZUNFNU/hjWHhzCVwk
pYP0m0cTupmePddc0Krr64XQ+hsmJo7ql0WSphzzXQgDmA/Lrf4wjoeqmdhOdxP4+JfCqsTvbjw5
kxceEvCxkx+k2gS17ce1hpWc+snN0/19tbNhNBM7gTROvPp/+5AchMWmJ3y7diuWjrj4/z59q4UW
zpOG20M/6xMzC+FkrMZJdipYsHKttBvpg5MbFPI4EynxtK8/dGENFo2RRZvqMJltKjnfUbS2agxG
efhNPe5PxE0yN2K8nlEOsrrpzudtdxXl9LeHTh9F0TuVbFMpd5o7IDgbFIiC6kt6a9T9ax2LE0tm
oygLXiB7wZlambEZCIyAUy3GK2clWccpNAcR79ySQ4DxW/ye7CbgdUriyBFkTyij6tLxdYalMd1e
9X9/E5W+Fn0G1492cDCO5pVxJ+jCfpZfGGyeZtjdjKcqUWtsNnVUoQlUTEkS40rIS/lBqUUaoxAq
XzYKrDy3gz5ff9fsF/QK3ehZ1ETyigVjAsA0Rp/yGhSRznEFlouSNc6BNCuyRZnDrWjZE9IsrLhJ
CzBX4r/2naqq06YO73yP7TEtxeKNvLrmm4b4JeS0MmCh3R3O7LaY4vOENgM5zFU4i7mW9qM3xCyW
Q9VtRSNXxJsNtSPB83YseOMEK8e26oAHUznqrxg5183p3R+oN6UCH2SZg1ZcFwgHIpcOgw5Dm6k0
OouNzJeaC75c21BTGObJJrPo7tfeqbcv8Kose6ymoCxZmFz786rpcs18FeiVTH98SoSldKLk1iGL
/KcyI+QxndfqniYcvWH9l3mJRG67MtbBzfjPaOnekbBDFYlM/SsjpS8Sh7KbMC3/sFyns8tSDuR3
MYVvAG8mK/x/s12BeBTx2gjOUKE6IeVUGlm1jM+gAOR/avbsGU6hIq3TrcO9IcMbVDyrB8RtLQbN
Tc4HlSGCOVIBogyKcVBVSCeL2SXaObp1rq60G+SJRseiH8GsGrO7u6iuRmPBCcd0vr2MMN2kqYGJ
onQ3MLHUzcFIX3Cfg/D3sLr0hELoGEoRSKPO/nLuM2vS1yhS62ZQUV16LZA1HAH1VPQ/vsZcgF8p
8Q99IJ1HH5mvlm+yUAuAlX2AUWyW74fwybWq2qDBvyij1cEb4TgkqvlqfxW9Mo+C4TCB9PoRfndI
BZCl4tPEySPayKhg62m/ABVvLNqM0+HsaW3qzJn23Rs/Bt5RHjKNUxtS7S24IccsBFGLrT7PF7Nj
IL02ipzdaqMlPZO6G0WzWvTgTDD01GO67xNqK9esMn3zOPHb0fjpyrk2qGDsLgjkRlYJhwWg5scv
UdcjouYDBFTpoqFl3KJj4IGGXm5LrOkYYIPtHMhwECZ+Vs/cLgppuvYhnQNDeen9AED3rLiz0vzn
NfxNHvS+sbNoM0L7XxoOKQFx9Eh1LLSXQ+wi/x1s1HmlGWRnvSPT4o4RMr+0oWrpjqByhnW87IK9
F2Qt0LIYkUGALQ5hSlFjhBH3huVSzA0OBQovsmrPkSzd9Y0u6SzH5iYTVA0gQKxNjSYR4RbQ1ehV
45I4Afhbq7Jb6GQIkWCAgMW1DOXZ5xwooBZgfWgVEHnctSEefMafX+jQSow39KhwrxyBvLRE+XUB
ySAt5aSoSLcDu+5xj+6fGdzy2KSC3A8VLG9alN5N0iq+a1ijtnwvx1dgCl1ZMAYRKL4IFhyJO87m
C5/C13zMDGgDNunfmdrX4JRroMEI+imFGzBu744yPBwrMW9YTyMlFQL4LPgdRsOXyJwKPtbt0UZe
QBdY+IOF11TWf1JdXUXl9daLPdrj6akcIMzrOWtD86cL/1qVcvp75+iA0PK7DdoowxmUUCSgXCa0
Yw0HGiXFcjr89ihEkE8Z0qAK8a9xDpQEDlDEWdqicJZO67qRV9bLwWyKA8w0PP24Vm/VfdNay7nJ
BwY/IaZjZn/BQddc+nMC7YvB9dwWTiwfzgBN7xS3MeaGgn36y03ml+5jBX/c30VZNzDlwbkCQ++l
E2v9W/bNxUK7s+Yz9wvy4x2vD3aaAzW0beTfbc++rdLjY3hgl8Mt+fGO6aKJrPRYb73+uLPaRFQH
C88YZNJwZl4vOWoj5luEC8O02pmmR2i78wblVZ0pw26ObETM1OzWjvUKNQfuUBRBlMXdfUC9L1Yw
+4QScLXD448+r12WOV6xxL29tN4iQupv0gnxCtkSqMOAuA7B7DuEwCkjF84gOIwegWHUJvGCOqzw
O7aVb9sRu9PaglrYieW2pva+1sn7zzQNPvmmZQlcvP4IiOcsFVH3pUaiZ2PSpXdzyeuN3GnqbIzs
sThE4e24r1MRCCj/DE48Hz9OFAIQPDzemX5z7aYy744dz3KKkKsAFkbPz2XC+TGOgtImTxLi+aji
BSvgVPmstq2qsLxUOV+KLrnQXBVlggECYjAO8md7k8r9kNqDxeLI+lIwutqYox6TXdK0PmClOUQW
OhAK+IWtjaarfN+r5F3TSVGlw660dRNSz01ossoOJgVLwFJF5Th9h7uQ0XI5mb1xYXHAk+6oeJgW
MPNcm57Ydxvp0KQ2ItheKjkzPCB3XiCE7m6udlyhJRtmurKp3CjGWbnmk1sgNJO5IrbOCIctcSzl
cLN6rMM9A4TdjBPzlsLHLIJsufpTg5/9talyEDYtTPZr/0RRwVK7bCHMXmvl20u7rK4rOz+t7deC
1QzIydclR0RN7/PuS0IobcB2DDPNkweIdfCI3Xg75/2pD4EQBEkyRt8ewoEy5Jb96uey9HI0hztj
+TSGDnyN0Uzh3YuirobdNza39yGBKj/fKy6BWM3Lf+P5N3zdYopl9QEd4py2dDEIcfTzsy32xmX5
NGf3W7mWmv5SkCu6jh4ESeAjuHbdMK7Pk3LeS1rieb4aQy/dc5PjyGfGjD3ey2Nk8JFS7ojv6PZi
osWH3nvB0MThDQnTyypigJ53+dPHmpqgi9zWiNp0rR6sCJ+rzk6Iz9LssMRjyK1LDIQYG8JwPtTx
64A7WZlynNV+UZw82nSDxyfNEUl9fQ+orMJpWSzoc3+PlKH+MIS2VquS/RLrdu0HjJx15DTnPKpb
9/rTmxFLwX4cIc6gI7xHv6g3qQjzExA3xZJ2/Bu5d4jTCHBAx4CNM1pfK7+Bo4udtbAu9BrKu9Zt
a6hK9Bcab/zW2J/m3NRHe605yzEh2HESrMUGGZyvEgf6oP6INM7K5Qx/h72YDxNxutEs3AOTLhlu
QzrSXhqIqdbxb035S124MXgcv0tCy4fwSvRgqmuFn9lXyBbfFgjkJ/Og6bFNVVn7iELSICycEKQW
pQ7VZRCwamJTzGf9gt4PMC4lrLfo6SEQx1jbMI1cUZb1Jrun37T/yB5QvFMMYxT8xPb4TxxTKnRi
MFesMPbhaI7J/DWZr1SER9glaBpPIT4XTPsZYRjytnJ3WcMl/I8vM8uIcerIUD44RlOZWKMURpjs
LLyNhwINTbAbiwPZbGYljeL3bGg1B601U4VvKqAhr65+k1KjZfgpm0b4SkvCLLZsL4I5f3gMpbNW
l+vALmmU5sV0F9tisBC8gIxEtcy/trtjhKRmkIgLbwqn9CmoNqtnEx27ukttA7DefZvFQjtVg/mc
9HBphLciNgfIWt2iD21GDE19B69QhexYyrhpzK9vcgCEbPovEyRRk5Eos1DKQpMgOdEKrTZLynng
SPueRU833q0PFQ3xTO7JEqV61Tggh5FvVbBHWf6cmpYisEpqyAOS0hBBFL4LGk656xOJ/Wu92DkH
OS59IjZblBhqecWHfV+iX07N6NN9KgGj23ya6hb2O1mLhw6lMPHKwgdQP07koPDJtWiVXkmUzrZL
r+R+9TdQTelDN8a6MNKs7TCsX7TaUoEPTK+g2356FI4nkz0HXqhO5AFy1HcNid8SE6G9khhHsS6d
NyP2iurJP/OfwII294x9GvF28fK1wb+gkY0pJJuIDBpNTlZuATOV1hlEvzWLt39cWfHIge0kBPVL
wnxIDiEVmRQUU6StI9gvZ+ZZtUXgXxP4QkTY3HElHDP8UL+Y4F+vxtTjfeXEbmUBeuv8hPAuP9Kh
86YV2/7lR8GrSa7p8Jrug9mWSY3D9aVQrK7NrAb3XMfgralUEmVZ7GMSR1UEbk/3iWckKZ8zqzcg
XyeCbaa1ZTkLlMSCFMOJC+p0g1QA3WDC9799k+L26pVX/kNnAHb7xRDzvs74A2i65zKYExEAU13B
lp0qDO7TE/9ZUoRIMNnTLaa06VELmawJZ4anZRZlENN5PzjFH8Vn4w/ZwP0PoQ0ma1NtxWxBN0F5
1rvjvz9DtWsVDam3668RJCPk83FSUw+2hY9+DcOdPnraCCbcT4UvPpuT3aYIKwhhCFPvRE9YGeQW
QQGQleW6sCT+CxIk9S9kMJMPg8m/OI5PCawens1xzAz7MJ8RgKYBTFLYJpY3Tzy4noCYv+j1OSUr
iNupucWKqy+ZDT9loV43+ZiO4otF+oJL5R7UZeNG0oVYT0Nbx2g5vd6+DJvaUmngcnPSh8/dxVwS
KsZWqfTOkEehC457YmpuXzp/YvCf+36Nzby2ODiKlBJlE3xKJnvzVBWZhh1C+anpSgsWiRg+Grgl
yf9pJOoZkgHnmqQHmKP14DrzwFwjXfdL78Y9ug4ebvnuuhvV7ofNqNNvwtHokHuyYVASNSCuxXnp
cYmrWfNmsHJfqDwDb8TMhgYb0EFWU+eHnXZkGg3iHzGaZiBZP9jOvJq9Dd3P3aEsIyw3hXlIFji9
T1V/xz/XLHYwk9GPB4Grj2ws2NvtvCZhEs8ibTjyjN/zqsmxhpKy7mqL3r3gnndbnNrrWSmw+Btl
BuZlW8R15HuBxPuwE4tmUfG64qhjD5ZSrBhxlfutatixBDKoYFRAtwGmHcIr1vcVihs5ddsHZmWU
hvsaGGJpRB/PO6FarfKoYDbbF64mqk885nGyLr2FCCmxosOHlgNusnYivEkWa3dfu8UKfVyaNvdK
LPmjxLflc5yaT162yQEsNpegR5MYwbK2nZazTTGeNi+iUiHfXWR5uuzRErnTWM4rdi3seq7V2MFQ
wj1OhfNvaztxTjRzfRYUhwznUXmFSyTd+qFD+cr0cxgRa8czXGaNMOqdd8zQ2tw2OLesN1v0o/NI
1bpzeFfkgEZ44Uwh6dhcFdV6ShxgqmNcAbCq3in3q+RR3L5FyYxcooMARIS1aXG8tvSZ+umKBm2+
Dq+Hw3O9MCet2M64culpEJdWRBKbRGZ+gBrv1JKbA7DepF2GcvPnOPxPx6sU/ABQpeMmdOxxYdI1
b9fXWPbmWa2BYPVMMQQuVAdAv0MSSBzUZXkFSsqulo/3zQP5D8GPX++pp7S3xExN0q1Q2EYOaHPO
U7ss7gVyVTNVRq6+ENekZdQcmgNFvnojxvREySYEVKU+TrLajnM1UBV1/kQAxe/L7S289s7Js4eu
6jnrzbAqapaIfIY5DjZj9VFON8dDfuIlEYGeoy/peUIIy+cZ5dwRE4qV6Fg9AkVVr5pGpkGTwAbX
BqfJj97yjk4bBSijC/Dmb44rO6YThrnTq2dVTmkXUOWdt1bvGtLSk7QjZFc+Z/t7kLG0ao2Fudvi
UYp0Yrn0sFOA8w3gIlYHSXUyRgfJUUAC+pp7sKS3nIlMNTc4pdNhJQsTVJTcgQsZLOOw1wHYgt33
8dYKY3yL65H2c8wvcXpDi5FxpzVCpcOWbuxxihA7Iok3FHFKk5WL6eYCtJ1iOaCpX21+1b6U5fZl
azDKkuF6I9vKURFNUDSGyuTZkaouPcusaTq52RL0NB8W0FC3jcZFG4dQBWEngnvO8d4Kh9gVDyMo
FMqSIs/1R8XrCGHG9rifRsa3oPgL7wa10ysBxpRvlt9TsyWLVAa8QSqVOEy+6HIQZQnvLcCAAuL8
Xraq6hm91tJv20cOEQ7JlSAXB+Ja1a/jG7XMQOwUNbSxu989yqO43WBHavE9yD9HAG86SrynTAga
FfF8l003BFV1sGjHWd2GXeumo19B6OHebfrMce/S+uopFiukgLOruC+q+asrZSfQf7gDHnpYSob8
kAjUKgurF/nWBrzYQtkCiZvwmM9cArtW76Kz+4S6wl8UMdi7c6vqh/odOBRfNpoMzg/84a0XGL/1
zmUU5BAr9vEMXCCHN2189HXxC3gng6Lar+RxLMsDSunicO59Jw3RQy25enPbsBQ8y9yhYctLV22R
pSqkig36e07AGj6zcD+StAsHygyqky0rrCzLqi3Lgn7tYEySDBgS6LOdfDDEV0PvVEHvCYnMAm6i
mZW1gvWCGHwAFzBYE7j2h5Py1DDiqfD1+BTqlJAz9fTEv4YbYVK9v+E0uJuu/l6sZpdHVEHo5LiP
ormZweDXtV2iX0Xfo1DC02Paju2YbBOk7eJiFlQjVNVwTa0reIhyUtWPXUDVyzYBmZi9W/UUsVDh
jJgDgyEQStVE63fh5yK0ZxddIsGYbmfdq/gFF4sTv5U0DmS90hIUbpFZ92iREt+u0/PWM4Z5aWqb
C++Md4qhKQ6ywKpEr6Dn5HXzzY3tZxUTv1aRdj7JdihcVqG4MbGXj2nV5SiyO0eKk5NKVE6Hpf4y
qupgPhnQkosTXDsHoW6FnztSlOZ5PlehJMcbHf68VK6epa0LYYVBui5GfcNu6nd26Vb4aYYVhljy
Yg6niokYpXkZrv74vzwbuBf7XP4Y4Up0RYay5QkC89YrBTYTA23m/7v49xEAKWSwZMR8OnpxCteN
/8HUXMf33JPuXFpzB2Xunrz6ts0KsBPaiLQhIK60R135qwpQz61MYiE9K7DjQEzblLix8uhwFeg2
jUG1arI8PBloiXSIOzwC2fchRtPfu+ALmGmej7GG96hGHYldWzJpQMnVZvLYa90C740VVl3kXHi9
T3YUJS20YlHIkzDZVi9TzS07XRNwwKdMwLL9CW0VAot2i8RctUeZuWDpph8IByPc6B+GHg0FpDYg
h6p5Xir1exdZRwtD6M5on4JHqzgsk5+2MGIDEvzNRclsPl4u9yVhpagAXgSZpHGLiBYx/g9EThB2
wG0jBcxd1wFFDrux4beDraJUJOMTV48XzNY80wAm8GCJCq66Qwx8kZ7JRIG0cO+k+ZEPnmzbxw3Q
fiyL0fN+ZTcAgNR1WioVtHT5IztrsAmIw5Su+SUYN51uBvd4ZHsa0sVbhs50KyrSN9eRsuVcNY/c
avOQA9c2xQjhXXzclU1RTj2bI23ee/HQVYmtkWlVAuZ1icFYERVd9Fwg8TRSapELkey4/ZWkind+
2ZUfhwubjOf9/jYcoxHqUR7DLWXf1vm0BU03RCgqQ0NGR1zLAR9ZOjepbrFCpbV5vzaFc/VOP005
hpx0D54BCr0QfZ9I4hcoqTIJ8rl1nokkI1h2vsKG0Je2H7XoSwEL2iVB1Ce5JF0Bu7QVOdw54KjS
fEq0rgyqtUaWELzPeXIwDsmpYeGTki5gdwotSxdMQAzDIr4/ppEZUrEB3R+fa7Ygaik43y14J87A
6g+S3b1+qzp+FPN6hp9xluEWUuvF3kF7oIx7nJrTQ6ejswDq57vPeQuXlFkWlczSXHRUoWbqntc6
t8lIRO2pkZk8egcyl5c3/vNrzoq05nzMZUpq4/5e1LLmallQaLmNgFyJI9BxXLkv3caCz4Kldwiy
3bN5IavAW6U+JqUpBA9a8oYW53jD8u8OBeCEE97Af0rDgX53C3HWghKAgdo4HhaCUDeJr2kScEL8
3HNYxcEekIr+gxFV5A/x79PQQL9zBP2u3sQVMArQyYDf8W30DK/U1lDoqVtDFp6L9LTQJkNukKde
+LA6x7ka1+IIlZtzQ2yd2QXx/2w2SSvPQtf7sT9A88RbV2tFrtiW6Bs6binznLAxe4/D2nh3Geep
eNeA1wMlkfFwPuHSZzcw3npmN2oMKi2vU3vXdV3f/VJ6PKgP3mCwE7Z6ENKq7FQJVzcEOE9O4TWq
qxKiM0BpBqqbRKSmnUo9o9aPHE6qi8m9fcp5l2tEAp8uCdvu9BhKnieXHDSSmOKdBdO8IbwWGak6
Y1114es+nJy3ETCLCXxIzEkAqvPb+POr8SO8VARP/namG66y/oL1irEZq1LUaMZEhB/t6GETGpem
LvBsmjSx7fkGY+R/yparlGODmEKDXpPG/PZoqtKutks+GRcRUiNZoV0f9mtg11rhj87/ld9GfJ6Z
Gck9a1lHd1MqPMhbgPygslp95KASk1jSoqhPugX3GkU3rtdEV5ICQhpWTtE2/3eKEuJdahIlfeck
O72CKlzkRO6xw69O29ZQ3wC06thtqY8wV6w3JqTMasB4SgTFXVL4IoTSICanGtsEtOav7cUbDvbK
1efyVCqb83nkD12WUkEdKfA5RqlJX89QKrYSW0YLdx/2rSQIC4uZYh6UTNZp2GZ/BrKpnRHzF1WC
zivPGkHPSHtcwbk3LTl0urj8yrbe2SMmFdY4Na0uUwDlWUv9CUE6uRnuS03RHQZUwt+ktzwqXaDG
jdrrT/X4Ze2VjSack3evqwVc5XX7AVNXuPFLiDTK0UpQkpxWlaooD7pyATPOpRPPbsTViv4Dlma6
X6Unzw2cdbuoRp0KbVHVkMywxLsG6Ej2l6o4WueUOko5Jw8eXpaVD824IJV/G753vZWorATx9d0w
9SKYuSyiA0ZElbv3/eOXearT2HgsBHGcRAAZBPMes4vhIa4vHX5j/xX4ksKLJaQfq0bQSlw49+xx
+DgmBZdd0DXCLG8bNlK/3saa0r6IWS9hEu4VoYmmluUSVkYoK8N1n0c+0pU2j+Q5wAIuZ/JymOsW
KOm1N1IflmDwE0/MRnNM3nerzbo/xV4B8gWB7qR6xVoQXw+Tmcd3+REZJnqcfTzycyPszyrjtgur
vr1Z5fSLVgyTtFbI5bmtAG3yqX1cBI1epL7w+FdpH91h0/WvOTI3JLICiN3OPxkG37oQJsuapWZt
6iWW0+Qo0BoUZV8Cs6yHjs4Ng5M9pdwoS4JgkFPsXeDz8aVR9Ftwj8MNb5ApdUaX8dLuP3J2LJ+o
z3k4s1MHnRj03q8LYXQxRQ6OxATqY+9AkW5wq0ma+4AE3GaG3LVDS9patAMWD18HCIlLXb1xD1e6
4bbUUj1AidslGHN1eLWtGco3UStg9+iLKgy3t3Ny/J/c8ERUKqIGKf8KSJiSrGjr3EAsSoOsrg/i
ysDN4SPGPfrGOUlCFtugHG+HptHZLFiETLjW72kjJUlpmkHj+o3nQCOzZqgNoae/XR6TswzlunT9
29I+8X6PCrmA7Y9rSzZT2ZniDtbKrkYJB1iQPGvqWQK96OIJ/eIs0nmJ1TfJUwju/zWlK8TGsCod
umZuOYXPQ/Hvbg04tphTtd00qN7MzVmAi1en/UOUMVTCCWVawYYSFT6UWP5y3c2wniOALqyJvP4A
yPEkmrrr2LwgLJK/QJNprA6eVrXv+jWHLzVY0m3GTSoMaiOOrnzX4tD6VFEeAlClxZxuS6Wqr+4E
NWhAtvAH3N1sz/0dsBnoj4NM9VyF4fg1tTyBiSZWQVInXIupwOt0YwpFagl/6b123GbBTVplxLhV
Q6PirBjCAxAERFlFp66Sa53xGNvt0ccJaD6gjispZmBS6KNTuU/C090ws/JP76SllGyykNznxdh3
KN9WfaJ4HYq+9s0lxV7sR8vfIcE4hU98cLsYN5lsnNIq0txcFDxMZh67oKO9YH4APN9Pmpoo9PH2
T2YMrBDuBqi0yieE9uZFhGn8SU27/Wa/KALmKa6FWz9oi4lDGz13HRFDy+3Q/R0GyvRChGoejPLR
kwC4UcFBmjsVM5goYJBBPJR50Vufq4oNwDj8smQxF/tEjE/9f6yEJyBx7YUrLuQvK44cN5Fmwk3o
cdrJpAVf70kjkD5LbdDOJYkPTmQ/4X3kS2q+P9TdrDk+33bottq5xaR/4ZzEVe475ERVQ55pjgf1
O92hWYEQhJleqw6XQd3hA656iT8BgWjkIUTADswpqfTajv7mZGydPheiXVWudLT4XcK9e3rPeY6R
BjMSwrFPYd5Hmi9+UeCq1GieqVHo+j5DUPFGoai0LyeyZ6RpZAs6odoZl0+7TfwkAywB/mixvRjh
RVlFBGpQAQFfoH9C+vzO9yyVpkVZXFMxDU79Okm5+4C43jh+Cg3juBZpCSQMuFPkvyEM5T5IDPZn
bg7EizoClzmZhqWHrYLMYthhidVd6KdFpY/e9LJujgm+bMMLLn7YvpR0jXlADwFtBp1UlYW/AVsM
mlfnJKIbhLV9wSl194F0agdlV2Pf2K3XMUIBxM64N+AGgXlf4ToWMD9cY5ffmSxHF0qVDAWyL1Dn
7CjoszcuuMw1++9DoKmbrb57EXjb54GXWBLsphtoiL8JLNNlHdw2glqA1vkiBtIRWGWN4u/bNqum
lH3BicWiRBsgx4yq33p3Ari+n4XWCMiQzesRf5R2OC5AvNY0y1D+ND27rINUyzFoux/EzymIE6C+
SPFhX5fps8I2Py2k2VEwvfnkWm9EgpDPIWt/g5uDg0F19d2pkQLhkfosjJDxtSff3vt23+nqI02g
Jv/FgtHjpA4lZc7rPQ2eaaGT7roF4HAmyeAYC5/6qZSDqdc+j+hG3bbqsV+bkaCp4iIC9pAt14EJ
CMTs8Pb+HZa8Ry4FTJBYFMauOACcWLrRfZ2lndnmgs/I+sgG8lWU7AirM3W1QPrgaf0UuVCxANT5
SZ1E85PlKm6w+CU/d116zKYFOhhEAU1AaI05h+m209G93j8mOEJJFcH+/8cIB3CK48TAwvM5wCOZ
HbwAsMatYvkfShxjrDEl9yx+hWT0Zt7q2lFUCiK21irOFkIZ8KW6kIw1i7D5X6v1XUj4gAfIwOXI
KJ3UsnRsPxAh90Yy41PPdvgMQVIkOAPXJ1XGYoPD4Bmyz909/wp0+6kWN+4oixTY5KCI8HdFcLhx
zLrPZkjiI65fOKuiN8xF0HDASvmyqAF0eG/hAWYT4gzuMWccqajn0NXApthTzdqCYWE+ABRk0FZl
PGdSTd8Z6tCzF0m/rug+F+Rjz2xSI/wpYFYOn4F3i7RX/V1XL/oKrh8xId9NXIUEqayxN0EAr7B0
ROS53fflv5/zF9k080JeqGL6/qWDJW9xPPb8npPDEUE67buz/bp3CWGL2re5/c9WcFeNBcX/fbvi
8KO5mK4izp0Ea8n9S6MGkYgmf9LatocxeEUHIlPyAIqBjZHqSRLz0LKtDa9FcefwaVl8bHd6Fmch
bgxElcs/1Qo1Ar8YF1BX5FYm4jmlmPaTt1WeHlF3qcG40ifWNnkxk77gpEVZqA2525jkOt/zfLWi
MrvSC+oqDCGwr3t0VLIHlgXGptQ9e+jk1IOAASZhWl+H5ii4LtrNaZsZbUqNaw0Ud5/xFc/G1ixX
bLI+9Lf0NUb5Q2vRKRQLWDP0+uFwCxJD3N1sTxf0rDAt9ptBczXk+YxeYNyk64Sl/zkMTeoBtAn0
BSPtBA7S1L+kpKomNn8iHI2p1NHZXiA9gRoPz4LMUxtSbgSqc+CODDcQsF+uFX8DQVWMbtpWsTyz
K+C56t5WisHFdqr2p3nunm/3oqRewjeSLeRvuJigICtJKGSjCJn/DhTCXl5VLZIJ0IvViC6uYWjt
yDqAtoA/OEOmqfb7TB44lfvJ0uSPiRgp19cDrdUEMJ6+bu/1/LJ7e5KJ0CnwChcRcgXnTCuQMc+9
8w8+tv5rARPO/d10L5Vtp9JW5gAVZeeN5B6KgrpQWzSDDJ0X752urDqpMXnqYx2N5W39+NrBlleX
yI8KgDWqkiMyrfAmfL82HeEdg/UO5Dj66CAs2+mn83JPgAX8gOAAUamjTq9PK5jKKXzPho1XzVGy
oLdnHlGey5aw0m4WlzQfuev0Rqm3guOyGPW0o2w27HQy4UnT+594pDTFsGozrv4xSuAczk6V7HIo
N5YSj1HykL0UawXKA2pvd50v4QtdPIN35xwFHdvUpb1I97jmKWZkNPSsPECdFkfclJrQ02NmGrfc
KhoD3Y3Oeep4NYN95fN7tLwztyqKjBf71ZxdhH8kWS38gUcY2UH0i0oZpl/zwh6brEuUBcJlarpR
0nQBjR+q8IZGPNiBVkLbN5uwEJIIbmPG9RiYGu2XkDTzNO+qJknKrWRhqOOmhySW6Iq1XTxqUEc+
dIwlw58EJq2nLZPnP+KQ/cIoXzzPISEn094JKRaIlULpidgbh7HHuqRU8A2z1MGHF+LPT2bcuWio
uRPp5Bru2ypTds2KyUkoFIGfHzs8A76qpVL9xiQdHIXV4RD5ljcZqdrwjr5QHBsJaFwzBB8XQCsV
bu3nR3rdeC6YgKM1DRO7NCPRvAk0UR/9srwlZxxD42xNpNM1BFMGjAEkiT9gHuFEH0HA76GazGZY
17dumiyn2E22x1ubbc7sGMqsMq0SGTHjqGW9Y+nTD9NLNoMwXMYjUfj4ApLJVPaWth+A+0+LyRn2
n8lIF3t5Kbls6vUmK0Ib5MVCgS5TiKAeFWxolqIxqT57ksrpgsn1iYKbjIKygYYoGk94AWDvFZ2q
8xZofZX+wtP+qaWc6BFHtgz3OSGgWOiZjmIPcFUtCVAmXwgr5ZHfHWN6vaEaIZoiRNag1U9C0tay
EnY4GCDIhyKtDLtvZ/eWfjHT753UtYpFQlI0w0kJ/ikOKlgl7LDgJtaKSB9pRGkh9RZVkKwsnpjb
r5QFTJNm6dmFIHXehRbjhMua8uCLJA9jTg21YlpOKvcTGhsBqtZTZJayLvYdwYibeJuSssA+ZqEn
bdfAznD6B8yE5uUwN2eKVI9E+/7ww8WLTDBr4dZzKDDvDbYZOe9MWzDBh2McYuZu8FvHBt1eiLVX
eNPFkpBGQv0CsXwSf8/r+Av7Zj2ODn4A0oU+Ea38vaXKGrSVafQqjyUZUZt5WgHHc6yay3tK859F
U2YjUx9gxr4Q0G2sINwp6S+h5ukJfEToF50hhjlYafmLQFWfmDWEi9//aDh9+oC334Sl3NBVYnv5
hTEC6ljqBAdldtZlrAt8Yt7Jf6uSFoXXRju+Y/HA7xnwRQL7If+YxFDgoRXkMb404pSRE9vKVYVC
jGmY5RX7Iuoh+3jACMQyo5mljtUAoHzrJPVwgwXNjq1HNJf69H3y9cdnuixyEJ5G+TJqyiNNHuWD
MC1UzgQ1lAsjuZRXAkctLL0aOIn1kO7utKXOVnuSwCSPWxGdyRbDSZdwI880BICS092QGD9Wza3o
NCYvykTJ7goeHO7CljTHqYduDXMdMN5xCcj/bT2DzVqEKplDgLwE4qn9IMRBq+3dAMkNB8/Tw70Q
l43kbOLWtfOVYJJh+FrL9+afLbgDhmAOIMGJgNCv3TVEy0pQdpZBJa8ln9061vdZahBfhsq2EUDo
2zPYGyMDHFrwK0oHWdOuAzFJ7zXOPD8ghbAJgqOWSDcQKG07JIjW8/GVqor2zplPrq7g7i/KQI5b
alSpJAf0JmRoR07Eol8oQc/KWV3B4imh6p7bNj0FPqtpgXshkBLtP7wnlwoax9Y5VshLDVMMXyvA
OwWWdPSp1SflH3iHwO+FuLabVIjBysg0+gWSwZuKBDWeg+xIveIBWEUJyyS8614vP2m9baTbbVG9
bG7+qz5GUnXmCzMWfgdIRe+pJHTRfMqFmBkr3ow5VN6h94BHCc2azimCpnTw6XFRDuFs1kUoUPpq
H1JNfe7vG4yIrW32GFkl8Uwep49AB7Mt/ewSD8xVFcuOrD0J2YaGEJ9d/Cq5uhHdUeQaE2tTrfwj
254ci/wRhfdC/bBGn+SpVUD/KKhJSUn9+hTp+Q6tWRxV1/4iA+Am77wp7KcwZ09xMvaNURFoJF6I
5AbKs4YD/lvVqbdiXJn3h3mI31zUhVcj+J5Tgbvo0L9kYPjaowYDABfDBiefpvODndMpTcjBbhGl
HHHESafBbedqRFvOj1nu+ImgsVGwe6ioJEHvrERRDcSb7NBvis+GjT2XrcyQNN9ZhsW0qiIFxZNd
9oFfRFOolyP76Wu6ltvqDFHWfmZZpU+K8W3aQXyl66JeTC9w6EnJWeaprMx4UEw8cmObiURwGDI0
HoRpwU0JG7Sv4LVgdYFXfvWMFWN1uVO+znL494nPU/Ye6KWWdRPdMWnddEoajLlxL6xPsOWyPsbY
FZztuBQH9RtMKkZs93sSx4NfgHSDOT1bbtkS1Ntv4xD6WdQKYVUEq0o4WEuoGCV8+B/uidJmPwtu
ogUw8R7dWXJV6SOuoD8zO6TCclTh5MjP4HRxCuKJlc+yzf0VEyJZ/Mlao6rB88CRpVE1pr+TYUbf
/kew1wkc5zvm+mAXOKHfET7P5xhBuET15RVpaa2ZW0Qij8uNkyZfUbo0CoufysS0q1jXTycKNdZQ
e8jn5SPr2YR+qKM9GiYRQa61RlP6iPPdmWPbm+Y3D6n/JEw8jnAfszgOBHMXIrdkXgr0LVNFDZHn
k+k1uHaxKIhw6Vmn6rnyYpE8Gui119lsHmXXjz6kHmDD7hitf2MuPpPhljWCmuU0gTbKal5dhNy6
DXkHNNqwy5d5N+sK26WeXFP3x+sjMXNRLYBA0c85TTZ1g/vnRcgLE3CW52PxWcyhHrLtisfkm1pM
fjBr2+9au1j5UsI58zMCniflyPcS8PQUsVET64eaVVX//dbIP7N70MeyYWxMCgcBHNrkcZkw8YIs
LF61amAYG+74sPuN9RA8n0OP3XWWdtIKF+huLZ+/XSstnJtY1uu3sunMrbN/oE1xQPVEd/D61iN8
8+U7TDzB5Lw42gd+UuOXBOPZzj8K+LceZUNjKu9/TH202dhToF1aRx9FzyLahHZDwxAJdIjKX9dK
EG/VHy3tj/b0wJ+4Qycg4/FW/yNAtSJtiPntC14ojctf5a52O1bSQFvm0eZxU5YvmwBIYltCadnm
iJFrofwVWB4vIJ5eW1zurpxVb4v8RRcRwEcU6HXvFmVjet+UpdIgi2QJ1jGFi8b6nNi2EAT9tcaS
O962WVID0B0A7aKiylkvDe40M8bHEL/cUmwrVxtPNK75+03FkwSPDLGu8K8RMaLqRAORdmvuRiG4
aarEquIk0EOP+2QfgITOPXbl9TG3XGZMEwizpEkADwM/3S9N3KGhqQx/tG5M2rJ/6T87bFHVO+BN
BbdqtD7Jf+Ib9DluVIqA442hS71miQAtzWnMTzWd2Bf1pEGsB+BPFolxal4YfwU6NhtenKzbDZqu
T/ZkPig48CgyWY4d3C+lQoQwXLUsc9T50Lc4fjE1snEOX9YVdfp8d2xBVF589JMFVlJ2tHMO/8ud
2z7x1C7QKaMecpEvnr8W1QbmOJelSQpSUgm0lkjIjL3s2NxCI1hZdQoUhLpmRykn058dXLy+T0rx
8jIndAuuoDIoANevNwUz2K1suR+kyPgtGAEGr5Trnwyl69u8I5Vqa/V5rJpos9mT2IpxGGeRTJb8
rBpUdXZQonh6hCziJY0tyJQCvkgHwSpeL8BdtRjUlrp+R/FrJy0Cdc739icUALQxVYd50HLGDgdp
h4xPQi7QsHXpcVftxKwQvrfxtlFYbd2++Y2AbDkq5yMTBGb3wT1OZc4+jcLHHW0rEQp9E15a7qCe
cymin9Hx3ZMB6HhoWg9ybZXZzjSmJ356olxwMMjF8u5Aexxy2NaVKgcoW8SmBe3opBkYc/no78ZJ
EaJZjO2v2vt4mDcm1Vx0vs606gbtDGdqh9/shpPKMj4vaBpuSV8GydkOfW7P6w5mWY2ZN0dQeYf+
d41E2qiGm1FG+L6M8cVvRjCjge097OMnXWh7NNJI/PxZuo+4M1TkiJ9iO6klUBpZZhQuadYE36xL
oJdWfNt+FDZ/erBSgdQasNWN4MfYBJlYTYkELVUecdCcTaFnlGszMSUEXa/betWZrTRYB8XGbHmu
V3zrs9DXt2D51YGZ/AnZ1WLRnMestdqpn9A59N4+lPZw6mCK5GVOMft9yjCDq23zUIAGuZEwzYz3
4CRE1SbGZqrwUL3SUnscqBb5khjZTJMS+xaf+Z40Pn3Ry5UkmCqK3NsYMffGRU7ktfuQeoyV5Vp7
kQBSFJ32rW4EDxk1X6g8/sjuPeNA6zi1Y7NCFPNcB60htb8a4kfs1P5fs5thBPHPy0meGVInd/dP
70t26JLK0IDleQxfaRwDxdpOTA/RpK8E5zHAAI5UnJboUp6d7JiezHOE4z/GMl6wwLtpNJQa0FAn
JqoNcAUQGJt3ajcb2hRpWkYPuAYRAtF5bFn/sI06XAoiDwQQUZjHY8c3/EDRGOxkWjm1VAZ5Gkrm
MNodAuS7+gTCYCgcgVwMlf/mqyEXj9JbifV7sLajAti+i8zZeznAiDnvg2kEiNNlaycb+4MlgzAY
r95XSOPhFI9iJUlHlY7V++M9vSGcMzRKA/pKoctfzQwyYcxttblrOpHObmq614ys2IZxm7QOltRS
rmTTWGimGDLaEAbQyoMcOTjiWfPVXHV3x6Pth294oFWcJ0R+DIrMcEPKcnAabsJwSO/mhwKPRW2/
VWeTvWb9
`protect end_protected
