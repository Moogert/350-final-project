��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.hq>dT?j�6� h�6l��h��u����5Ag;�7`�}�0�b�MC�A1D����4P�c�lz�#��l����hi�[�`]�q�7Aۭ4�Tvl����ٶM�NH!���q�+�:���.|�����X�z4��<��#��T��ɜ��j\��ȳ��'��mK0E��F����p V٫�p,�$ov{c_n���Wԉ��jׅ���<n� TƮ	�[�^	�6(�k���PUz�zXU��&�@PzP1s "��Y���l���������e�T����{��)��v�
j�£`�\Qd�9�WF����{�(�7����Ru�[ѣ◪:��~�kݹ ${�BO�:]M1�R$��C	M��b¶g0���n(4y2,38O8��SV�l����PY��7o:}�F�1n�鎞���3q�}MA�uO  �JCB^`,�vGLwHSP�`x^8��#iKF���pv���G�������_z�7��@Jf�חk�t�F�[��7����w��i�g�d�H��B�{��*�n���Zɿ��� �H�
pD�5�N�O�t�QM�<[�3o��}q'}������>H"�D�p�C�9<�~jmŝy�f��y�$ �� �K4졳�.��W�0�>�a��SV` ��o�%,;;c������4V�2�k
��-���SiQ4T����"�mÝ�Mhq�!"�R/�V�gN�Vȋ3o�m��qǉ��QAFkP��d�)⇏���
��'�8�Q��m�z��És63U��_���;�i��҇�a�" "f8�ڠ��=�A1� �_k���zy	�o�7�{����?�m�O.�A�+FŀX̪�T�W_i卋8W��ll 0"�ѐY�fXI��L�罃!R^����Pg�H��yȢ(_��g���G;�Hx�匆6q�+5�)B��Jz.i�̤D�',��qg��� �*�I�T�?^�k](ThoTA'U�MH��u�����\,QT.?[g��XN�݄�����!�	/5�.�93�<�
 r,cſzh���'�$&�\��$75�j �l.muţ�_�?��>VpY�F�U��oP��a�"nʛ)��9�W�6�"���f�q�ݜ�H�׈R�[^;/W��2"|�\*�kQ���0��������Y_���g?�J䆈8<oϺc>�82�@�DBe�y�y�����7�>b�hp{:Iq�X�GV������5�'b�o�GB5�d$^�G!?q���J7�p�f�I�h���C�t4����M���T�݈��-2�3i�}��ܻ���&���e���0�v���E��o�-��)7�u�֤ �r�ϥڛ����u�d���;}��Z�/r�^��rr�e���Kӧ��
�Gϒ��/�ּ�q�xD�r���K���M5��ʆxyT�l�Ug	���'����Љ'���FU{A�YxJ� ��G��;���u��2k  ��BX=x���ҕ �����#T��r�p�Z6��]�Rj$l����R4=���_&��l4^6����3��2�n� �(sKs�骐�а��@_��H���4�;����y�'������ ����'�����G���24��T8P!۳����f�(2��ZN��Ėj�����E\���n1���,_ÇW�P�N��aӯW�DfË�Z�S0Ѧ�U`��b���?Y�kkt}�&�x�Ѫ����-���
}������z�T ���sŎ��r���?�����ԬՊ%r�ӽ3 �"7݃~�+�}r^�":	E����ְ�x�-�u��	��dA�kR����4s3*k*9^��۱=�CD�U`;0Qm�շ�C��<�s�Q�3e��Ʌ��
;���+��+��\��P���Y�
f��+b&4<�*��'UKyUA�8o�o��hf���H����E�]�/��<�LT�]���/�Iyo�IHyTƁ_�,��mU;_�M �'�`�6�P����x�H��~��@��ވ�ݲ�rl��[ڟe;�_���|��8!���[��o�,��jo4��テ����M"Q��6��yjl�6�zl.��R�Eh|�4��eH�u�PHb^���Y�LF)��a�/K&a���)�x1� p=+�,0[]5t����%(�<|dIDS#��&�+���P��@����e�OY��X�!i���*�)�W�y�u��|����^��{��.lw��'��,1�T���q�_�I�WTJ��
����{��$���թMǜ�>c���d��bA��W�l���S�N�?�ȳs8q���2���\l}�bi;p,x֖�%sz��θ9Ny�a�}�8�B���ZQ�7�����Ai���f�$��bK4�1#o�V4�\"�?e��L�V�O|��2�.z�s�'˜���t㻟v?��6 ��D���!C���{HP��y߼#��Y�*#�'�*�Jk&`�]�$|5K=�U��@�ɋ��iU��,=��̱qJe��4$����\���&�H�wD1wCiF���|���O:?�<Z')��-Qz��.�V[%�k��0�-���T]�x\yb��&U=�E`K�3��)E�(|V���@��v&��[_Bf�9��f�0ɪ��z��g�e)�Ғ�nÊ=�	@�V��nQ�h=_x+0p(K�I���&��;)���yI�1��%c�]*	 ʏ���24�����O�R�]�E$Ä�m�5+~�D, %|F��'���B�`��"Ɗ
��)�&�P���2����BN�W�i�c��&X$z��h������Ag�����4�������M��g����z��@�pm$b|�@�a	���~ۃ��6%�:B�ʓ�}_~�0o�wh�·?�2D]��ՕvO~��B�	�N~�O�$��#婛y�C��̻��V��/�GK�~]b��|!NE�\����w����|H�y(�I+P�gjcG�â��Rx-^��M[$
�(�#߱&�(�����
A��"-=��4Q�v��Vtur'�H�$?� �P�j����w�MſnȎ'��t�E���D�(3��>l@�T��Kmb��ȭD�2�ޙ�19�DO���)����(V��J~U��	]���J��&�-�J��KƲ|��|Y�Ԩ�W�Y�E{7�}�ɥ��D*�'gb'�ק��WXD"g�[n��,�����K����J9���)��{�b�cΣ�PH���&x�:����M�:�|�q��Dyv�;~��9��a�:��y,mR7}�Y���ׂ�|��Gp3EJY��&2ƪ��Rp}3�OT�f�3��֐��?[�,z��ׄ�,T�+؊=��[���T;�\�iկ��sx%���Ol_��/�yku��,���	�t��RxC����_���&p���^jQ�7Yj��8B��0.����{|8�1��рo�yWOթ��=��vc��q�
��������xFQ�湍��]�,)��	��iS��N ���/������_>K�~J�y-�M0�85�QU���c<��w�F����u���w�od'tA���W�څL.]W��������L�T);d����|�(I?]ڌ��3e}k�/�kVY��:�pF%\�b��F'*&N�	�=��C���s���^���q���^���EP�4c��f����CE�<)���a�é�`ԩ;�!�&o��<_���Jñ)�C\9��e�0�����qȐ6�K��M�	��>��[����~j ���saB#"��0�o��Mj:Dr���yq��O�D��ՙ�H�̍��{��{�^�����$�f}ޒ<�@�3>b��ܩFX���7G�z�F��B`�������mH!���]�C?BsWL���VNZ͘�nS�2K�4�9�P��u��q����d$KD�f���,�t{�l�{Qow�Y��L�c�P�1�ڭ��w�fUDB@����/�w\�i7*�ࡸD��ۉ2�*���O��M8Q�ˆ͢:_��s�XN��O��1p�\qo 2������E���on.N���n�?�cSC���|c���ѵ~&-rm��Vg��yN_;����Cʼ[�r��(Ё�*k���v�U�ǊΊ�e�8��۝b�*��v�qp�:5�c�ٙ��WR�-�#��N]�t�vgi=��c�O�2�j_a��m��cx�� �lK���?M��2�ޱ^���	mo��1�Z��B�E����L�t��@ex(R�x?'�}hOX����:��Oi��ÈcW*Ciʛݻ�&d�_�ty�ը�	�����Y��VwSrO��R�mk���,�fs4�%vA8���� �[-�'4���J��_$MqF;��:H�Ȅx��0)7����0<]>G�!qD�z%�59���l/�e�T��&�s��3<��� ��j��s^�p$pzh�D2(��4�� �$�Z�[ǠY�]	�H�Hj�2�n�B0���8�N�� �VGT�<�"��a� H%���us9)�y��V��S���H�q���l���)�nG�T��Mc�Q��0V*E���×�7Ev}�p��rn.�����C�ɇXU�0�P��(λ�딅8q(B�m~/���Γ���Z�n ɱ�e���)�@� P�`��A;Ll~�����!�w�d�>gZ���'go��Q�����?8y)D~���Eȅ�S�/,	+�C�p�A@���`S��a8?���|X+�L'7�B`�qڶ�N����u����_�L��x+4*>[�E���Űl��d�23G���F��,��䈅����~��T��~�s=�;Q�dq*����,�!��10��5��ܮhq��󛟬=�Q&W����P�=�l��@}��&�5\�_4���<K3��fL)R}�?{%�Ev�lڱ^8�Am�:<t�L�8�1��Ж4�44�|]d:�!�خ�\ �����{���QN���ﯺ�>$[-�.�a<��bj�썯��?�~���2g�٣�-�!�tߋ�Lϋލ�����-k��ṙ��s�@!��x��ȹH�d���t�A��yeu0�t�e]�tEJ�0�kӌ�)�AK�J*�ǥ��P�V���?*o�&O�fL90�]�����uyt�̮k�s$ïhT��6ه��aW����J�*���띞`Z�KN��6\��R)����?���y��J�[�:d�X.�w�����\`G�c9�:���_���N���d�RU�!.��el�&H�40�zS�uzZ,�Ĺo����T>R�-U%I�BT���[���q�p3A�*~���D5!Fp���H���t�Im{����찹Й,��1��};���e,��t!��M��롭0u���v��SL Ye���r�JAI:�����!��;��P�D���m��a�U�Y��C0_ �56�o1�a�G��f47Z�R������;Qz]��������f^�B�(>%�0����6XY���"�0�e��H�?�2*\�䘔�A����9o�������.C�D4�0B-�yxE>�N"�~��ᗪ�W�d�Rí�C�q�����c,��i�
���aEA���Z2M�nK
M��07�J�-�B�Jf9H�4R�?[��r �z��햼�FO}N��N/-�X}�M-�`H�6���w9V�E�\ >�ޘ��T�������&����Eγ-�E!�C�k�ߌ�ꌛ
���;yq����9R��r��R�+�M���&LR7S���=2�1�U�i:����!Cp�ғ���y�iwA7����f��AY���|�Ja4��H���C��<Q�e���uH�����N�!(�Tr�-�8):��Oq�Y�̉����s���e�1��d�彎��ڊ[���l���>�z*ux�&[Qm�A��J� ��mąX�NL�Z�������=HC�oGD�7u;9ٲp�4�F��aHO8@� �[��$$T��N�j�G��8�����/K�U!�3��__�Ai���5�/ki��e��3qk�8r�X<0!G�{ه�n<sנ�"�"�&tt9Rw��>���>Kσ�M�������C�� 3U8�u"���XG���n�+�2���#N�tC7�'���п<s$�=���X&(��~Sw<2
�����]�f����.�ۨ����.A����h�8YI'q�Z��"�ܾ�����%��!m
U�������.�>�'�Y�r�d��өl��1_m��<�H������m��U����=}%.�#G2�����W�����V"E��rz:D�I���R�%�@zߴ����(T'4T)�0�P�1��і5��V�R4Z�H*�	�O���:���8�?��_'��G*}�̯�a�t�Q�b{�Ų_9`�[��q�q)=�K%@}��ĺ�����@}�a/IC����E��B�B����^��Qrl=3�c<�Z,�7Ae�u��7X$�X�6��SqH�}��.L�<�]~�뵦3�o�ז�v�
��ڛ�O�T�<�
0ꗮh�%��;+g���Ǫ��E�P�޴��!���H��myl��D7^a�t;N���s��W�M�T�{M�7+͉Fnt�H�t%���!!\���F�N���Bh9��te�4鼕ZX���aEș�ҫ$o*Ū����DVYF-C8�hVS�e&��韻=!"?� ��H4Z� >;����i�ig���g�薏ł���w>��O���s'��l�O�x�튄���6!ˎ�J�m��Ċ[��g�'���V!���)460!�C��A�bT�G.�L�`��Ht�!E���yfw�K[��Fpf���Mhh��Z�[ے�wlͭ���T5T�ۆ(
�X�1�M�q�F�}wB*+�K�[V|JSP^/���,�f.19T��>��`�*�:����"�|�	."��R"\�L�XvXв��/��G��o[6������jF��z /�k�kf���!^�S���5;K�|��B�'��R|����������ԉLh*�.�������ݚ�l�X��֛�� ]E������)�U��ju�͐6bȿ�)�^!�x��Ia�p��u�K��@9���i��c�1� 6n*ʐ~�Z,$x�?�UB�w/{(bP���%��I�T�iV���5fMM"��+XI7^I .��Z�5U��om��x��{~�4�(�W2PLq~	�ڋ���N�h2�.�7�����`�ٝ{9���(}��;�
��"����|r�`՘�3/M�4«�]S8��^�#$wM\�Ó*��'��4���F�P��X�;B-�hж4L�9�?/�#
U΄~*R'�pUq4�ֶ�\}�2���Ŭ�w�ot���׀�������NbHj�f�l�G�x��Kgqt���(@]s����S �7T"��R��2�����c��E���Ęi�.��!qڜ;�J����:��ھ  �Ֆ`_i���ת4[����1���ϓm5�"]�5\;^�v�9Sơ���ø�}����7l����_�7��"���?3o�s��6is��k�6�	���,�P�����!���0�d򡂘��Q$��p^��|g']�/���;�Wv��Y��htt�<U�pCbz6f������0H�@܎�K݄G*����#X.���;��dV��d2��"~�-���Id�o�Huzfb�y�O�7��=+��p�1��Q�L���D5�)��a#Q����>%12��%��e���ـ�J�n2���@�p�u
�� �������>Y]K%���q�T����*�9��\�/B���eb�K���8Q�=���\j2Po	�ὢ����0�mߥ�8�{���!�����pUx�8� �Yu ��Zn�ڲ=�~�C�~�|| {Tp���oQ�fc��,�o�F�<�R+|���j
�R�"�(.]���r�bm����W�B��i�b�8�Z����O���[���J� �_bΦ���*��eRU�&8⠛���&ݗ�8w�Cd@!�"*.���d���I䆁��x�I������d�.�����
>�uu�����2��C����lcym޸�mrG���$OnB
��$��`�|�������E%C���Tb�)� �N�.���v���_`h�"J���F4� Q]R'�����
/W���;&���~*�� !�:�XOZM�`�$��?��tH�;oZ��&�Ӽ�������*��u�� �a���(m�1ݚ�q���w���\T�@��$�������u���x`�����"�������C�?DiݩF����fyy9��]��Z�}�T�鬿ͣ����b��� T ��Ľ�WܚZt?��N��:ㄨ<�qz�Қ>�;T%� �&Z���	^�a�Qi��,�"/���Zi�����>pv<��%I�k�s�ԣ�|~fwlM���bd �Dr�.H��W��� f}�4�['\��G ��.6Hp��Q����oA��C����(��52�U�N-�\�����#�8���v�r��S�Q�.g�E3k��_@�W��u���/~=��ƀJ��J�.2�v*C���`�a�擋0�uJ>ԕF@v�c&]�Nx�<�@�Fx�㦂K/_���f�'\9�Z27�VsyH���6�S�(��S}�@��/\M��.���iM}$J��Oc��w���.����,�2p��������ݵ���Z�y�R�:��?wz*�/��3�k�F�����i$-6�Ť~�5I������X�
8�z��D"X/(���8�(�0�-L6������^��ߌ!e�ښ�&�/U>L���X�R���ف�Xۘ��rz����b���)Uu�g�1���jc��5�q>�N`�U�	�-���6p!�1��8Z�t�5���M��:��l��I{V8�؛�?���Tjb��'��E?����M����U����Sӯ)x��!�y��l-	ꂎ���Hh�<[�j�3c��ou%�َO�3�����u�A�j�RF�%���lR2���d�
���7yL3]�<�2�����jڅ2�&F�}L��l�p�+�+@�E�t2a�Bn�]qdhj�@D!9�������� \�D���Ė�R���c߈�Ou���j�vt���q�Q����.m+ڹ����&����xɁ�Z�n�x���Y�C�	E���,�s@͈��$��0 t��3����$��v�YS'p��9�.�1�gtGr$3:�#�{~���i�>=�*�5�$h��`��8��r3�$d�}��Y�Fab�K�fh�чψ�<�3��p�U�:�)�N��hbDp<g�{y*�T��A�ܨoC��Ǎ��+����pN�a<�����8ć��q���X�reЃJQ@��oƨ�d2kI�qؠ�.�
4�&�F˗�saBb|�;9اY��N�y��D�{�5ň���g觰��y�TR�b�ɆWd獲���4�Wy���V}�����j}�]2�� \`�'�T_h��#���m'�:"�Ѻ��-�LJ�*՞�8���{���)i���?`�I�'�qR�J�7�	L��п$y�'=l�v6�ߋ��r(�k	n��*��D�Ц��=PܿqݪG@�u,��ϊ�7Z�3E~�-��x���M�й��n����:���w�y�i\ӽ�0��Z��̠Z���V����S�_L�I������i�k�6�~�uS
��M��zQ!�$r}��B�'(	�`�Y��%��&�䔗�:�]��� ���%z��y^-���y�@Q+a���~��۝�WǬX�Z�kE��,�� L$k���F�����Ӟす�JLMe�U7V��d&�pN��r�c�z7Q^<rr쥽�;d���"T�������j�(�S��Z����c��8x�����mMo�/Г����Zj*�ء��M9���u8<ϻ����o�d6@�Nb/�=&�K�5��N�**Rb0���1�����[��n@��i�y���~@t��K�c3	���&\��z��� vj�J\O�	K�8�Sr��جt.-�$ĆN1pPy�u��iw���H��&.Q?�j�|�����`�� �H�y Ԡ(�Y�c�%����GN0���5n��-,��!����*�+E�QtU_r��%��y��ƌ����=B*��W�nϕ��5�����c�j!�aW�!�(�X�a��m˿�Qڨ+�� �����#�.�Q��3�2q��i�/���}�oH��"ڜ�^��x@/ ��7/\XW�f�d�H	����0α�v8]�to��z�A�i(�f�'�����#1��<��Z�n��lO�Ʃ�����s8GM�v<�\p�D�l�814Ͱo��,E.jR�z^�XK�:(�;�#�[;���0�����h�w��Ұ���\<o�]���&��U���#�Q�֣�	�����D�,,郬�o��ә ���7����Ӣ��ߝv����%��l��E��+��NE��/<����L�'�~��S���@Yȃ"q�����9�a~Z�蟓`<\,W,&��d�Z���7�>���Ot	햾�A
���CCC�'�Ua�W�R�l/�3XP����A�ד���v-���A���P@���8zػ@|���`��q�#��J��=�,q(�+��؊�t��M!]�A��r�sC�o�͛���n�9ҳq�^�y`�<\c�+�"���ġ�TG�A���k��{m��R�ѥ.��r�Soj�,K=%?/�t�Mm�9���xAL<Uj[��2�E���Iz�+g�CO��{.${�up	+�u~A����y){�<l}�2�R�?sT�ͼ�����SE��Pýt�?�z8m�:�Q�n��D�(��f�z�ȡ�!t�a�R̚lƟ��+�5Rh�fBN,{Q�0���>ݬ?��
]�_�*D��������A/F:�L�}��F����hO�j	�_ν�&o��
�q�z�t���-igMM��iSV{����x���G#�2A-yd��7�M��G���A��->wB+l$54�c��a�n��w˚˅�g��ynnW�эz�Y!	�+z�".��	аRO��~8��i����TY�v�_b�jV�X�X8��ukG�9]^,�z��pN��O��J��Q��s!�#�1���Ǵ����b���!��MJÆ�g�_z"<}yg_L�L�q[��ٴ�4�I���>���$�LyXdL���<"S���p�ھ�U8ِ����fWË�|�I�T#zF@5+�m�pN[ǉd�a�:1R�;-H ;=IW��-o��u��-��,��D����J�@��S�P��x#I{��v�1��&���(�r��g��k�mh�l��R��7�.��@��2�
�by$��ZL�ә5-?0o��V1��@����+6��a
��-TZS�_���֌��5`
�"�P�A��9��e�;�������*nw?�vH���p0sܾ�Ho�s��㌿� �w5������J��/47ۑ��e�M@|����}�A�B/�@�bhe��j���a
�_1w	y��kr'�\TN!|ݸPh$�LZUB��8�h3��[����ZLDښ�uΤ��e��c�I�!+��(Y�qL�}=k@:��!_%�/ӌږFMc�I��^��0ފL���I����	N����xF�W��}O�@U�� ��Y&p���Mᦿ~"ƫ�p�A�c�ED�/zlTj��\#��< �X���XS��N�[�����ȸ�}H�����5OBi6},��U�t�DE�����6����ۇ�1���e*�z������>�Ƞ��؎��,c�1�=<4
�j:�;ˀTי�L0ۆ�8�@�Y�����v�D�@�����:��r��B��mg��7�Xؕ��:�zx�A�J;��߿�B��B���W���T�fQ"\w��eM[��Mor`Uϔ�3��=NZp��C۾Kۆ����.�L��F:��O]���_R���-k~*��L�m�5��;`�߀���}�38�KC,ܖ�:\��J�A�J�֞�>�(����,A���@���n$�|@egPMr�>;t/�b1��m�`oN�"R���ڪӢ=;I�����1-D�hA�������,�As�b]I?�~��멎�"�	^� ����Eu����j4�ڶ��~`��56�P��'�2�S_���Ӕ�"�>>�<���\`L���g�z���)�Mf.�l���Yu5~�h�����@�/'}���f�$^A�~N�T���0=D��$�>�1��W7���S'R'���#:a]/c��7W�����Q)��>0��!짞�g`�C*7������k�1����{�����	�*�
D�L�/Ƒ��g����G&��D�J����[*�P�	o/Mŗ�㰘�]��4sҿ�8-�Gk��U��^�/�Gi�@�?1j�k"�Ӯ����_�Y�뉍 ��o7�	�N�g���]��*�kH[D�=��0|F@.Aϯ��723(W���;5�بY��⣛k��5����"�#a/:2��uT��MB\���]G���<�T��𩫗�Lu�2L=Y��|����+ȯJ��bg�g��.vQ7t��CwA@��&_?bF3�z�i�˛� xEjG�v���ep��m��1�l���db�'gc�1��'!��v4�����C��+ĩ�9�p�!<�i<�����T=݀�����7��W��ϵ�D�o��K庒��t�$��Ѭ���2?�x�Q�'�5n�ķ�caP2�^���I���<Uw������=`R�ɕj�9�V��L�z;ل��-����.�i(d2���4��R�Z�'��������mq��2�C'���
�v�tOQoNMKޢ\#β��D8�lcْw޹d��<LT����+-��(�W�I�<��>`� �L��I�1�ϛ��x3Jô����8� �f��x��ՠ{��~̅Zր�C�+��5-U��^Jټ��1���a��v{�5'��%W-v�;{�I�8J;�� �HĮjޞr݌�+�NyM���J��J�q��7�@-p�J5�mB�/(��L�p ��{��Q��1�J��ԷC_ʭr��X�'�ʦ��f�W�����p���������+4m�l�c�/��.w� k7���o���$�Z�AT��5����r�IPا�K�(^j_r)�S"�����F1�=bc%���ߙ,C����w��WL��T
�zP-Pg��F1��"s�/�P ��3����%_�]!�7�;���L�NK
ĝ��wd�I#���sw0��o�V�6Jg��l	��oS�%t����m��ϲU��0�.�nC�J�3�{�w3v6ڷyw{�|�jV�b�vX��|	�	H�|��i3�L7)�*��/B�AqY+�����w�޼}��`E��~E�T��q�� �cf[�k]�Y���3S3�Ra���@��E�@�{;?on����IV)�BSH�$�&P�����/�$�����ʖUt�[�g�F�|��l��0�b8ڻï�eh�d�4>\Խ��[��>���v"�#�6.�1��Rk�?KM��a :�и�6�t���@��=��I,Ս(_go�$O� 7��\i�^)��\��=!�Y*d7��n"0�[6�' ��)�����x��DAj`�^E�9��e�=��{�$^ ���%�H����ᜤ��^�R�n��.�H��XC���{��v!�ǃ��\�0k������Igsd����*o���F�B;]@�t|&}��d��`��l�_��#�G�T�s��t2���W���c�~��3%k����F���U�X�i1}�.�����va�][N�5�ȕ�s�a�h���%H�*����Ez���ۉ��|p�+�xTg��L�Z�s�Or�|�S�	H��M6��>K�2�;��-Jū
5J�M^r\���Q�,)��>B��.�����3BU,ړ�vu�kh� ����)ƧtUE��$�l#� �d�&��E�$�_MP-e��g��~�r��c 2tV�]*8!FM���vǩȟ\ ��Q�����)��E�]��Kz�L<�g�!�˚Y5|�/H*��T�S��_�8���y��T�[���N���4	=���zj�ϵ_��+�1��K��'l!��M%�L�iN��" s�����F��n��WB��� ZD`J�I7YT���||��3k/��e�&����~�9��r��}�&z����?�D�_U�P�E�m�E�A��E��nt��;�N�����N0����X����vM-Rَ\B#x��"�P�Kb��X]�#��(C~�1]�3�mB����b�y�.*��n�T�q�_f�[�#Dѓ�l�KN�/��cV=��-ǁP�Ϯ^[�8��ҡ��G~��F����?��o�*h����v{�Q��l���C�:�ݶD�d�l�oթ��e�^'>|(�&�x|t״��W��F�:�N�x$ם*
_���31�	����4���}+85Z�,�q���%�8L��?�H�̃1?�&4�pYX�^p�Ш��6gw��̻�q%���=���q��1�A�{,��E�+���Ca�M�?��{����ؕ�v�	P�I���M�i������y,>��5��b҈��l�����O"�\V[����{w�����t@R�:Ոl��#Gz���px�o|�������A>���3^��O`�q�e�_�Sϯ�C��9O�Q|�D�=\�Xy"����3v�t�~��𤰱F�U�ݯ%O4��N�c\��q���ԂbZ�lQ	=loB҈	2*vV�
��,,��j%1Ku���t�j/�	ΥڎI�H=9����u�����M�&g���m?�"��0Hъ����G�܃Έ%�
��ά׮�� J��(-cL��$��̀�D5�0DA��CE��c�N&_������ޗ>�bf~������~#WЄI������q�˺H
H�&R�й�E)���3�mD�i��a@�Ӑ\Dz�S�{P�����܅r�|�}�u�/C�H� G_��l�J^����W$�\5����5/Y;$<��
 /qN���9г�Y ��s��np�j�V��.u�Q�t�d0�CW�W��&����Jv����C�,=�3'�|����$Rl{���X��S�'���S+�dt*c���(IB����ҏ��54 ��U�\y����@ԉ��]SZ�}�'��$�iO`)u@�ʄo��ƾ��9��2s_Wy�U��:��@����UR��O�gLɚG~�x̖�̯x��<<7�\i�	�u��~E��>�d��<r9���mo\Aد�	�'{@Q	�lJ�~�������1�����|Р^���'��`�m�ӆ�v�Vط?_�ub�(�NkCy�;�'���p����N��<y�EW4�9t�����}����ɗ�=���v��8�b�j~ټ	J�7����<{���m�����ư�!���-��ӓA��O��IMaj�Yab��� Ϟ�*��\�=N�E)k�ȟ8s��臠�(怞��v���{�5���It%�a}
Qn�]ck?>O[��:Ź�(]wa��{f3������#�]?��j��Ep�w���������h���jX	�3�SːH��¡�g($<Oes{�-�L:6l�* 54m��f��RҢښ���8u�����-� �<�/Zy#�`�e�蛕t=$P��I\��Z��E������	��� �rZ��q)m�1�ΐ��7�s�u��dg@¤�|QaI��O���E9 Q�Q�v\?�$���z���0Z�	���s��T{����UDkt8�k�9�`�=�q��YxuPj֔��Jׇ2{0��z]��߁�0�։��cP���y�4d�C �`�R>̟�s�k!O�B�gW��ca���'�<r��<&4#í����}(ѹ���b�4hE��)���t�[1:b�$�F)X�T:E����04ۦ�ƌ�MS-(�l���|@����GXT�~��,�m���w�z�E��dҸ+j�:���f[��&x��G��j���uy���ֳ&�y}w`z�ۨJp��Ef���sA2��u$gAaTs���F�\�p,���uMT�[m-��Bf?��-	5��f�be���WӁ� '��P�F�!�d��Fk������)F�v1!$k�̾���l��e;��5�*<�3�r�C,�Z-�iM�.'�0���˄��6+�7Q�����,+����^7��pR)�l���1�� db/��M�ċ�]zr�P��ʁ+;9�f��]���g��K�me�X%Q�T2=�B&2���O?��ā=k�<�~A�v���-Uj�4a�\r>a�<�����v���򿅐=չdF����D ��	[M�3{v.��4D�o��=y}�W�ގ��>��� ��\}�����KY@్%M�>�u���Ҕ8�s+a��G�o
�Uc%i�ٺu{Q)���W+�rV���\�:��Y%%���!���"���uv�^D��#���S�;R�����s���,F�ɨ���m��qI�$�v���S���u2<`l��R Bt߻��b]���̞dn�N���A���`J�42ŀ��|!xj����C���y�]�6�!�p�a�
|��=h�[���Z�ʩ{#��T�s��.G������t�v�b��(+\�O���%J:P�̓���e�:.������Y�����rug��{���^�7M��������/��3@t.��[&�,��u�v���9 �x�5��������+���_�?=l�ݙ��9����3�qW�$��{��!��pD�V��#�A��^9~T�������Ǻ�j"k�$�8�g-�$�+q�kg��2"Q�����O�|�	�F ����!���KM��@�g��T��i.��?�Q��i�P�&�u�|%k�0{�Z;���Ñ,�����sr�" u���3c*~gצ9j/O�4~n�/�̰r_�*�
��&S�q `�6�?�x�
c>�@�������E[��v�쪮0l���ڦ��<l���Ѹo"7OnQ/v��X%��(�#>�c� �d>z���0Uټ�y�\�]����]+�F��i�\@�8"�b���7�uڤ �}����Y߂�� ��0p�Ο��J���tA�B����I���xZO���o�u��!�b,��5D��O#��&x�q ����u���h�@�[�"�XT�g��$B{�X�yE<��7cGl's�O%�a�!7��0�#YK�&�eL,�6��l�mG���1]o!ڦ�FX������j� �R�VD`���<z�s�ؘ�f2���X(�0�+g�ޟ����Zz��p���B��.�?����lˬ�z�n={�)��~��Pr�q��f�fdݘ�� 25x�[�̠m�Uk�{�{!91o�c?��V��a&�~�i?�c F?�z�aƤ?����a�r��+?�O���Ͻr�8#��9��oP8vΐXJ�k[�k�&��MtE]��k��:�����82����?�K<&NI��#�5\xe�V,$��Tك�됨�nC�ݷ}9��+��q�}m�i�zy^@o�΅YJ;:�!G/�����z��͞Ҋ�c�ϔU�Сy��b]��fD��c����t~� d�	l���Z���|�Z���̈́��q�� �Ϊk2RmV��ۆ�A�C���=���`"EQ�~�Ԋ�v����>a�o�B?PV<��<����7c�Vq�3�
��G� �
 �p���o8����nN�'�ָ\������ºD�'=;#��zj�O��PJC��z+>!XU�yG��7����UY�����t}wX��QO��wWė�*5#ˈX��3�v����?���W�ƹ*�r�*x>��RJ�펋���O���I�%@3%��gcS�YF,���?==g�Dʤ�4�[ԢP]��{j�"��l�Y"��+����|{7�r�8XQ�I�aӵ�"{Q�R`ҷV��W���P��Q�a��``�����[gL`����^~Ȋ#��A2���c}I!�Yp�#����c�4�i֜7��n1B����XB`�;���T���0�)�qS�vC7�CZ������&D/s|�l�/\�����%F�͔��������B�1:���	�昘�����7���V��Ht[G��r<�#e�p�Є�#�\�讽Q{�<Y>KC�����]��'��2;3z]hZ=���)��И��i�Q|.N��/�����8ү'Ak6KV��XGjC���
0��v���O�1�sWH�p�\�-����`��U�u�wz��?�~t^��-��驅T?�=#��9�U*�U�B����dM�@kji`���t�4ޥ	x�^�?�]'�'���2���b�Ȅ�`Y�O1N�&7��9�g��]���/�bc��9��+X����c���K��0w�d.�"���{N���.�=�QT.�U�M�����sȞ�"�2�N��M���a�p�@����1�)bD+�(b�ޡj���<G����� �ÀǇ�99^��B*���:wQ��~��i���52���(���WMOd�9X���v�
�vk~���#�O�������k�<PV���I❿���hP������w�n8^e�������-�X	�no�����9R�:���!J%j��}ob`�+zoL�Pc*�Ҳ��GN$s � 0�7:���4 ��T��X���F���� oX5�5�'�	�'d����-棗C��P���/��U_۽>��̕�zt	~��(�p���N�W�Q�h=Oűܲ>�Zx��5�!�H�^�"z@�ᆢ3�Z;Z����)G�;�l��}�!Y
Ά�.���K���Q?ڟB@o�1D���r|ڭ�.�� ��`��%}�"��ۋ>E��R�j�%5va�O	B`v��:����Z2\p�hK_�{f�e��T�v�^���B|k'C�~��4N�$��#�&r�
�!���"����$>߸���kk�V'���|62�šTP3q5��BYWqM���1�/h,���X6��3�h2��+<��1�D�u�}3���`jȗ1U��zN����\q�g��e��ePD�8��F{��%d�rCB��G]�_�ѹy#�<$���<cz�߆*�mp�3N��V�P�Ĺޖ�e�3<�زB!�'�B_N�A��.-�F�'�Wƹ����l��{��xj�K�la�Dq����v�U<�n7�(,����Q�OB��BO�kVOB�#p5^O|�{��O|S�@i��i؝p�pmj	����Q@Bt:y��
��c�L�{��5Q�������h������9��y���؀��>�0X���u�Q�p�?���+��TEQq����,�o��C}Fפ����d4�־20e�����9Ο����n�A����Zɭ�LD��tG��.�+8v��T�O��VW�{����T<#<E�^r���E �2]�������0��5�AJ�N�z��4$�gA�[���u�o�c"p����<���,�R�H���o������e�xൗ�Fq��d4����5���U�F�zm���n��3#�̏k&C���A*3'pX���d໋*Ѩ/1��:�&��W����`���Z��-*��?�)
Qw�aΟ�;�kT�R�1�`��\�g�����!�ف��WH��R�5@�,�� ��tn�@$ ��ĠB|7f�y�z�y�6�Ƞ���Z�fp���z��/���ԁ�Jb�P-O�x��'�K���MD�'Y0��@/Q҃�[�z��	�Ǉ�Y] ]��M�N&��6OٞET�6�v����ƽ�T�k���\c�N`�{�WJb�R�ӌ
̸�����C��mg8��U�3��K�VlnO������V>�r�� ��fF�s����gu���B����i銁���8nCnk�k�W�*3WȾ�����^wsj�0���Qݨ$1
�ȍh�2Șg�1:U�6�'3�4�e}�PB4�'/U�u���O<��4�M�0�ut�����!dt�162�9]�+�:K�b
p��"I~ň~+�T��N�N: ��)��Ff��E�Z�( ��bώ~+��+��t�Ĩu�L=�p�"8'�J��00�x�c�����e���=�ۊC�R
�P�wSLw(���
�{>���\a֟�7�/���Γ�Y����U5l�����L����?�T�S\���|-ĎF�S۟�3�sn]�.�(�E3A��$�"�ȧ��qi<�L@�YX�ʤUI��nl��֝�t���w�J\xi��Ɩ��%#S{��͊4ۢ� ��:����C�z���=,B�q/T�t�z&��]&�r�.��Σ��rR?��"Ow��I��2��9��x���;ĝ!/��.s�X�h�e�����X�x[`�%�9�B�%S1��r�v���?�U��I��%��sԪ�[�N�F�xWC����aY7Ƙg wlz�￑$�Г �R!n�zyR���I|�	�3�$Tj�u90��FƊ�5=\q)cm3�%�Ar���ۢM=7�d�'��W�f׎&$K����%v7z�����Qg�g�[G� K�BP��0x�\�
;�2g�� <*!���;�����ђO��T@j�)�*��9�ճyj���hVT�h�18��v_�wv�*x8a~x��[!��0�U0������V�d4E�~��6ڜ�zr_F�8SM�N���h��ȭ�aD3�#�������8	Rߝ�b
�����Cn~�0�_%���}e"q��n�]�ƽ��ȑgeQB$O�,R�U��!�]�<���!ʖ�����O<ҩ	��9�%�i��ko���Et��彻�I��2�5��	b�Yq��+G��a�K����kbj�(�K	W����m��%������2�������
NܺE	ДN�o9�!Z�owj������r�l�Ķ��'sy��]�C'Y[��ʺo���!L�ʑ���4xi:����X����`=��;#�FbP*��2�P�A_�+pL�~���& �!��'&	㜘A��#���TOs��M7��.ȭ�M)ZM]q+�4��[]�y��2��(р�Ҁ}��C�\{���?b2�3�!LֆW�9M��=��t�0�d���_������ZQ|�ϴ���*�m��:7~f�n�W �,c8��$RԂ];�k�)"~����=�{Ʋi���A
����11�k����E]��w�hJ��L5㏿��j���Pn�a��/�����=�6���(.n���0*Ez4�r5��&a>�jkm�|avcD)bVHFꢬ�"���+�ލ��`f5���A
6f
�!���ܪ� o�?�җ���ۗӅd�7�]yX]�7��i;�p�ߨ����dhه.�����I���=ġJ�|Y�k���Q�	y��C�)���*�Y6�:�ƃ����{���~$��W�f� ������܉�i~��#�_�/��м��z��;WC#q����[�� M�����)^�������L�-��?���/!�I� ^�T�ݙ��3d�9*�(����K��{�y�&���)8Va��1 ӣ�z��w�>���q�}=D�co�^�ՑM���@轒� {?V%���5��.���/�-ZH�����+\���e��'�f���""�`u;= 0&�CΞ95�!���
�M̤���_�x�nY��H�w��(���"=���/x�Ty(��C�ʹ�����:c5�of҅n��SufƔ-�7�&,{��lse`s�et���⊎)�()0��f��R>}Q��}�=E�j!�4�dj�/�}$Hⅇ��z����2x���m��S��9���F�N��hDq�X�L"�|���)@��^��'�0=>e����t�^�����Ç^��5*7�X����8�"�L<�>kN^��_Lx6ئ_�gv��5�<�Nr\cIlC�=��
����)�
���+ו%/�ʂ�O�(@���YU���G׳���4��o)ܵ]�{��ԥ�סJ[#�����̖}C�M�&���zHFe�ԊuDQ�O4J�5&^��tQ��s���7�b+�'~=�3�����x���X)� [���c���v_�9�|w�z����A:��Oiu��=7Ѭ��#�p�ڱ)��V/i��
��_d���9��Y��I�J������j͹Y�¿J2����k]z�Ň���36�[Jg��������a���=/4�v�`#��U�~�w���jb�!��"UU�>�)_ߒ�@=�J�z����\1\�p�t)���P@:Z*�^F�뻧#NB�4�~FBc#q��i'��R�I<������=���&�E��X��?��%+�xK50׊-�ܡ.�¯A�b���<�V&>�WR�q����g�Y�?Eqڦћ/|p�������st���sBTH+���:��+/���i��K�D���0n��'�PX�ߨ��B��t��6�>?;j}/����[���bZ
I�#JP�.�oOD!p��H�&���ڛzk��$�e~�4���}�Y���e�nV�/E���r������a)\�W��������wQ��Vڞ"��O~xq��zE��g�o�Ќ��9�k쫣m���ɻ;QPDJ̥w��u���s
�R�E򨬬0��Գ�`(؎:���	��/��Ja�V�ȵ����'������Z_I�dԠZ�xg�ֺ6zeه�@��/�ϩK-����SF�5@�Fxv��hZ�	�w�g��r�w��pT�=�	�X�^�y��D���:����kLY��a�`O"��O$����~1j+�����M��c�D'�R���ŭ�0W«���H<��9:^2p�2ܴa����ޡ���蹈��=�?���\��ſ]	K vy�OX�>��_	�i���^֡
�дG�\������t�
��[��BJM�Q.�5ȁ�Փ͹Y��0x!`&!J�P�@����@��ϧ��-;Qx��@�� ���Wa�Vz2@Ϛc�9AMh�u	���)�A����b5aͯ�-��K��`����)l��3���z��	u�h����;+gr����6�=�������{�~t������3).z�z���
����hMā���)���'�{uR|��U�hW� ���Ĕn�m�����V����Q�_��~���
�[��]zZ���2`\dB<�4�J�By>/\���	�Z�v�UA������NJ��8���0j�q`�\E2�%*P��.(���h;B�ϻ�3*���?a��q��Il�� u��)6�`N�E�k,���@�e�0U�M��\m(�g�Պ �O�@���r�L�\�����0h5��B�'vs��X�5�������:(�_v��~޵�p���!�e�F�r��c�����c� ��#����5)aw�I�R!_*����k�0��P��2��>�wG��KD�h���sUo�6�#�T@E��	^H��FD6�F�A,})�'�^/^0���8��Q^����[h���8Y��W���1&F���Ш]1:Iρ�?�a���<!��X��81g��Bn����h;�~�j���aUvf���D�p��LB�CwL6�!�����J�Gn�DZ��1�g�'�^GzL�D��4�Y�UZ��R-+���!%͈�]�s��Z�$����Y��]տ.+׬�KĝE���;���`�eQֹ����^�#��!���%2�N>B��CPœO�F^:u��:�P�����jP���RٟX�������G���I5��W��[Q{��f���m��#���d�Zx��5�^���s$��|�n�[�]�4'�FW�-%� ������k�s�Q����������.�N�(-�O�>cb����8���f���Ϋ�5��B�E������8b^^�+�(F-�l>l3\[!��`�H��?K�!��8e�Jy�<� �柷+�Ii[�k­���Ze.��'���R�[�7�Z����Ǐ�Kn�����>��g��Z�Dq;XBz��[[j�)~N��ׇ�!eȞVL��="�^6�}[��p&�@5���Lfu��UjfZ:���A��7*� _Ң�2�����Eh!u�ȅ�z� ?�8ʫ���ٳ?e�e��=��bu�����ڞ�W�H�K����.�����ϗ����l�c�S=����[DC�Q��]�����/�ϫf`F�"ro3�,�ů��F��ɭ� F�x�`��T�PGAa�+�3ݺ�����%�Z)N�@6�5˴���t$�rc��O�V��`� ˫����~�����㞃�Wco�
W.��'Y�hθ�Rռ� ?��F���	�#* c��;|!� �=۫�Ad�uR�
���|�>�r�֖���U�y�6�|�S�B̎i���5�07��	*�C�!�[�\1�-��aF�nY�ߣ?ծ@M��^��{�r�@J�R��i�N|��bzψ&xlE<�R�K�~^Jz�������8~�FŜ?��ڈ��>Se�!��5C�f�Ћ!��f�@n/e�����v���}�-�;w|�4O.��
�w&�ZU5K��
$3���F�]�;�P��# �	;�vQO��+��A�C�E�C��`0x�;B��S�e˧.9,��$/�.����-l�$o����O}d�lc�X�]KeR�z�����,?\�2mxd���GH~>��wz��� �
���zcv
S���l��-Rt��Kˋ�O�zt���w�D��my�?��ER��]�Sɇ�o*o�������k��C<�|�XZ_��_�<%�%eI\�Z[&�u\�>A�4�F�^Yה"DB[v�4��}�q����E���X�%r�͡�"]��Rˉ��&@����P�lIL�?���E`��aY��\���q@�F������Lw8K���ڷ�lwh}L��Hpb�3b�:39cӫ2;���ѝ+V,������g��C�����oOlBqA��˯��"�����{ Y�%~��u�}4�I���9��GZ[����/�ܾ�k��d��yu�I�D�"Qz��x5w�b�Clc>ehb�c�Sc������^6I�J��qp$�?�"<���Ĺ��(�������|�� �� h�����s `���!����g��/����T�y1�T�q�_Y"?P�'[��V�`�NCR��l��)�A¼K�����GX�?��<�A�$<���Ãӵ��J���Tj�G�g?Eү/���%�x`�U�q�R�s�k�6�]d�#-ղ� �A�DᢻU��������Ub!�l�~��RQ��2wC������� "��&wa��?�p� M)�ã�����]YF
�S���N���ԇ�`��c�n$����T q��b�F+��,wy�uF�9����I��p�^SK�ݰ�M�h�g7r@Ǝ��'ur�8��1�P/#���8�C�ʶ�*�A�mƀ���I���T�|�{��I�ƕ�xW�T#l�K�;<���9���W
�ې��6��%�$����|��}K���^NR�P�Rx���(��n�G��{<��5�t
Όc��_{4)�aAʫ��N�
x�R%]��}�^4�K�j$�%���V�����I�3��Z �J'�/�{ls�7�����7,giI6e�Ӫ���]�1�I����;��gH��^��$s����?J\
��eAh�ⵥ�h���W��p�
.@N�Rsy�b�����u�`��È�M�Xrl~�֌OTҭ�,}��2y��Ɏ�����o���$5ab�LAN� ��VnV�7(y"?1mw<�|De؜�wݯ2�o9�E@b��%��x´	Z�&�x"j���b�s'��FK�rݭ��I��0��C�����:��6�M�f&o����/��D���s��ۥ,�v��Q����9��d���EH�<��;|�?\�Ҋ�|�Ct��<��d����2����G��(�jX��^_��F#�����.�pٺGma�����@������L�A����� �ltx�B[Ԇ�2���&��i2[��m�>bo;؂<�Q�4Sϑ#���5PQJ�ۻH0 �R��r� ��&	W2�'�+̊7���4�Z�z$D|�~����U��e��L ��J�Gk�����@:Z�LˠǊ,W+�C����I��P��Ս��q<u���m�M�ɪ���
(*�MQ�;w�DB��o~1�^l��*(�/g]�D4t���7����>_r���w�^��L����$s�W����v*w�ƚ��`D�!L��Z&<ڛ��n!�<���J4��ۗp�"��E���������?�Y�bs����J�`�XSM��I�ϰx뿜���&� ��d�^�~�&ᯢ}>l	�f�ua2����Ah�h\�s�#_l�TO/��R�Ou;j�yMrc0��IY�ɤSSo�ϻUcU��GLJ�=35���Wn��Ѫ��C��V��淨иq�^�R���!cf�X������޿�@��%d�:�]�2G�CC8 ���޻��=L�N�6��-��j�M����h�c������-�|�{H�b bA��"lP������ޖ�g:T�D8��0?)�Z\tP� qXB&q̬o��T�m^���qU'�����4��]��T�^�f%��W-dD#N�F�t���>��q���ď�Qf����e�x���wB'I�}%�Z7��'K��hC�UT�Ĩ4ed@���>�C�ă��OL\�-���Qu`:y�gU�v�x�z��[�XJR�A�ۇ�aґ��L�����])R���a�����Ɛ�o~��\�lEw'�N�l�3o�ǃ���a�zc���^v8dF��n�+|ֿ����f��=%r����%��� ���
NC�'!:�`NTD<M����g�-yF���
��>��Rt�,N�_k�}1�ǲE��@���`C!ki$�]��@<1\���;sP
	��Z�3XP�Hl���n����W2Ƶׯ�{�uƲ0�9�#<�Cw�j�:�T3I�6�1)��(/�Q�0]Ҩ���&̞[��!�u-~W�^S�=;&�F�����y�D����Ar�"z�(V���fHA�Ք���u��N��4�6RP'�SC��~8��5��j�ks�3���^g�E�2}���Ш[���?�~>���5��sq�)ǡ#-V[����@58�O���� ����2׉M��۽��Y҄d����b�&�8r�]+���FDQ�~@�i�^|mJ�����(%.ēVy����<K +�~������+��Kny����3��K�ꆡ�4�$�!�ٹC;��t���'zD�>�X�A��5S"�C�K���4Z4l���ق�[- 5�T0��pt�XKs-k��������>�`*�����������춣��{�~�)���r
�w�7ɱ8q�^���z(*�IY��f탱���G��ό���B/�!��oˊ`�y��u{����?��4�"�j���8�aZ�B��S�?[�Z�fQ�p��ǘ��c>,�	�L5�
�M"��5�\}�_�(�T�XMJ2���M�i	�H@��)��LL�P)$JٛxS&�|ŁZZ�>)��q� ���-b5�MCr�)8�*O�z�;�O���/,�.�05��!�;� }}'=�9�<}kԇ�B0꡷2��v%���K��z�����P��L��5v	���M���C#�D�Sʉ���tm�_8N���qg�Vf��<o�����F~5�^���f��|�x~1����e��Z������U��2$�ª�/H�!(e�t�1��..z{�B�"���t]�7�h���]@l���\������^��g!���ړ	
������>r����k����fUGJ+��+L�L�&� x��-��u'��i`1bL�jY4�I�Kn�ٻ7�����@�Y��s�W-�^L�UY���
2��2�J�Сn�o3☼m3s�ԅn�t<V�l�ǐ��Fg��Wg/�=�Հ��aV*S�"��,�\@��#�㻆S��i$��a�ɢ��N����AsC�y���ӓ�;�K�1OƤj���I��p���UXG$�GI��i�I]�R[��U���,���=�&��&o4$���)�s�+R��g"d�"t�G��´����~�c��"��E�����ɷl���dI���&ju=|1�"�rv:��h���Y{����6��}��?� HP�Cy	���}*�^|�v����S���7�����z2�T����\zzo@]����'�y*I��_�\� JQ�:$�GO9w��m�8Ի
t���c3��>�5�盧��c���<�p��Bt3G�$���,a $��_�!��m�KE���(#�__\�M��`�L�M� ۣ��]*�`�%��5���I8E��M#�����J��Ч#�{G^���o��<���yj�=�}{VG��\�۠B�iŚ�!x�7]��/S�y�����g5A�my�� �<<7�"���\LW��37�a�N�z�����	ےP���c�	��w�F�>�	(����X@�_�!N�i����a�X�� ]dV
��v�C�t��v�G��k��&檾XQʣ��q�h�0��i]�0���k'��G�tOI[���˦��ݣ�����+s�j�#�&��u���3�ʬh��lt�1��K���)rpo���&(�c%6,�"`��UI�踷[���i��C�W߿�����O;����!v1��	�fd�2���o��BVI�I� ��{r҆#����	=a�<P��a@��Z-)9C��2�|�A�[לa躥�# r�־�[��d*��pͱ�M�8�G{	��������4�O��8DO���Ig�W�q���n��l�4#�����Q#�q���s@�p�T���]�.4 ֖�'j���Z@���wEZVŌ��V(
��t��kP�||楟\���+�G��AY�}���Z���_�4��}��L����Q�M3���Ou�CH
.�jZ���߆���&��$��Lj8$L�N�Bk�{-�Y���@��y
N��x
���S���g�,�k̿���R^�J�+鐠[��,�I�\�ݗ�̎��+z��������N����}穇ä�[q����4�Wꋑ�\Eu�%��զ`ߧܠ�
��� ��4 ��X��'[ԟZ�ztȶ}�l୴ >�
�g�	ɞY�"'F%J�/���R~HXR�j��q�(��4_Hr��˒��-)>7���T�������/9���w�e2��ib��#��b�� �kN�-i%��
��8���i��)�ke�%�[͌�8g$͞�7kf*�,�/��&c�Gn9��d�|�=��J��j����`:�f��ih\�/.���߃E�4�'����
>��o;>
�� �,��Jr�ڸڗܼ�>�l��q*�!D��!�
��Tf���Nw�a(��ʔǊ�� ԛ8�s=�~J�,��tg���K�*p.W]�E�z�m#���5��&�����e[ܫ�VLE�&�6���������XI��~��"o9i�gO�$�ǹX���dkJG�T�"i2��0�Ab��A�:��7%s)�.�ʝ� ��b��W�)�*���n���Q��e(1���=���|��=b#k'\i�57>�p9 Q�Ծa��V�&���a�"(������Qt�A�R`��=i��'�%P����P���A�W���	���JD�K2��b{����7��"_d�������w+���K�������搥W]i��`�U�{�3$���~�_��t���
���n��T���gz��ea��r�_��H�9{���c4�]~�J|)n��dK��W��_O��˂���Ⱦ[��
j��WRl��R���u qA�U姪�)��������������B�Qo]�n�3$z�ĳ��!�̆#�����|��2��X���[	�<�D��8�C5Q���~bK�%�u��%|�J\#5�$�r�<O�*w>]�"U�J�H,Ԉ*-�i2�%����
�!�y�n�|G�|x4��l��$�B�V�^�Lk81�_���5K.*�Y�'1q.����$���`�� "��$xTۇyٽ:�pca����"���1�~�M�.ȓ �RRw&����Y=�$��f�H�e4D�F�w�e��m1*��3hn>��Hjn;�:�od<�l����I��O\n�����n��t�O����} �j���M��[%2�r7#~��2��:�B�-XG�`B�S.|ā)�N����	�\�)�N2��������
kj���D��/�3CU������P�E���ٹ��k�枊�+�W �煇��@�ii��w�E�`Ľ�U�~q���G�U��ud 8�]�M���w0�FTi ����6Z�Dx\b�A������U��jt��ḧ(��w`��@�'B�٫_'�����B�8H�Wǈ�&z�]nj]	���̟�T�nA$q���P��5loh�۾�7rS�xk�����̂~���j\m�����;	���ev���Ǭv a����u0i���&���2��̢��o�'���y��4a7#�������Z�L$�� �'�%)����6����\�Q������{�q��^T�JxZ���9B�(E�Y���!zy�f&��/ᯯ'�!,�	T��:xSL\����
�e���Q�����m����7״NY���O��UD7�A���;�gb���F��
a�/�:�^ॸ ��Em��[���R�y��6,�he�C���"�Y��`t�+$�"Y/�*hѯȫ�e����sЮ�֮JM�'��R_��d�gy�*�Ύ��q�a��y~�bw����lp�H��U�7�Ɗ��H����f��T��t���\���׷3�1�����/�vQ�鲾6WM����I�c���P�3��r��.�oL//%|XϮK�--#o��-��U9QOIL�Z�b&��3�\�51����DQ� �_a�+
�70�Ľ���fV��&(V�;m�I���<��%�d�"��<a-�ꏥ=��ܽ�[w�u�Y��c{�$�t&�<a��(I�Hj.?[��N�fL������D�F����$�c�49,M�Aݰ��v^��8`D��rLKX��'LG�D���څ�L���6T�*l*dy�I5ƿ!:OLj{�x���>yJ��Z�U�AO��v���g*� 7"�D *�g�Fyp����c�޻#iCAIlg��C�)���B�`��>���3#��ү�B�@�0thݺbn�3�=}�@���
�%�w��sĊ��o;Ʃ.�w�R}��n4I5�Z�D��� �Oq�5��
]a��T	J\FZ�J��^�1��� :H�I�ke^I���'�W��-.S"�ӣC�0�>,�;A���ho�ACg��Oj��5��^��1�4�?[���_Q)���9�s������~vA��a28�� �\����l�vֵw���N/m���<��9:E�*���Ί���T��Ț!�\c#�6�V�(��}m��*S��Cv+�ݠxW�-�,��:�H$LY,J5:he/��V��H�A��͕Oyg/�f�>B|;�j��$PFG���)�+y�����M�nu��F0�o���чt7�H�+�<*��>�}�򨞳qY76���_���������[�-�}C�K��b����&��%7��
�ko�ɟ����,`�z5tBt�
e,D�Ɨ�N�~��8�wV���8'��h�?����̽�Y��o�)Z�[9������SZd�*��Li�Q�N�}�0)�s�=�--L�+���I9������У.>�`{ �=�.�|%O'���sXD�;+��5@x׼A/�&�lfS0f�Og����F�Gy:�u:~�s�FiD��66|8���j�K�9�|����y��q,?t���"����C$Æ�J�����Y?�N͖�y��-�i��$��=��X��R�5�����@��b��B"�]\�4��	����#6`y� ����u�Q���	�m�y�D����ܵ�P�uy�?�͟����R�K���HK�̿�9�\���o̺�H0�Ռ��!~��c�њ�%p�mf�]B�'�V�8E��$��k�&@B�7�oظ��WT�ڔ���w����^9�3�ؤzn����?�U�h�p=�Y�
�.��y8��~���e���fvIJx��H��)���m����-�<���K�x�c��DN%o�2�E҅\�Z��t=�[ۻvB v#�T% �7Mժ��QC���x��7���j={�/,L���/���@�Lp�gB��,���� �(߾V�#1L����^��+�NJ!�镅������ �VW�m��/��Ɍ����"o �'aPP�t�*3yi��5��h��F��>��YR�sd{O��E�U u"��Z ��걫5>0yLd@"�j����ȗ���(����m�`fAX7��+! f�{�����lbF-z����U�q�\��E	�T��W������B'j�k��Q#��6]Ǹ��iW�2���ԯzA��f� 7�N<�"����xw|�A�]�Sb &f	��Glƚ�PI���P1jKP�p�^=�6����d��c�&u��!����jeJl4Ġ7ǡ1��B�'���.�mx:A�Ba���@P�-	���T������m��m���h}��N��;�q����v�73}Dj%�ơ�x�O����Hm�y�Y�W�25��p��vc�	�;�V��Ĩz#o\�bPH��(NQ��h�x�ލ�\���{@<�� Sy�#��F����`!�+۳��K����K��|�߉mmH�=���3��T�k�ï�&a�(��s�s�'2�6��k�
A���.وBNS�jfeJ���D-�E�&�+�B5��ު��ֶ^�R�][�;%�"@�L�pϙ��L1�e��n����3t��͟��ӄ�~U�U,,ds(�������D�c�Ơ̕A&B�=�l��m;��S�3��|!��9�TQ~&�����F���u���BWv`ǎk��ˈ����x댻n"Ѱ[��p�%,Mb��F_��'�5���|(�X�8���:܁�	�d~U8WC���W[�3�@!�3�z�w_�pr�&�t�nu([�:�yŧ�h$�;�&~�"�qnR[@^�A�j�/���2V*���)%z�=��
�n���c�VX]夃	C9���̀���8[���cS��u�$w���&�ϿDs�����6�����e��Gm��7�L�z�bJ��<T����՛<L�אʯT�d|3���K��Q]\���3��+@e��ब3c|�]����.jW��B��j�)�A;�Uq�ҽH�ϼ�R�kCr���V!��K�h|N��cA�8�
8N��w��Q���8�N�7�A�"E���ק�4/����{e�HK�Q�ՅÃ#��x��7��5 o�3��T��.!N�F�#ġ!ydR���9��g�H\a�w�,�]E��mx̦��.������s{�	kKX�[����J��N������5�i�Q�1� Ӌl��W�=	�\�������c�H�\�$��I�i���������2��*�h.u�p�Z}i�����~ER�}i)��?�Oݿ��"�:���r{��;��|�A�quY�q�n�ݿ��'��]  �,ܼ./���4��Vn�l�vn͉cvX�{��Κk�f�;S�g@Ǔ`������Q
Ͷ�K��X��+[�������L��oh�aK~=�*��`�(
�JBJ�ϝ,��/����aԼZ��b�>b��%=.W�}�c�I�-���������6��P�"=ù't��E����z4XxD"����4�0:7�MvH��S�q5��(�ϮS�d������lH��;{�����%����r�ݰ�<�.#@�G��;VΥ2�d{BCN��S�aaJ���n���>�J�R�5�9�S�/l�FOyM�$M�F� ,�/:�֛b�^�Ji�:�?�_Q�S25��p�D㟆�r�2u�/Qb݇߼]+� jc��.@8R�����}H$�`VrN��p�����hy�s |ٺ���l���g�� ~l���@�jz�A��p���M�V�����8a=~'����1�h���ٖ4r>�،�jN����Mȏ�yd�"��������q=�)?F����n�P��:t�q޻����+qW�}RkwT\���������Q��c������h�)�G�h�\�8lQ*�:sv���d\߾��������;c�?�Y�[���]Ͼۢ���BS���^���y�����6G�i(|�?9��RCʜC�#�����<c�"NO�?�h6qh��� ������
q���M�:��Z|���(4��j�ϝ=Ϯ,�)K��{(���׼����\-�P�B�	�!/� �Q�����	?AK 0�Wm�J�'��H�gES����C�x�����Kӫ����d���hWz�.B��B�2�yW��B���2m)��9jS���F��q��=�ƱPB���u����'�݁Z�F���N�5�N�[���'�7+o\D���H�'n�J b+O���ce��w�4����+\��(�朴U����-y`����vn�}1�����9�)R΢�ZJ�E
���V=��$�I����$ sgt`�+]N���������<�Fd�"���p��������(�	i��G��(��+���дw^fF �Tp,�rgR+5�ҩrW��ܜ�$�cfjE�oЎqzh_��P�DGe�V��Q��v��e�J_A4�.���)�Ʊ�f1s'����<s��e\�~Q�,���]T�`M����a	���#�<$(.��&r�a`�෕����	B�(�Q�N��ycs��5�&���ʝ�y[�![l�w��͖<)Q���!��c���{�y1��l���s�)�3�X�� �Œn����3Bc��8�c�������j<�����0y�Ź�o�õQ��L�� �Eq�q���bNز�߲��I�8�d���W� �M /�%RQb�=���_����������L:�[1[�M@�@�����-,�[yH���q�_�qP��%�IJ��^ׄҐ_O+S��P��Zu��V�߂'݈k�������f� P���L���6�UX�v�ß���o���wƻ�r�(�f���Є�PC^���I�C��� Lv-H��0��^�VtA��uz;�mh0~Հ�R��NƯc�fT�<�YquaO軼`_<#Bnkf"�R`S�p���u���8�@���>�Q��i�IS�L_o��?�����Z���oųQ�� ��T�z�T���L6���ޯ��d�!��I�_��C��{�ɓ�~��`� �T/���}re땛����5ل^�l���We<h\��z���<�H:�p�la�;!�B�`���}~`� �uoL�G�	n5*��c�d�m�&�j��)y$��Ɔg����QK�וq���0	j�	F��:ͯƓ6�*��c�z���Dz�K�_�D&(*�kn���#�T<Z��}E��<I�P3����S0�&PELo�Rz#+*ʮs�!`,���zj�~�nGvאL{?sW�y3āS9=�% i��#l�ݻ��0����9����Q��2�}���/�֪��#��	V:M<Q��#F뼞AҼ;�]��� ��T��9�0��U�6T�,�g(H�å4��Wxf��xiwR;+�Ⱥ����H�!�»~�e����SR��t��|G��@#:%3��نzI_k�hCx�PL��k�L�v��M{�җ�a锉�����DA$郸�J</��=�?����`�5�e̕�mԶ:�ʁ�W��I��q�$�Tˊ�g�,���~Nl� �5+�p���U;���drg7��U�Y������	n���AF����V��0�p
���i_-D�W?]�M�BLS������B��:%��U��m-��"��;FE1'���������K���Ku��W1Y��
�ەHYRd��p�"�9��Zȫ��.��/H*eK�ޔ�����~({�����I����o1X����W��i���h|���ʆd=S��J�o��j^e�PV*:�� ��[���'��&7�Pg�W��ׂk{�+;f'��$�|��pj���Zvbߩ�������t�8��6.b-��*Ke�`��'S]������{k-CS�.K�H�i·�e��i�2bZ�X�
ۏ�'|5i�C����q�R�vה})�_:�cS�N�K:�S[��2df[
�NAw4@��'
��281_}��R�n�)5��������?�j�z���͹ms��eT�-
��DE0"����ӱC鰖+x���q!!	�a��*��Z�A/��5	:a���1f! %Pq��Yeg�"򳀱76@x�v�k^����Ys2�_C���1km�~�����x ���:7h�H�g��6Gf��i�}���P$lm�\�7�)��<甚��}�YT��<��#c�+�&3+��4lI��w�O2��Kp<
g�Sa��������ګ��D�ʿЅ��G��0�\�ZM_���o��r0��S��9z;�v4e�����t���,�AyOB
c�t2=�S$!���B��ف�^���&��_��7n����F�c|���ji[:���by�@\��H�SL�_�M�A3�>$���>��_i���+@��g��FE<���p�ԟ�&:���ݿ���I|��r���n�P
�v���8T�5"%�>����zg��R<:�\tk@�)ʈr��*�)��$���f���h����.�8Q�ݜ1����j���
�:b�R���Z��U~|������1q?>�ԦS��!}�Z�	:���:�=��^�|�O5{�ޫ����%s�|x.�^P�(A N����t�sV�l&�d�$��D��ׅ��V�=;I�эi��� D�T�h;��Z��� v�㢇�]�_�p��|�ϫ��.�0% �8"s�V��W
\$S,�� �+F)#>G�����z�B��ZOu�Ͽ?O7����(\���F��Rl��-1A�A��¦'���~]����?��W���6�lP�{ʷ�h��<����CB�Y��ӿe|��No��]�坚�1â]�}<%W�N���r�Z���Jђ.��Kr�&�����ڗ��e�)�@�4:��\S둅 �����3 v�^�
�w8y�����"��L���QZF�BX!������g�ر�M��kߗ�0p��x@J�87�H�h,������>�ro�'�e�G��H��V