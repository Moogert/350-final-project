-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pwySr7E0QzlMDqVXENCUJSHyE0zmCWxQTOcktbIXEIHpaIdA4yasmZmFzHjT5UbyN6MDCjLg2LWt
0LXgm5tseAScQOmRf+cgLnibwbTK9/MhdzIN945LHFEz8Pgh86qunt9KG7UrTKm+Udaeg1Fz6+z6
IoXeMtj0Jr4blnbZHsJmPUwRNX2RAShAlutZLyDTvPZeR7Tb8oUYbl3mYVtWajM/zM0iCkP0KrwS
Mwh8jodeUawf12gW4KWjvi2VJfy9entPt4J2l0UIOj/hiMO3Hq7sYmmSirr1/RrASl9y8HYk5+Vw
I4ZfPthJccoIbwkmh2G4R6yVNkHhRsIGGzc5wA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
SZdpKT+Xh3H6SgJboWLkIhUU1KPC/KMKx3tyWxMMhGq09TNL4CY/NdN5oieEhphFNZhcoDSjq16l
DtIkrNGfRmg62+y/ZRTkfb9VtD+jx/5aiqQZvgjrBLN182Y/BysV20RdyVJZknIzBk7foNs14iYW
gAMiem5ECwuj+cif/yRhH3N3Ctajt+TCD376m3FyeQyB7Cf7D3WpBchJILyifAJQrw6v5LD/fd0M
maSomH9pefBKDPdj8P5dd7x/FDX7CxuLrarBqXV1pkmf+kxykNv1O+FV1rNvyGmpmusJYdLALKhJ
J0l9xkLyRLw+Ntn5/H9bD9CircG2IyGidJKd07BI0Av+Q/pBA0D17qrsInQ0O9g7Dsvrcock7CIM
wnyWfJNJe0NXfQuT/a7lhFDX+Pd3J5LG7b+16znFJPTG6lOfTN/KpYCE70ciGxYENNCrDSvH3qYh
OrxD9r8nHDhm151pHhrPFiS/fJQBgLgDhrBuUhjmzFJ9G76nhsl+XobBOJl05mVt+eLOgfy19YLj
f3vg4ri4qgTcKgvnHB769r8V6JbwFRg/Cle3vq+tkABT8jvzUxoTiVt5Cun39pruM36CjtjJAL/J
hYEntnxe6Ivh88Z/OY1iWc23PtmcOhw1JXo7dJl2HKWGTppnkrLv7O2JA+tGygSYgd3Vq5Qgb3TD
ZYr2Wg9Hc6zfcAtB4VQWTVItBGlSit83Ds3hlYWULv4JBJGrCTLT2fj5MT0cdGOIPVmJegaaypuN
5WJpYkJlVoWcDJQYpW58Bk2G/eOp7IGlgdjpaZUWsfOI6yoopqLYWmIOL9SY8RwyP13Oh0s5gcZH
Vhc/CMXSNVAdCFo4sH07/YM92I4TeNWQuYADdsEEFc7SNZ17RqwZ1BLH109QYgZoJ9eZk+vKziGa
U0Sr0RWoQgLIoRwVa5VCnZM9oBHxqQiMJONuGLq/cuimDjmYww5nADcn+EczdF8/5NYV3TFvDYwL
wEE7YOnjVQ3ZUzUe1v2FB4OT7UKEC7r8I+31Ms4wyNtibKt8Y8bIIjp3QW0Y5QmM5wJpZ7LFtmJ/
elIbMjSZP60KdIaTk73UrOgFGDjIj69wurFYIuap+jUcERFw9j5tvsrEQogFh9d2spC+kGvnvQJ6
UZrVHCsOwTc4AZcUTCQS6R+W7n/aUH30225MYqEClqGNZDF4iHfw+cmYNdRl8wMWxpH2P8tk93/j
42I0ft5lGj+qGO5YgGQlKFCZ+RnBxBF4mcT4JHKfl/eG+WyREF1hefJdG4kdUzW0sBIdysD4yEJF
87wy74nPe6kEkih5dogj7da7H8SLvILE9Wv/UbKwOQxtoYLpH1BR6zxKY5BW6DLn7NOAWPM3azU5
1jTyGwbi7e+TtyWdkjD4NyBhOY9BCD6TH1PpLgu7zX+EtmDki3j0o9bxy0sx2ncmTScDiwA4rKr9
9cnLfxGpUwuJXJPhZ1LTmV0sFG9C4mEuNhxeNce37Z3CKoSK2P+36J7AodClItyyqybty0yZYVZx
6DC+W11qgdFQIqBotaIndh3N4UF8Gk8VoF6bgBtiurBAfb6Ivj8FeiI+K4iRsMchug2SZ4RHoA9U
povlpX2Q7EN666ZnR6ZlDI7bQzNU8jMzjNXjK92ESouaw2uEqGXsHgg63wMHrcOYE7F/4Lp5LvW5
ep5wjFw3LCoeIzQiyzXAZlUL/ys3L1g8kCFLEYi3KwgXiO0SppHAmTf5bXAmDC6v16GnG2t/IZ2l
eM0c7Xk0bd7OfYeJ4b9F4/Ke/5xMzzTC4awo9eGfhFtVs62Vpgfz8T+vMYNySjg6lCpgSQeoWkpd
SGUDB2HAiUfNg4nbTiUqjFdmz2lSd+8CdPgRlOvrn15ASPBIxZ8ARXQUwnKk8wH9KS3D0d4isbZR
IKR+CI8DsZqfGBHGUSACaBmfsQbajxDHVFpKJ3XdW8PZIqVXE4SRMWI9NWGNpLVrgujT1oHrz+VK
F86KVxOm3gOkjGgQONLkN7+ZlLVeUqTluZEJzPjmne6ZwI0PUjpFq+lCLO9mfh67jOVBCa8zpDMv
HmYKltq978saeNCVCi4/kXRE9T+mJI/sTuNEadC1eTBdZ7V02Zi0r1/+E69fk0gxttChvPrxRF7f
Xt5Po/YnrG8c2+AvnRj3U7zm1dLZ4W2MplALpr8NFBeGixx1dldR72KZflU4OwjoueHvEHiVX3XU
ZRunkvBJTcHMk7YfJTPMk6XsjidAgo5A2X3PayW4cGLyFw+/Trd1Yus+CEpE8A+PrEfT/g9Wo6bZ
YQ4ewPly55+ur0j1AphAZ9cE5BSu2AOOkf4yAvmZpZvwFQqaMaJfm3tKVg2WUK5kwcNV5Hj1BlBH
iBvXr2xSrLqQ9mtOjtrJ+6NTI+h4UA2pJK884nWGqyK+vuA+lvGIVCpmAuro4dEm4O5q+ofAu3H1
9bFEvOIeFDsEs9yCL8PYfH3gZvC0t0CX1ZkfFJvS4a6dPkHH0SBRaYvKAB/uTlnnFvM1atjGh3Qw
RTnO+9hxNtp9CUwUPzt591HiD9NG7xEzMFoNl+0g08M2IKtdDzR7DpJytQN7Rw7rhKC7bVWE7ezr
XE76m0J/NkVAhXKyszNFRkMEn7F+U/P3gMm6+bqm8LiU7HgAz50bT6jP2iij9qnEpZCI+7TXDHfL
LakGWSBec2ElbqjOLQvLz0uKZcC9kbrol1xRLoJYuIZX5OELj8knGynhkf6hr+FxYn8k29s2MUD6
l58OWLL3ccMR8+uyuwwPv2iBDCNsnfovOlW02DM6zZdZJjQyt7QvAlkg6C4j2nm8NvktAX5itw2l
nRI5pVyT1ngUrXa80+Ug6Q9Q3xqDWf6J9SQppf69mZsqONSVgDgULAFGmeoTJpdX54k+Pgg24vf1
M3g87ofr7GB6UdnliHMczTZVyxQh7UyeBiOiCi1MfyL/Nu2FByh4tPBiP9c9Wf4+JCSNtr4GdrBd
/RRj6h0zkJU4Vt+35jTbxTKA3uT8X/eMCl6ZFZvSd4sCEVHYsijiZ8vW09Y6YkqoIkCnmbRH0c2+
LEZozzJWFZs1rh53iSWV8zEHJ1Q5hCL5kA/OXD03qk5lbP8zqzw+FOMAroArj/QxNAegCWmGiVrc
vJbIiA54SJiqxUzEFSCrUPMXddaWwgaKHPyOxn7zZ8QzLo/9Z0y7U+/JQYGAfBIFZbIxuqY78zUD
5bkcy8d4Kr7GxxRTZOj/dA8CJteAt+j/j1iqKYUI2CEB2KribrygwHcwbfLuGd6hJ585N5D5dQ1+
+x3OdUqNHQ8LKkHombbZ22v11dIi2km3nZcOfOQfiakVHQoHOmIrVf9KumS61v1BneLLWj/3EcZc
Q9LjSvIcRNK+WdsNp7Uuqz/PrHLHf5/gjsLeDJqpZloG3UHemmzMlqqXfvIc0fho2XQbOl/f9t3o
vcSpp74ji9S1xpHC6yw5wM3WZJDm29YADDd216VzvGytDLvXknEBNIj+0Q4t3alxfGwvj1zWa2S1
qmDp9v/KdKOysfSb75A1BEZIKCLnTxlrCA3WiKQ+QNsco3DyKg6NdqVeREhGunOGUUpVwsdqzxut
1HQsVmHD0cwBLrkiZZWC9tGYtSGSIpBNVG7U+cmd0p4oSTT+d0eSiJVbeBLoecsc5Lf2blOWfi50
vjxhPOOhrUeQvTzBq9fegzCC41Qbg3V5tQ4b/C7PGJbnSi5NoqdZBBUxg4fAJY/K+jt16xsiEFn8
I7V3pYyhqy4HwHk4BKVCjmwZxOl33TGJ8PIhM6vx+iiHY8C6atQ6oe3hocf7+wOt1KeKX31h5Y5L
Tq794rMnfdchMDaIaDre8WPlS14JR52ahhZdi5TqpK+jq9q+G/XJPGdYUdCfP+P4GFvCnujfbiUl
3S1X1ftJ4ZpPvT9d73udcFgWFKOMvXLqXZzX8+mNGK9TK6zpi6V+zhQ2ldcgDZdSYlfWVqQjUDzA
JgkYyI1SkfWMlAI8auYRoPP0CFHK3gJac3ifPgnoABWWi1z3NBwetz80JC/HIkpKRaYhWwAX6m8H
2C87oMm/5+yP63/yiwlvC1dqwJnJ8r1Cxg0XBPmhNGjzQrlVMFdo1QdvacQVnaiKPFFVjGjCw2OJ
VkiKqGLHckZtqsaTtkEp61Epo3TrM3bDDsPMFTQqOGlseeMOKSnxdDiF9OhX1u67VTXyUVjx11lb
JJX3ZWbFSIakpdwlO240HHe89UCd9VOAWYpdPYRrNN5QAbShf6PaHiBJSahjnsrW0tbaRgeX6Khw
W9e/eJag4qXvxnBhfodtBGyu1II5quawPQKPPkX2wM9p/nRI2chccHeq8Wk/KyOAB8l/okOfQjED
37igX9/Bbx95168dpZOBX6dhSpQzJzZwd7/Uo0epyaMdESKR5hft4AJng9aLdBqqE7TWmzQ65WCa
jpBgZhIPoUf+4RT8Vs2XkA62R39u+G7bzSKTDmU8i54Ufe/hOTbT+ejTg4dhO8qyc3n5HoyclZhH
KkXaJqGJPMeFvfSiIFfI0hqdXjZD9zKsg31FyLZdp6vUAzSnhkMWXBwpmi15wA0sS5Lzct8e39YC
5TZRQnRrlEJ+n57bVTdpl0yHQd93804i3gR4qOQLvOAbqlVfz5NBBVMV3KAjaB1yM7JoEZatPR3j
M2w5od1ysk7xqQU13rCufZPVG1J+o9RpzbyJ8xaOtQ+s+1yqvTubtGYuc5sRMPxkxHR7S9JZoxun
SyWFb/E6oa6mxOIVWXt+DZSrqtZ69X/08eb/7yS2vrsoP6E+5J49rRpGpPSYEkoI/PsM36EtemjI
IQ0ppghkXGhsljLuFVFuedS082n6k3OVXDH06Bk613TjVp0j685o8fpxnwD4n1/wXhUP8gfr6+iX
TsxReE5SI8T2KwNfiFfbpQsQntVsiUJtcXEev+Bx/roILxv83KF+dA/8Mpm0JFNE420CbK2ujCJw
bSLy5rk2Oza0D1soGBXHfsc+KiE3MHYnsCZW4R+FK3zCwRBKNBtHBHeYu0pUwjT+/tadCl8ep8/E
ZD7yF5O954mT9IP31NQ2G+KKgAmtAFFeVNdp+3zFEuR8sstrydgq6lutKHiw5WMiKcDXHV+3xYl2
LFf7qASIT35WEECEiJaFKGyhKJnsOE4buAUITTV+mcsd5Bo7+su8FWLHE2DK6ntCRjh+xZH/jMt0
XCouns0172fhnu+Dvg2wy4O1MTll+iCKDGQ5N/gvxZoNSAd0liKhBVpXIGvmJs2IgUJzDvu5Hqng
bh3okZ3gwrvhmT2OUHXO7SawLKCRV+4yx1ZdUV91meQO6u36z33ichAlq2TPIA286amsYYBt6tGO
s1kbyqZFdHhXEQxOfw8AGWjXfwSdwzGIWlFc4njLOGiP15/8ISoo+TKLJ4Wknb3cn8XMn0qj194H
VSCS/7y9sX4YVEXlSiQ8H0UNFLZXKaAPoZiT08Ahphpirlr/DY3MpoZXUeh/z1S154/3d/VKpP/F
Qal1WwaAkzFFDZ2qAKSwRl4xa3gvzsDNfjKxKW7gEPPXwNPYRCaOmQtvuiyvPP3Vmt4NKJI7I7ju
r2uNGY6koAyniyal+l0kEroNAUPydHW8EGaz3KI+RFZum6djrA2l0dBMxxk079HuAZQiJmhNAxL+
/stdo4B903GSZ4bvw/2A/9Gb74fsZj1/xIi/7HkztJt/GPYn3OdcN7p6rGTLqWZO/BZGmtJaKmta
rFq1CKadbO2sVv87QXQ8a4FES9UpYdd87dwD3TUaRDyiifJXOqlWkQKrqHNFMpyyF6B7iLLusMhV
wuzhr/kGtuOH5GpD5Ua5EPwtRDxiXPO1pnKOsenlt/H6uJLnU7HRZSCDhcHbDDhMS7mEOhmeobYz
mdQgw/KaQqTyz2oc4KtVbon5xwBFiDlXrFeCjnRbU1vaZPNoKFdam3XdYeIJ2M+gve7N4yFamYwa
E3RlubKrA+I2Y5jXf1ksDkAvikJ7Wz5DuZPOEwrzi/FRvrXiUzLyL2E53mcch4Mlo2r3J+j7WovI
RlNrOwwn069CIrnHbBU//+EowdozDdoXWmpiJAZpQFVv7nJe6u6cqHoF7T5ZKbN7yuXwAn3iLHaJ
G0KbDV6Xf5wLrI8+62ppeJHeznxe9EY0gaG5XSlqEaueLqds266SZvnU+LJVUmIGzDKJ5bQlZa5l
wH+Vj3ZU7biGoiiIZYoPAPLpIAORQ8mdgF53dBMZNkfjqBR2bA1A+GpX86nYJNqXLOf4SbJ4uA4g
Fi7CUQsVW0yNr/F77I8gakbsbYYYli+7S5xiHV4981yTRKAer0o7RNUkLWlHNZ3ap74S2NY6+/EP
BZwDL5E62R1v0GCfwtstKZdtcJMZBf+A29P6HzkQeZY+x92zVtZGJ1XU7sGI92srK/7eJwSQs8IN
qO7KP36UkbeNa4tbT1NBm0HJihufA23Y7swezeYGupI25KmmZM1tl6OGje0A3K7AgTVaNZiGEe12
yUAqvwirHlgjZTgNoKDV0IEOR0x5GEr4wHMj35g8c+vgkCYdHJ++u0R916n715/3m6Tv7wiJRxop
FeHACAl2A3kQtDpldZsbQzYSMG2K0P7qGihSJfKEG9zyUFs/rFY0SfiOLQ4AZgoaHw95qFt+QTAC
lPMUUxavJH6xWYSCf6wFQT25wK1ITGNAWH0sgX8XPOMC1T/cmRWrwAsrzgjdXTmU87GyhQaZIcj/
ddifBcfR3bLIXjXj9gwRrFgu6y3/qtlychs2Np/wUTqGyYlqh+vzSWESIxw5CKQgPKaw44npI40P
e9qFacW/kqavhUGJtoBnrd9lL/QvO44ImJ6zCfB7KliuDkHG53RBnPTntLCNRBjkER3BCB0/wRWD
ED8qTp6f5zfIYwfY4Eu2amEMZyjpMI9WLnMPHOq5jb0VZjLs4a6tkhJTLG93jb4DB9eoAEe10Fu/
WwOuBycTQtjcv+RoGvpvo/2MEo23K6RP77T+Vn+GUcll/EN8s0Fcj3adFi0VMNQ0W3JJN6iipJ1w
9IL4u301yk/LPE8S8guT/lRYHTGQ5GGeWoCcAvy8GDLpHRDFNRrZPrPQ4XeSJ2dwUN6+8HeBvS5O
37ahgebwjTg9A2VIz6wwwYif7yp2dIyeLKL+y2+vX3dvHKQenqmgHgiHCPu0446ZE68PeVCIapMM
3SVNOpe+w9a3EeXP/QPne+0iHIvxa0Vtg2VHYKMHaRXfz0Qnrvy2tDvcoLsLA60EeSe7XVK8otvT
I5aIPlyy1hXfEaGUggb1IRydp+djvTG6IBuP8bf7tEn6XR2oNwokFEaGXxsNpaQLHKSoHAeK3BTs
nGdYAzj4W5S9m0nHV//ite+99Mpvvbr0aBVYAs1ssNwMSTarkIcSXv9DGro7nEZAucIoCOAbv7L4
mvwOsb7Tdy7h/3UzETlwMIdfc/xiu3Unso66rnAQSHxCxIrcaZdwgsFfV+ukG63TwxCfZLIwZu8C
Bb7/6543C83T9/QphLZ2B0PhYL01wXs66GLeYgGj1uqujISFNGjRd/FjfUrsrcYJYMl4QHlYhdwm
w+MlIGEotTNcdqLftLFgcI7fazi953NA1Hk+WZBj72jMmVGa+NRNnSqccYg77QqJ9IouBwiqm8HI
dzENHLiICuu8tpyUzYtKUv+ccXzGlQeIaRvb5P7k8mM1e/oT2lIdVJDsRFAaItSxnnros91GPQpA
a2LC9ITEyfUGyaUc7PqDTvPcJ31TqzDt6l/EBtUqu8sf5E+q8IMXzc6bVSCvJENOlDJ6X9JD1bV4
pP2miB16FmP28Shlq9+V4/svWPG3b9NEX6uvi1ExsGC241t8REsy6AsjxlWk4aC2zpEb3o4NtVZf
jI0Pr5eGcq0qpDz6tQAcEs5nK7UHhIhZvl9xDs7pKkDThOMQTJOOb9XgnWrbEWdcHeDFx4LNxeKb
XFIoUnCuSfR5QVq9MSHnrIFrsqaDG7Mt78/+sD1HvKBSCjMr4O2e4Q9b1N9tLokb8BiiSsRcOUOM
wsoXZ0iZMeLq5kMcSYaOUaIlz25RZTJl0eaIy8SnrRlPH/eN62cJK/lWzdoS1Xyak5puYjwlX4RU
c8lAjJnFzUHmqJWq8cpuM5qcWgq9Sfr9tVoVgVwSy5dZBuleMpMRq69fW9PAnPUjOdPwo5klPRuf
5BAFatkeIEYgM/vPhkXJqPPHPaQKGpnfpF4kxK699tqLvzYDWR6pHvzXuRKuuVEfiTNyAndUUUWK
C7iVbnY6NmlKT2pN0IbrFxynQtbc6ZQgZuF1XpU9R9rqnY7+LiF/5gDK5c6u2C452VrH4ypuDO8l
LNcWKVVtogz/5m4B2Zw3l7ZCqTjdUGYtnw0fq/dD3iVTEjiqqNLsjgzoLYMS+s5sY2s4NDlnly24
YrO6L9AmA9j95MFVWkyzlQ0YvdAR+6U7PPwKXuQC1rgHoi6VApnsDt96tXLLOloCq8xF5vu8sS3b
LZbUTuDuIcwSSZ6A5NN2tB1oOxdqzIVUwrFyQr/uUwT3ndTz77jbzYt63PJRNNjzgmkH4IaA4eM2
lMhMf1namm72C9j+t6M8bnlhHI4BjnmU3Ko+S1u+wKYSVCBxraGf56WkudFbMIS4sSOgrsOt3kGd
KCzPM/nyaHJPMwUCL7mCm9JV28olaYcfIPnF8+0+WlvfFxp9PDK7Jka7wlEXZZt/tY/B4+J7onHo
Ig34ZuAs6pLSggfjrA6AFXyGLNC6Ys8Qcqs8UGjWKfAqn7fdFKY+Uci73tjyai/3zxXYx2fjge6+
s8DsEeWoO6pqikKM4nn15mx0cve3MbVy5bAcNB5f9iT4TJXKvqgtkw0ze1L31jfuLCv3EMlajU5M
r8y67Blo3XmEqGhD9LcY6fTjH2YGe0ewh/NvkApgL64QvUPCsT++N9rCorPJLkav/5TbaLBE4hBL
drK8lQnkVvzfgBEAmGVBjKux9SYM18LRtr5FmAFW6c+Vx2A4tX2eAvYoFvhSq3fLLtpQ8b4J459/
wlHC/WiVxby8pBVoJ8oAdfAAZOVsNi91QHb3tof7aZ/ZCHJZJwmInubMAkTtNaazAESMKOysWfXN
J86PEQHOtuoJ2jmSX93MaUHBI6hZfAnV8WJQnSrMbseGetblz3QtANh/7IyJ5U/dfQ1QWkBEjHcG
yjhjpQ2J3DvDdASxTMC6t3y7lQ0eD9cZ1lfKtdTam3vkJUHph8jZESYwK5gMny/yutFEF1Nh7vj1
hF3ICbLkF37zlYt3RDIEILiWMqlvUKeCPMAPJVgMXcfPjoF4Bf5iBO9LUQji4G4K5F6tdjxuGzwF
ZQXY4YecTm6Upol587HQkNrb8CnRk2yYJ0DJZ3apfwH6HfR+3/V93oX+VF038rIZNuuT7Houuejh
h6pFGDG9oZ3I0P3e4DM1/2swDtXsDxzS6yZMaVL8cyhZfBl1cyC74NRz7CVfuylxGTjG1NBnhNbA
NNGTJI5/VwA33ekTQAK4SPtRZxZ33hwNwSUaH7tUurPQRxKMGAt1/kySfcEMMFtZArvPNU/zHG/P
k+O/ocvA927qUYfDPWqIr2slk8OOmY6RHDcy+GQrJ4XR8Zg23k6sRVDwiPJJG4e3unRuk/JZF9t+
twJB/connR9GVkBCbnU9wIoLEivDqTFAhA4QWwDSMB4HFZLVIEPi0yJuTjF0Ay4PC/IBVI1bt7pI
pSwXM4bZBom9YAUzzlFvl7d8f7TaPqdzArXci4oUyP+NkJnMMkcY1LfX5OKajXWJKHh+4yiCbvbg
hoEwg8Y+8BUy/y4tpZKaQaPUNZVDQNF/Nn+RlFSOCSw4ZnAcYI+S34hbZlzuX/05BH5LYRdVBp4T
7D/dE/G7jbtnN0Rr5Z7NoefbVWPntEXN6HKytXlhVy/xvwYkdctLbAwSzZlTkQoTqXx0PD2MPTYl
zYZg7YpO5FMoMM61eRK5TotnFDQG1wGmPbymOlSm4a1tIFkJlUSoFAqiFTR+Q0R0B1VzbEeP8f+G
lv2uXYxWVaiq4Qxzr0F08KJR1PUEzmlfjwLg1KRnNRMBDZTHGof7CYlot22EgChoajJvGqwg7ECr
5dMDerIviYWBsPSGwQ5EWdX3ICJbbdWCP0i49BVERV51a1ohpr7+LKX7A1pGMaYO1c9e7lmL79ZQ
UHOHNnr073eUZ/siFBpEC5417aVbfM/i278d+bjdLx9uosuK6REQlS0T7p9bmEbNob3249GPLs39
0WDBVITxhYzGQu9aLMokqbTZPq9sXgncpdzLkBJs5gcqsnk9kjlFo4TFYr3pbPbfOBuDpvpcSyIG
t3qanc2sGL7kduvDaEPy97Wzm+6PZw4gnYwOt7H+nisULnIxR6r3OcYUNOVNtB+udfN/vZczPJI8
PvWPpS8a5TlH8Y6liUApfFKJbzDaiyypS/89TmFIaOa5WcZdfFx4v4jgX6UVSITQI3wCXufOAR0P
DMRjuo00BO8hBH+Kf7dPCSN25JubbHckTy+nCsTkLx3W1ekMgCZHamsk5YE7Baq2jyMzR1hGWM4t
duFPLQy8UIkA8XHcmBaI5Ep0SsaK0pa3d1qRPZbIuTIJR9DPoueTIZUDhG7jplKqIwi98UcokV7r
bPgfxAbOlSmrrlq33qG3SfpRpWUKWFP0oy4c4Qwm0oZxwvWVYuQDD1vMzKNp5vBaXzA1XepPv5bQ
WZza6S74d0tfGkiOZNvC31mlGVc9LeL0QOvlMGVrhdEQMI1B6iYLTOKXBsur47Fm6qS8Mo0gWNPN
iBJiuhojrFXlX0fSMedJeJ5M5amQsddRaIDq2Nvfc/Wucv2LnLmLQBmzG67WVxAK8dvELmUGHK31
sVO8TzkYcOHEybVwiifL16FlaRYXyZOk1mvdL/4QX4ECqlHkSTu3LnFLVFqW/dVZRffwAKad5KJ1
KkhO3spvQxgxyNJivN0k/HMXDg7X8Yxqh9EkfEYHxKQhaUyFDT86muEceNegJVhqkz+aZc28oCDv
f8PDeE4RJCyK8oLk+98BhMiDfLAUP74e4xN9WnjseNU8GkJJrAEhaogrwOikxguM9hZ3kwsJMSJM
Niss7TTrmKkW5uLxIvyFHeRFA4+MglDXSRtzKj7B1yp3irUxL4mfGiyZDMgd6lfStUAwkhJLtVWV
MsGXphU2KnYkCtU8WT6u8l92LPk3f69uQDcObvpL+EPj439b3Xi/R8nDMaWj0kcEzlCAy2Mk+x4E
0yVkokRshNDaJG6vtT17PeX/zO0jKP3gOlVZQOTJx1M3kNwM6hN+WkoQ9XpoKPjwGT7myUu9ShTN
W0TUiK/o4a9smwAufK+cFtw6WO13wElYwq3A1HrSfWvK5tEptgLIVajP/hWJFAgWEx3xVBMOm2FX
XB5MbLSj6mGaHs/MIUT3vPP1PfJtZ4KvbGbBv9XvUPEKcn6DTkWF9/5caJSIa6N7fW4FczMDY61S
eh/Z01N6EcI046g48/JyYi5UaQBvwk2baIcP2HRS/RZ4giiZ1UvKblo01hnwxtNmY/I8YBQKQhg+
X1wEafulhZmjyZGoEUxesotVsVvCpznjlxQS7kVG59pjXom+YpIWu8G3NzHmhbtBVHrHq7M/LJ92
k4+uubbVuZn3vprnNJLXRUC7mvPD8Y1pcvw1WwLAqGcsVv/7F+E8N4oVYtv0FmR219vGMYFsxnGv
UvUV2/AJ6OdGaa8pdLtOIOgvjRMrvZqSBIkRSiIRXGqQnPkyzRwpUBj4m2zIi1bMLQRJ+/UN1a6O
uPEVR1vwn4zQLD5kNyFf9791McbY32+au6WAqy/axnOqYQIzDG1ZJZa2v+eYlyCIfJQUwqpBnfQA
LqJzzUKA5gpvW1WlPy9fOmt+2gsCLrG1APp3g1qJVw4DBCIExi40i5CWT3SJukGjkT0X1GV+X7zX
b8ntVCBXXBFlgXjHFJ0P6NjQvlt/iHz0W0Hoid+07iohbn8hAxDQyZti7QoiPfYfTJCR2LdFQIC2
Mq+vyXl/4Iq+1UoyAyUh53Y4WCpt2gIbPc9WNZ50ZQUQLadSO9v+dtBvMhfzf+0igNV0OJavOpwE
SjnqGI+mwaHe1J1/Wt0pdVnTwYSti0eM3iphnG/mWalm3ZY123Ldywa4nGwJm1IcKLs4YPhj578s
4U8ZkwEFrYmNGBhbGvvCqWJpmpkc9yTYXh27BQEyQQosQdKy0FM0b3MiFGXIceZNiqStU3dFh0hI
F9bITwcwM+cTFwWVfmELBrWC4U0kvzcw4OTDa8MBD82+lNN1AH3wgKvLFZ9cXKNv7m8t6SJTl3Y4
Jd6euyLoJTR7hE5sO0AafcVR6pxMbJKMESLZ+lfhjgJl7EbqW2R59SgDrFlm+CqPobHETDPEOIgK
wClBwoFhIIKy6Mc1X2eXMLe3b5DUymnDUrMV1+Kd5ei9AiWJslNW1rop8Ikv7TNtv2DJFP6tg5dh
2uvTBp1tcoNVYoXrd9laCv5y62DggragBzOfnF2zMSJjXUiiQncm3nzQBl8dHaTr1Ll4rMQSvCrj
SfBQi2V64j/iYwAR23Vep1SQHjpaVn9giesTGP1/lzow1r85/vgIwap9xTxlTJn3nYxlDw1KT9YH
P/r37HGf44wEbUxcjXOAb6Jeon2Bhs7Tsgz47d3BehutcdrLS09FrisDCjK6ECIa7tcMbcMW6wsC
f3mjyTP2F/t8wf3tuOxDZbAgD7QO5kaslBq+rwkEWKxWpAK25nTCkklaoFB2U4gkZhajrcjqWJcC
Ce1cSDu4jkABqsY6joAZC1dOLmBwltv/aXSUcnT48kIUiWPYtVDUbKIU2W5X2bjCa1zBssmnrT9+
2cmwsDfwzWSiUDBZ4llw0SSDIBG2bVSxjo5Q1kD5IF9eREMpIx8xekR3M5gjXMGpF2TfrnjdlGGW
hBKvaDe2GtAk3OMfg9gJV19CaX6ObMHbg4byHxa0yjyZOL7AgCzYS3IsmcSI9KnUE80TBuSHDxIc
o1HfZIs3cwJlsiPeU83FPwWPboddtZDHOj96ymwgL0g6XaoaqT8NJ4WAWaLodNYqbE52IUzoKYId
IukAZXaJ3AxvvsTSBXy7TYpK+TBsMbwzitlpjShRYVZPvCHD6KTLy8dAEmwukJtx7iPNPY2amxlo
A8xCmg0Iz0R+yuWGBQJFWxTcGkEo4rHfZpTtPT95uh0eZYczs3zDF6NlExN+eEP2VZ+AJre7LuMq
Ij5aiu286J8NQcpyZY19rb5JryI2++XcLwEn+p+KKVPzo2jEBS9A4p3AcM37985guF4ETS0J6vbz
5I+040BewW+03e+0emT4991QhGCZAKR6WwX0IjlAf1T0UO5p+zEa660mceW13i7WZlrUxXOFCB+f
SGc3x0taAcf6rOE7OTeL2VWyKwqNi/Vh6kcHNZJzkhMcSdyxF/lnPJ0ubmHRf6BDwDPvAxI70Gpj
PiW/PDQif/WPrsfX1mdKTtR1W3OXQVUxo9qNF91Wq8FmXY09x/F7va1BRul4t0LYloaoXkp+uCFZ
Y/RNJLXnTVGqUg0loZdktez6YQ5tfX5NCYqDDWTg9q/GB3uCPOqVB1v6znjEKRef/OXSUIfBSTTv
T4rwYu8V1SeGFjoU3scn/RD0tIC4ys9RaHPRH46etZxtpkoH7sCsgyC8w4LtLkei2HqdE7befX0J
bvUSyHAW6u29z63BSXqjJSi1FrbvOWDa8Ux8Q1MimwiqhxkG72So7aQaxBdnMWh+zh6O4RzrDRgo
nhctLd9rWM8Cz/92Nn+E4+sXw0gJN/BhrXpzvN2EQ5vEXFAusgfSEALyYP+NPbObEtrif0moeX9T
Nhrcr0J8/rE2GyzgeLi5Pc6LCcT1+Q1w+f9vVqrT1kDE5JLIR7b5yslw+VDy+R9tJdH/KieK2CBB
WxgxBIqchQ4kOJvDUC0KjOSHUO9cn3nZSXyttZ5MTlpOTXX8BQ8hcUollqBbkWuDqSgs/BJPThq4
rvfaX2jF5/9y6NL3mWBqTyqMdmtn3MYJPoDY2pQlfCHhvg+b/zKckh66cKkEgBn27mWpA6a5bLLo
bAh5Lmb6d18IMUqGXq/0pOX35zCf0rZUvnUI8bQn16/RTzIt0ysDQWFI7S3iBikt/Mek/BYFUq0o
l2SdYpLpe/SkbcCQrOcR/Yf9b0FHpR3xc7PAxTG5jei4/B4vrDSYdO902MgmtbhhqzhaGMfRkZG3
yY4TkaPWN8GcGRDzzhrozTbCbgCDEbjjGBAq3XdggV1hSc27XjDtivwU+PJcwTtgCMi3PtyuE+M+
eDT05lc5pYDrDIVrPvcKpTwMGYuaLM+pU72DZ/GaoLHRVsbZ1+ryPTi1eWEOcuCKDojABPByFPew
72T/VWC3jkUQzCmQMeUAMrh/G7aBlCxWRD8cSkFr1Au/x4BM0pgUIbLajhBa+gf1hPvxZFglk4Wx
su1sD76LXcdAfSoMU53EbBYVOXnxnR8e1dljfmyAmakgtHaCc/hnQlafLrbFJsmnp7PeEe0R3+la
X+JpXniEvkQDnVTGHgjiBqVGJ4hZ3DfGGI8rLTfF2O5SyxNtvAgHZ1SDNJGSuGld8GLRyVNj9EbL
D5UGryqgTFVxMFhiiaGl3NPaXDT9RefeX1XySf/CCX+vwnXw80J9j+QUtK68SOINhWCFmTp63+dw
l/WfbDqK6c5qfd3kdYJg6asKc3L9wAQzgiaxUoMwPMcFrEtL0yx8NS0Ab2WDtXsHO6SojRAHzSdd
vgPq5lAz4TRxsFZOikhmGtHRyPcgO4SD54JnhMcRIwKWZUHWAEQRJZyYDWkNVo3Oqr4lJH/Gqs26
CLoAWIMHxf7aGPAK97J5nwruiCGYOMwGZQe/p5uwo1tY3CxYbWomCMiTcFb5vZfcNWSVZol93oEL
u4bCU+42ZDWyA0N0oYt28sufcoBhfSJKc+eiN/FrC1rzQlE89iQMlX+brulkRLcqR4iU85vBXBgG
CtoDivNWNDnMNl0r+s9ptx5MgRlovRatTFj4gegKl9JWfNKH6weJBPJn7d62kpjy2DPUclxnRf8p
ALrMi5DqjHXY8VE2e28J9XLD3JIy/3ttaG8IpxhwEjdCpfH1MQZf8DyoRmO3Dx4HJE2icQA6UEJj
Zvw+cM9JKVw6Y/rBScFrg3zltUs4CjJ8Kyf1ZigzesMTxbcYeetPvzguuZDIA06mVcs6L5W7Cwyk
qI2GHxsUtXCiCWH9gVJGYtsLFrnHsSctuU1iz3VjKV28C1x1hTBedLeGlACY+shPrMwIbNiL9RPC
L+vDtWoTJpEKuCFp7Oh2iTNqnOlD/Vs0yvn75X/Y49Fx8mvbYTi0vCqdpIV6xrzPbJ3zsxZVWIoh
dtYJZo6Zla9tGYW/T379rqlYR1euvv7gRKKUp5FhUFZhn+8vpuzYPclSyE5hgwAU/8HtTure9SVY
eHDnkvyAbQkAOiO8lseYsrN5M3TphLAMazgS7EDv4EODUdePH2se7yooRsYK7hk1IGHmDKHxEIN3
FT/bFCDWw3I7pa4ELR5H8XW18OiZDzI/qY+NA8N7T6u+nRxd8Ny4sfxyNNGnNdhcMlX7bmzgfpaw
I14Xz+ELnKWy8zPDsnGNaNDQLO4jqpW9Tdht4IyOLmj7pZjGFgi/FskzrSZsC7xrCb3xHOyGlpdd
UNBCvk4HTwo2eXwa/VCcd4bXQJ5clXS/U253nrgCoNpF7Q2YAMA7UgxB9qdCHsQJXOkAP7Kj2Q2N
bAS0QPR+dZpt7H4aqMTTyPL9IjS6CW2LFeqRDZ07LF2l5XMgdItsIW3k4xTcdLgCRBIzaDNHzXk9
Dh38n/ppSs4uXP++qbsftRViOku16K0NM0SEuCBZNvbzgUTLMOJTPIdlnmnD5ebQVpzoeyHsXhJZ
oGYH0oz8zZYYzYsXOeJqkbIuaxygZnRkBb4Xcw9eFhMMNJ1dJwTst3oMIKlmEnUvnbIdJ8kObeXS
GV02SiVuZdGMPxbqnMvrYbKPvD3x3EzWeWHOjvvtOsAiFpTvJk4p5M12FovE9lOtTZrxB8qy1Jzq
Jym+9MPKeuof/rJnwhsuX/DIfMJSDbRrAnsWCxZ1HXKV5qyTQOrdRhGdImg1+OzGxEPRdzqv64RZ
KGuIXoKRYuRITTtUHcdRyl8g4MF3elQUQuUBxsWPBge3zfmDzoaYixOTRXT7Q6jNVY4HCqQsUI3F
1+LcFUCyYRCv4fhMI3tKAfr+37B/NsBDY859LcBo9BoKvvY9wzIH5E6XZKSB0rqgGO4dDNgHdWjG
RbOxRsb9wEnaNX2ZmH3SIVB4oZnyEVlJnuuieuEezDfz6KCkN6LN04IGfZbwpOKA2JRvUGOW71oF
Kq4UtRimdVaJ53w62fCgKNxKFzq7OF9UOq++8uFEPX5ZdIB0xVqA3j/091zc4LQ/Tf0qiPhPck7Z
7DSwRFJT9FP/uJII274J/ec0MJ9gYk/8KSkllj2RbjlV7WF72wMF34aTv9hFVTDi9lF0FQgxnOdF
sTITQaM+wTkqRrv+El1cUCLXtUYJHaEwHfzwtJtP3es29/uHTLwA51XS8XLG69VyhZuONYCfwj25
stsyDPD9fivrLTT2ZahRWjF98DPU3Tj4Rs4v5rf2po8zUsSNyaim4qJTUPMQ/PcMNNBJvQ68PrNm
TlnXS7YnVEZCpUlmzmEE9mNiD6JjJiIq6t09oCsC4kd2ZguidHMdC3lNMDCyvvfLim2JT6hoWZtm
vyJIq/jyxW3Yi1Wj7a1iuYjCwDQI1WSXaFmsIc4NunzX24KKfuvugxNuFeGGqngf+kfG1IBlcChz
/2KjowiDkhEeBKv3Cw8hlX8cgOXgOt+wjZvgVWeGsZIAdZUajJf8MJwMEp/9IuTdyxMcWoTMejoz
7dcilLCJl5femc86MBMsBn9MLoPArqOcW8nBQNWKyTiBY5FnNM127m0e1AqYb9wP8hZbAkDTDohW
qjKEp21twY8gz61iiYvFajxV2TlHdkDnZJCoLINYQddkYwsBYwVWATew7sHERuF1LMB7ERywpZTg
JLNcJaoGj2wDbgXGtQOoFlXmlXlXxpAjA1in/9b7RimudfxVfFIHlPzrAHWmW2hdwteU0YBilIQs
VytHtO3URVh8ROAYVsWB7cZhXkIrYkChM34VCwyg6UK1KizpcDyklhz8TPwiMG/jpIGE+44/X9nv
HIrrSmZhWIVXsJ+YWk6FpYOlNqO962Q8k7JgAlDij+m4r/VYuz7XzQRuSaQ8BtVflCLPVAa5rzWD
leCNYlGHCtEbej26pxihNrwxc0uCLC1RKRPNtq7VI/IWpMjeobAQj0vs//XHMTWmLSOY99gAthHD
sbrEfNEhnZTPJ3MXg8208Ym4NMdXo0tlnCAuvr/bqiGVcnwfagquFXItJDupY+CXb72Lp6xn1mL4
15xtyJqIKQ4zGKF1OL3BN6qtm3YoVZhh1aGuhv2lajveOwZ5PcnAifYC/iTpKbrR1nMu9zI3Mgew
rkuZ3tZ7qTn5hk5defHBvbwSdQQpDd6qQygq+LhdSGnQnbSVcA+iflMki9hZqWDVDPJNAxq2J1Rh
h8G48dsDKA05lXm3oyVCQIqA5/uC6vy8tx6dyicDlUcx9N9ejGHBqjBtguyxgi1I9MUwo/lABgom
iTnwwZ5Fj2Pqf/2mZ0IRKtusOO7nbrKMZFXUFbG14vwDwSv4lh2vQc+3EG1vnfIvdFWAspIKMxj5
LbieFUQNmLOFIjNOVhOEx/Bw9I/bAAm4ep2gqbdbT+qGSoalnmhRYFtI9du8lTuBF1Z01DRE+rCw
16NJpARe4pgxoks7y9dyV4QDFYV2PbC4q3bvZJIKnNiun7HYUEUwrlx1HeO4XTKXDdYv0+Ww18x1
/WiN+GMR/a1Nvp5iG9YOqHEXjRjVc7O5QUq+AK1HUwplHFrK3Mk3sKUpksgzW2H8iTsKKOXDK9XP
aTF8T+W113REhBO0JHT8DoUi8IZvNZOylY5uPmO9bfYwQUcXlSIzq2EbeBu6EN6XyrKSWI+1skCO
KOdz9OPmPatyKyfj7FVavjLu8IAbja6zjeh7GJGxKVc+zSuj9ozQFfhtleHfRt5gFdiI2ubpI1my
3liuSEuHZfq4wGzCqlv3ZaNWWZ2kY7kek2tOYlHx4AD9vFKMyWS8Bihdp8lGM2lrLWqD2MNm0Q+6
bSZ/tBrbFOFfPj8jRWBWJtVmtb9vqbL7BShvP0egYD1uCKxl+kFZ5waBl8vLnf0nqTiE5fSFps+I
5wBw0w4xdh/qCyCyLVqv05/NZavkyF4r2lt6OqttLaruEPbw6wrA9hX9RIsSlQcOD0/MLLcDO7ej
INMDGxlNlAs4r+imyq8frhPx1XjC36hFXecosaXb3705GKeRSFVH5fuytFOTaJUrOAPKZFCU2wB9
YDWLpsmJZw0YvpB/4cWz1JY70na0gCUOEKGTQM+Ozbr4j95Wkar2ELCMFSADEwIfnaXZGE5PHpoH
t9wkc7+TSyAll7UXowS8WOOZNCYO5icnwVVocc0FqU4fRpvMzDzMKHVkii2CcRGxly3jhaHThj0k
XkaiLmRlnsiZZ0eQpLgxdzwSEpW50WZZzCRsuSh9kg+Q/Hx1NnRJLhrfoHhd3dTpaDVSGB7RiC91
ID0LMzHWSa9nCWqWAolc2pTS1eD61ASmaImvfmNYLlonVq/WivQ3FmPBRcfwTpWgIgH98iSuv/bB
KyQ4Tt4ET6EPHnCtKqGJMciEqOe7yX1qoDkz3jlf4MIpjy1FRPWGdKXQ6oFFtz5W/7WpVCXBPCG5
tux92pxcKcCqovaxxUn38q6TLk2CTZODj2sOKqpA1CMOYw1mqgt075U8pBZJwRE/ABL+5sayX/U4
WLnRHLUg0nobTJ/y8udQdzqktobQn83A/lCSR2cFEG5x0XhH3RUuUyQToINiFwEM8DHvYp3MkltW
+YY4DSRl/SffeHg4y/GfNcNhj++fWrHV/NGPdBafvWy8dVA0clNrVTmsgCzick+SIrmBeXStk5Y5
V9YYKfmc8ZIGu5bjpbQup8saM6MXWWM6KpNo9Dkkr3yGUU+V7tG6f9+sFg5gwJpnaXesxf621nz5
d/yhaMYr2woG83xRX0JyoJi3xdXHLredYg5Kvcaie8JJglr5ss78krU87Dq+ydpLP2N9ZWd/4iwy
eqepCwacCY/2yFSDu2Zi6bGIDGjUxIhwHqJuCApEL2TXAg522Ld1+sAfLFWVfjQlufWMy3fOM6JJ
/wz+wSjRvVD5HxZHclwlHb+/Ia0FpUx61dNMZKhKGNfmAvNm/HVcCCZ1iZFMfnBg7rS5mwOgzC/0
ycxt3W6j3KT5NuUO7vBbKtGukOjAKlNr7Im05XDt4sf2n6wDCMexezMda5hHC0BbCaZb9bIeCqFD
CesbPh3vihjZrAtjYiEcJsUz4JWQ9G3TA6t6+0y78keaw+ftLoSRZRj72hJsaoUa4wejFfQ716qC
Xe8nAWnzvPvG8MwacL4HR+TGMCZ/RZnyykoNhN7IIy7BNGL5tqka04PynGclo7ySKLkysha+jWQd
/Ks4TTOADZ+O2dbVAJXoVyCgggePaw8V3M3abkjgcgALit/rWwkPZVG+7LoxdHg70+V9r5bl1t2w
jIXB5Xr8EMDd0zKTQcwDuCtMkOa9T1VHYmwY6iPaHmRinHyeRQz1fLXfuHnEzvDYmTk1k7QWmhZU
ftzImvJ9IVbHI+eB0oysYbmuGN1DptlMZCdv0G7y6xYXtHdFrtUdOipiRF46whvfPufx/Agi0Osq
XHNuVzDszBgzD76wxU5gBiMfjteVSevZP+CLYm3sKud5+3kbR+s54xN3YFlGCbaGOeDl6Bx0KWaT
n0XyhCAM9XK49iQZveRfzB3wjqB5rjlXifhqy6VuWEbE/4OtAUI9UZM0pGXknQQnf9jBs3CBNyxa
5XHMgm//EacDYLKP4IwZIHg2vABKFcuG/kP+WH/GCfKN23YTTBncZEvb30vGy8ZBI/afHRILz/Sv
IZFLXwsxh8IpaxhogmdQtL2vnuJM4X5uDcstq60EzqKgc1LHFQQlxMQNXyFoi5nms1o+/IoROlwW
DfMEBQxc3j1gJEZGRVLOHwsK+UfNNr7eyKaQGOMV2BSRHSr3vUBvsoIG9RoyifRmX3gzPMxWuibI
5MhpB3x9c/aFrvUCFLP3MCA1oArbK8/H2CHBbRvUBJHc7mVyZqG2gvdTREbRoP0iEqXKf0+Gq3Vm
wXxA+Dz3e3Agw08zGtZIXUw5rqTWGqOz+8xHU/ZoYQu2jJJinynG4m3PRCEkDzSx4N1/zXvXKgbp
QWjE+92rsbT8JerBqXV5GK01ccuv1uaXDj2MfOjdHtxUoeQIREzBq0S7voHLtY2gB0ASO5mvrwrh
BPGH6IIfzyBI/W8ish4srrC9XnBscv96RUxujqzDh5h3MxG4cJdMgkDW1nlB1OyvsMSV/2br0VK1
aY8Epok9mD4155VOMYA68rT9PPi+AKZMmn6h4r/awAKNUzjFmRjeoU8+ODFX1BAfBsN1AspjRQnT
CYvV0Vdh7qjLfjTZ5hCoUnNwrRU6xUbT1jRI/RusQf7i3q33TPhOadcZ/86iyo5qwthDrGQb20gw
uvX+AcFLXPdsk5pNgHlolkuYIXo+RK1+ytNOsnZkYTlAVq2TguuO8Q80UrzgWDPTVAuFeVd81a+n
OllXBkMHTf5ng6Duta5oijWnxKgMQBUr/mPeAi+6gP9CJf5r1qoCaTr4GDUSGu5Uq0oMal7Pnapr
rJDbMjJYrWP4CfhoSPckEm+rRlkERz1/98It50ckhwUQHvTc3JmDwnoa7IUVa1aNtQQVnKblaGoa
j50I0UUY5lt6pyiy6CYfNdnLq1hjrmf7CkDwsR9/ljMD/Tv0b6jwri4HZi+vkkX0GueQHAzUgtp9
/HclbGAzIiF0jRsFQOY4Qgta2V1p/pBtAsRqhTsHMMz/jjsBJ0gtYMHZ4ePkVxLSqoXsE3fy075Y
xN3nhrSJgHHY6oNw3m38AHMRhU9IpixrpGWbhREiuKrs/LlBe8YF/M/UTTPV0PPynHIDnIVipz5Y
Z5K12W/mYf0blRwTcuxEx75V2SzwMYfuENBHazuyE4xDgeUIcvUTQB3ZdL8WotkIyqZhEJG4OPfL
bGuNoRGsoZ8eAOOCEvvrusgEJd149WRjHaH78eSLNjyl/hMwDFfVywfFLYNWfPzX9y3WYYO5gmSF
BIkI79W4e4zqrGnPUHbcfKumKrw09BAEzy3EAGLM1kD+7stayho4TiE3DHBB48eayGRxKwYBgAN3
PUkeM5vvpeKosv0XKz/bITNcbCHpNE+lhJovd5LXGSzyhf8XyqnSaOUAVm9hTAybIgWKN0NnaDez
qKSdA20Mms4tUOzMnLXBIzNYsYufqyrC9FdgP1NSY1H7RnCyOuj5ndfeyreN7wS5bKrSCyz6egaF
9XvZmSgJ+dChs3rtVPACuKq3V+sO2h1d2QckvO6K+UAoCFHnEsK1ZZGkq8Xjg3O+877TBtMh+FHC
YwD8Wa25DhgFNYZzEq34m1hXQJfYh9HDAjeVvp8AC2NTQ1bmlEwVjpwXhZTXWWxlTb1hNRVXDRkh
DCIn/wYIbZgQcOjjavvKvbp10mGFjvXI/tmGN0DX6+WPeF93NhCCkEshDSJHJJGmI/cDCGWb4YB/
bUYZcma719wTr57DdajAQwufrtVkm29flwLh8d2suIme22f1zHhdbjgphFhYDEtj6v1vbkmGXmhZ
ZPpENXG/AI8q5foJkpuIrUabN1xy3Qj9euEmnPXfFuEGeQysjiO+1hkqDVMubyA9X/8aFgZ91DfE
mPExLlxrBFki40kxC9Fl+edXib0IgDlW+gpZFp8ACq2Gvz/9p/WK88wlLpZvLoi/jLj3MIEAr+uM
mGwzSO3DJtmpnJnKgkZn5eOHb59FjIlhutTqMvSE4ZBcuITxkq+/sH9ZRcRZTlPTDv365QBCCT5D
bOdF7u0PjXFA7YIKXbsul2R7RS7IX9Gifk8gScEegUi7GULUswXTYPsFQ3BeC+fH+awbt2MiMCGL
ZVUGz84tOFbUVKzGGEzuluhI1vZ1b8JyTJ+Kw4J+4ZHCYAxkDjf8f4ovhH5JMFE4OjA4296lgfBO
Y+5ljuhDTyWN3fpOKxDK7W0WMd6pE7rIy4zv/mExa+zffybgsnGhqNvywWGFhzORJCpusrT6/6Ao
MekiTBUyJIaFds5IdldN/M4Noe44e0NgEt6Mh7GAiSa7X4baablxN9P1idBiK4d1nyPs1AhmRX/u
wm1afMK1llM4X37Wowc7eeRMPgwbxNbgOWeejP5I1MeC5eHCfBvgofPp9pFvGDUwCDihQsMHyaR3
Z2e6swBTL2XU5ysPhown1BS2iaWKBxxfVoVszN7MEJgNnSanksbxkRrB5LX3w4Hz4+4WiNm9Us64
v8sXd2W4JI6WkLb2l/nmVa12ZeW6npuYjlZigxPvw8DWGejd8YAkGi+di5Lob2eLciA26T2MTia4
UlooxJdU0d8h4RQUySeknqzz0DoC6EA+53OTE1lXY1vE1IrDn5VTIp3zEVFLd88N5q3yPSxP5L+L
H9RSSZVgqq6thYlOetKtYOO7qkVECfpSwYkCgTEvEowujSUEl2DrZrnD6CwwTPA0iuVsm4M/9D8f
miSEjNOgyIm3OF5raHBWg/J4ZW8r5/akpt0f8AamKS4MyBSBWg6Zh8trpbNXYHtRaimtJfEc8CYp
iXyBrsqnStO0f5a4la/l/z6omDmVsYAsqpZ+LFHhJdX0Q+F+OjFU+yyCnHWGyNb7MKCgWlEV25jH
y+/OPvMOMeDkMofuw01N+R7lXxcQmVL6+cQGjAZOl2SwHsSGiOrZXJTBXr9LOj858R8MF8NeU5F0
DwcFqKnDz4zi6H+5N9Sqb3c4AmcJifAzchIyN5lGkQEdHrW2qpavaclNi/yM4VdKNbLd+Mp3vcv6
u4FJEAi+4S+RcHRResB7FEhiOR7G4e7TN695oA43AqA2VupNRUxeYhKpPdk6HyoIToEw1ifbs9/s
Lo9yXAuQam8kZ5ES9GNmAJNwZEER+ZUsUoRlFg57E6BhAUAyWPJ8QjZshaaN2D0eX+959S1sMBbn
tUPXNepcaDTimhQ2FFmtmErsFIXcy04pDITtv41skHWEUsSdOh3lUflzx6sreWHccrj4aK2v5NsS
yYeC61RSK+mgvbCVctAuUiJnq7EdEK5xUUTFfMj6bx/koLO4IHSV3O4keStbgIQ48U7UdOHtG0DS
j6XeF4JHjuv6Du73QvySo8v/iD+rVEeZCHVUr7BriREVbJj5Ldu7s6/5mu5NeSCVptkLir0Ax8tG
2Qt0BWn/6kS5fNDvekCBfJcvs9kE5V6eQrG0rBNbFuvMef432zAQ5hh7RydgrNP6tt7TK2M/10wK
lSNxi3f/ZnzpF5QtM29RSofTCS8IvRIAhxdP5SyGtA6ZJ/Ns41Y7TNlQotIPswj8nFypOIs6ouqd
zoA4sQ29z2kOg8fYi7XMdMGstRGr5D4jh0qBL6ulmh/qSnavpASXjrZ1N7mfY2S803gR21EabCWe
Tsd+HXV3t1keTxIDd7UXGPU4zjH1AXu1olMoXV9ENgfWo9XEpj0YXJDEUvzBc4r9w7QIQJxKU28t
DEYDZeMt9BdyBomD37oBrhuceS/428vfBwt5VTEN3TK5N3Ol/l9lUQzeHjMpCJUBhTaA7+Whv0Lm
LRn2r4/KzgN2x2VM2nEr7/2+j+o1E+Abw0mCwXwsPEVo1LbAo5wJUr34CBY1OW7dtZjFYwh2ICgf
Z+Il66IWTwQCN8SpRLYkQ3KGz0PmqHzZiQf8SI+FOxj5RLczefJPNfFwnpNjH4a4D5CCuaMrjdXE
IFKgL0PQfMdpsCWHTFN9QOFFeDtJ/xR+p2BujStTqGWe88AfyY2tsrAq9jqjVdz5dHn/zsJl3XOI
ySs4sBcb64riuTBr2xtjR0E4R4hgAoK0UsT+Pyi/yluHXplSsWne+iMCo2gpCLtcH8ik7YncyFEn
RhDbFA2oO9nzn9zkowXELNngm0BX6lV1IEgctCqTpX8T4x+mfh0bwY1tF/QU+Qib54yX/9Zix/RJ
LDCrMev39FV2/xx8LXkkT1M0AL1eeL9fUOB5cQr02fvTEOmzP3/N9xxTMl1Z613OuQRxI4UFYu1d
bOa8COidzCW+/GeNa1l9hGPMYl11qvUgaWbfIdPfcPIfIPXGivWIQkQfnmhk/BUh2bFsqigmn1tg
hUS6JFcPdcOVs4ccba4OSS7hUFsinc/7DVQXLg8C/HRD+nAgbHaHA+AxGN6onoOLMfSMhMlsM4q0
DMnpJYu7rIfXjr0iUSOSnIJpZCHrQiM4eTwZztJvK9oc0O3vo3uBnPx2XQZWOHh3ltigpX7aJ00d
FDoahODX31SO7028xDButAtCZU8Sc1Mv58tAeR3RAYI+r38ldTZHtE4GCQox0EaPJi8wr/eTTvhl
FgAGKG5MvvyqKydUrgxZAlLRQUkTy/HU35HicJIbLzg7xCy003bdcrEfwg1vzj+Kh55iItVMrfCZ
T78fDRGktSsosTuzeTxsy4H4CXbpJ6u2GFdOQSW+NiuiC6Gl7qD1h6g6H2reSSCUcc9VVRQQr0uE
IGSTLSm9smbmz0PpqsUsXKXO1WGibu1GVBqQKfwjmBdfW63ybmRicZKZaH2SG3NAgSyewQmMD9uy
puTlC03TipyVUwCY76e5eP1yrX3/VWO32pCdY9cz2IfLqqpnssDWOMyRRbORZwePeuPdVYmpleGX
FiPGmkzcBpxIDEzhBggpmA7w+X8gU7TsUEvxXpT4W4B4zb8BxF5uheXE3X3lrDCMgVzMbos3wemI
wh5in3ksmwfymE2mbmUQlqDl52bLtGQwMW8foBmJ9wLiMn6BlzYlOZz6BTV4VuG+PGnM0ahJh8kN
hej/aflZ0DuPlm0TFPbkrBm/XdTLNDoZCYpWF0YVVTpXO0G+9xZiAl8YbWYMehgIaHY0Y2I/iZ+j
jduqR89CjKD/QrhhyXdldRMrhB1MAGRk4diiOVyVCDJDawSKNGax9rRyRTWfAzEQI2AGnP8nWx4d
wAvNbdco1JAeIY2/pLfxleL7bx8laNKMucj/v8DkzXK6WBXK1MJPYP+IxHi3R9QbVAdU8LQ+0A6i
KN6IvMno2uz2NqdztiDZL6Lz3lxOpED7SE9eb4frCWWV8fu89jZ+TE0aTKz043Uvju82RSrMcUBb
fMgCzPwpQxCCZmTU1R8qQeoqXpY9fi30XzsPIS5oaC/3DyVzUlD9JhPi+xhLD0Mp5FO0Uh34Lp1J
e1joyWXoTPGfggod5uOOgx6JSfBeaajSCPE+0em/8o1jAnJAsXbIFK5xt0C4WDqDhLBcdFr3dhEC
vhzsUDZtJgtrUjlVH9K9JZvj/C/895DNTSy8zp1jCwYFIuYrbqNBbns0B0qDGXJz179W6XihXxcH
Ebclyq9NZvfezO3o9tbsggzAb8CJl0wULbomauQSRXbjJYrwcbQamEdVHXD+YNrPKtE+9ttjZgiE
6PGKSPkk/bGr1/d4Tp1eByYl/vQDwJBrLEI2v7S/PE2qz0I/ndaGmARXpOl7aqyFBW6sUmkWBBZy
5Qrp45Mba3fDKqDsANj0Lj8m0q4vvhq+s8KmhmmofJ9qW7xqYBBprMMf3znrh6MikIVZyp3Ikag6
dHXvQVlljEKR4eiKcx5cPDbOTRa62B+qtB++xF7Id30Ar1jNZADiG8U6m2nKZAJQI2kQu6uB9xiN
gcoUsULr/PEFvK1OLwAJbHugOzmO5foALwcD64s13/Ec7XrnlMgC9PeHT4DzdAEaCjJraD/4f5Kc
omIaTkrCx4YT7RbhXNgrQd8aDW4osCjpnoS9h84E/tP12nbtcIJWQuEOWN2y1E12207kVZDIUbvd
DR5iKKpJRVkaWUYUzK0xqdqqO7NPwnXAaH1V0iEfZUnZlVa1BVPQOjBQcxYz4ibVQAuKn844qeEy
3o+pUDtGAmezO7FoxdgdNkvVBIymWiJWQiw10vIije5fLLyAMlkUfAqGiNuaeFVoKMbEkBzYE+3v
6s8eE3YDg8bPx+7pDHMR2ASYHiMZFuQ2nddYGW5QwdqvtNdKOJvDvqbNn7BcgZx/7+Swio27If66
5L1EqrVGzKhHllOUzRq/Cg3NLLAMqCfU3tb8W5Qq8M/o8zzcELWmTYOsgERZcFZ1BeybAo/ztjuL
Mm6eiXcHwOfmGLbmTrQekcfS4DCTrXcEuOeMg8P4n6hEqZy5zgQXbSoSRPEhdaJjycSX39zSVZaf
VUT03M69SZNlge1s4M16hXGt1uE/tbaqbmBn5+lOykAQouSIGOeeiMl/ryISHQLkK+SmtcbgGP3T
/Uwh6fSGhkS63PTJ+XwAZlF86ekPZHZUBe60h8Cx0GVGERH+s3ds3AfLoB0ZR+luoCAO6zwBXqf0
oCCHyskZIY/WM2CZ/IrqoS1m+L+tauHNl8Vbiznh9Mr06IUhwKn0PDmfuSaMQ8U9rS0EO2+H0SDP
S9dAYNFQMF/k091MxfoYvdR6MzX8fAXPmrWJgRswEZZqomCaBL6lRazHRpzq9pKXCHm2JDgtQ/24
upPpJt6foEQSAEfETAOWfR3WAGQYJhthCBfeySSBoDgAVsKTc1vCfFQdYl8b3JRF8eLm6LOvp1F4
hBmhGOGG0Ouxy71X/mWTQs6hnf1THF9rmaEQPuGqZQXj88gr/OJUV9z1pQybs7yfOlNF87dBzEfE
fWY/TAsfdrRFzx3UUx7AurRtjNdLrTZ634JBQPbVUV481M/7qVqEZSRXZbKcqulVo+/laKpVrlLR
1gSq1OsnSpDEBm5NQr8bezfNxiA2aW7cV1IQILBRg7zgWf1AdGJzdMpb0jRIT5THkFmBTrxuzq+2
YFs0ODJQiHsQ5ia2CSGxnEAthurOJmHI6yttg8kStN9O4dSznHqFGtoXXNWzMctDHVmq/RcqbntZ
cZWqLZAjBoWfw7Est9kDDVKYXHSB7WYxmo/CwYDokVCN9cR6dtv3puXXZxb+BS3cUdPO/759w4T3
Kd+dpdebujW0Y49NWWcvtxdf9LF86LKGiYtqQwfBPpJCIjm5lkyd1Sw2gYBM+4+sx1CJaNR+ljmC
BhAIbHbpX99KoGHo3ZJgglnzXcDMMkmT28YovCvnIo58EQqCM/zst4aPPpvdLSBSn29Ur7cougD1
E6drUEmHeeTVPCmfdfjsCVwN1Lzc/eWX7JA0l0kkHvKJ1larG1rxYnvDHpXwyhQNboC6ihEb54wG
AgOVx1woPFiWlN8eS84ZuWJWoDpycjfy5hfdJzbLkFVIzKl41wN2ZhsXE9F6FtiPU8jhE5uFZUzb
n2aUxMrR18uBTN1N9H3VqoSz2CbBk0l4ktIKqtkEXVw/WaoaAehM+Amjb5fqlhSXJgcLjrkrFPqz
yPcMROsgfQ1FTF6og0f6+k602n9irqxolxnDclX6lkBRcOe5MWRTZ8Z0pbY41uU1nSuiNyHghBKX
uNStyxG0NQ4OA8cDPYoKs5aNrMCUfLcym/em8kQkp2xYi8/Gcmfq2c5PD06f2YqSCIpRAYq6NAbl
+FR9GsxneL72gitFH4W7aaj503M8Q5oNrScKld1tGgk7K78XQlffXmt7MyJEdIWhntUG0jzTQl/l
L1eqHkQzibsLTvaUep3uylQbUZPF/m8bv4gaft+SxCSb0mnqE7OBGH+QIwbd6oNmeFP8C/Vf9JPt
zE/e62dsgS9a2GWOpJnS7K+0ZBomACe0WF0ebcO2Jlfe6ZkNdjElFWAG5ho5D7l/8Bc8A8TDXsRX
eWDnghindCDcaDghQfXNVQUa9cO5D+dXFnaxpIs1Wjmd3ijlzHaxy4R0NVVyT4JQmOjgRvDLm2s9
o98ntOCHSETM4EqBwdW7z3f6cTZdFEm/XwTRqT/5KDXXvKWEjjxuuc2t+ahLQeVwGXiPuqIWBeP8
kcd7IdPORvhcdCzQtE9pDQyzkJhQgVeHXFO/4uxwoRn49t2wlM1+J1r86y8dmZLzY9P6lHt4h6Lr
n9CJQKqknrktJKreEvCP1CAt4EjtiMHDGC1FrNOxTLnDzEVIZgVXaOF3ar2hfBeZDoLqM7wxkyqn
mxuXvkjzfNBJhAHBFQpVGt9ZG6D8oN/1Rrj72gl5eyJW1+4qzC2mQ5anMy2fIiijL8wrtVe3ulqW
DXODFONE487++NXlUyPtmM0CWtibZ5bxlZr5Dhbc9PW9zfwyVnmeUQLs0PX2aB39DH56emwgAoN5
pnMCsQBLYbk3BXV47HdH2UIzzpLRAsKQiYEM2zcEjI1td5vflaYVON/z6h9f3dYMGCtauMmS5RuM
geEW4Kb1v3RUW9vVS5vzr8uyMHLuy9qnKNL7PO7aIG4ICvnHbZX4OAqpwKg67LaxvacQ7t702JdY
ybUQQ0RzqHoAGMG5ClX/DoL18KdRYTcNdhX/W/M9TBf0PKUd66MMqkLJt90PULHv38OmRmo7r52i
35a++gRiayij2Jco14qM+7I7nW25lJ8mtWJQF49m2Ti3ti522cDALYjP36CnhV5Fz9eymEO9fH14
I+fRFUvaiaQHGJrJb9dvc/HZAvylzwEk2MTyfkA8fyhikQDdJdX7v8ZjrpzuAExqasMqCA4jm4IZ
GAmK094UcNzwHco/IjmXPEseuyLcBaDDPp+rjI4ph6+DEsl6O9JaQif0BzR5DUOGpTcmuR9fVKPZ
EwEc6Z1MToXZ5p7CHAx0O0T7Nrfp0TL/Ea/eW9gC4KnnOevAktWjz+XMOFTWlgeaMrWEX01isKgX
vHA04C9iiDAF26yPO2cnxSw0WfHSSTHjzXsRtcTGaqoZ3WlADdgZLXb/EetLfH0GwpTd+V+YmYUY
v+B/VdlzGk4jATiwXUJKRJMoOiOG4yZe3AEMMT0o18QAQAOK+HNMRbv2p/4x78NDKksE+n4gQGVe
TQCCMWJYi2t304whPviR9Yco4iS7ORyrHbDyhrCi4ut5ROe5ac7jsBLt06ndKIjeX2LTesvlyv/D
uPEwF1Q7pGibO12u+Yv/Cy/dI38Z3dRyS9Rb8LNCnEc1Mrj0V1SkO51dlTJ3he+l3tknv7TdFI7L
w2myO0ByZcH/m1Kdj5XrJwLOWWJYcSwKRDz/U5pbyNKu/aePEy2TxtCX5ETgL1wyyYX/c0ior6Ec
HBDUQ7k3YTQaxQj+8aEXhpBkLahubtPdX4jNtk707R4yiNTaaBYScFpV3uX91KnBuxuks9CvEQhe
E/mz3C5cUMPHQTCoHKON22Rl0dgwTTbdH1AT7yomaTfIeC0KGrEbWNUzszeuVjviWIt2r/PTFZYy
TQ8cXsLMZVGkwFknao2PPABEU2fAqdRMAO8kvzL30CLgf370geVfI9L1uLp66G0atcrl0SHuUE/b
qW0nPlKc7OAdC9Kq3i+EHrvzLQ9ynZyHxmt1kfTm3ulRAgQskDB7bFYP+Kz017phoIWtHy/cxJ1w
PD5l+dCaz/P7IaHGiCWK2b7C4RcR/sEKTRuQGwKyMg1nX5NG4SC+eviOWmBPsVTyoolEdPuTV3uN
DpNik1zdgHzUtca3kTMxdu2Tc63m/AsJgmVmZHeYl6+xy/0DqwluNUnikVRLHAVOwsStZKgLAqK+
aSYAPibW+0nfQK5LOiejFnWw3zsqL3a/3bqur1lYJSpdJSi5zW5MxoK7xy4ngZSA144gGIAPPLys
kbJ66AbgORzS06QpQRqJQxtw2YtSFywRqXgAwgdLXaDTr0+STzTzKL4oaa//s196oHq5peFJeIBn
ekqeXaupaP8gwtMsOrB3NGxbk+DV0IB/LioAKM5Xm8+1MKPLx6B1LFVQP7KXqL0xnMB+NltR4UVx
6v5SuHJvx7wWE4FEuQj4jp3tIrBTUlbvPgEiNtfL/59GbIVoIedFup6ydZnIeSpfDFDrY54VX2qp
7gEKx9gcZGhOYJIHZ1dzvIgKCemTS6lTbrJ6+Q94bM6Y21EyoaFAPsIKC9/+YrpfwvZznRGJunzs
T75FjWaSI8DnUYUp7MjeVh71aA3uMNNyaT/yJWqiDirI7GJsHT5WWbFDK8mQdaEga0AN5UPHGVy3
tTy7liUCkb9s7N3iWlllz+XS7sfhhSO9Qdo0UZv28X1FpN9kL4bU6OXFT26vHHoiKz4nXoAF+4NL
EuIOHTZlYeY1JDo705RKrQB/9xWxxcsgD9IHQnMPqWZWTmcEi0aWYs4/QfusQAgiPTQmOVfyuK6f
B5YT2XL3Ro6pvg1lB95CmUVMuwkxrV8IvDta5pY9wjQlIRtojJCCtMwcr05K1NR5Mz8NXHgKr1iX
7nL2heaHxekusHqaBrqy3P/+DJr1i/b6O479xdUdnp5pLk4Bv/Y3BQ1k21f0Fxx7KjLIEGs4Bxo9
c5dNM0zx0ngp5x004nMIgVdEJSX2n2G0TEKGnaezM6db7XSl81fhTi/hLNjVVUnrz8xIrhlys+rF
NLoA7nsE5Fwo2aNpr6tr7xDKM0PhySD0iCLbf29HZfNDQCL5LW5ZY1mhhl0ua6ahubPJj2Edmlry
qJvgS/pNzFOs9LhP12h9Edjm1nmyACRqTVLow+7fiSW2E2ddXE+MsNuiya57M8iq0rutZNot8Cko
0hixLlg84YtsKqUFVrP8sYH5d6J8J7b8Sz72yRyWBo6jINrNJ1OmKylAAggOLkBIBDdh0bXs07nT
AHlApDyDtX5HCkO4zlNEie9V0YG/O1C1U2IZ7wOtBj5u2iEvBJsWFf4mMtYvzZ+UIHSSabhiEUfi
NI44YswfO87+fxihoWYvYkPVkzbtmPuEFAcH5mIeUc4LsBeaR2d7sMNFVsByTOr/QUy5TWeJLI+L
Z+3ep50WAN39+2MxgcRYcBV2Tat52vNqt/qHBnuNiQ/AFfh5PUFjXoDx7bNRpyFPJWwNJLaoTNYf
9sYhX5NMuPtGpT5hqZAfaG9FLKUDArVcgBF3VjZ+hQau9rpSqX2YDRPHgIB4SLsfoTBoLPPkBT37
mfh6JM7CBXItgQkzO+IXjXXxLkZ4qFrEU9d9UyuGLIq/XTybEjgVUeoUs+OvCQMHJ8Xt5advmu57
9BFi3yW1MTkpmgB+9gaMzWQ0aBpfFoSF22FiTpFTnGswuUvVzoLn+bAlNkeAIpEsieI7+w80h2Hp
mlOVKw1to5TTjNCVLEkUc4Lk4KokMOh8uPmjYjRXdd3NABNfJNxeVymBTqwKKIJvZghcMd9zEVWr
PB0x0+BHq7o6vU7at2Zk0saTv01EqXwUyE+fsW1kGPuk3cGec2HhtonLlT1IUkuqtUp2tRqs/02S
7OLKDNLWI1VmLGgVSY5ehkxgU8EIQitp3koXLTEEoKFJpwtr2yxFrBI216mEkodIvUKAUR+Smv0m
D4a7BAXle3LkBHQ1b1RVanDiwfNh9SEHqfk+w7md0KJ3Ek13HRAKc0qc3qWiHPj8GpK7plrDR82X
HmHOvM/fCiDDjNxq8T1e+UykzMCP+L32+aFprtQj6/R+rELOrnvbwuNAJGYWnqliTckScPkBzkKf
ST2OWbIDn5QE4wWjxRc2vBN1Hh8WEhAgLUW0N8D+cHUkT1soNsofvXjdMyGBHYd87SmDYj8fe99+
Atz4YQCWMJ7oSkzpCvA8oQYr2Xw11ST4gnGIvIHGDWvjKsHnBxySVmiJqYkYjMJ45IIMpqoQmZIQ
TRYg0Jan/CZQhHxGaY+bpj7fKid3FMsgAvVzgwqc114TEpMNSCIA/67mMTNWXDpeLXmxSnYG7SJJ
L42iyBpYPYkXIw0l0wpAETLQ4pFa5k2jfqniVOtBAI3DsHT5M2vLydXJ2Et2qmTRxZ+coq6LgOv4
yIM0q+fvIVGzb3qf6ViM8CPdJKxlV1rRDNBBK/Q6bpK+K0juGcbhK7BV6QAEydRqT0fB+Wu8cOxU
qCf2z8YeYaMCnmt88vEQHWZQ2a9+nl+zUp6FY0PLvf6UqQOPlq1O7A5WxNFYsSBlwvm2El+3CPBh
D/sLRTPOEg0nEBMHN5FAEvN/QF1Ti80q7/KsptwEyTuSSq2wLRWiSzpIzxVxK6R5dYMLTIW/WowH
5fbqEtt7kxmSEZwzXPeys7SsIoWeHmt1gZkvurIihlDtDTc5UJYDzEz9iaQYWu9/KYcdEAKOJ6dv
olJ51jkv0rQgO0tBTnxwDch9HiGZN/35k4hdUgTjiDWSTdxe9gthKMQ5nP8cMsDVoWgekK+HZ8aY
bGgc3w8jQKxj349TXAGHDGQDYH7L/M/7NYQgVCREGPUPLhzNYT99oS1kU1fa76QtZxbp23oN8M/h
HX5QsSCr1vQPy0QUumBWSSBHG8jr9kh3M2SDCZf5r1zK0wAh5qzwsPLZi515PU7Qo6h5MAMiAsuj
uURN1aw02QxR58w4guq34NdmYVzhL6MUKo3jekgbuKhLEpjdkx0ROL/ZWqhDAPDmrh67jpN/THUE
iuunH9T2ZBUoiEee0yiWwiXNv+Kckno5lFwqeT9nFh5CIr0KgKzJ6U2w826Sl0Yx0ya6+jxr8tz4
bMWwORQ5r6C8RC03zm5ikmqTjiUEAUzMPv7Y2YHrj3xB0rK5nWevgFNMrVz2j29mCY/pndvqwdUM
9ydw4L95YTBR3RZc2HLppB5rbJ1EOj9S2nWCjjDsMi0aF0v/LP5tyxpD1bDuxnV6j8qRVVpnob4S
ZNdOpr16crOiB69NTHX+Q2Y1sPx+dD1bUc8RqPrkqNI6sHI5takNwmJTIJYldQn/Gf8E3niZJYUS
tiXBadBF3IVxfFfNuDy39wj/j3aW0lYVXuSmZMCG8h7ZJOTB5Uq6Uof61VBPY9lnLrgeWIfw6QyI
d6qk9wPQlm9fP+YpWJWLgLusgY2c7vTYMhwyqTv6FCV0TaW/KVlT9iev6+WFYdr96u65CCLlCoCk
j23VpGq4DV4IY0vRWt02FUazX9Fy/CJKHty9J/0MEKXnyoxh6xXmNAa3Fx+uWyjW753cjgh9qW9r
O8iFdfRLui16fX78mwaYMQWvaiRHZ5e9mf48BghXCbV8YeskkuI5YFPDsGrh8Jb+NuIL2h5A8hLt
2o+/EtsCoo+LiFNcWi4AR5pV8LO9VxMY+jknutJ6S8LJUgK0xYd1PMaT7tilSnxRWKTmj2CUeK+L
N5KCcGkJ05My/gRvrHa2mYLC6IKfyy7qpljejDId0mG4Xs/jmXbuRAgpxzyzc8OHxQomAO7UVkrd
JZZdpErs2CMoLlxIWanIIU3Cv3CwttsFJxCC338960sZzOynlOpw6GFyOJZOggl5uNxMzEggeWnG
nPzcFLG7lWIop+IoFAkIndjDJFs6OKy0fIPanmbtC7WHiBtniaqH1EuKDx+LvnnRhdNeHP6keD/W
Vj0Jb90GOgr4DfodJn+mYOJnbtkHX3i0DbPg5/hQLfL65XI6QTcqmV2+Xym516w56km6GbBIkYoa
gWfTl0qW1mnq4E5MLadjGFtUhqMWn+vXYSnrZ5+zRMr+hRWqmrYOn2F4Xb1wupC4F7Uev2+FO24w
mPl6Q/hHVUU3DeoPj7xM9Zf4H5iIbJKwtKKZsV/3VpBtncfoshULaYR2TflCBdUcH/LjLQQfgyaf
Rl8eDS+Byxu+2W+nG0Ovryx7QZ6yB+VbrkAUqP8/+9rzOcN8SW5mpC/1D7HaAtsm04GLBAXZ9Vv9
B8MTeZiHaKOkSeClEurTa+qScMIcPb4LxcCfIzrX/NmA4St/cqYQ6Z8RBxewFr+1pR94RcjnJACq
pVmQ/SIqtiJLdlOjetR/5wTwcL6qKksOF9pNf9J+kMDUV1RigtXL/EyMf7XFGvIFWmzl1Q8QXXl9
+0OfyXfbS6/2FNfxgDvH8hedxwVnCbeLL7fYZWAgmYObvpktrx3Us/rOtg2g914Qpv/D4AinTJvQ
YbwLzeO0Sz2i1rzlTVTD9ps7hbmSkh3KM4/vVHIk7kGPk1ZF9I1tuzu9hklpvb1Bfp317ponRo/Y
jVzOOSf+o3dO4IofxMsX8UysP4owlPBmPqi0p1rRiEutEn9jU9RKGzC11QC/y3V5inSaKBUgYdvd
4nNeiU/7D6hVpWf6GMQZVbGT3kJwsWsyouc5U0VCzdU5BhDQ3hAF+XopD+prRVsyPked36HBr4x4
MlQw1lXqbkl5H6+SAPnMPiJR6KsZyV7jAlhjPsVf0mh1akMqi80DhwdrrE8xlu5owmUbMc1pDZ4d
q3FGbawwOU5zcR6LETUvmsRvYB4fb512Suz4VZ0JK/0DZOfUKPK66CO6O3XvsRZTVnce7Z4GYzP4
qzVTVbBsAymRDfwNmWcfmoyay7Ds9bmqbqLttQjdwOJHwPthDB+qm9VIF6bOTrQoLZuV+kx0Ifqr
WrWenh22Km+0wp241TjCMjXz9O39aEI+WNJwkV4NxCGvP9wu1qoLdyZA1IP8ycH4CZ/qhxAQ8vHn
zQaxx8/Lz9nMfS+nWuGJI6wB1tR8pNRQkf/mWZ2L5kAtruuMx2wM2Bg9TrdP5m3QRMgVZykYVN71
ikM/xzadiEP5G5HKyjLsjCzlse7I91c0NJ2e4pcsz+zyukbFcwdGGVMVRpFQCHNpBlO3Eghi0AAw
HVXWHGEo0fMbUoLqd3tLWZrKDmlxUrzFPbSPHoDtg0MOeJ6PSMrr6DgiVNyAEkVg3HzTXVYWenpU
esnNWp7r5nOsZIYFg7IGUzrGGCP76jzg1haOqE+H4l2FpUGi1KzA0UHo14dcnGCbsIgz/EVEZKNh
Bkosaq+KqrqME7VgXwWBZrBhlKae7K4NXbAthLETGUNxhQLuitkCpQ1GQ4c1JXQC/tdeY6JYCEJi
jtLriO+ZkJA4LvAmLXyb9eRp6hrWN0QgP/Dy/ve2OUS2gLKGq8rL2nXsuQxoQefQJSTslRpzAd85
njoyozPJAvst5zEj4zkWm1akSLUq6qF0U+3ozbqwCfPvbpohGFu9jE+PYXkLXJmE5kqCkqIsQJ5+
saEWovyGtiqAV+LY9+K8CMRX18JaQLdhupb5yqp0+mhZTR+Ro+O4MMocQdsDwJ418D/fukMCD2P7
Zp+iWRLxjySp0wtk0SJRZEDfFI5OiYwYyOnFI/gYmBES2qrhuzNVZTR7txBaj9RIoWculedKe8+Z
k3+H5IiEmcfr3TSmipd4iVNpJcqoOjrej4TH9MqzGBQIExoNBEQNBgeuTfg86nl+UUKC6rjFiHBx
m8ARnyq4FZb8FeHoukvSAR+pYQiWnrLD1PT5JicRXRcq2dIX3VOI49S3wT1uXULJsvGMMLwlmxwu
Px1VpcOScjVU3HJFOR6RO7EdRuzBgoxdLn7Dg9mJ0hxldUJoovp3LPZXMwKYrZ1OiXtYTBocjfus
bJ0gaVbn8BXd4l10wYOEY4AmgbPWuyazYXiChncJ8am45a2swXIoViB9uW3IrXjg9UEaPdUhjkwA
/RfqqJydJbfj0WcaF/31GzsUbW0/JRZ4/iffY5g9ryL6ezVD/kAWl9NyDHdQxSbu8uefXhX5hR+h
6YzbG/QUTtNwZVvVnrd3/lkQxg/Jp4N0ZKSF0YaVOVs4P7viVMyvBilWniloP+n8Ul6GnV8uuyO4
QtRzP/YzClFt2QPpMT0NgyWcm0JT7UDyl1IaaZf61juorK5qz4O1/KDk82WEpxqDf3aw2IAgjlla
YvGeHLryotZ6phQFsmH5Lu5XuQ83Ojlm8ymjWiE7d6i1mQ5ZiV95ZFyALrIEKtfvhe8G7B2q5DQg
f/BYRDNp5zgT+p3fTPAv9Og1aLR2cNw8lXObUTXTrW19oYoVYNHApTfUjp/j3TrcEG68zTwQk/f7
nx6UR7cTnpOIdINjl8DfurWabUhSRnDdO5UKJxMDJCArZgfuXU/aRPpB3rZKYlvXOMVAM4V0KxL8
oLTmGKLydl+OVxIX+iiH2Wa9s39m/d8ictDFpX0N675GG/XluYNDv+dg62GZ6xoAwaSozLTbHe6S
6WcDA/nId47ETo3Ci1BFTlry09MY4xGRFBgemriXY9sqYb8ZaABNHpdV27ILqT0IQ6X9ocpSf9qH
DebBmLSqBY0XpUXp6auuG1SNZMva2V0FuOGzO7Jk0g9XjauozDMcdeRafaxUzSaLX1iYK16d9Xd1
JkzqOBlJvkSXqLZwmW109MWK8S1Wa/R8zhXdH0UC1uwNSdZa3vTqx5c94ydl+PzL100+Tez/U6ff
yH4GpXK8RAm5abGZTLE8hXghm10WSYepirpgC4rTm0F1Qt8CTGpT0cgjHZj5w1/Fdr9BcVzk1dBz
0ycVCK/uJHWPivc6n0Z+1vRmLKZ1DZunAAEbiIsnFq37CrMwed/YcLle8saMUeZAJ7IPRnykk+BD
Dztpp7uix/tNwxntn8u0cqYLcP36EVLXxjM6IJJ8+n6P12+iq+OqZoU/CGf+FcFRxQm20/DLtXLU
O+l6eREZ9Kc/lHxMBggDoQsOXtP1Wi19xiCXxNxqWLHeGd26sWXQkNbuavNU/6RtO52K8KK2D6Pz
mw01hf4i2DpC4J9HDTaSemhIXaCtHGngb56RbHV6VNOC85j3HPtp3NL/KHdswom4D5jBaY9KH076
Yk9Eq80SfWgdqGGw6cg/vqpbDaeHxcZ3Oiccu/+h7XbZZ0WyMpNHef/RyHkfb7W3KIbxx8HgO5wQ
e1KhGslJbaQ1o5DdNaYkWEPaz7rNOu30QQqdyv+ggF+Gc4tuqnGF4Gv2YJNACOQIBvRpB1Iw7zoy
PAMIPfOvNxc1kmBUcU8K9IN2FKkz5AqOrRWZm+R5+MwwSMM1dFvzHAR8ZzuPD3rM0qXQcv7dwsDM
CXWOvlPl7HkCt13OrZZWjluXnlndmb+ZLrLzrj3VoqGUTWKqFsJgCwPr6/DGurWuwLCSG82P8jm5
pDe9LogOq5a+lHCKacLc33obJld+24YP7vcS3l5fJ+pT1PYNQmTyLgOzxu4ZpJbPANFUGZGldj2b
SOcJYTazFKwfHxQAs6bQJhU5F8kIlY6OEYFfO7AOHJA8EvG68S1sc20PHAqVk49Rj4SW/B4Zd1ad
bQwhpZRWUjwuY2tOhfsAOlAazgYB3XT89glC2QMuAVS1oxdR4AwiCNzA0SAQ7Jj4S7NGHj1Dk8lH
X9/XtSkcyDue5ahaA1t3l8/pNtm+dRgRog/uw7JGOWnWHm6ZFbrvAKQTVEP6niLfUXLNkmGKNAiy
4UGfp9jb8rQKueK+LAikPvEeTsKqaM+Ek9Ktg2RH9Sg8hn2T33wZde4vDPEvA6og+qycSk3hsBEH
Bfx84UZ3TI4VlUWx4H8h1OutptjqZsQhC1S5jDodVk6fec6udBU2PU6uHzs7rjEF2Vat3VmejRQW
mo4sD9abes/Dl4FU1QH+hG2WovvmBD7chB6+V39teh29TTCzWokCEErAzlftN7eCQ6fkNrgjjJ/5
VOBv8LOxPUN+4q1U0Dvc8xKbiR361Gnk8x9xaaoR6UF8wps5zlaghxNhljzdv6/dMui9htfKc9ek
t09nOwjEY8y2Vg21j+RmFAChsJi0IzIDHYJ8aD8G/Ss3bT6bMHWkmYvuYF7aWuVzu7YXb5vWZENZ
mA2LeBudvWmcOTSojsOf+CEpB0OYAV7RToKuuFZMlqiIXQUhDMThnWRzd+6IBsCSu1GOxCrq6mqE
nQatyGSsXBloSulB6MFzRWCLpjoat7W5gI7f1BhoGDuwmfK1Z2WslaVGW2P9Y7aoorLL/COfM8c2
vmkF5Atd3wxaurNNAeoqIevIItIaTT2318UNfNfC6N3BVx5ihvz08XJLCp6ME2yE8GE8ESKtRRNU
jDeQ0U3Qp+Ifyx22PhZge7992uwUXdOJ3qEPiXUfQ531F1s/nSN5UP6GceZ5RgbzeugdMdayIciX
+muqfaBjB0Suer3+NySrc2FwgGbDqETT+tlFag9HXeAWY9NoQDvV6RuI4CxHUA46NYYxvIVtJm9k
PR+pNK/0l6xxQ/sKI3llg0g2lT08ikPiBt6X4DkTppAw97vtN5H5tsrnug/poyHRpzG3bTJgYm1Z
bKw82pgELXVV4gVkDNfErpvyooECxaReC9/gTMEd/G6BVu0cGr9I+4Aam863FExPzqd+zzPbmLgl
zZkqvrvtUFRGgemPy8A4zRGRReXvhf+CtTSO1wvGDqd/EyVL/AnP/EIaYrnsivGqF1GkL228qqH7
atnyE0o9i1IUyqJfpALt6E0rEvxagkG150U9BZZrVEMsQYlOO4bTslU0wRzfBamVJJah8i75tMwI
Kn9+zeAelFAnz3za19ejlJuZTBOXF4GX0FENgVdFv5cnjOZHmbse/H/C2gwNhDdwMQDce45crnMr
d9YanXy6SBV/CgilsqQXPwWKgfvgForsHxwQTjk+WKrfiGpmU4N7S05bpZaEeJoKym9yUwxjOoNp
Glr9RhbkBEu6hhMtVjYvyNRMqTz7Jamf/M4FWQzTakKAmFRQEgnkklqwK1Zs5eG+dX5VfNM6ec7x
3WIdvTDflWL2Xsr9tftNse9CgsFx2MtdFjEJii7RFuDgQ4ddWqGu7VbUnzBrH9lHhnz6C939cpwW
BJ3PeSjN5nPltRBx1fB1VtYNb9GAarP6sZh4NeeJtfwSCiT4z01kAyTlx6mZWx6ktMHn36S6vGKQ
GVOoPQZ16F9BEzhYbEbSEBxqEfCTA66+tqnZhGnMEAr+uUb6lyk9t8FbGSkufj1Bs0CRFPHQ3B5Y
r7OHds4lRucpe19RGqrzT9zwAbAioSJFBUDEYkaBWMDywh71ddInwGx4Bho23WG9maDjRXCpn+gQ
VDUUG/8tuoJHMNRPnzGrvEsQpBcu/fyUuF7FP4MD5TJwJuOY9Us4Lkfg/jBhgIkWMdhlwEX/3+il
PCZVjXAtw8VZg/iO1jGbEWbPxX8tt0nfO3xuCmqqFqSCE7Fb59Fp3a6rFHSsZAVh2PkinJMp6jJe
xASbKKtk9LfhagLKqSbzIV+a7BmTghL2alXRjIGs7F0Kx/Fa6H9MnKgtqf45k/ggSFN91QTICEqS
1AXjQljkPkKawi2LjrJmq1mcf2lyq5DNTJzJeqHQOK8fvcGDj5Ujwr8UlDC9hyrIULM1Fay8G4r8
4CQhGir6SuZv8fW8JhyhEUH6T9YsbFergq6BVqFJtEEdM5CINnQi3Zn5KWKKRvXZgJApptGVFMiT
v6k0yu73RactIWDQKzv/A85c3TtpfFosK78Oz0hdVTMr2AuT8UxN1idYfilYJqurh6LUUdcXGHvL
c05ArTPkwaOg+jFNCis3KWiKiVW6FWKx8kLtB3bgsu2J24bnkyEs2kCDZHatGGs/LD6Nmw+nHosm
cpIVWrlXjoqqDT4LpqfIgPwcJGpV/TPqKbptr0nloNUyV38WFoAv/wlWTnnPGY6GY7Fi/y4wKMJQ
cxpXkbuH8kiGlGlyHoP/iE/PIyf7VaSB8DjsO8HPZt5ND2BaApwZXk0o+HoNocOz3eOE/reSTyKG
d6NYw4BjLq9OsIIWFcnuxkDyFWcs4YSmOTrzhy5gNG7YJMqTRGM79WCVeV6J55U5rfI0zAHhTyH2
hp/0JkxDB6H42ja3Nn4aViYRewi7xfgYbxbD4JyHEaTbtSB3OCMM1+GltrOwe1snrvO/4xvl44/D
El3NcGFB2lSE0WN2tgFnjwOKQA6cTXRyMryentSopBOLEl9eUcsSTmfjVn+mXNuDyiy0jc2oXuB4
6e9QT6KLAuuKKMe9DYvFKaqo3K+1FJOACAqGqwqNA9Rcpp/dr1FAeAwN2IxvpaxYz6kgQGVsv6+c
mP8S6jOt6j8HCPeZcZmYSz4Sx6fsbSCgY3SXV8mVz0xsF9RZ9MeGecDIuu7cLcrzJ3v0vxB70apj
h/z/eK1Lg8cx+XhPQDL2xLRzOiXJk/ZAklu53PEKjIKRxN6WCj7IHJ/rp7g9Iixcm0mKVl7kopDT
sw28v+F14LffkBBSJNBKahbRurABLn8sC9McAt08osDoNLpNB2y7Tt8ZTapVAG/vyqDl1G5oOVGK
eYgAjVzZ65vCEX6wYacKO0PlbTnO4Qfb/DXdAxLaTa7/YKDna0z2XV7EsWAUnTElLOxwUtrvIS0k
Mt1Nxu3E4mO3Fenh2lG/j8xDrNtSBnSb8MYX/tqDbl1rdsFZhDbeifNfxn3sdFmAVoMXSKyIOuu4
QRgzfFzon58AEJNV7VOu3dwPaK5od+osnvCVgJHyuQIX7o6RXaqfIR0GsjAcMuelEkAVTPG1Kp9B
Phe6/5AV5mYmIok0Bus1j+App7O1pxCiKQORXMT1AYaLsrKOXWByGQBV9RSCsj131SYOF4UzASMn
PL/2A8LpjeNyxHBM5ILhZKrXW/7FvwKy/C0vyEeaj7CKaIDNl+cvalwdkGbuOKUr9/2UyGJ4aJ/G
o+pTIkozSnkCME9UFtkPnyFGrhQeVkoC670t0Jm3l4XWVEIuesIZB1uHXTUuJFjkWpOpKcPr4hQQ
15tHhBUYGOOu8XqM9PY3BXJb1QAYAl2Epb2afgLsMX/Uej/3n0RpCfMwZS/0aWx8mGNnVEwRmals
muaemFJ3iTYsf+tTVfFm2NKaWc+RCzGZoTzp2QRXZbIb0EHvMjdbejIOxnx63u10rjzw/gndFS6/
PIDkL7MuypCFxTjonJ6+5ud+ep14+gEItq4rFVUv6GjsomYCF/AR6zHmHuIYppDqJjAdvfUvTLYu
H6k5C9fgP2RqjmYWm75sYMxYvyC77HMc475OCMIyM3WNdNqfucBP1IWY7GSrjcUfMgFvtrpQAESB
xzWd/iwOSIw+7HDG4jrBatjuvdUdFsy8O8HFgMLq3Xg2HyqiA6X2UQj8eZDuklq/vlX1XNNWhkQG
I+hy1X5iubcwkRfk8GcrRbNLcRYGg4eB7eR/r25GagCFPqVUlZe66fVYG+YfwuKWe68hiw04wtll
mXGpHJDrfGjXLZtaNKPezBuKcS1pNgD1fjb0zIKM1FqcY1uxJU5xsGhnk9Z3n8jc+TsNAaNGZo2i
QWpFz/K3WS+0B66x5PeOyc+hkd2Axb9NzDLPFCIqmxrlqAAEev0clxNtg92mlfZ9wOGcF3/8KPBC
G3lO8S8bom3kOyIWuPeGqOpUZFKAG0syj6o19FSDUQ3Jfg6D+EQrean5RE3TPG0O//D7qm8ItwOC
SMiBNz+LfiFE8SqpyljlWCg8b5EDwiNRnPkpOyQ8bTdPPUqd3v6pg3AHQa1AbZBHiXhitiW/EdcE
FM7Js8rJmQN+6Nj3oCAtTndxPE2BN9QP41K7JfwgspY3SXF6+YCUL2r7iSVSyIHSqvNkFYMEGQtB
TmE2tE29LXfiGFwqyVtvNj2bZ8e3pauG5ZnSofGV22wjE0RpbCHv8xAoUwvqrWP5g83wLcvu8TOu
vOxOAeIf8hFyk0B0i/J8PdJkk/c5NIswld/OEPBvrp6FSpmIn+JeHGUz5Fpw5hYmBHkhR/fPOiV0
cG05H+8wICvwsY7JJ+03qAms9cZny7a6a8foOFRc76LgRD4HiZgZSMDMihRqhWeHsH4+gIQmFLx6
YzbsG876oaN+2XliEhC3wNHHhrswlht/KprSysvRMHlQTnYIwhQkvPDgiHTM4bHOdz4jpW/LN99R
9+20Ib9+r3G2u3aAiesoUJ1jE7vl9Hii3N8WLKZzLhIDTd3gAgV2C963xY9roLg3qtoPhPGK/WV0
XKyKF7rFv/zaeVAvJlMtfJTfLP0Unwc/g21Rjb3RHoGuRRepXlQQG0bJe5V1BA9gMzkIHkH7BoFA
oQaw4bqbbJ4ukyCew0lMH2aJyb2thf1H+6/PxbM3d6KJr6rxh0vpFmmTXnyLe9HULim3xzDXbZs0
w+H8LxrbR/iQnfBHDeoBIs6eqlOXT8I4QChgMXVJCsAXoWv1qEqdRQLtkG0PuiJtni41ZYFpomrs
xRUZ1KeVbTo73lUrI4HOYpkQ6qYE4gLYqFIpZaP+2y/1mGrj9896Dd/VHkIhkWCRGOtXCw176iQ9
tNl1qCx6bvAW4Q/p6u1PIlkEEr94HXcmv5tbRKMCuQtZgT6LxbL7BBtDTkd1Rmsuxkvi1lBGpV/6
J6fU8YnHDkrZcvTT1CeyobQN3o84HFtyLRWLB865WZSvr8M7QwrY2yC/ejSV0ROmbHIp+kEGk5X1
yTWfHQXZh5OjsxV+Nla/Xuh/iCaUmXdVBZWg8vXHvO7prnxFFGnPHbmVI7bA3/c/PS4oZKMtwkdF
Y85of0u7XG1zuFa1HpvWqeqn5WNTZjBvf+LbsSVs3UvBu666W9qMMTnsXkciUTX04www30GUyG50
4H9ByUZfxVvz5sMO9uxW3Qx6aPcf0xyjATuJ8NwGqmcoE/cY3zwcSf/VuBr0uW+T3eY87cT5Tcfy
4/X0emWPD3khAIwbqKT+GZvIW7pL4ODE2egNwgUI6bnoWtc5Nwegc1CzYzZg3hRPWAyAb5w5NYOv
5sLHE+YdqzUe1COJN1Nr/oNR/+Y13zkzLhZFWseRkYUM0ugj9XfhpasdqP8nVfDQLVDM+0Dn9sV4
e30jCCon/EizZLkP9t0GDT5u5qyBL6m4WfHQd3zw/E6XBFjYgrX2GX1oSmCm3nUjgrAGIU1hlocT
XdBp/GP3fvgtdlA4c2RpYjvu6raMlC3gcWgsMtLRjVbjkmkzVCmKV6vsCtotBQaeixjzMsffz/rE
1am59mgbXe47PLeUOojl4jt5XXyjUUmaTC7T/jFWOxnAv/u0MGm3XQ67nD9i5TVsbSyRPtLXnC4+
GvGswmLnbpA8DduM4UhKM8pWe/9449i83MciHWgzmP833vMRGARuOA0vqfa0m4I2G4MCGY6GbkAG
KOY73054broFrq+O6LsbW/xVk2tlB0GE0JrapEX6z4dlxyt0n8s0LkBzTrHWhnZLPXNSMucIwwq7
mxeZlVKRq46II21b1KYRLEly6cPx1DDe3XVEk1wDq6ea73Dz+L9yR1kTaJtaLNpICdJKdIX1Ot1r
p/zyi/1PipLAEf/IXD5I7XMopQ5Bdox7/LWp94P0wbsIjmYEH0733aHnS8K+o8sY4vTQz6OzCrZY
TZb+tBfq21HqikpWCoc04iv48nfbVGB37BsX84G2XvNPzm23LoR8vIobSqJ5EfRAWtSwoCwG5wL8
7HAa/7bFVVwzj1M6fpwfpSmApvoCbYrOfFCfZfqVMXLL2+3lK+SN1mbBLZ3YwQnSfMMhkkVHw6P7
7Xodym6uTJ2TmbPEoN9FGGaLG0C/fSf2W3ztqHkkYow2nsPV8at9EH9w/8cfsiG8SteAKmXvL9fe
7nInxvfW5WRVmRg66J7YsHHxgYce0VCcYr0H2G7J4vWhjn5eKbZUAfHKTKsYaHJSSHCxYp+tIsbr
yicS+PYpgJBuHzBj2ADtpLDaIVc8egi7FC/aL8lohHI9ywaepxQDjQfZS/Ar6jQx/Zp7gseYl4FF
89wWEBIXSm4f+pKWCKPzmz4PCn/y05tjkzSAcp+JJz90JBISdo2t/VR+/i9bUwfuSL6pNYziJ7bv
UXVjoMLr3cc0H0yNRgQW5Hg72l5xA9wYn/VruRzhJCQ6qB18XhkuINWs/6hSSDYIC2T8j+Bzbioe
q3wAlrwCuTZIdO8aKD/6i+ysRtFmFQJOzpu0H4tcwq90lBlCfMnZdPBAmMymV2qWZ6u4VIZ2UZSq
5rYAG9SNnigNKbFG9Rl46OL3AqOD9SkMyXrQvqkEe1tz6ckpJXh7R+7mUBnWZSqMkjtIfTgwIjYO
rpuw0XpTVH49yfcv8NgY/SAHCCgw1/SLkEmrbyHD0LcVYFzYJjTxaL2bKpZB4AwyrOo0De7u8zr9
XwbA5VxZ23pDYTfVrUaTFVYZFPhBwwWorGbcvUgyR+FRbvwg3y36WR2RRdBq7Iy+6fQHPHTFpPP8
c5Ks4H6pZDQpCaVTWOS1ZLRxiFfwo9sy/nVnTM4dffGJcDqp9nZUW4yEM+HOkQEcNNaaBWcQn9yB
GO5C39RgLJCMMqyVlta6mCGYYlykw7ucrsQFEN2eMlKL3d1imw5eLdfBdLZY34zBC129VWg3ZUuh
dCkHfxZCv7X2hNpu8QYEcK8IQgf7NfsSeKQ/BytI375NXx0gUmtGpQhq+K06tzOx5afAH9dB9N94
AP5N6NTKseuHt52XhByLZAD2WAQ9qMILkiwEF6G29meliNasf44BB+nXhIQQ7aFLRleXomTM9ww+
YbyrNtgokjuVvV/Ghg1DPE+1MsnAio/EU18ipvcVVALyRl7YnlynJXBhtKml50cAgjHRc45JYQRN
JF3weIXNapXUQY/BvO049VOS9tqWeYN+MjYLg9ppFzEkT87VSpKTKLdeq3a8n6VyLwCVO0tBpsoG
cHbNsAx/gE3Z2lUCRpT8eumXp/z2Np3whhVLwUQVrNB8E2mYe+9/aoDpDph3Yc2EzArF9Hbd85/0
xGHkP9PUNQFvsjANXYIUv9CEHCtxjdWcDbVaKC3sv9FhVpLR5P3bCWFtfELHTRu9G0hv3XNTY1VU
QFws96/GOoZmw3NfU6xXqPDGPjmrBtbEwK/f1185JIU78tCcOIUju41FwCQJ5cMj/aZ+qqOmXvQi
y47pd/WAu3zi0sQoj5ZvVZAPD/N1eY9z0dtbCgahcbfnkJV6d7+36i47WhQesChQSN1cTL0iADjD
FpbI32OgIfo/cACGmglGtGQWRzQOMMyVKyBYBGsF6Q2tZzcSl8vhx6QKYzkUEJFoDKdb6Y+mgmI2
URjGh2Ue/ww/42nkyAuqHCd2hbXWApyR3scanjDJWoLp2NrpAGtEthb00rnvWfB3PXEii1B61//V
nK09szvW8XVMIEd3rJGVM1D3bU6zlVixuQiZwLZwgwAXx1F4mpQwxS+lpz33Ud1U/qork5zp/oz0
U3zDCErgl+IQOBPsFO7xvEDXZ+v0/9IDwOkgbIvDXg89oBE+9j/oDPkjZSNxT8PdqOCJCUJ0rpbG
FbJPj+NUS189BEXUi0tbR/9JFrZm1iZuuZUm0MJTEqkomXk1qiLODh5pm89m0wfdgF5Py/9AxMB8
eg2MubmSMTn0cky9CyBA9nC0xf5ujcl5M5PtG1VuVc42mQwBv+8x5qTE8GHxr+rh9UM8+cegxgyu
TBXj6zaumoEx+jLDtWCMIADtmeXwwi7jUFFJB0FdSeHc86uJ1xRl1hCCF7XhPZ3Bmu55onRPzCez
6RSQ0Ke5hYD8gBZfM4ktvBxfKnn0X+D7KEPCH4KBSbfp+68oqRrLqZsqGlJOvPOOYB8KYi2EnLa9
huSehgPeWw6nagocIXAzm9AHCJnEiWzuxriqcSL0vbsPibG1b1Ll2pxl1fj1PdBaBTVNnUUTp+pg
efVkewbwd4nxXjavkbjdS+Z8UM3v4kRoIzWSFYC/n6r9ttbG9p6hs7/YQWAWwdznMgr1Sahwhwh9
5fqyIgtbuYtrzgWuv49f06yULcmM0KAHJWKCszh10ZcCPtzSQblFCM4ncz7f64YOpOefkCHxVUiD
n+coIoD3pDFGhTE6UTW8fotdwN+C9lCqy6cT4w66hCPWy2dvlqncfy9aELEc95aAZ08t3V1W+RCH
FOtxxmXGqmICeCWlOOSR9tPNCHLSNM10NrGFmM0wT1MItRskP7hbK5p2n0jVmX8l59FqQCGLmXAy
BdztRCm/6FBxuEW7uqaGdxU1M57FGVGO3R9L/bj7Ud2gK40t+Fq3HoerlXpIs4DqbwkGUEv6oX5q
JQfQvmD4fC08JQ/fQt0S5+xxBtU19Zvx4zJAu1xc9WJsbHC/DrjHh1Al0a3ZnPGDPdPGQoOSxxc1
A5DN6BGx8vo5x1FXAlVFaQ4IVWI0STbWjfOsQ1OGXQw9oKgNwrlDG4PbddvkoNBOQQT4CBqmipfW
ZlxPen2zO2t/zw/HQ8QiMeGTMJgoBTzL1mU97USMhb/eec5J4eZlrA/11P04lFe/h5MxDpaNsIYi
uLF9GxatB3z96qcFdpWbMrLSJsVUm9Fl5wG8xEfxTytC8ez7hCHNTHpvqPswZA6dBi8Sb3KDicPe
cu8MhRY55P4PGymvNulTcUbBeTHsfn94L4jUB12f71JMxgZzkiYTWRAUIcpvr3/mygN4VCWR8L69
ovLlYjNZMr4LnJdGnWhdpb67vaIg1gCqg49DMptpK2p+4u2StcbQKd+22THBIZAfWlu8LXMfaFRc
wiHvexNR2gXF0KZb8QQymf2sHMQ3kSFpaFnih+JOnKsj/zuH1Hypk+GInMuFnGwxeZXD3ccM0GeD
3im1FaXTX7PG5UyyQ1eeManoBpSKUXtVvcIJROlbltsvWwtiulzQ2a3XS10DKP932Ro6s3Zn5XIi
sSDl9W6BizPvmFZqJxJGrVzVjlXko9NKjm8Rrk036GU0MDjAXUA1oS6pi39sPHNVVCut/HOxJFYi
SO3gQarujg1B5y5P9CTpubpv4mDksoDQKw+6dDkYd9lHI+/OwWVfo4OSVTjwFcvl1N0TAdklx4ZG
mwKBm9QHb6KJEpGDqlxBCUdRKfg84mW/3oUs/Ey3HQHLi1NHDliTExUwEuFWu17qU1jXX2eHhgjZ
Ek/BI7vDORzGJoOpcV/hN6Ai1Xi5V/q5CcDflnOYf4fjQAO2KYzg8wI1mWdp8URQLThSEIeHOKzu
M8CD5g1sW+4tCV3J91NXAsc2AKYvoRj8nWV8UZ3Mmg6dUP4hxt1gXfC2LD7vgmpX7utsvQQWTmRT
RuMXg4FogojYr10dB3R9sxr0wl9WUzXO/m4ZLU9PZSbnpN8eqgzZ8T0guN3U88TKeTrQfAx2T74v
Tjos2opQGn8EIZL3JqyeThrbmTTW55nwaVLLNZoTFzziHVf4BMMWQwIYSrNjpWaPa701L11fCvCv
e9CPZ8OASbYWhfnBU3pupf3XTTJT7sQ60zxTGjXB0UNxAxLmaj3ojlMZvGJthiKK0+QDJy9Wev8O
4imedU5uloGkhAi5idVpLXL+KaKFxxsBX7QqilUdDtt5eobGChJONvsoz/5QGYua1LS2gVoCXWed
/c8srIbh70CJQMqYAGBF+Sp65Kq2nJp+i8QXBwgvCb3uDk+7FxcKr+SaApTR+JwQSmzO1k7W6CKI
lZEbt2ajqx2y0zzSCVrnkWFj7yyxBb1z+2Z/XzP+uF8J3rIs99xC4sMLpRMfQU2Bw5GBCIZ/rcAQ
6/2tkKuKElduKoN5l0QXsVTeATIaw4hAEOqlgawTuMDTlhJ2js5IqbxuAWRuUCLgj0T2rvKa06av
VGARFLHIcOPUUkPV8JELpCKHI9QR3uu4tU6LI2KNnyxv1DvEHDlP4xFdy70Q75AQIH0gbJQw/Xu1
kAeip3WxkYG8BJmFWP5ywwoIOeeYJbZthHXko0ib1K3thpNk1EXDaEZErZ2O7D9TE6193rnvBaoe
CdYJhsRI1qLe/l2G3IxgOsLC14SEba3uA7WKtyAFWAC9vN4ooAD4NwZJd2t5D34wWDgXudbdeokA
0xrB/qtu5H/xu/lExpVPCQOdGX2WJwGvi89Da5PrpUATo9C4aP+Stlj1ksqsRXfFv+NtM3b+og0u
WZzC1LbZzKTVWeN4zXn8Wx4718aSEqFcZCJOnRq0/ORHfOHJbbZwRUBSCRcvml4CUNwruth76UHU
uMjeDHdAg5vf4rOPxJlhEBVzvlDTjaNaiQwPgEyjCn+6wKgDxs/QwXJDQqXxYTsgfVA80dbMLJOy
UllNoVmno7SlFSyrxi1pdSfvDb72SFRxjLtI2GN0mgP+BXCTC5JE0Wr74EU6OR6bA9eRPS7CH+9o
pNm3InvILFr1gneqEbH8p+X7i+HNVPIKXGyWF0qba22U2xtW9gTxY7FXtzDvm5Dw3HsoJe+kRMtk
lPcFfoIfogvYDGc5bYNTEt+kQNWiVXchEY2cZq3nvvIA0yeW+RGLYFgyYGPSBrh04zwoop9WHac3
3tfrZXj03Vo+KolW4GC3sRmEemXEr6lYwLgW1OQ3sbuXHHGoLicFoLt+D4eC/o9xieX4ROLATuMS
MYz7TPzY9uG8ppNISqFoNrNN2acyzYjKvudWzKA7fmUfg0WMGl3f6EBBe/gVuZSaDjFkg0K3RVrk
b//vcWLidFtefiT2bsBNWdq1CLQkStfe1IscPNCzuoOF6+jyWNRNm5mKHmHHRvR8iwcPBqz0rrfK
Bfn1Sv2QwKaDydsNMD5bv6fwEn5eavLTzWEPuhh2mfIPQEXoYcxFcWnFpDGOmpFYWXQImSZ/tvlK
6NDdb/ErD4xeqoUpiuXJ/5ZyQjk9XSTsaT97lRZdOdfkLjAuYRQniKBx4kscv52e0Jw47RlEUkRy
4qq0FwlYyCP+r3GgDkhj4fUpWaNWyCygP0U9C1uU/AaDL8GQrTH8qWOnVXr4wh/b5rrR8rwQNZoa
r9EH0WbvVvNV0TBgy5nUHWKBp4JvIY5ObhUS8PHPMvR+iHGtVP3OSXcvhd8bVqAJCSUo6eb3+rCe
tsJi61Dolcq8V8KaSc8XwJ1NOn9TfSKruTrgHW4w20t9RlACONSkkV/9LebarHgiTksQ1GxHmgB0
4VbWjCbW6Wg0N9cNMIgQeXqejPILdf3U+HLT+rHO/nuZOG8if1XLN+keLy+m14Tw0aE2BguDP6V5
0mWfgBYI9Ep4EEttGMrljiY+O+PGvO8lunfYFBmA9GBhSR0JSnfyzWj/16TbRJfWgD2PiR5yLfVu
yvMUQ0pYRwtPNtYFfp3/a6/hWR8CjgMDG7H/j3JgCdJU36gN68VzR56axHd5/3Vj8D1SvIfLhIx0
7wvZdCGMWyj6S68t/sd4O8hqb90yq2t1tFEbKRP4NMhAekkBziRA1/4CSxG4H/nh/aERhrYRMdKy
XiRT0CqOK693lamdQQR5eZI4ovM+suKZGWDZY3T9xVlhYqvch2kaKWvh/rTJV5M4H2sIQ9vtKJFY
BdO8HiO5NpWlaeSQ7Iq7fXy6P0TLaKZgOMH/cnOk0xDNeXMI/HY2Wg2ohb1pIKj7RyImzKUlmKdy
2iHpGm5ct3O1yi5G5sa/bG1X8PYB6z6mjWwer5THfCQr+897Z1O/il+qdq/iWq9lb8Vs8Bl3jQbi
3Wwku2B9vB+FrUjwe1uZ3BthPndMcZ6G71sjFuaCaLki6nnIfEYWCprqhGjeNNUuGBmPgzUQ2cwS
f3unbUN+kHR4/YdKCIll7MqqLlaDyQC/HCpVX2vHN6IJSpB2MCHw5kP0xSXMpsxaXEpxH+JdUeTl
GkczY3ZbyxA936R25DugJNlC9o15CcKcFfT5e2waoBbvESiIbSipNQhBiOlmR2R0KRunwQ7ysxBg
d8/aIQhRZHxoswlICLp44DlqqXQ7ztcrgNOP8gY4De/AgLMzswA/sNfa+QpHrdPHhD7T8lgpm42K
W1vTyQ44iAtjQ1CTKxqmWuFPOkApneRDBeA4/DxrDfizACJeg5JchOkD7Oqw8uSaPxcu49XJ7hoC
VotYDhb4RYUGVoZaG9cwJ7vK0M2NaAJhJfH9vkZ9sKdjud451H50A8Cw9C6Xw3HsRwMOFEL4Fc2G
AYNkYfjgt59nggUetrh2gsMbrsJcpGbwgmCZfw0NebhVLy8geyPuia+4K8RSU6U/i4QSbJgefATx
koibnRB119pHXg5B0UmKsi66fAD8I2vcyDJ5tmOwa+wRmzSVC5WrKm+rRepYmWem2a4d4Bev1Tt2
iDH2OFO3QYsQ0hNtPxDZKHfJES3nUeSWypkZTOyNUlbDF3giBzNwwSNqikcIYLys8ZOYZp5uXaq+
OtMHeH99iDHVdVCOdpvWzIy358cUknfyuaGKlYT1QMaZyCqgileZMnZ/FTfK5NOGXCSCa7K9feny
t5zV+7QryRbXA3iqT3b4P7qtVBbPXcZIcd1gtiOUbbocjM1jKLygNr0nH7IkQ612mZRrE0TqPcvA
s83a7UGCP1B3BrzKyjNyMm42ZoZA18rZqOcF37Irvc1JE0a6HKCpCtOp3yuPYuczy6a5jTY937zr
2ahFSwZBUGLcKtwKAiqKpnmNUwk0Fs4Pshl4yqKoW/YIa6pO95Zj8fYyRkJ2WZxO6N9BSLHjn4zs
gvhT/uKjW2JxRCJE96EJVFjUaIgwPnn09VDQitPXOj2rFdNS9UK8gtyMKzrDo2emJMeRyZmSk7JY
vYMgpeyWGSv3Yc1xODzWvj5cCgEeEnFJgM1vomRLTT7idmkPTdrG26gWKUWUIOBZQgZgzbLsBkwI
yPBSNlkoZAUZSfr/9FthZd+edrHUf+TT7L7RiNb1uFHIpSBCVUrtCfM0LUQeTbriSTpi+7wblxsq
Tl1qsDcRYWBwbOlkV80zUNoA50nV12YqWSPpwXliAoig0mTN0cWagczsPefygBx/D4IyX/q18N5q
s4RKJcng7mYdh1U3+CdURGoASBQBXa+5xSG32Jh9/oixb3qx7bt660G67m5shel3YOE8VjR5SqqX
o2LtJfeHBrh2nwWHJhPZPHs4oLAB6cYbhfI0Ny5o+hhtzhuXxmEt7oxVzeqj066bKNZ8eCsVp/Xj
9YeBZbf50QQxdhE4gItmzKyI4p8GJsMaugEndLfG0hXYJzdXx+Dm05Xf01pY6wYbmAbfr167qce2
vFnYkP6UnqirVsognmTebh4Kn2yXOT+2iAhDZAJ4jZO9X/X/AidKLXSizDmLooIvehu93lA4HtCP
uA4XFqWSRmJ+q1WrH3IdZx+c5J8eN+tn9GHE38Qdd9ewOZHyvFcsLEkOtBrvrCnHPlL1R/LzjsXE
/zp2pACv4FuQUa3Uo4NIbtSH4FGbvCiQXio4JjXOb5s6UF/oOnluyUMVBw4hYKL3yhRnCClbrKoE
+TpjKeuWWnZcSws6NpEBR4jnpt3RhuCajS1mB+U1nP7ZTsyI6OV3d7vjT+j8UH/MFOR9Y+Ejodxr
XevR/XF9LZsPuLwtbhd1I3tx2KkcXZH7EVw5PRv81E6PmX4B8pflQgiFm+6e7Gl+SyTc2T3zryo2
M3ueMbdqHz8IMEfsQyiLdQ7WuRH5I4vQATOE07TR9ZNN1jL4DE7n2znkXieSnVP8pAbdVc8Zk6Sh
UKBCzFBA0vYWyELobXuzlEcm+Ylk85I8ldosRBaMNDhr6SXPBJA6jIj/Yr69nw9/JMq9PrUpLPwi
vvpGtRKjF0iVA73qNkoaR8nAgmVXJVAYxgG7lXKUpwE3CZxEv+La334KUAZLl7fXx1Mt2MEeOyBU
GLoq3JbbROVZ+oC/3HnU/CDIiHim6PrLP/i+8Bh9vRn2n6zq7tECjqQ+3y4M0ZYJlKNLP0ldn9hO
pghVD/iYyAUSha2eht3DP0tnvWnj6048wLf8+0wXh7J5xt5SQ93SH7gMui9syadfYJCzwyiQyZ42
VFK2qABW09TIBSlH0SlMSUenslLdweGWhCr22UexvflJOSQFA5/Bz07XIj5cLHKulQ2bi8yfGtx/
o0LJ/wliE3T4XOuZfJ4tIdxnX3EHYoP+3cV8kWVZep4/fhFo4R3npeI1VQ4IMKt77qnMrI0BAMlS
/RZ/6nqNmAv1Rx3IeaKWyIsm4MJ105xriKjteahZn+wIJ+SM5l+710BZTkQXg67kStw5El0rPvXm
sStOC5e1P1mElEbrfibiVQrd6qHEQ07+szV1Kk5W+AeOt0quhZ3YrtVedE/BO0v0VeStv+pNnSpw
Dr/fL9joY++T24qmGKGCVfVgrFrMnBJODk8aNO9NjN6Ayw3ookBxrpuh6N+0R27uRAc4R15Tj9ih
K3BTZEIHAyqNaXiiJZqyChlatZ4SDKgPw+pnWfMIhZ4/ZdoM0VZMhyAxHxcjAKFcpAqkwg0wUxOl
rwBNRqo1yTLfl2E1s71p1hPDFjloE8jVm0aPwlZEZGKIFGt1J+9KnUTRJFV5ZvgSvRE/VNrAZ8fB
Xc6hiRvWcMAzqi0NAhyaWwbklgwLTz2p2B9VlgTZ6lRp786U+uJadwqrRI5IIgEkmgvb/1kD1a75
Cj2xt+x0dAF7Jhy7ETre/ygMvpUhpfAqxuwmECKH4OAh609o8H3GzSfGznxVxYs3kNGBz0a0T+J+
uvE3ksnO7EFmOueci8g6YO1PESXsp1dNIxAouPsi2KOIqGZmMuC7Y1axZwvLxBvmKRfHLr/g/KKl
c41JR25pk1aLR864W6g0lqHw+9EfGhRv9nfxWCSOxArvV5+0opSkR2er2cUt7/f5j5GAEdxaMAQw
M8/qRPZ6dOWPNdNmPsHUaxEbmkdl8fwQIuEoYoyljNI1kGXn7EFdt+N+elUqHUr3HdyKEsXMnOwL
DGwD4+e09Vuo7a1hKlIktnGqugaN/GmfcwM1d5qpNaq9l1CSUAeIdiCS0JT3NRdSSpT2MmN2TIie
M3y9PDVeOzTivNTZd4LpDEmhlXKUTG1Mk/3LJOsXG7yHdNDN/6GfBXxf41ESaScwkLb4tNTgSs3r
SgrNRjWA1s6+Ior6igXRJtblD9aG/PKzbGOOxyRXSGnsxMGQxXkW+6aEt5KRTvJ1g8VEJyXeew/c
dhNsXG5eRJMOfzsZ0N8OlKHUVo9M0q15KeZX4kaTvKH81dHy8xA9kv/avQ79HiVAacXqDOZIv6UF
3tHOSpY78apWWXTCY0f0Fe6qHKQsDVYRLbddnPfg/gkAVRRZeqf+rFkC4/aTh6FTSsAlvd53XLEr
JSKrYNDUdNOPlbRVRSLve6WBz8sexa0dXYlbCIGSaUCefcgGRYd3+gRLGhITD3Yb/dm48pRkW4D5
LudNNASb9dnYcaL9A6xhuGsDH+A+znka+qrZMHvcYABPJhwsTh4MVXWlJYrRsHUlwZ9GhqajEvXr
nBobLsgiPvaEF2cwaaAJ/CnFmIb0d378pwsfw7ryDFJ6YtYJKYM/OA7+psXvYmL5JfF0OWWD7sA7
okyL6DUBxLXz2CrWxxsHid95wB5KVHs4YjQS2AL3LY0k6JVW5r4pLWFPPTQdIg3NDQbFbQxfIYV3
AMjp+L9ze0sVEPxzRGEQwcEQou67RXvl1ETv6JkQPZQ5YNjcAvtQtiPLhABRln5amUkwyayXxtS8
cghf43V0938u3G0hin6UAQ+xpQMW+FPrj4JEaZNS6DnNMjHUOpsKOK+yEaAVjk170ODjz5HfmiUa
93Fx8lhDW660p2JMndoTVed8QVae1PGuQGc0kofVmlrJmsANG65lgO/5JOKeQVpXLX/Hm6rSn4my
+Rjcu6p0oeI8Xjf8HIV/aS3DEIxCLNO91Xv0We8BxHCv/DBfZ9rcqZhParruuhpQStKKfKUPpVvA
lzRTrY4hsSsCj+xThrIS7ctyIRaAtRUw84ljB78FBFVLj4hWQtc3a4zdy0ZLfOio5Km8o0+26VI+
NpYpVGByKnuVTPxMPrekzKXeKlT2NvyQFuXj/kw5sQeoByPsxSyvgnlwW0XzIWk6rkEgmiMGrr5q
NLnlX0sfwzQ65PNLkxXbQeZ8L9AaocF4SQkgP/a7lD/+vAEVkUJAjke0a7ZblKrM5V5UWVOpy1fn
rrGex4m20p/gu8B+gqyUotkjjhBSQdWcFTWIjKlOjNjcXF8VSCjbUXPk4rZI8vu6xe+pcenZF/bR
pCSA0/saSvPCUMIT8o5opDZRrIvezaGldmj3WuQrfj4XVlZkz1eiwIE0mZCaX/1jKySyGWWrz07i
1g7sz5trDwv8nY12+yohlCMzlicCRAkIHrGPhgy5K5WUH7934lmWAHpxp2q00AqF8Qu0SYgJTTPF
SCyRBg4Odll3mmwWBAQ9qmdTmTKoE6vfbcRJkL26ELdGbUhycB3GNY6y7fJCE6c5v4xvcD+Rlvfz
bU2tZNSI9ev+fl/nEg2EgXobpehUSI0YSwx9rMbV+Xt3OwIivH0Z4tMg6kSUBMRM8swH+JRv2Gp3
iCYe1zVf+7JJvJQi5bF/NAL+gMpMrZgsXoBzttnhhCcFFhA63ImSaqSqMYkNaXUrrEhDltOHb6jI
1DJ4tCZnObeQRceTXSVRIUQcMkAFTfWullP0iZ3Gt8PUgFcNj/+UGF1BMpitWDlbzKnTFfhevxl1
HOe3+Ht9S2h4h7Ktc+D7DLwPkDqorouj7rQcuXGGVqnhw7C2zEIIIAmOZJLnjID5GVADYAmPIxfU
vZlHyF+lVgWhDc6Ttt8LAErAPfWjoufICerbmHjd6dLlYlpDAXLWI6rqIRgLzTgXq2Hqzm1ySprj
dIxZiJAPu5bo2dedRqN1bDQ06XiPWIQCZRNCnyL2LpSv8mKByhRtbMJeNUvJZEcWUchbz2TnCRXl
AzqPPTVS3AEjS5Gv+0B1iwO1UWnuWy4Ujkg6MdUYaBUgy0ImOVaPrU19u2UYzvkCck+doc/Joic1
Q1R+oSLg4fhokPMqSeZmThHmAE9g0Fwd/WpIzsjCEi8jd6bz5Vj1TX8hPcQyMmQnFzJ+t9/YJqF9
w6FD8bdg92HbAq10/QQBZKtUaHazf6fzNInBdurX7h7soiLWRb4WhHvGiSTdQxRM9yuGl7C2uycv
7w6JoK27z0uQUDxpsRIckTQ+9moDH54T16aMl60cJk/1gIMvjt/3lX5WaQ5K86XC4c+RhTmSv/G9
CiE4NcpWKmr/eN3ugk3hd4qpNc8YCfndGnE93NPoqdRogeIZPLH6ogkhwgnvaeifrOBRuZxEJxun
n1p6hVjwB6udDRV7LTs2u3BHdgEoO9OZPlFdVSwF4L5ssFc2XovbGASIMPXaHL4ZjAIbSVJpQ/uC
E6Tvvgt09BOsL/qcYgCz4213Er2znyXMSG0Q6TNyAJhMfeJdTtrhhqzgfoi/JqK4fS/nzxP4JcrH
aaQmGf45TaXH3I9CUgox2VrJIVtRhfg+ppfzwQLWdnKE/lPD+Wgd6Sevcxjy5BjV8tuQN6CvO7t/
AZF0bvg23LgF98nH47EbEhavoCj+zSjtw1qO6lpNTFN9tfHBgQWyul/wfj07KGbKtEsaG5BNoCWs
nz+9h/fULRJR4gMT7xGf1ZUpHVAvPoRUED6VeSKLXz9LN0B8MTdkMrhoQHIURsm6YOvlrQydupfd
wEVPQDYA/aXgqW7bNsS6liHg38pmFSNkYppaHmD81dD6ELd0HnpZ6F/et6frVS2WneHa2KjFEu2O
V67xYVQmZR5YW9n2hJHqwScwWH7ZR3YxPmAAgpb2tyZeQYVB3GgDuyueuQOuU2iG0cMd0m0DWxhr
RQUBmBzDXxAzzKDMw1lGTbeTh+vdrWngkzD0z43TqEDl04GwzkP/8hS9atx5wwew7wkQi7ubTlJY
wtUULIbzYoOYqaJnp85DOre5++N/Y1IEb+m9y3z/M/851pK3EoLxBsMHGjMT3dNET1XZjZqTFvnw
DWajgEgZ9zRYLTVuw7faafyHF/2HmGD6EvtLZ+p0DGTpuFY0EF23DgfsPQ56g8x3/l+oZiUz9lSY
DA8bty6i0RVA+lX2aSpK33E6LbVQ1yvPkp7RDQtW7GkPFvBusDTX1l+9DLug42J7cWG7lDk0Z9+K
uiYTrzjwe9Z+r8Sci9tUtiDd8nOWN94/yGG9CY7P4cfLCqHYGS5JecmbsMhXukGDG9HI6jYnjUAR
BQ8Mk6vie/Cx2Sh5W2vsZOmP3d6aUSnhiLD/sK3mdDS8PISDVDdGwd4lwWkHMgXsC6f9aQrUkCha
xpPGjsexvBTpauadPesjSAJZXPeWjz9cZA4QebumA4DJkF0Xjd5AA6N2XBWD/yd+DAb7BW3tKuWH
eEq8Ue712ma0BdQydCw9aHchz9GqoqiV4gmq9Upi0AKAvuCwDpM5e4XskSO2saqIvdudG4Mv/y+Y
2wrRufR3ARzq5RORH+7alUMN+sszgtz5JVOiRlfJlnpAeUycWS8138SbJe/udyj+g88EKhyWv4J1
iCkvOo461+Urdma5yQQtJKzpPPnhP8TQ4viONqNZnn28d/846I9BD/ALIcv2l4D3H23+VrgJCwB2
Qhmu+PCaLNlNfnXz9a8OtFnx94R5CytCXtkhoJusn7tWD8lXA102F+oDizM7rXQS+WAB4yNGxfcE
ipY/xhVZ1/0+/E1Mce4DlvOmZtXARExof6GW32myR48lwm+84TRjaP0YqVCrlWnngv7cRImuNGpm
uO4c6Wr4SoLZ4qOugGyDRGInHnbaMUNEbdxPcNDBbBG7Au07Wo8iFMka5295RsbIDIHBJphxUiX1
8XdCtnLrd2a2tbK9vT/Hni0v6a8O6LnMGVe7gKPK6lQnGdAbdwTWNwaiERZxSKvrau+VGMYBNaUu
dzJSVo0Tvi4OBs2dvzFBpq1QR14sgnMJgZ7itu0EIIb+OhPMkdunnu1yXvUhSS1nD64y/Z0hozus
KV9lrGd50YbUXURhE4YaFvOfzv6DBejiAQVe7qMZQKbSXoxVw6AUtHoWl0A4FwAJ4CRsMv223I4N
d31LvAhH6fF+NISCXUXzq/65cx2AAVmpVdsxLLWSqtNCYtYrhxon2D48MQQce8IZexSg2UflNbFW
MPbIev7a0axNkrYks4qlU7nVo90hcpX/faWxiE+sCtaiY0qvU7xatR65bbWOpdB6+5V5sAj8waBN
ek8wKqTG6DLUeKlwZZBlSQJVROK8a5Wk2ZzvL6L5rMQoOExThDo7N+CTdDMl+QaRLnqqj2Dg75F6
OMmeaDul7w/o3oikGKjcmXLwAIa17fjrCqKEsdbmFYEa8Vdda3bwDP9YVkYvLn8svaht0kyCZ+yw
GW/rEkBq/Ccn2X77iSyTh1Glu2w/a169ibnuxAuIcI6Krcx/rOEILuVNS/zrff6daHlpxLKEqeO3
eol0+ouSluWUdcWtjfwFgRAFGsDtkk8kth2iWqIJVxI90vtn3TBE2cmjEE/u2FX7lxvKX8HcoIpC
UM6R52oRLiox+7ttznIOxE9YwG9D8BO5EAvm5PWlk59MLykmz1bqBCZQR5M2ATytu4qEVOjKBG4O
RcpjOA3Dq0OZK5Fse4TfRLnPWwhmJX0iOqicoDP+V1BD4HJ3TLpzabKVhImKXxK1IgkPqs99D550
1Xn6+b1Gwwna4NRE6cVeG+mbvSnT/a06BIATw9jHUK7jOSz3WUHoq1LPuUnCWkplLp+apff0x7yE
s4XOVEyZPjrUmtDmWS5HgsWyex0N8pZ3FoGD6zWpMU2hmaf3XOVTB3R7URzZv1IcjLxyg6JZ4t7G
ie+iCbJQKOlq+Q+VzAyI7jI5/hE7j1Vsc5lADGjQ5rRY9H9jhQMEWZ2RbfDotQcygwKLfCf/Eg82
QpMFL+rt/CekRhsCwS1RxF7n12PUF4mxVi1Mt27j8t6lIl4tCYdDm5JfQqE/oUDxKkkfR3xJH5yt
cUYA8hllG+wHb7CsApf0veDbgigXeydLI2aTsh/QqatAY6KSy+sNxYjmKYBzm+KGd8pBr8pttaN8
hThxLIK6ndXZDC2FGxPuVWCLcZiRuS+oy9hlJceGJ0HjhnduhvNfQdkBX3exUKvXdyOeZSIX1is2
XcVxCajBp7a6fxSVfWDClT4avbZS/6mDUaP0rHZnKt3Rx5NvkuiGkDPMlSIBs4KqjCxDHcPylyHk
7FN5YW+gxkUAxetlVvopLbqNVhWSOSdQbedwdzwdkoq/69u2qu/ul/kvr32rAS6iuO2bcEdQuyoT
BcoZ4lMKXapPx5WP9rsuowvzrFNe5nIefBXpeqRiHrj3Sl+XROcfqq65EcQqmX44MlBzoHIncA+/
o+5Pi/I0SPuP/o1Io/kA1/AF3/UeHn4RQYU+wY5bKOg8PF2OaOEvnI1tucsRsdKAhfX/XQqMDImx
mqIBY8MUHZIBpstH3TdQ/MU+OJWGRx0ALconr2AEwhFYryui/dTahvO/Vejt/SAYoTdsXdq4Lfhp
q80BIgXsy+hZ+btYeV+XZjgixuL5I55C/SZOonmvrVmHMqCcLoRNOT8JhkXklP5QbC6MeuBFUDc5
PGMm5OYpPXPGzPnAvlf9yRpg0+iGOD+cyzlYnmUb7PB5lNMwNgrXNIqD3DXOC3n9FB50oOYj0YHm
7zNh5zBQ85XU8HB+usD2g53E5p3EbrAkn9eDSJTwv3QR6RAJ5HLrlvWU6qzbcgH5wpVOlz5Vga3O
CiqPTtGqXThRksX4tbrnTYnz6udeDu8eWfmw0nEqU4jb4W8JwE8XlGS1+VFAwUCxYuy+8qdzLNFL
EUjm7yhQOQQvqzqZmYCuO1Ac0lcmcl9Tl27AKRWe7BnYVjB9d+OIHR6wmWMJ6rfpG7IGGer81WMA
g48pKLIVvIljpoJn0u4dsmL0Jre5EC0avnNb7m83WLE9NUTTyVQFSJ5ClvqBVUDXvfsJ2jbZHvpv
VXP62cqQIAfSUnMR45Q+m3/ujCRAid8ads2BE3z9O2yK+fA0Z/qWvEYuB86ZXVFCPrt7ttoKWvrh
hrETcuqnkVzLzkR/pJ1eIWCrhmYC1Mlxcp09EBhs1B/KQYSO+FmPgZCfn4weSkZeDoYGquwcHbvq
f+YGS00/vRyrzjS7dU4hsNYeuX4eNaF+KrWu9WUz81GCZLGWJZkvgAw0VLVtQLojr7+7Ma/JfZQ5
f7ivLr9oKHDI9rcg1UfMMMyrGtjM11RMpTduMXQU5V0u9bcrehC74U73Dfq0EPsdzecKrrNWiUqC
vhKebXQUmpodaleHmbhHXSN1adYC2n1zZnJaDIER+XJLxsU2ZGsR6LRcNcOJx/jI0uDzege4Lunk
emwbYfd1sXy+CXOouArbENP826t2jFqJewEoXkVsLPU4XI/9i5NnhLo7S12jlN+Uj/Kohe4GCG60
BYSpkmZsksiJSQMDuSayNFqLonh05PPhgaz9RmZ5o15tariAZQI8GBNvjs5IhUjA2QsmXU0Dtshd
HVazha99Vwdg71ZA0KlaqUFih8hvNwG/mbWNL2zXieWo4jWnB8mwS8x9imbjeg/w4i1aehQ+ExGq
pIfb+8i0k3Ift4y77uCZ4enJiue1h3UrzhlH4aT9SLO95+8urlGioPK0ljsxJ7k+qbjxqRIj06jT
OQUmPJbgH4IkoP4JWy/Mmc3orXvVDICSbfFO6njG6L/NamgF0j6kQtsj7tlNA8pByhOdMUjMiSPo
s263IqCG2/MTWaK0HjC5NIc55W8HUymrNo+9YSITk3XAdsOiIVpXXnXK942OQHT7BNY84PH7L9ee
sNAlb7LjWyRpSx0kMcEW+LV8bAxcK9EqogTjTjkTz18WOM7x+HdND3doEyVfYgA/UBUUFVUlEiv3
RcH+IFyTDaJ3GIJu9+AIFgWfxewaq+37sz86Kz/6iT7S02oL1LglZ01l7xtjRG/7mljVDEp+7quT
XbaAxhQ3WR+bg/hYKu/FHVsjuMQ0WV0uIN2mb35k1wFmFgxqNR+KLa7utpghszywrnu3Q0/OKhOv
XBjodHWEF3rDiGpPWjWp51vA24Nq3M3URXPydKdoyGmapP5/KQSpp+NdrrnYy4KAe3E7uG+bkNkr
DibAt12JgK+UWJ3AOgPNXJvULaBZ5cZm40z0Mh/dnsAlR3s63hCROO35BuzUVoZMu5F3+CKHOW/x
Rq8BZjYRHeSFNYJS84F31oGQo/epA/le9SunJfZX3k3r5KoQx1Rs/u9ft0oTu9bvYQxnqtoMRXO4
uTJdyU45GnPw/zGCn4xeEI3YPjD1ODyl4l+E5Q1/jxy6coyNlh9zbvmZ9mnSJSOgGSJDOE1yBSGK
kn3MDJ+ON8OzAVWAUp4/11wAvz0bxh0j0xOmYcZYIklxF5PriRbdjJO82HCdI5IgBmFQ456TnENh
wpitC8bal5sRYyJ3XOvPNPNxqXJUkYymweOx/9go4c2YlqgzNu5bWODnpw/7D+ZcMxxE56sU7Nsy
/e33t3ff8LqYf5ZNlNNQ4ZB08TT/2Cb4pXfHcI4htefUHId3hgDIrvDohVMpw1JGsb31z4UcdjWd
kNaET9FSkhJTV7EpASa//tf+oFTmLt+P4qygXQTtYVLntoR+agJQo9U91bs5doSYgshTGeRRSL51
0RoEnt2jtlEi3ZMl9I2kqwO41M+DtFKEBvgjYOxp9zP3V8degzyHxi/L7QHoV5dkdQHhMg2Y5Vh3
axfbzALSow9zxT+da/bwxw1fPfMs4ahZlWcAYysDBYTdiV0BTY+OM5gI8ILyASkjEu2aLbJeLRs7
vSoilg6bZaUdsRhwnYwWrQeZrf8X1YGxY3F4Oqy6eTImU85xQ2x6BAd+lZLJgslPzJVbNEDuz1jL
ornBkU+wGnpnzpu7u2hbenDWkZBiv0FKTMwGXp6Etv/92M7CNbiGwz71QOafxU01q9RhkbBLU+oG
XPfb/VrOoEEdqx8m7qIEAXKDiWgzoJ88XCgsxQNuuDe9qXZS2Xa5WKEb25rzXr3u3yyR6I1y0ZGo
3ykYlSUcinznDTYHwu3uFDCdXyynHGgZp7jNHXDTl1WEARPOyDfq1kM7jWssQBJ+nfHQ8i6c6Ngl
IVNGn6PDXR0aCOrQvF4v1LO+AJRcsCCKchfwHKufc3wW2wgMae40+pc47tODBD7dsPY4WZQkXCcu
TQX+nErYMe61Tr87sJ0PHsOECEVTEB5U1WbE1z2p79A3HeOCy3dCN9wnRscRFWt3fixLLy/OA8fn
uRILbyJyrCXg+6uF+CE9cPPqEyEJhhqV7ce0691pXymIO2X6BuQHlbtTnz//jTjwp0U7cE+hKoRt
GUQvwWBHsMlw1j32omuk3vygb63jv5tbf1iIA2Or3TROKg33oiGnsD4YsJbIpnTGkWv2Q28Fl9sl
aAVRkixkJe/wUn7dPMODpQLUwpJc3PXm0qZ+9RA/jY/v0Ab4u8fdDGEGqwqrUj3b1AKKcxEk3Fkw
TDUrJFytCd9ohp77BoVa6gvWbH6yj3dIZMJjwbQklBXWxEPSW9L0CHKsfHDfo+sDWJ+FbX1RmKkt
nBY+WUcAa33aePWLuzK1MArfePehicDgfF1IUjlvGHpwyognTsf0qMnJ+qf3pvx0/rkeT/sLdanS
0lHqoocNnqP+jSp59StC48tyGEDj/OGsy5QEFLcotBns/CC/OE8HGmdS/kh0SK4t4q53OdDFJ4qY
WA6sddESku7PKs8eAEJ+HrE7uVpluCekzdQGsCPPNaR5VN1RBxMvm9Wx5yDiYLOQEMEzXLpIUA4B
+ZSuiFRp50xownqeNIAReZUvlNlrDQfPnr97/6UXSj0ngI60jx4jy6mn7kcGO0++GoDRQJCPLYu4
fYNDuxjf9wCZ/opDkuCOUREKqYqkVrvQvcUNi0NR9T6HdyE2ROo6bJ13/N6XTnMwJ4EF4rKYJAcD
t68OZVt7I9tAeDWtE/WLJ01J3s70aIIijsFQ/NnWSudcjqEeBiJLb83q/nGu3CEJcTQS4gHXNCOU
flUnWzIf6taIBnFiTfe3+uyYdCH5AxFmRBVAaFe3Bz8aHeKiF817t2fcf5iDjo7KOaZDhFwIWcoJ
JdEx00jh4zNYmAP68xdg5M2CyVLrfhRo8P2dSzPWWPqJCQpdPdcQAdIforqMkl+QhtxyfCTyzpB+
yWZNvir4g/mwab6V83EODV+WCkp8SV13vcN25PV+pYCZN661q6t7rlNMXUHy/vx30e0+D7aqXoyn
KweJdJ7QtUnGRh4hRognEYZXuxf8WnICb/CGFzMVQA7qDJx4zD8eZ+F95op48ZABgXkKB1SfJExS
vBb61dd/Zpn4F2R2tH3rrIFQoalF3FvxCZ0Jpb5hwkHRa8NcmNppQ/pCup3Tqe6wv+7XCucmYttz
CCwrSyB6inCMJ75Gnd2fUM9ofjwKCTLjS1BE90MKG8EohSS+9CaSI5QZ60NfGxRqyVMwPqon2DU6
EqVenlHjjHeS/L4H7Qb5zwJK3SbMVWxXBYUSukT0RRQBJddECsvjy5Lgse8aGTqI0FrZqLgoQlL+
hgbqA5C9Ih3U+RRRZFcrIzMEzqx9mfN4aAYwtSjFSj1srGvrvW+QeBuWGZyVzyV8lfTb/Yh6eVUA
tctw/1FwU0I6CDnNfpw26dFEPdSsLlNu7nLd75PjTQBkZzM3Lj9+0aEEq15Q9P1lKco5XrSdUoCr
md8YJ7MKSWxMWmBEKCINH67oRPJSqyWujAjDcPEIzoOyVovwgfqZrrwPo+dGXaF7wW1FMkCdUCVe
ga9d70mN5Zuo7rA+5Nibafn8hYmYpA7jvMSMCuRsaMiYLTD6C9G1W+I+C53ktEmI3Rdd0Bn6H4jC
t/nAdc0QmhLV5FqKEN8VLMTtv2VZX4rOyZd8ptH6Eo325QSqYaOA+zJarepf3mDvMhwn0Vy4g+LK
YbgDQFm8Yr6p1hx1yQ9UI4LBhdbBIDjGVerWJFlZkpCrBquzvfL8g0Q2wZR34tMiT4aaPjyVRXH6
OLVOGNAPfDa+ZII2SB63Bd8omSHos1f7NRZwmVaLFOzCBal9H7bOmE0tl1bCm1laoBXoyVVOY3BP
FjqC0PXxQRA8yDjftkohq/CVo5b4CREIXbF3rOspdDRNalpXb45NZp3xrBJwYVtRsnEHbNITLzpn
T+Xsf904l7rZ7FeARtC/syLsJq/mafs/DrzNWAarxOpignFA7oJ8emV2i5+sq0akmKdSKSUQzpVa
DYSUlO0RSMbWd0+hLAdR37LNu7s4WRUwS+ILYeJEyxxBTF7RHJTmN+NcG2XBzEPIVmI9xl4wNqpl
nidZAywfBg75zbBEjwTRZoafWQKIMpagqEZS4nDZnepGPYs0XOUrLHqDd1TW3Xjm+InNgKmzF1Iq
3tZiToWVTdXzBbvp9RkHYM+1ttq1qllgQI/i0Hsu3C01d6gC+9scA8NwKZXQsfWNPCd3T1SAL6N/
PBDFMkxRhnnuEMbnCM/BlYmsjHgFLBxeZ7fWzzy2xn7YzTl8a6NUWziJfJm5YhQ0BYcug5vMSmXA
2fAw0NSE5V+MG0P0Yf1D11iWLGuHgUdpayi9uvqMQz0HOY6ZTBfarK4wLH4HyDgDG25lWTgto1zX
hGpoO0pFpL3Hlu8wgXTC2NbVigARCCAusnVH2ri2lWCCD9XlbaOoA2PILhIdROq7BypGL8RMTfms
e+kADytayloBmL2SlaSbroINBQip7D0AEaLIizjgW2uLdFrkUhHoPup48i3EAIbRLvlWfsUceHRH
7MU05VuCFJhBqXaQHwQpvzao6ekvi7sVx77hHgIjuhh0lFF6oc5JRZi6e6xhm+3Kxzr0s9fsZA7w
TgAYsUuFG22/GLw4BJd1HNOvy1E7ZLmCt0Q83OQ+rNzT4CG6nDNP9xpybTfCCIxOxA4ttJZBYN+3
HHhcrNlS36zvqJ3FBeBreXM0j6lJdtyvQvQxLa+gRZU2CEAWnaqp+yRKMp/oSGKIh8UVpecGuIfK
Msz1XPolb99a8FIxAWQeFOI1k09z+16V3Zg4rS7DLNad5tS/NiSDhq92O+nVKkjfFLwlWhWM2+jd
e2YcRib2U/Pv9SaQkwfvffJpMGcmLLuu1kdyxcn55+pyu2ObPsE81Gbjd94YmdcGaJK82evM6Ud9
SZD8cir7/eqFmEBHZ4ZjoJTXR9Zpwy/cerZNvQBWyQEwCWDbmcXGJBJ1TEPtNgHicDVe0oXPU4xO
4G9i0SnXcut3BiMU4ZBJusbj602cm7X+8T6wVywY8e6pOjmNd2fYCtcPsfauBGZNoRkSTnVfly5l
cp+R27UmpG1Bv8h55piNzk0dFEGCmynu9oYQK1LfkbB9lXa8ODrMeuKCQwCk8rLNp/zonLWzAvWN
1Evdq9ZcURTZLYs2dksNrCQIAZzvYSUv6XSu4jhKeXGVrEBnQlD0EYDmJ51GuD4oDLXy03vRY+Nx
j6AtNz77uvqj3+WOwx93tw3R5w9FSMMiw4d7YgsjSUd6irUbiD8w+T+qWmEMAjLSEVV+YsnboT+L
yq1ARr3lRFSwqlPJ3EU2qsgXG9pNMuHbFu2tyF1yj34vB5SCaK0MPZXkq7ufLCzGcbrmJKYcplpg
u7yEe3P9/z/2xLKvHcc/QCGitsuzposQ197CJz59FIxrqDp3LlK2yKcVx5W1XAw2xFCi4Ql/at1K
67x+53orD/oNnbfYwBp46MH+0uAe7dJHjM7L/2Y42CupT0BAS14tzT92b0jf61AAzAePzbeSZypo
QfzgkQ2iV6WF876/9Hgt86kJqAxijjNMWhbjRhU2ImvSYryfsAfGW+/S/9HihQBctBIYQ5LoDw9w
exiBEGtx+3x1fBy1F4AMUE7b4/cnfTSEesjTQKbJ1KLOR0PM4QOdfJnjcidMZkhUjPJbI5tb7el5
oMPZwlYadpVzW/APQsj6zFMJ4ypI7qvttZPofPRHF/nULWcf2g4jYZBzlpz+CymFSj4YZM1fnMbi
y0h2YYQnyzuP8AaOfHhAsA3H4DevKGLRLKbKErC3TmeRay+yeEan6xSU55683hY/22JyH8h24IxC
Sqxw9su7jpsGtwfXN8t6jU1IyVdBoM7M4Zg+QWPz5ziKjF3CrTCWx/5MEO6DFJMllluKX53L7H0/
RlZ5KTnzg5+66NBOAIpVo3IU/zK8mQQfGHbaHgpw7HBDFV+gbauiRzWlQ4c7fLN0M7J2/TF4BFKI
EIaLaf4A18ER49qyhgymMRnKrsypxwR+Gpnu8t22+Ro5Lty2w7Ow+yzfMtwuRbSbyaRmM/lgtP38
sfVByh03zujF7th7ShNXFzXgsej5KCyOmBXajh0qx+AKRswHYleDUUpjw8aCRMZc1SCwuXs9MiM/
6e801XSx7+/QZat1MxODAn63ntWb6wtSODbE8zESxZFApk0ne2fgUInUtIp8JdXn78lI7Y7n6QvS
7+10pg3R7YP5PK/ucLq6oGL8mVrC4hgz+3AAv5YcOdV9Q4vJshQ7L1pFHEu8cDKK3X/Mr2hD/NIk
rKAhnK6QLdj/4BBbeWmj2WE3TgiqhMyBFaHG8kwxHZ1QkKSCmFI6vmJIkD3H5fC7GLkoRXompgUT
Yz0knwOmsEU5VZmw//u71FoOCHgbSKFE/YJHB9RMs1d6Zt74L0j1R0FTVb66gLrvHp+yon2W8bgO
C/IuKS1THRPxT7NRtES42+ELBQ3jIkF90mrv3Pr84tBSzpuWX1r3ErHOwql5ZCBDL93Ra0cnSBRk
yAawzaRyBMmk7y1EXEgshigU3pguYCcpLYhYlEGtyIKCA+avb0r3IP/4Wc6uaECq5+nA4oq8/Zcb
72j48V7LOHil8fyykqZR4HJLNSTe24pA4uQZJPVsDGLdSOqkUuMaxj8BeO/9ELTzl87b1txYA5Bt
zkAH1PWwVOhkVRjXw64GtprsFAXSMTxI46Z3Kv7PawUCAGMI7BHQnx58bhzKBDtAnbzZcgHdenv0
OAIlxYW7d8o6b4AHS4VhCMhrRzbzWV66h9cCUMMHZzPs58HUjgNvOPLhFDGLf828ftIpYkoyrfeU
wOVSGqmAhSG7+1L4dPPiMAQJ4QpVFUIkNcmO6qpLdZDMHIlcURnguNQv6Itcc/WthZqav5rUJvqP
PiCDMwkU5vgj4hY1McjxBEAuodMei53HokrRXHSwnUHxOYpX2LkfYrqo17uVDkIaVyGVYCu3h+El
hBBdO1GlMuOW/dSkR7DMtBYbZRieG0Mf7uxX/+m82cI4lW+Ri9+W6EzR3OBPiSyA2rGRABvc4ReP
RLpbn0LOm9YBguH9SNtwwQggpE+go6HayOSr1HsMNhOzC0OCw92mWmKAxgT3yb523LTJaF0RgKc8
ut12pyMKm1hxY9HewwmmmnzI1MRiWNR4Gak/WPkUVNI/9RmdkK/m3sevG5DVW83oGTWkLn3YCklk
N5ozynNARXnJLijRoI2460aIJes1CaflfukKqEhLQU1Z/yur0GvlLvvW/gEq/hFvLBc32m3VIMOt
rICsvuexTgcT9EMcGHEoWfE97f7dw4Jk2yNZ1Diei94u0xO9jD28sCW3NQjTeRKrIE6v0V3QiGYz
h5rKPVL7yAQFTUlWzA6sTeH67Yr/0dS+lUrVUov+jNgZ4B5/XUlewALUvNKohQQxQybrIwsVDC+x
mUo046c/4Uz9HZ12IyN+K0dk2BeFAVuNEEDo3tOyL4IF/JSXvgCHRKanAnMg6HuZRYvJgNS4yNGu
EPKdw39eA09xcWfvOP0sT/SoIsbz5g7CaYfkx3IjzfnLcc/SlGq1La7mY4AwNB40Tz+r+ZtQuzk1
fIMb3Q+iPNwCt2mww+1C1Y+5Q+pFnrc4ZhciaWkTNX/yDWREJ6vc/NfxlF0YSEh02aPurVa+8PBI
F+YgBO8m0XYwRdLuxGH0aEprF7Gxoy4sfwMtB+PTw/btgCkPOuGKmxEVp/xY5mVYfNpPSth0Ykly
naulmDwEk8X9QR+/gNd0aEWOebDsZD/pacsFxVuq4q7x66GNVdsN6c86bHVolzacTuUU4+zwIr/Z
CbnvDlbRrvwXRFiL/l8KMLKxQwKDznhv79LzP/Hs4Oas69WRTXRmA/kQntS3hH1qyRuWPHkM9FF3
h+BZn5fSDPL6AaePwejbLeebC8kclbnxIBoRXr3A3kHhEWyMtHCxQzUT6u5jawyqrMbUASMq7mUZ
SVnIgjVmbLV6cPgEA986QDvlWlr1BmwpjoaoVj0qEPsKZyrIKm+0wmSv2LaWpw0n/3OXIZD62t0c
wNlj39wmbmEYo1yPOM3myi5LargSVYMEnv7mhok58PSdoFg4mFqhc3qpFGH/ymKrR8PyMHvD5gdD
GcGOTi0NUm9QK+qTAB2l2nH0qKadyjKi88bmJTTmD9t0DsDrsa7XIXomXYmVe0oEcnJYeOhFrhBO
Se3qMLaFvl4IxNGEfRuo85PSej2oODzT9iOS/TeIGXdk9AVIARDzOL4tit+TqhGSSflSipJy4t+P
0qLuzsVLcg5+vClzlu67VOPQpqhOBX4wVVY39thtLg/GJaTTTQS09vABSk/Ee8cfOXRSRiAPgjuB
9Xb6sMibVGIUpSyFY1W/RtfX000KRuGMoLOJ2F0/bHfiLP4+QnBCraywR+RlF3OuB3tpQ3dc6yj9
xBsh7iqnQIiILJKjOjg3QKFpB0HFDVfHiHyx8/Jx+jo3uHAJh8FokBPotzMjfsJ7Km6t3HfPAwKA
XNXi1idckqliVdtxH+edxL4kPeeOwdLQO8RniXSlRio+k/q1Z9t/NUmz5boP2N0MUhh6GrGGPfK2
j1GLeVehEYsRm6sf+7iYFyBYcbLTjNndbFIinD9qGHjJfVRvf2yJxLaQudD/HWXfsCGSc4E4nNk5
Gimrv+Dw+TLQIOH2rAst048P7pBmbNTAJ8vjTYMruEHwOgmJMKQeTpXYnBGBYF5TUVByDOXg80IQ
IkQeQkyeCen66bQWCMZWOUU+2WxHDH42s6CWrcsCtrSdAuWBOfQ1jiUOeuPgRDDMmgPwFQRjUSCn
RTuaD/bj7z3DNhr8uasLfszo8rp1Cxj4bCt3sS85Eq8TFRl7x3+Qofg15uW5p+c1xYBDKyV9IvZ3
p3/11rHhMHH6N6ZPTHVCSU7FtT7fqGA75j6LZQz8lV68hSPw0cOI0OC0mbC6Z8y7DFDDslDgiErK
I9Ec4Bvg4ZuIHAD3yQiH+mRs8X4s8NTol7acV4iqjvqBnFsNiLvm4SRBtnhJHQS+RPdKdQto+xe7
V46TiJIwTS01N0llZa9hFU33lmIowlTYacewgj20mx6gIu18pSde9Kseow+9dgV2bHFnIUDkAMHK
kof8I3dLpmiQHpJhqrqtF1Uvc2f5uYGt/GRxqRYP2hlaVamBRkhakfbXZL+n3shGmWeH090ht395
WcxsNpFSPjIcYbjoj2PBNJ/zyWLdud0Isz6D7VKfw1k/5VFx4hQGXjxEoz+kwXRNs2CsYEooOmKn
UMbUzVOmHwfynAnBDsejc9EkOExOWh6mK3y9JnmC054f1C8PjQoaKCUbCs9+TYSyvN1RN31dlD8T
/EGsL+DrlnOAGWOOI0A35dGNICD8PfQsrg4d/qvUEvwhR+tRbcgwIUC+/TaK6VqKBKmkQGkSdcW3
MVablgKyuFIX13+rwxRwftceY4gq+JbMVFqQfsqVeVydplCZAps8PF3UdOhXm3D3+gKugfOR12ty
/cL3TtJC+iDwaAlFpC/MsiTnaQnl3LHi62VDa2Yw1MKuSBzD4KBuxo+qonlgUnHNhfeiBZdYHk/s
QRMGjD6yx6l6YtN7Plj7cw5d3ZI0CgsV8hI95x+8icr03RVQminTSJyitNRnFz95/XdrtAtsrsOU
tbYgrTR4t/1bSYqwU4DGK3vuhZ+7zDeXeN3yoMYzq2sA0CsPWYUl0NUy7xYoeQUf6JeZCKLHE0ne
RX3S2nu71U4vQp8gg7pxOW3+OaV0shcC08GUmGQlzZOBrxw6qojosWx4Gr5+4siEMAXddeUV582q
c+s9GExhs4E5M/O87eh3daX85W+7S4f8yupvbMCdtqusSRCbZiEuwQNGfhRnYk5A4w1YQocI/nng
8j/BE8bVRgAaZpxzw+XN3qSKt062mZAzCJDQGqu91apA36aAvunlKH753e4zTfbjeYo27LdAYKqB
RkJUfGFgesLoNfQA8a4hDMcUxBkRqKwTe7P7Z34O0o2oMpG+FmPXKWoirNhuEYEoqjnwYlespZ8d
U8EOPKk085x8v1IfnCQ3X1n+ZpcEpfLigcZ7hKYedzREuk/hdo7o1rAPUz57jhFZWzs894HadMxq
S3AUfCGdhR6sOHcOh93ArRSTYsAj32V3jMV4nhBVXdG4NVJ6SlLLv7L9GK2Ke/pJMRU70FnXTIuW
UP+9i3t5lF+borVjsBzxJBzzlhZbTSl70Zmu+A58w+S/nYmX6GNST4srUDf73ZSUkEgoGiXEhGgL
Qfb2wWfpdCNEE/b6U0BEaan1cX6FKnIlRcsGeX1ILGFYMCtMjCKz5HVZ6g9DXSsbpnTYkkNxVd9l
Ruul6MtyYSDnNx3fIBNfOqO6NZwY0YVixWcfzlQccTK8d+qWpL2g5s7RIpvT7vS6VntLUO6kPuzn
bjkU+Vg/DUqzoyz9LN6r0DUo9oGhjF0XW9xbesFKnrWNsJuyccofbmT41cu8PFCKTjNItjwZF1wF
IInH1/73eSqpjqppOy7yrsCrRD4qGyY50U98UH6y1v1CQa11wB1Ou7BcXmKF+eZtpwFcW0a9Gf/S
khxW0SOU9maINhlGuelqbZSFjxiiVJH4YXt1ZOsncc7AyRP/ubXkgQuAMZKMZyfZYhHrEJQ1mpOT
4j+n4nR4fZBmE6TqrTW2REordDgC7oyvCZVFptZQjfxThNlLRw0mOI8f7O0Uzi3KL2RevSN6lx3W
RyVH12sAZPNdTPH2TPdjR/oNvmhAVV8uZBEmIdmZf1ZBiNvYh+8ZE2kVRzP9kouKz4IehWqbEb8m
yMa0b53mLy0E43Xw4BkIBAppsx6QhfE4w/NrXgH5tabbpnE3mrgQhYgeFfqDsmFva36p+DxfzhjM
0r/0Kf5DbT1XmvaplPymO6SAR2mjliVe5C4tj/SCiDK8FdLqU5ajl7JLLye4OgoG2jDmZoFqCoBh
9+NwWGKA9DX0GnNLQkjN2mNoWxmzOtMAC4493jdcTz+wFai9K5gSdO/vpReZhmttkGBGM4mNYc9g
8JIfFsNf3x70jxV91m2MTxzmvM4zK938ig7T61EUMVw7K1ULqWl9C2xAGqvPlhY/h2iUBhbolaSs
PUzEn43nPERXiw7hEK2oPO2VtdjBLbZITwsOxQ3BCkS9B2ib3c06Qn8lonpaD9DE0lkQ8F7Ueeo7
SKKWUv1y0e5VKwKumL5CNV6L83nejekSgBo+zxobd5Haz27nPfCmbhu4Gd/9gIhz18WpVLl3Hn+O
P9BzRLOSRkol9ur7qdNSEa4uKWea3I0peTfCxkf78I+31NZlX+HPTqaIZnVDB79TIJfg2UgcetaM
mE3XS/zacahysieffE4ZON7Hb39B01e8IhO/nxFK0ulpOMC8jVxm0p26t5WBN8RF6gEC5D2tU82T
bJgDdXgSXae1jEe4P2O4wgkXrg8UTRixOn8qqOE4EEcaLUkWphqXN/zNFTuuSaYncYrnrN4uk34v
Zo9+nU9+7ZjgMAKElv3BCmxAA+z5qxotvExHHQpHZKBEOOX/Sn5sp+zRnycZtsxzPefavjP7iSaw
Lz0YoHrMXoIcDJWbY5UJnhRHQtNAALFfJ5kIbbotQmC5p6E5Baz1DR5QtDwLbrinu8PZZj9sXe8c
nDBCDm8NdX8r2ZGEQVRrTrTdZvZH6WiVrjz175eiuR0lOcen3B9KR21IBZH2PrY+jaOjU07Hxbkm
3RkJS00AOJ2PfWQ3hAretKkdjl/YhTue17aVSEK+zbwZrKp9y7yR/Mwe2mD5W0uJhrwaBN8jqrDU
0jQtF2+niS567W1bTY+jqakbr2Ih0fEomUe811L4ewZP+uvYN6yK5CWLC9ljnp99iRY8Iv0Ncw9+
ORSzWACfP2lEeVhCm9byYUdky++LvUdR5Ef50pZnxhRBqrzwKWjakjq1reQPxC833xpaLV+t9uFr
PG/kVDiGL7mtnCiY2gALKNTwByZq8oo4sUUuO4n0jYX32AtWl0SIBo4ctZ0DtXCqsnpPlq/sESVA
uvLJWh4L68mchmf7vd3ZgP5h6SIwlHqaqFkjFsmE8SFog2HvSmAJHtqJB4MuGFJvn0vTy0Z0tnSx
QRLUusA/14yDcdsvLTOaG8MHaPdCK5ltM6gGTZSSgtyl+saQmqes3QGTObZaoJ+lnDsjMP6KhrlW
qR0HWgDHnbkM5ykyETwX019J7ehhIBXu3v+slE+jCHwyTw8x1gInlCPgF0PgYwWTO1/ijn5Ydw3S
HX44kf3LunCywIP7qykxQ3ol+E3yXAMTvhbC1mFIY/3TI6X5+vF1msHQUobQHKlqbYoMIcdmZusQ
KJhht7PULDp6Xz4XWeQauysfXkMbHgIsbJ+XfsK3ckQ+NMf0hw42I50BFxq1Iheflfq5S5Vy1EUA
KWbq25fyRsb8EFCvNqLvzuMankjGcBk4HKCESKSFlZ3huro1IriJzgTtYAqxDpV4OwnNzAtLFmCE
iI3EdhIw1T2Q98lwPHOttnrmml/BHSEyXdp/rWU11PUXR5dOA70/GApHDUbj6cSMqCkXc8B32Vpv
27wy5YnRn5YjsTej4yym4zRw7gx1HSsZpMGgxxcLM23MPAAHmJ1jpmbMimIqR/KJaMF8pbH3HIHd
9t+m/6Gy619AYJK9HLZJmmm5r+rqXlRqL/YMeV29z0d5owGyxr2dMWPO7O02KtsXEHIprh34KkMh
h4iXKDmAFL/F4iCQbdZSassGXJYe01VUNTTgUJxEAaAM2QzUVhCfuSc+QNIpr1E/plm8fJNern2n
pRx2wFYsXrCRDu0eNcF8xHXZ/php4bZCI3lH4g7ds3taAOhjb0PuDqlaZOs1sAwLlQGP+tcR2vXb
Am44BbzU6Y0/6KUdNXMDb/pyawOMaAOKaczNIFv6ZXU5AnHUyj+m0vfcedhFiXcf1HmoN1ms+EuZ
rpLpVtDjsVhPsVpK5DdWMt8vrlPq5bG41aAs+2XCKOfNl9hcrlfOMa0NtMojnaKnWB92mI/uuQWL
UJ2x2UWR6Y+umMbZK2ac8hDmBNavVPCFGkk0NZqwoELuNMI2pmq1vS6ZVjzQzf0WxOU1fmX68zMo
kFcs8nBc0fhAc02e5sPqun8C95SGDQOBAmu+wLM//IW3/EKqI6thmSlkLd+4Aaqe9jCoHq2d5Zxz
HtGL1UZdnUiKF4yMnxjbCZ5EMMpy4Pzkx+X6QI8nUBJV5mU9talV0PGqLJt/Raa/6+/Al+gav2Q7
7lcSMmh26ie+V8Vh/P/kcZraA3CxOU3Aeo4nFv/m6MJBQRi45w8oapCSoPyqhR8cTCMeigFRa7y/
24uNZUlEI8ckf/PJiqMTJkWxvLeCC1ZwT8sKRtxKrtnVe771aodJjTINk/t9M0MAgWBmc+BVbfiu
Ph6opaqj7jwjd3Iee+0MNj7s7RZfl5/4hvp0UwHj3BH+wDoqrzqiUf9kCu8LBS6dh5EUfLO9TRA7
W7IKR2xUcuK5YZs66gONXePBn+ndWZUofPm3u3X6KyNdKdBclfA3ZNzmF+sdM1XE0IK593FvHW75
ojaCxPZhLKDY1VmevOIXSW20/qNh/YmVuxd56Z3lJkPBKJgCi1rO+MTrvoTZXASzedBQ6uaXBeEp
Hrsxzo7TKBR1GgL30YfIZPO1lmIcV6SJO3s9DQfsN/dXs1K0A+Nnngg++cIXANWVmKKpAAQ1JRhu
rmoPUOsWcnMzD3OT+bmJ+CjbsxtkHDM4nUULuxX2flZolRvCBD9kv5iMBk5/hEDXUAYSQW2ezKCN
3BOkc6HGUYuNK/UA1+O9LwCOmBV2Bm6MAW0eezcM8lhdHk6wfz0I3xlhLl93tneZhrNoSEhffwLl
ydEm5XZXw0PdJUvuVl78fNq/OaY82/LdYd/Cnm8UNNOSICUdIaYcqO/bREjHeMsF1vF+Em93ArHT
GZX26tx3/O0987DWnHWsgLKenL0l8AiJACFfFTQi5W1HssO3pJ0RRcZeNYKj+AjUeyElZgX2Mah1
sXzi1q8mm3haBAMz6DkiOJ5re8fWEvWEXOC66RnS647z/jpwS+7hoiyGkCkcyWN85XColzrQveQc
DWKyfbIhqOubADjniAgJpWT8JYUHQD4tWke26d0RvKC8kAjI3x8cvxc5ZPoqG/quEKZD59071CUv
OwpLeTNWgUssARXDsJqDEfejy2X6gt/mC2n8u7lxJBc1ug6VHuCikMFLPQqDTK5Wa6qWlAMrP1AK
KWXCDEUqGrISf/oPj/0cSAfK7OQ8t8jClUc9NpVa1fg4g8YSorryas+3GpTBjnB2VpJHtw8I9NX0
5rUlFzR5UyNog22Koj+d4lBg//WRoJuBJ86gwRuJMqORgGw+MjXHW6FM4nhHMSCAlAnca7h1fUbw
/Rsb449K8RFEJie2DJUG1mmcULfZmbKGTm5EEip10rLg3aYdFZCRR5iHORMc+6+8GKHqc91kWsrZ
bY+XJsLzz7cx2lwFLOT8u3ElmtpJ0oG//8jGfUKrY4NI4ICEfrJXwOexiSbXv9MNBX+Y1wRaGDrI
4zoH64RYOh6+/rzR/ElLEwkzuZyGg8vVJ0VEwZdDWIeUCWaVaU2i1XHUaVBNi+Vixgt7+1zAnv0g
y4+9YfIt0a7AG0t+LWZUIz5eSCz2FNsKwNvhjHXYC0Ajv6xyA8SRyQJP+WO9gsqnw/tG7GeKCtFb
1MC3W5Uybf8tKP444ahmvvJda5ulNjx/NyAN6peYEmbez8m70qEYZCNQDEMAqoaOIzp6noKmsY7x
2X+3uHvP5G3qt897VYk3YZz4Z4y/LtLPSFy0diFTL+4xnPGmxHfzPjCIdZz027P7zTh3ZvWkYg0o
Z2c2/4v8x1goNG2YEl+R5BNsf35hM7qxM2/sMsIqJnACvly43QGh7II8XycgWoMO8PV6+5XsvoG9
DD7bGLtnHTKkGM9nYkJrxFr5WzWf9mdxeqALfsCchLEBCjg3mKm4E+F860BFc6DXuVdQ8tbUVdqL
AxnvEZhldlWVXUNcvYEfaqzhvVBnBbcScb4PO83caqMXxzmD6Zs9b3cSb+koCphOIrpY2YQuA12t
gZQsBcCUvDYOKTvZmCaFQqdA8n0ZhNFZWtubcJ76xFSXIgNWVi6Vju+N+Oy8k3B+cMYeBFpPiMeS
xAFT4OafHi4PYUl+c61mztWm9QdpSphSrWlOE/X5O0C15szLbaSySKDaBq1SmJLug0N95yT1iQ7a
xhuBCZXeMg8MhudxFDodZ+cUwLVPihOoppBZiEVJqqybsQC0Z84YQDCE/pZHx+VPaimzdK6bbrpH
mrSGpstaUL4kIceKdDPLEjuTR7P1qupeahrz/iRLPgEIbq77cjjKacJcK6GJfaBredoN4vcczy9u
Jo0QLftYT65M6J9gk9HNw7egmxODTvrWe/vQEI3ZuXMS6h6NufT74U5tM8q/dNyrSjpJ6jrx6jIj
S/vwVBgI6UVq7hOO3h/8w616rXQT1ZbFT7NGooBNnP6Ky361cChoFczDnsDyFVqXmoxDC/n2dLvW
PDdImyos7iajQXRIDlS3NylbZnXocCwSh+LXX04EcxNx0hK9208DFKKy0j9vad9xEyISmJrI2HzW
OpoOUt15ioIj2OF5gO1hKvBeFEMVf+pqiYqrJIQLYFbW0G+gYQK4AHtvbpXQxzzLNeRvLA1VH7iC
3qC35n2ije64JblFs8QuM6jwFSeB04kmAzT67GRBkuUXVHH/zTgpY0TF4CRrA2KFdk/gsxpUYGbU
DnmWteapTO8M2g+eA4keI6BUZokp6TP5nJogRY+npYkhl/HD2LtWwZ8MkcWWLuaxiSbqoIMhkvOm
wTAVVjNaCIfpzVfk7GjDK7gfgq865qv50gwlcriJhvkrU7AVplarg80XrGUzJIQQMYu7zm5f/HGp
vz7oKqxbMSEw+8xLB9QG05kPV0EuSVNA5HANRX8sTC9zCIMvzQDcawnbRbJpoIF5EnJL6eFGjLOM
dxnKYioHb6g0WBVpe723vAjCs4mvxm9rH/rSCGtwykScxsjNc6Z3wZ7t0SsKtxoESv5i3O5qwLPz
aZjoode2KktV2SV7q3DshEMAK3jclp8cB5DsLVJuVs5Oxqzm9uhlOHU/SAFmCwvVBQfL/TMWPWxn
ffN764MBm/xx/SbnfC0TYl6vyUtftXhN+HucuW9MNX6+zYtlG9u8Tj8Vv8JbVc8woZZtIViD+/FG
rP5jTxECki/lroZjx6Y4aKvjj/tMehrriPb3Rrn1wz28FUGvFZLFS/OZjUXih2Tm/PEz8EdLh3Pm
kOmJ9ik+KIVMtRp2h14JY/UvoJwl8Vvk5gDa7NPv1hBARvz5WXd/ZL9DQz/2IH1l6ChRogNw5wYT
M10920n8E3uJqAvoymSZExmTH9ONb/dGdrfgoVRVEqswpa73A0C59NRo+EyMxjOzzpa3ipd38mtH
CFLjD69SWmL+RZnGHLfp4PC5lESDIqf8nUMALAZcH5GD+ojT9ib3zAsINwMnly6baWCd6QWzz8kt
fC83Jk/jhDi+AJ13jJkexCs2L524oqFtPuf1Dn9x9H7+rWPQdVIfbobKrx+7xl0hKmVamQPJAT/l
m9QmtiHgr1SpPn8REf1IX0LiOz+iCW45rQ2AXy+DmSd4xe/dfr/jFaMCtfFfPMXu68p8hPnT8FZK
7188OpYee6MMllfPTp5f6FigUpQ6cAP4QSRvsP6iFBuppTNjRIFGRePVT4egH9/ybd+jJYFkaMJX
CWahGxjowtmp2hRGSUoY/dD1Y7wICs7E+O6pn6+qZWOEIUSqYb6YK+Ii8xY/w7z74hBm0Ml2sup7
JIgaGcgZ1/vTGJVuZOux3wnxaeUetLequSekf0kG7EBMgLRXy/8kNToaEQ7qmunJzyziyoGMCGer
k7WE6ivulM/JEruub07tpol+7UF7Qlj8W/+u0ZgpEzgvLuUhRTnIMJ5OZ0D4T0npjpnaXtK1h3pu
sV4rPbUMs7c5bfLN1EfSVN4uRkuGutT1Gpe698boD70f9JWqlUf931t4uEGk/ApLD6/5hFIqXOZk
HKv5GlLWxVDUjOV4LggmSjYPZ29hZ6wDc4VQoym7JCHE73os3FbjkVxC7UMWHek8LRjo9w4ICv9/
1d/UdJOf+/IsK42FH9/zCue020UoX930HEpkCm0WfCGjRLhtSVVc2XfdqxZBRUIxfgLkj2kmUZFu
+/+QYS/f9leytMzl+1SRz0JIvkVYkahadnIHkwIb8+TkjwCu/vdkkpxIP/lnkCTVEBzif5yFKpky
Q3H0vcY/uEXZxtI/bBdZfzw7LpawPOJWC6OczLQZKh59ceKo1NYmSAFBI055lPgUBnbwvkfJQF/q
p2WIZ2FitKOyTZEvT0iYZiQuGWE+6Fv2MeNpN3WpZqw/JBbf6z7aA/FldBGKg+oU3XWNEI5DxmO5
aAqwpoiaXQ7LyIwdd04p2U//XuA/p9y2NQjW0X/46FBxcpZ08+tkzlN+2ed8k+xZmoQ5WAc8wetf
0DEnYkJbRfGXTdst8pM6CWSE+S0Oah8lHKXs9V1UXKSzVyZcc0gnACf1w73nt/3HosSVOszWOQ2v
xAh90Z8k/ZM9VCLjuDwV1axnkGKO3WNP0FjXJ7VxJykDWJVY28/2t5zg9B68TOpzmG6lvvfx6xKr
Ft+oJfD2Mdnt8x1m0X2JPTRiVo/bX0Zw+mauNst9/vRtsR2OKo7acAz7FoZWHp1y7p54OtEhEvIH
GY+5pDJybKYEy7k0z31JBN8+l8kHIw5J9RiW9L0gds3+fSSG+nqcAFe1h04Z7iLfkT6lQe3ub6Io
tG3lmeW+LMf1qs52H2QZf5G7e7CHUibyeNAXqlcVxk2k/6bnAd5Vp/5Q9wafq5V2EB3vhhc0Ete0
ytzso6B6UTOYYQGXumZzktZ3yU4IAp0qbrNm9hNftodWDjaauwmIkv467pxbH/0OB9KJBcsopwOe
s8UJoXTUUsdWml8z7LtR7ZMieja77XNYQq5Ud8RJv/2eseGf6HXrSDS7uuP84qTBGHTPaPUmDba5
Y/fSVoZnLB3YDvH/06SDJS2yTdh+iMJRdYUQd+TLYWrMinymi9u2vPhCQIHHKCqaUu07oux/7247
Vl4jn31bxsDlVtfdLWL1l82pTez1eS7K1b6qikYeV+AFTyKdOyJqCjjntX8Q3OaI9biZ9K3YI0Ny
SzcbuMXgMEfsLkvXMW3kaGh33adh5+S9USAh5DOwWtIP6Jxi9csPSlPcdjgjJkGu5+HDY649JoVO
vie6EQG1UefxD6dWZQi8TT6onGmoW0kaowTflOz3SEw42bILD7zgnA02qr4XzBzoWIOPMZlQYQba
yF9lt25vTGf345eWAxmHnfBsP9Ii7eZJTKn/UIqLfBETn/Sg0+eOMd0u9q7f4zzgTyHGuHjwXP8K
WietdHv4FixPbRQkHOh222EsYuhHgJ8MJSp79ooQjXdaTb1nXcpi5cGz/yIZe6GkLsVWXTS8ZoqW
VZD3BOiuIvRt322MB69onyu9DoPSzPyWTu0GRkKQvRP1olroIDasMB9kOjKsl36O6IlPYQsCS6p4
Ds7LFaaxVWHBzBa0sdiXSLAWW271z/0eToF26z/BLvOhTaObwghZE6DJy1Co3s2mOZKSSRUGszOK
jM+tFyT09+1o2IXPrS5bTfBft9PdwXQ20eL5D1efEEyMKpfDyToxcQpFPlPDU8jNt1KK5qUhESjt
javgTQ5XILUz72pioKPl5oVCvsGp+emPWU7CrpNU3ao/lEcClbk2UWgyN/CDBUZIOUgIYJKfSf3V
T71r8Of5emwO6hpH3+E92QWOVcQVKUN+3BVwXagt/8OLrpguqPa1wsls2Zyt1iVk8RwAkEFgaUWb
hN7mIahumgxmLh/ziSrfkyNajxrSIMcrb2m227agT39lFw33QUaaaui+GFa8pti0BII4zx78VcbN
CYFDPM3YqI2ndHOzGI11oAwklBW6ofdS5t+qAbmrOp/C4zHqDO5ybfYG1dPs2PeP+hWXjlbneufZ
5saRQ3csG5Y1nDxme2FlZa0/n9CxgtXA7adceMeJxhFdLgdenTYQvHdvZJLushg17FDOZcOpGs3x
Ug9XYA72ppFgnxE9rKx+aZ2PTbjK3KvIlARsdt/ZdVYKLcEcMHt3npB4VijqofJf47zx65acmOJ7
4vzpjyk6tbOFO+icWX1uw7fLUXXOAC5R9+5xaH0SSP3jbifLo1rL6mS7LtVU3S/z8YkswaLoaXYm
VzABMCxkDhnJndTr0t0a2bKjZARCTb062213Poq9tIR4WHxqr5kBonNhU3U7lLZB13eD/XZLBkYE
8aHCBskonze0dO3DoVHX2+FxKWejfovL+fLwT6MGDGRxVqseC7/BVFU1f7b2I55nvjYqShOCn5SA
7ykFwpX6LhCmOD1R3O/GxNm+Xv1jLqr3B0coYjHR+pib8psbZ7TlB8vlnybHj97tVZm6U6rys/tE
e77jC9JnjSiA9gmyxuJPpYf2xDyw6VsGrlZENN9YeVmWuSWuErEmwlMlLbVNRnKQ3dyxVsuGHzPh
2wsoz1fe2AVFp7yc7ZgfR7+k2PXt0BA+yonPgxYAER/glFWbA4tjI/UbnAgGH/mvmkLztRJjxy1U
WaV/q7bHxVsY102te5BR/inn9a8XN3f7lxySiWGXoVe3X3bdI076PVZephIyePUh/96jxHjVoo9D
wdSZZeWXcqW2AmQyM9v8QVk0tMBMxC3+rFttT5nh9DNswirJysa8LF+CpZ4AeCvg3uYByBFd0zsM
BWwe9oXipGAHeAKU4ifzbPdzinbd1mXmjsSgHmtRGK2ebRXDOd0ArYxS/WsihyWobkCOS4qGnw+2
KbnmbDKwDAg4TvvkrkcKDTqj/M3z9f8TpiEbphSeq1o6z7p6NGNSOMIVacL+6Z6SXSRAVYis8dif
Kd4fct0/t2b/KGMWItBTUO6ClJlXJ+leIAI8dypbatr1EAqRozRNUssfr1tFmjZlw2eGC1hKIcX5
2IcwVqTZN0GUMTaVtjL4P4aTGs/Py6BLYD1fe5HJtTr7ANrwQ3H5ZVQ4CEJXRvpXU3k5I0NnzJuP
Oc2nXBPLFNrWj03iaQL5L62aPsf6sKbqzDSEmeQoURCuMRmNO+gzW+GKydD497oF6vTqyf5WzDM2
MWQzxvLltcNpgclT8VUMxjO5fcYUGhc3o0vAeyDHKDPQBBqU3SpYr4J7UwP9sHPGJ1iI1sHf1D0j
zcITp4x14mLHyNzLKhfYL2yLSk9/pV9v3lawktRrIbsY5W2iSGr3PHjBYYZJsLR7eNPJCYPKQZR0
ZTvR/GEe7UQS8cdynk+7BpnzGxxUrdHjYQdjYOLYYDpu5OCHmViMYb8wE0hDcpdP/I3a+SXcZBa8
30nLsd4zshGczThRsHCOmz8mz+v38s6g3Xo6ly9xMteIGUh8mi9WrHCB290w4JxIr/6kOU+gSlw9
GltPJ00B05UOyule6KjNnK7fsbyH8Vbf55y/tixsYFqLGxWxld5xS2hdYOeiJDg4XkzkfczvJnVL
XAi//fWsKUMQMY6bMK/WoaSqckOpoNF0lxpTMxEHlceaKtMr/V8+T2AU9h/EGaHr/XbXFTJu1wRH
sStmwCjy6Fm0RpO+haq5Pf77D8khFotQGtgbvK8eZn5pJKSjWGK99Y4jzemSZlpraiDttGcVmlVX
IIXP3O7a97D3IXXdXfNg6W6t86t33K5DRrXSum2oVVKuKq5oGE+fNLkof5RSLVvWtgxm7NO64oTj
5wZClOIOx3qz6gmF0m6NXvlL1obmPBClRHM0U/IGa/BM8QYP7mKV+C1gQtWEySvNmA/bs5R/+So8
qkXhlQx6M9l5J8GnqtKy2X5LljSRVuxGvT4SpnGsSit5ybppG3JmDYAf4tzWnriBK/s9Nmrk9n76
BirptsKl+dfZfCUOY500YjlXgHSZIna67MrfGvUiIJXVwGOlS3sUMjSEyeiEWagKs4wH6CbesyS2
v3JuOhYyFgcqop2tI7duiQRMxET0oiQ+r2g+R6C2hbhoIzrdRiKYqAi815JFN8g6apMSOlbKhJ2Z
9hZcf+PEWDyimjZrFT8OXlplCpFtLqbWCe52IkIXGN4I4e2nDXLGv4mnl8VyG4JnUDm6UzKFyO5c
pTaTHVR8+YAcRrhAh7Ah2pu9/e0S+VCn8cJL2KBb2dUs2le6V1Zu4MkYfCsP1c9XlZhaUixbBFuP
8NysXNIQMva0Mv3KfXGd/jkmPnPxfWDyap9LfJfELLvMw+9yHwrORbMPuRtyulKRUsSvu432uioJ
iyuJL6WWZsmLGrXwIgKU1Ph9ONZk44JU5imLooJ+BzfRk7pycZew4LRThMcGqeB9aFsUaPDIPMxk
n4oz/QdeC5jFFk7YxVQhpGkux6W+i/NTEuOTPJ2LDUTl7u+I3lBcQzNQ3VmP1H0wWhS/PC1//pb5
Sa6vUKJQsel4L5uBvqWkxTbWr+9sW36/AgrbUZ0eqQtRi5sI+4JOQh0JRoewP1gQTBpOVprS5qmk
OoYP8UtgcHmreR9C1RffC/vjt5xwM6fy+tx1kRhKe89qf0ZV2NpqWciEgUfaEm6oIc46XCLDRYRp
wqnXA6RAZUAvTiy4ZCe0Wnh4bMBq6+jSCA9Piaiy/XZNXcrswATSaXMqeyFX9Xue9g+5V/OczqM2
katH7YWjfaSDbWc7A/heHnVplrxWeLuHyULq+yLS8A0gF5SXBBHZhlcg4r0zg5ntxSZeWNsWcoxJ
iiJ8GOPDZplUGjbCPP5NWmlDGLFqRwUSTMVR4IS/FFuuWPc23H6omcAeV7raFXIUfvhU6U+/0aWH
CRAwhMgNbukI33eK/aX0ukCYBBOz+9Quc60ft9fgSlyzTgRL9FEXhKkfDyy7PTDcmwL95wwrIebO
kl1ihj/Gafzq4DkhdkwVc3jZVTENTBsVEq8u6T5pA+lL16hTkg4dAv4k5JfDNRA4p7MQA+KGbU6b
6Zld3EsuMeza2mTUqb9IBYVl2aoYENKCLPeRoyVhUPzmkpmDLqf9yiRdZGP5SFPJ3l+FBpHuiZk2
YYHcq91QjZzDU6GuCIvlkIbBeNUKRbjHauURtvqDXb8WV14z8ZEuD0wc+xFzNESXXKf+y/E2+Bjt
688e75tUwhh8inHomttPr6VekfCoDsq9chZre815fhzvtsH0eeEvmUkogOWDZawRq2vIacjaIpQO
MWSyDcjlE1E5pYHlxqbA5tQu597kDmvDxqkJ84776AGVC5kAmvfjFT9YrBQ4EFfDMFxRnEvcw8+I
NGkH+/3DUX+4uNma8X0V+xzR+4nzu589v6k3gx2ufsaowxHuUhq5YF/7MlPHatr+ZuwOrQmzv4nk
FwaXl8yPSCO1sSol7efROqXcEmTnCCfN5+f6DH0wWh6/U9rDAiindHixiGm5oBikSLMM1EEPoekF
F2lmTpHKBMKFWOXqxO0bnoQYkeaOi5TqDlpjONsjD8wRJpOF1jb6A09v6UVi+B9DBC9AlVCVb5S6
vgzUz9WmY83hB4g5OtbaEHdthAQFk6ESB+YdwitmNbi6n+4GoczA5MMpV0oowURRsQsYhB0zEJWj
PHKiJ70wJeVPYoJBnaFTK5R9PS/pJZJTBdlnR6uFEM496npaLFEE1WV43FR4Yx3tpZm0OgvbxmXL
AsZeg0PLyU6TskgWA12lUQx4ObFXoMmaHVBDjWXqThvW8Dec79M1sJ4zqzKD088BkInvl+J3yoVc
FXuX4hVBkmC+CV27u5t/aOYBSr8dOSfQWJLdH0fPqRq5py5QdQfuZZrhDKZK4Yh2Twq0M+QSDXW8
k7CniVbq40vYFTz5trVc5qDlkgP3dJhc8PndvnMpUSLQMNXFFf884Xio6NTWt1HEEqUSz5imu8zu
CG+ikgfEQOq99Z+2ECeJLDYW4nYuJGV+9Ajjnv6s1NnpR4nf/SO5RS7tJC11SwslrszGQbMKLwto
mliGRdKc99KKMQk0TXx/jgpJaQTEFoWHKNTTRVrrUzO3h3Afq7u/xo/idCCh4xVV7Bsxj/vbHJlF
fEA/UFEy2lio41evKRXDOvBuWr7Gw0eS6MxCMh/Gqek3ZvoaI4S5+Txv89MvNmI6RuLYxTWvJXOZ
mRZlVvIt+zRcQrCdGsmSGC351prVQHza0VIbT52Af5lDTUEfJWWZDW045hrvO0dyUJy6qDB1yFrk
njbdUSjinbemIex5RnIgXyFvTUfIEaHEtckqPB9bruT/dmZVgblrSDw+CtmzsjIfvE2r/9qSqj5P
VQBfrLkN4Uyk1JiR8pVMxJjq8FSOstwRYFFHGuADRhZZjvXdDyQ0f3fbPOdG+QWZmt0yDAfnYrdy
RijWtccIbvJhHxbqFshqkmqjoprSk64vbmu8HHe5dcLJ5DZJtb2eHgR2eggy+f4NqOm/ACcXkXyV
0Lr55XcbScSMhAQ3SsUsDJ5UyLizPer8f6+it+VsX2XhAn5ZPvoCUEkD9DmxFURqUaM7CAJqYsq4
8vtOPyQwzcUKiF7sRMuPjsh7Kwc3UQ3jfJ3c+wNd17gGk6BLpZmEZt7d9cQ3UaGoXqbYRZ+4xD6e
vLf4OVtSt6bys6QIBYVV6Mbntn8X/+Dqj6HhjwHxA8vNz2hVNDdPNxSBXsChf7d+DRXDrGZPinLW
q7ntOtxmf13yDaTqUtQ9lgxA/uXeO4svLf5gDt4uIVlvoh9x9VT79M0eFr6MgF+panv7G/QTj4Lv
bVgpJfxPCe0NEw6COiJo3USHKdeLo5eYtqw1TlJPL6TTvv3zNjsQIMXHtGYGldk25HgSlqDE+Wxs
sUos1da0+aZuHJEcn9eMeUIgWaVyfQEpb7W1fNtpAG/irMqIEatObiAAYb5CRFmRDaWo6ESMWvXl
Uvn2dgAtH2/tuYkgDolI2TLBgGB3sOKrcgtXtzCSSV2AtNAVrzbYeJzRnkjW/ysqQpsdnf2Ggh2F
XY0+vfQGBHVDhRxObelcI4dgMV1GffSdQrUjjLZc/zOSXjhSRXTxanCqkDaRcyftghdfzXx7YQ7B
QsX3mnWzkptJ1QfxrEPqpZAMEniHygGjG9/Dzv+023inOfoVhtnJstA9Cb8/5jKSz60aMGYRKIPW
JWopE2xYgE28gMdRGUS7g7+BuOY/W2ca+s4AAOVYltT82yGZHNh5qruqenUdg1noTFQt2QawwjFO
nK9oT7ksPcRxrf9JafQ9dzKgJOvf9hqeQvSpUHrEG03PeSeqCQfYOpQ1JktxlxWZpS+ac5lwmWmM
eDQNYc3Pa6PQbd/0yqHB1uZf3JGXERE77+OQTDm0+W9yNTkjIFTIaGlYEJCeWiDmnUcxMvOddqga
1p8WPpOsA/y/+sQSjySvFifpkC6qxxkdt77BkwGvFEtUhwWh8yi3goiU2FMsvL7MKOQ+A1omg0qo
pQIp+cD9dL1k+R2H4u9iVNoxDi8M6EVDrRhkqa+wJHCz3jKp7LfC9cVNLMolV9CVLqrUHIfwllYN
l2v+imTUk3RLv1n5YtuJs1yXAq362Nxw0RC+cjSc7PgU8OQIMfZp0DFqA4Xi33/U4TpLI95jGStl
SlKhcTItOnxQuUZ5AkvtRbl68GTkNYbOewO/Qi3V0CfGiK7TRXg7Bf22656Bx4G/tycZyU+kX6sh
bC80NAlA05cKESmt1nfBh7ICzPJ9igTvO33gyEABjLG2wqn14izxiQ0dKxnALPk7rKYTefElSoMN
Q8QlehBPWpLs42NQAkD3k39Xf1LLHRDsfET/5XL4GFVrWMqOYar/AYFlBbST2d9CSiP1fN727gpT
45hgSZEns/VjzntUutKpYQ/5IJLcYDORujyMFXbZYcs8ApKmEEkOigpCsvKEwD3foSadp00RrvC4
egy4I83GOPncb2XGjxCZEB13fTfQr2aegO1n6GXKJEBOkPUJdD6Q+00/GvcowWPaUOHL00Uy3aB0
/1MUcW2AiUQEXJH6r73C2fVVZTK/ffkaJEZ3caqEG4CwdvCCQpdXxehZVDfegymlpuHXyBse8i6P
BEpm5lxyuXngA7sgnwzp6dGMnPSOXQ3yfN6/LpArVRS6NwLV4lQc63VjyylwdCdvGf5vp9iJ02Mo
3ux/stJUNBNlvnCn+bYv7HznxUZPGRi/fxIwP3HWZLOXWY4UYZYFemMYYtUb1t9CevSEtDAblUjp
ulxund63JMP4Bbn9bdOop3YD/UhE9XkXOjBu9AP8RlpjMfZd2dmo5IZ2WEyl9aY5O+Fx59PjA8tD
/q41bPupJUstfmvOAYzzARCsAT3RK0mjVo05MPXBCzEIE8y0qlBm0TAlNUwM6/TUHW2s5hre2z+g
45MWiHoO7oODK6IADckE/u0Vu7Mgawy0QA/9tmkDLndoR8XwXQaTteyoofWdXV7NU68eIjcx1SCv
VwxBVdf/H4mSY9+Ki0los550meDcV/hIL8uZ5lUw5CVscEf169ILYr5WAUEkX52bg46YPOzu+Xyz
IuZRikCAjfGyMbpF/+fNNsTaU7eNYq8LK4V/46Ig44iunbbx0v6N0XtJcU0dCGpqogMah2fQvlhR
F4w4py8iNDicJYq0inTlXVkrXow6aYwHvLCVYOx2Mnjl971GSyR1fi69AW7D19RSczsoFW/da5mK
vWU/aXxyyBPJAFY4dNyb6f6Yqhndqj9U1AxGG/oQ6oo1O0qkdQlUQkT0Zhexo0OaZLjWleRmlzG7
mZigB1hekb8cr70rTxen/U50wttfWnUZm+LIKaYT8P2W+FWjASjPmOj54bLHRfQoFfrD/khKUnkP
MqjCDntnL8Jc3ZQzETN89Mm3HtpygN6zq8x6gThE/bbNpK/N19FMvJp/5/BfMGecPysQVpZAgT0i
uwjpNr4IeavR3Vrd52XnQ7YIr7TtvkKjasRgkd3W9HdQ9gWn4CC/qyaEhTTGIXQwAzvmxY+amRjb
/8iBe5vJnLVZ0KipCRywlEfslQk9k/cOykJDBhd8/ERNPj0YG0Iv+fnogm0NyjFuMBEUZl/jp0eI
+4X2cc97XLHYH/pwQsTj5Rg8J8eudeQkyGsJ/JERmPqNnJefd5ioQTQox0fkB18w6Bpb2wvWNs4+
vvcyXHQvCvD6apaTwwwCa5UobjEDA+tbgfsVkHlsWnt7/iMs8kXwGyvvYKuLSbii9ZOuMUHtYiT7
gvG29zMY1KysEDjGU32hijKQTivT4Cn+iTDtzD3U7+XG4iEXmOKk6zLIPagm9hNR12hriIQNHl26
rlCq8eSUAe4MwfoG2pn0v+mWPdHduG8CbUo2sfJPdWnMD6YsBH8GiSkQhoGQtdGqIfUS653d0E+i
ARyX/tLpVkdprQf84DmU0dqN3tcUxNJocoBu+RasYFj2s9rxhxUi60r5Iy1SlLFg3Afgf7+nPtNn
as7PJWU/j4pW+xNicVsDCU/EEaJJDKqIQtvckKjHN7m5wT8pXhum+1A6t7Q6m3qDrk1EEjhVK8fL
wc8ILWooqfIZhxbPfwkXOHWVGJTbd3q/rU6oDFp1nYZwoIB6xluwn1QpKwIhUeV9tgq637yjMS8s
XrXm3xvielQl85al7oJF/iE9fWqnDTM6hm2ZqHIgCMgyTCBAUAR8rnWxr86gngDzrsgGGq76pWqV
Resx6iPjXdEFEXzW2FLbqJGaZ1chzxADNIUcqX+Td8piNLbSWatofEOlJbdDiml+3WwBjYRErwLs
rV0cO7HO+vBsBPO+zyEybeaF8qwwbHHNZkSUL6zM5SNeMZ9dF+wcM40JpLxKAIZDnsHe3Cz4TKvl
FofB1X391sYvSPL7iVeh3tZZRqLFiYWwV/enhfzur0u97Y/O/lbT7QRriAfo+7nMe/nmngNpsxYO
q8VhVERzaGzXNWMf/pPsJn5/thA0VYqE1ygoxOIpGPUJgjhAp+DiyYuhNX4HHlCtvYM3iuWhb5dq
Yr5EBAwNBXLDdt5ABhyTIPIkKtmqvaYRqeRZfFNFLuwZAbtIemPfCthx+QqD4NC6LgpMG5kOf5SA
zFfA1BA62h2zoFaeL/ukk4nOCrmF47zbBqKkCMZcPFofJ0RSQrSMv2TfQw9tw+8xrKMCw/xbtsP8
E54O7SIcFJM03u3NwnlUlcU3JeCZh1HsOUTPMQ+VxSP1ubpKSaq4xVbrf+Q+fEmimUjMT0PH6eil
05AQi2yOhTKdDD7HjrqX5znVHIRm2wT2ITucdVcWAWxczeAtnUH7wdK+tobStuuE+L50tmFfzvhk
H5Vw/TTtVKkUwuWuim29B4KDcsX0nnTwd6rdK7JSMwOpf/jYtIKdbb1+Nzp8KWJ8ZbPdgOzy5U40
Nrd6nr6mSkd13EIzErgMLttNuuh2T0eUvMBs84mKmfVh/SLypx9KHHnbXB18GpI6wvt8ck++Ln3f
KsOT8A7zoP7fOQEp25kSjBo8QcDi1VLq9S4VOmX/4IU3um+VsIUFTA3/FgMFb+UB+boL6iX/JYcl
50QeoTJ9wTEVO0y/jN5BKP42BsWb9i9ScDpd3m6qhyyq0Mf/FeVqMBMyKdM+yIvCPpEqDqpEAGbJ
TopvW6VSZZ350T6ttZsiuFifKbqfFcAMqirGF1TVME+hB/LwffsXNrryhFQt/sK/9EQN5oEPtRf5
MLJu3wEe4f8UV0DIrIECY82xAgQ7GU8gPcQlNaVwWI36+t2XwLwTu+E5a7Mk3iVK4X7V+W7n2cCJ
Zu521jET/HFhK3gvkW9cL83kC2maLFh95lgNBvk8liJ99WrB2lbWnBkoeYfPEkeVayhhcUQCE8vr
fSHqSnm2/D49Hwvr51312smrJ95D0zi99TUduiibWAa/FW99A2vE8t9ASZMfIbEGTtbo68moslVH
vhqLa1/1f5LACfWOXG62245M/scsxwxMbBXF8CwHda10F4Ly7i8rro67E1x6o+J/GoudQruUtlgu
oGRcgn2EfwYFrieQhvenbIxfZJsO/R1tiX4sfMPxLbrZqp0Zu1FT4ezAJAZmaJ2jJJCLN3ovjbb6
0oYNCeDYfVmVSnFMMO1OSty9j1qHqDeAE4RTxjtx5qipS/Wo0woDkvOy01Mp70i+QyhPEaknFrfG
skPzUX5uPn7SFm40SvWoj1RDuqj+BiHx0hqP/GjcHM2gjAziaZLSJkUuMY6bsj0fkGInHwlFCrYo
9dkilRDTHSpJlrfUSbPGKbBe6NMKCjZykzKOsNVYAz3mXq3brjwUtHlFgwOPziQw9EcHtvBshld1
f8wuVB+2IZ8ZpQPMAAmK8xVmyFp4yC4WkA5ccM3L84dMzDhDBzFknDPkRLfxUj/6mVRC0PCRkp1N
X3FrO1z0G/qrwpiE3Q+QiZq4JIsoNBRtY4FN11/CVoPsgGN6DYux32bt6hYiue/j9xAKwlDK3Ycx
NWpsWVzpSNbfVOAbmU0nnoJe64yyWPXNCI+8MWQ531pL1bX9nGUSWvK/N75ALrsx0aybfdHlciAn
Mj0FIKlkWIY9VJPrVpDFTMEkenhCVGsIUgXxwEYViGvYOmGWZJUpWKZjE+KESCQAat3dWy39wORR
1F/db8YHRZEdP3yrgHxgXyZZANdNvgrAUMatFEHSd/4hpMTzjCdFfLEr9mAzLWWA2XWVk9CT0q5k
syfwqO6l3ljN0xvlnstEdQA+3QqR2e13HBJTQYihMHUk7zVD1kvn+9k+g3q8WCTBHaeqF42AV7lt
R/hOd4afCLCQRDTfHSvDPn7+5yhRT9GGQOpY1ddKiZ+mg3Tl1se6tXd8XU/MuzWPDkHwPdN7Fc1s
tYJKSBMoXAkKgsDqB+jyzlE/b+rCborqgSr1n4t4AWLcrksS9Z+idXyX8vWJkQn0fHbXw51ytRii
KUjr0DyshX9iBsXuwh3iwxCA/ufcwmf5pMxqCiH+yFelB1/SrGq9nRwyFbUvMuRy9FDpRuFV2CZ0
LR0z17xSpu3vQjwAw/7TSuVlZj9J2VsIFLcElf0KgA2OQLE/IMbj/+w9pUAJx+KEj7ga+KcZgNXl
6HGpXJ7dfz2u+/D1lD+Y07D3UvU2V6J8eNrVHfohD7vhb6oELIAJ7i3BwsfTidPmNDwqbT+H3KoB
3ZswaImbrWdhx2hA7EchJo8vv5umm33Lt9RFkeswc1p8sdmHqtwnAas726BeJj8yVP16+ykDngYz
h1QO4868OlX0IfOs+BX3X1Glw06TwdeozpyHEY9k5/A0zBwbf0beVIAkcUxzkjHf8aRb92fXaYrS
P79IY8zPMzzQRyIxkLVrxiisIW/AYM5CmhXRiogt/g9vT6wnMnqZo0qZn0l2lOr1Mzf0AJNj6v4U
ZaDgvI8lAGUqjV60fmUtpB2GZI5qy5uON11sjOKD/Uv5QAPpqGe1wthpWgYhvlHRIb3hNECagwAq
yIsYfa4WUYFWJd+eQWUhpk8de/F1Vi3H2HVxtss6KR+57cScvSNyRGtsH4TBAf5tjDpze7/6Tdu5
cdHgsp3gwIhq7jvnUwHxtOLkUnRSKZitVvPLGuC6tLfFm8/uWtx1cU+g6zBzhcMzMgS6XKmMu8g3
dlXMsZ4AenwqKhI/9UZFXt1YQEdMKcOVEzdTgDCJn1CJabV5OMm2PIl/vh20HQz6POq9v703CNqk
mZvaNkjIMqzUcZa3Ge169+7VZFbaKqlx8I4mNqohshOHS4y6W2U0yXAVV2oc/gkSW81EdgBrZVh8
3Sctbh23I6I0bGxel7KPr8GZORpk0cXPPZdLmxBZ6NcAEKScrC66PINtDClipfkzyxx07G/ccw39
wZYIiZQg7H0cPm+gA6F9I3IhVPL7r6dYDqM+2vUQfZhUCwIm87hhyS6Aq8BWV9Cx76GxahAGjEl8
OdtQrOTKx+s9g5+v1Ys/jTlcGOS1GpeLhJxBniQZWK+tJnvOkRUmrqIG3F86ekbq2EbG5L6+u06v
SGwvvVx9/i0Y2OophKD9CD3WmwAuudumOr4sMJr8FcEj0frBluFbYKt4kM9Fpc1uyZT+aggzZJLc
tFZ5HBuyr21H4O0ZEjweAn26807CkJ0+Cu42i6hWf9OrdyWxrwW/9fYp0xMQ/SEGwoWVn6TKfSk7
udNvJzUZp0VqC+AbO18kVvaInFvGYxkbmvtAAJOvTvhZCb6tqXfe/McxrqJHO+G63dJ5BzPn1b+F
b9nx1WN+XU9d3V4S0H7A9ABjVbEbvOacfSIp4k3iahdBcPFDoFUHQcnB9FVZD63bWL1cOVkMM5Vk
Z0mdKQ08fTk+zEvPL0//JNeK0z+dg901ns+gMjdkPgRq51YSC88ExPzu7xaGMTKZ1hUHvZzUYiJY
lFz3lBIeIQzRda3hikz8IJ6x5ktV0sLONaBFBItMnymdhCawBSViRqqShzFnVAZluMaAwJMC3sXr
lmNhhLRXDtdtHz2q5Vy43zFtpEYs2wjMcnROEr9t7F+NBJoGfV5edymRU3tGxNldL+7Ejr479Sek
6FQ5QRJDMbabcwqVWXCwvFmwUgIuPSJ8owI8Ur78+ix0vjzZHWWs8lYnIVfuiimgejDCS8Wb47Dy
eof3ygNz6yD84aRvYKkJILNA3d2hQb0P5Reh0TD0RSxKBDFbtITYbzhVMUYCl4gOgBTcyXENY6ai
ZjotGabixdekLTV+6eiTkb2cJjXTuTUX6dhz07VLKvvnJnDIUvJj9WBoCTjozSeCzNYXE0QdiUHR
AfIHsrbQnegz4CBQpfqfiY2Ldwlv3IkicKeHtyQBORC/Zjz2sRZASXTGRUnTrNgBEwQsgXeUsyZB
e47yL4misiF/5YF1lGU+/p+8u4gLDqNF0YCTR9xtXpnliWuvCsLR5otW8BsAJ+kipCzRzox1Aysn
yZK9yvQTqv1nQ1GzlWO1ZYh0ZAkyfOzHT8Y6B2Ct9MnnUA+8E1lHIALAYe8M7jva6yBm7SM1pzZk
x0Yxa/gZFPW+RDuHYP6ek5lqWUKg95jPAiDlGyQ1ArV+YVma3LvmJNZqsbLZe4IF7PFb9JU+dSF3
NHXz/xTJfjYsykNXeGnHADiVZY8AtdWKzgbvdZ/zHAmGF6SBuSe4Zo/XvE9FfLAA7HfOco0dAQej
2y3e4KjeGBiBdprZmy2FAsp/9ct7oY32KSi7KDG6Cksv1fw9jhJz6TYmThS31+vzdy+r0ifz024t
Nmk/QtD32RHKqgj6L5eRNcqJ7Je5Iqva9GOQ2Y3Wk2PX8mT9FRd9iF9+a6F9s+E/3tN89GEQxj1d
FRXkunj3iCocWKhlY7yE9Zr6nnd7lIfLfrn6qJBCU/GKWqFaN9JC045x2KViegWat6XKi2x7hjb4
ehzqggf02LXy1C+odty7My0/O8HYEz047T40xKB7h8mcwdCNmst8mW+26fl0Bzy7bWqlZfq62f1d
ebWLmZP0SiFHsZ/AyVJZG0GTqZIKDNpX1Y8L2ME0tCA10U84a8tegyipyn5fXJih24h9l8B8z+uh
WvPoXB54UOduMz3x5coSP00IwMFAqyPa/8KxVBjiNeylimBCcRvlngsx1OubqN4svUjv8rgZP/28
J4SXrzI07NPjfkigY1nmsJHUUBrwWNEHk6EIu4bW9+SJ/+JOC87heeXVlXoreuR05WO3Mux6UAU8
4x+YiKXGObi4fG3x8ILlAanitkDMdlq+ZwSVIqw658BdMt7dDzdzJBcAqAONm9Ex0rsmNadVO4+P
WLLSBZKpQQZK3mKrUH8kqJgH2xQRzwr3L9t9FCbkOypDP1T15ABu5PkwDCJA+Qa/HSoldntupJWM
Hmioa71c8QpB3DBdcCn4B3B9LvwcYcav5mYDLsqB3ZATZn3MfSxxPWwbjs2eltHsx2JLDkgnrdEG
s84l+K/XwjnDcGeajSzZLJmz4JmwWAs3LK+Na1N3J+U/MT1ttTMd/ETT/q9+Nx9c6hyAsB2P2VDW
HbiVLNiEMhYUfivDfbyDq2CuilJanY1ntaa4Aa2BeK3yVEzEz2yE4yi/L+6So8+Axw0s7Fi2pR/0
HPZ0pN8cmuoDYu/xTjDlXrM/MfC9AQnmPguico1akHAhtLXBevuoHdrTVR3rtjGKqnie6TxwhJzw
td7nRKu552jU7yG5Z2EQliMyc1QKrygrbKbMK5rhMx9z05fgP20o5Xr/gfXtF8ry/SzSKw84W9q+
itgOpR1ljYwCTqAA8ti3ugZk3d7C+JLw8orN/7rwXb6Ej+1gRbsOPxKugLrgQfYr1gFA3YWpJLnH
Hc5KIor+eXrw4qvOX7YoBSoBZSbNn5lN1YqJT0I1lThkAixrQdehYMe1KX2MHS9igSIu8BvxZdR8
aQhQeUODwUQ0CTJ081gQZZpEeCB64ZeQS2ZHuz3z27Tl71eYRcxmEuiXTjuGUbCX8vhS2Oo5ny4B
d7PjkBpB5OeZWDk03iCLqgko83Mg5XpByMsSdabiT6tjW8KNbMyrUnMzPktHGrkbzre0HOWbZ+wP
6LGpuhihY7AtbTC2/xj3SGlXzXxKCtz2yc3J59wSWX/mqs37KMuwB+sdsNW114jXrKl4JJb8smPX
s1+zibJxGdgbk3VH5pWVcvYLMvTOhk0Ps3kS/3aX8DATct5XlkA/jOb9NGuaLdtMvHbh2oh+O9zW
9UB2u+msrNFuhEoJoK4ZRL5QhJi7fspfxMFtlZXjWMzIAx/UsuniYVChZRTL1h957iqUrZzxaMlz
FIhClB3GqzcD9QexXJKVShv9VKYnElqpoz/LuFVdVF2zFSSE4NYtyG6p8Ri7yEMpYmHAqUUzQCbH
j1YrTlQ2AE/Z9StQEjJGjHlMx2Cc5kjw27zebIjzpu/lrlQO09nDFt5XqBYAGYQrJMLkiyu+2f0P
xSEp/yRY2ykkaRuiqc8BV2L1v8Y42HWPlvu590GBuAko/KhUdpXPt//vv0zgdBrWOypbjdtRArzD
Gt9rRcPS0czJjZl76plSY7HpQB3SzlxEM686Sdk7Rqxsv+mxCtmLaFRoB5q7ky8ixlOXNamrvTi0
DmVEu9WHaq6r6I8BpNx3jPz3bU5+PJQY9JdzkqtoYVguZP6o+YVRDyspG5uI+fllpp67D6CMHkHg
QVwQjr7KLnnN6+So4r41UkdiEkLRH2bztma0kdk7Y4rqe+uWS10djynoD8I7/pQVprybhFIFJqr1
le5RwnPSdhRrCUfWasyVjL/zjhWPHiYoj2QhcBVFwXN6yFGahUeGd/srbC1fRauSVtf+oLRCSrdj
ncGmi8cEFJo37tqjqQGFA/5shjYmynILn1ikCGUNsHYevlejw4BCHnF5ZzcwiFnluVCb+oiKGflW
arVALiqF3T7xgBTZTe1oHKt+DV5DxlB6hfwt7WvDR8AVuK6sZPf42EfyXWL2tQfsVkdmOJ/hT/FI
j2ktU3MbJU7vsCpjsmKNa0Wlt/oAfQRSLCh54Abu7zJJt/yxOUlauUPcO/qZUEvUolgWY3VbvZXy
4AlnJWaerq6RrxPWTnjI/YkWcFQ0akJam/3nDWbs3vW5QlHwGZbGk1DFL12nh6+FjVW/w5dxiNqp
bbvrjQFiuEdAkQ2zowLeh8XaHkmUUzHcLvWu9ExtZIPXStEBIBk0sS3kdpDME1uOEjwN8pfWuT7t
s6qNyFHGU8GlCpr7bx9UhATYVloecQSs1KFiwmqGLnvB2WewWwyEhTlFAR8pKNgswX5cufM3zp8Z
oNljXhT7hKBS68J+AvLbisC9tLkha8wrf35JLEhnYlvZ+YXe2nXbO1K+I4v/xPuFFnPZ50aT29sM
3Rq15Lc3WPtulfhg0PyS57kz24ZEwknOy1VvUOs6NFZYxf4LjEv8EQUQ+Hnuh1V5+OkZ8A/nGZf2
/SRlIXFwqTVXUNl54MXYN6tIuy/ZjwOtKZopBTJeauLk7hIRuU7wAOIIneoOje73MSNBVYPVoD7T
P/YW1p6PH3WadV+8qH9+jPqalIJN3VYudFGJLhval29i0OY+R39klKrVx7ypV6uRfFSREe9EN+mL
E0UQwtXbA+HIEbtjA9hcNVk4sicu3FuZt2KV5UblOJKecgN2oTf+W91wPtJZplTzCMfHVdhT+0Rw
fsw7f7PPOoI9sGXagLz4Vjjfeeo3txwe19u4zOimIsnL59vyrhT4vRUcPSJsq6vE2TSAws9WjYtR
elVLo68j/WwMHsCIPAAkL0/BeyaPOrHQqQt7+Klule+ZT9GGVCVFk0uTKdqmeLC1+gB/0msSCkup
8EOzrCDrO5egBt5TDVDj3C3n9+bxgvSP2o1FiRFBBP1SonSxIa+vBzVaGg+5wwiXHXsyjYWGoY3f
4OYDgL+TeMDT738eEPK666Ih3edJ7Vn3HotQZGMCJyJHP/reGaQT7ejAZQF+QiiEkYgiXM9wIufw
ICe8CHYOmAFkLunOn5ywMQtGOxinFjN6wI8yLcFRGzb2HXu2qyslCqnSatGX+qCfISb2YSfhXXGA
rlsPGOhnwgqsIdqQLFb2BfBHGgDQKwka/u9YH5pSBAmbbUCjSWaZ34xKdKzJC6w3Km7NpYOw/Ads
qvToaT/rBzTUpklUohqic+8XC4kWxq1kqq0zE5Q9KK8Wb/dcQPDN7YDvSVPbka8rmt/rtaIBQoCr
TzcolMUdts1fWNCuRYSahNiFSKaKVPKzxb7E61bM17+smV6l01cFWehKM53iiu1nNFHxTAeJ1vnj
pzfpzYmuLH+2NktaHuUlD3Tidw19wApLEBU2m+7zK7HOA6JomIp1nDaBpQkiwbCGFuiXCxOLD0IX
oqdbfVFFQTCOf+Qk8AqZZK0zzWWd9GtBDuPM5E7fKQNUDBNap0/hN5qgztxQS2L86qMXqo+B5bMw
s8jb1Lk2mpT+/mBK2kvoWU4K7VyhVYSCCn21/nPV2LOJNs0n1A05URrwkBofjW+jSefdS0w2WPgt
pHU+o3TRQji1iyqUbWlqJQ/I14zImidBkyh90U3EuKW3z3i9Tt0+uB6LIxAcNp1RhZPQulRlUM7x
Gvf3tt2HUEN+ZfSGnPwVq+swuBF1sLQm6kVWZXU2WngueeYElRyn7RX5btt4Qh2T9W61A44DRB2J
cgPSElvcyRrzaX9UVkxWKseJ2Zoq6NQDw7adsDEihILSIRZ5zIfuJ26g9BIruqemiSzSJbl8wp04
9JgjUcTsufx5oCbg3t4RMy8xA8dRdZrrPMj8e20Crcmk0CETR+p1JVDaDg5eym7q1bdY8GPWUyd3
qcIzkNcrBkDI8WgzyCimMqjmMjjsZeHTMozCTY4a2euCtu+6c3dpwb2pEbnMq3qVK0mnpaOPVRzl
lBY559y7vXzub9F9NVhVq29x9olkmyJ24PVrEzrs1oFTZgSfMtkZTA5Esd3F2QUsPsLftS977cqD
RGZjZtskANtH0BvN47FNJqOADAIP6pId/pSaiueVqqOkzosvxerae9xSTaZpoaKwMWeuur1A0BWX
xHi9Zgz8pnaZNNrIsYDqVE4VjtSeKc1GD7wRNfYkPgCKJSAwHHvfABih3yCK0xJiSuIpa9cBuE4V
7GMBOvX8iFmBHEc/18iSozeq2+6cpPXYSqOyreVblSgrgPZ6bt4/tBjLJ/Ie19ICmAURYNCuI5nl
w6Jiu8ti+IS3ebluTzxpjP4CCNYGBUtoRkeXxyD1Uz3vgBPpkkmes91s850ks3c5KZXBCdqExB32
+CMVZTayv82yYaTqXpKJgzDyk/ypZpkUEsqgKypjS1gGTVaAOx2nfj/X2dD7GBcjDMKHSI3Dqlqu
bgXiTxAz34tlFjX1ji6RS99dI99KLudHjlX8lBt5ho+nqzlHfXfJBnVTGT/IiGu+962gl2U/D6YV
ieUpCF4Q3XB130QZEf6cEPw51ju5XT0GZ4EtRer0ooZxLWlMe9GcIMNPwDcvHlyYFs4xUTJgR4gZ
d34J1J5rSEle1OH/sm65wLzGB/PbKEQItPLi17WB7l5vjnciRriBGhoK3HN0RJBdU6jBEaX4ZV+Q
livUgCWUJP7UFfmCNUCp7oiB5NRP63gqQok6cHg/zEgKBXAO6bIl1+Qhn+mJiiCGAwlCQwO8Maes
nisuVvbb5RgV0EgXBNpeK76DKuNNbdnhyYU7nnQNeCA3feiD/CiXmNgjZU571WdzB8XNEAkelO7Y
z6Jl3bxkQxRp1ktEDcq5ni0bHbwcwelTOYx86YKXW13SUTI/tkUJnRU2ZZm++DFTepm+4lnizv1g
/E8nEsTRmp9SysWGllqMofsdP8i2PdEBG3qvsIMrsvIXRd04wmD4NB4r1UA4CV02mu2AQKli9XSt
yIHc1dDPhQLfU6ClqcTPn8y34h4nxit/RQR0vzzzqSmDxQXvB4iY00+cbLrFHK8M6TTcwmH3rQET
MG3HSCPnBXRIfGQIe0F6EWJU7Pr2Y6f/xs3BFj7WcmNHAeXh2QwRMSZ2bIqCFfrpR/YZcb2Nb0Ib
wgx8/jQc3OXy1MoyRtUc/NSd/6XxiO5qOY9djwNThz1PjOYSj9DZz63Vulzo6yMhp8/itnD69IdY
x0DbxOfqgfbKNgvQM8+F0Cz5wZcPuGAQLuycRdtR1A8df6XfcwqYqTiigSMBjlgtoo4ExKtRso97
b4ELZZNknqSpwTYY58dt6bbSaAYU12Tu5SP/bRvU4YKmX7V0K3VeqQnMcAWnIYbzV4yCK4LZhJ2Z
iH7BpyiMFF/zEOhHrMTckjMyyzA4COhEs/Ei9A4vJ+X51V9JRqk1GphHhjcUtNK/p6teHdzIQ/Fc
fIXw+Elj9C+KP0S+7ZDTLb7pu9QdhTFpYfIuqVIpr/W031VuzXD6DodiIwakVOvf9Uopk9X+7BLK
4efbGHLxX2gxULBljRZiSJWZ3hcB
`protect end_protected
