��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g�҃�f	��m�T���ƌ��"�C#~������VMb#�X�f�����|b���e���rQs��~����2����؋��&���K��٣�M�*�h��9�1��̻����d5!`�S�o����@Η�I�]���<N�����%F����0�8k<��~$��~!~��dV�Tm���s�@����Zl�U|{G�-?ҡ�(�K�ll9:߷dW��'!��ܗ��W��w�#W�q��ܬ���ݓ��Qy(%8jZ��{5�k.X*g���zۿ�@��S�k�!��������e;�����l9�&�V�����(�0mɍX$�II/�؂�A�gS��*n�N9���RB��#fn�n�����R�Q�V�y��Lh�����G�����TE*��k"���d)���lH�%Ѱ��b��5��3�~ۙ��>���l�y`��N�PG�[X|<;��F�/���ɠ�0�"O.١'FH�#y�$��
��wv�8��+���C �%dفp{�]�Q�f��ו��p"�+���VN���� ��7��������%+c��8����QJa&E2����|�����7H8Ǝ�J��'b\���",`�����b������"}�­���x�0��D������I�O�	��?���e�.��ୣܧФ,N�~��3*�+Qn��k��ĺ������>��'�(&���iӛ�Q4�����-���ؖ���_p G�d�@���a�7&�a�T�a��V'�E	�7�!@F�i�r�o4���^���B�q��*�#ߵ��Rp3�|��L���2Sìx�k4�L�Q���~oQ+�{W�ð'?��պ�JiiW@C�UD�S|�]�7W�,S�u`�t�1�+��ݤ������"�1|+Y�e�"8�����H�z'�����>M>�ŗF�="�>]�Ed}O����{��|Dd|0W�]y��mV��vcE�~̫J�%t�~bJ>�^$/1wV|N�mk�w�'�[���N���2:k�{����T�ڱ#�=T�h&l�\�L�1A[�٩&�����9���=cr�(6�8I��꽖���iϗ��ҝ9�z�q6�������s/sGo�Ja�j�O?��4�ǐh��9���F�g⪸վ|5�˃6�r�;��x2��A.F�d��Zk�)��;$�j��r�%�i�мCp�u�]:��P|q��`?�E8r��8.�,3@��ϓ{G�#��+����E=.��q�却nS#��H�LU�B��i�9+�PNCΞ�V�E�Ֆ:��s%��Z�&�'�$8�����ӡt�/�-N.��dY;C��ZE2?�T��oú�^o��
�}�q7�vVd{6P��~��4p��!	t=P�=�7�z�9^k�+K����XW��Ë�9�����PqR��}t5јǳ/Qw�(���!�u�X��
˒�ػ��u������j�<T�Y����9����c�Z-��������vϠ֠,u��r�/�	��K�sL�z��,����3%܇?A�n?���?�)7�jtUȈ��'��0C`��'5p�͡=�5�
bK�H2��ɷt�³��p?��\C�j@����Z�郒.�[X{������}��L�q����K���	�q�:��8��WC�\%�|y��0� ��ч~3ܜ��C\&?�I*�)yIs4d7m~X�Ts�NN��Vַ�P�4���*o����iD�4"�����r�݌�h�C�'w�����I�w��6:�������4eG�
$�]T�C�ο�,��YRE%��Y�]�������:(��}d�W3ն��f8�-N��	4rc�@��gq�f��Hln�Fs��Sm����a�+}�f��~�fƽ�p4�dM׀l:����?\/�H�m��QC����h�ї�̻�9"��ڒ&�Ǎ���%�M�9���f�]k��X.�×�3OO��i6~����L&�J��#�}`mw��z3��l�g�"cZ+�+�9|�0�tn̵�+_��C-d�M�А�*�?�E�X�� �a����L߉l��m��&��gJ�R5M�b���Q�/�Y8T+&����K�pb��h��$��z�كe�����E��nk�#���L�NB�ײ����#	Ni�p]��st)�K�y��������L�F�������(�Cj�H+F��< "l���n��`����ֻ9om��]:֓�ԗ�@X㹮���Vd�%Hq��]�_��q:"��Y�OH�(�s8H� �A.�Hs��,X\�D˓@��Y�"���e,;���#�4��&���C�Q�1'�/{�r�L̻��?x��;q�1�_�����j�H�߲@>��#cޜ!�F~a����D��-+u�,�7�L��Q!A�#��l�>����Mw��nj���&oƱ�wK�I	H�JH$�BDޮD��1�E]��%���%I'�pM�qL��7�&�-�t8���w�ڏkY����o~,��#-R��G�W7j˖!�8�>;h+�a�}�v2�B{�ޜ���㚪ۖx���2�X Cc��p����qҮ����;�3�gk�G �$q�D�n2@��x�7��%��3RƁ�>���]|�T�#�LS;����Q�%]�Q�M�ds�{!�F����2i7=��@s?��ԁ�e��`����QW~=�k����?�0;�eR��۶3) �lj��tB��k�=��S't��<
�R�7	�W���.��� <^���z!3�1G���Tu	b���.�@ɦ|����b��vz���|��4O��J2�M���\����W��w�{�]���1�] (Y9 ���-�u7[aq O����#HFqƃm%�Ž1$���T	����~�j�.���@%<�c;���A8����k�K��J3�|���dR��34	}s�	�4�݆���]|�'�}��F���\R�+
ߣnisM+�ոiذU_�T^��堙߿L(=r�܃\���j����|7P�>R屭u%qX��?4ή��r%	iF]��O�z�BJ���Ǉ\�/�.�ސ�Y� ��W���{�D����#��:��ܔ~�3C��`��1���Q-�{���P�͐�ꃹ|j��WZ!�y`�<�G1��8~�9g�OG�� /I�-��m�k�Jơ}���|�fb�#t�c6ũ�-Q�-�n��7��} ��'�ԕ�0(CY��H�_��	��T��~^Of:� 3�6�F/�2B,*q��P�!�TmA��W;�H\$d�b۩���}�pw2d;�8�B��.�f`I%FZ�a�Z�f�~3	��A��٪ttI�����_�nF$��N�]�v��?�gb �I<��ze��������ri�u�=���A�7ҍ�����)�7@�Ն�t Ö�i'7�ш��snp�Avfw�h�]7�m@��W�C�8�(S�}KC�����~Ȉ����2���e���k�M�ۚ�&O$�?j���wTwc?�tܗ�y��t�ɵ|,���P��X��`ݒ��&�ח L'%��T��N�nX��z?�|I��#9�U�<��_ks�W�	GI"FĶLe�`�%X��2�s�L<��Y���x��(Tz��-D�m�}
Ӽe�7'Sg����V#���#a^�����nT�4��}ha�\�V3����r���j���3�JOA]�&��;`N����f(6+�R�TN2�����g�u�٨��O �u�~i��#��O�V̈��3�"��}��|F�S	�.:N���z���'�E�y�M%��+hH&#謅��#|�w��%Κs� �:�E����3BO_~b^��^�$:�U�u-:}�>rU���O#M�����}��Uv���%��ш������n�K��H���:#�y�܉Q0��/dK���'Vt�3�1��E�ǡ�{�,�<0�9���6.S<��^�B'�rq4��I4@�sǴ�_�D�ǷYu�`S]��mngd�"�fݥ }��,���Ba�@��	���1�?���}�vĪ_f�vf�H6=�A�Rkca���=�H���O�ƫ��3�v��@H�Q��roa�g<�>�ٱ�`[�2���PGO!Jm`��w�_�X�8<���a�$���J;��р���|_�]�����هQZ�r��!z����h�LIl�/�z�Z,ܒ���yU�P�Z� j�Y�Ţ�SX��Y�P�[|D�0��Gm^Ş�F�.��$ē!i�#؎8/�����'0)��ϖ�7A�-:瘢��˗�|U_�,?F��y�P����j.2��ܾ���~!n��TC��8�&�������"]4�û�0��2q�I$ߣi�Pvm,ι<m/�;i�pt��%�!�&n�=��fƚ��C��T�"��^h�����'R�?���k%~4\�T _i_���1�pI� R,�5:`�@���a��vk1��6u��\�Qݭ �Z���,
�i
�Ĉ��|�z�0C��ۧŶ��t��6\쩂��,�|�WV,u�����	I{A�A�ER�I���[|;�����7���'T�M~��+ռI?����.p�y~gG#���'*�q�8��Hi�!�Z3t��b 
f�	�z<�n��Bk�j��u����L�Ka�Y�\㫞,��Bj^@y��ٺne���%��q�>���>y}2�l�m�u��������pY|bU��%}_����/�Zwn��r�3D"��*�s���,ִ��0��4���W�p\Q�K.�K�~�O�_�����s�R,Y�@wpv&e0vH����F����d������y�~�~�\��oߪ����R�t?��,�������]�A� �{ �X����˒o����b*)�����,�אP��j��e�� ��7�A8*����r����(��)��0~��~K���T�E�z��o+n�4d���<�>N�}$�6���%Oc��S��7�f\)`�n&e�B��B/Bt�em���;�hf���fԹ=_�Ճ1�2�c0�]�%�8\�}e|2�)��/�5GJ
Y�9�m���Õ�hE]�K ������ܯ�X}��K���,��:��ϝ��$[�[:Z�L{GAc���h؄���S��[���7����S⹡E�4�Y�s����\��R�����>vf�*�����0n�շ4ԮI6�5=�(#:�0���%;-�{��p�(����GT�����
OA�ɀS�8�!���{�a����&��͏ݎ�����@�C�`,�)�{�H���t��`�X"B���H�[ªPj*�!�-��A%�p�����/�4�-0m�c��;���:��+3�=u�tD�ۚ-Pц�BL����+�LR�<܅n���I�LWT`�e@<�wβ�Mf��{$2�m�n��9��W���3�ĳ��a��)��9>�K)��B8oA&�c%��:�l�d;PV�����;�p��S��pц�1�5ƨ�{�I�ש��G�-A��a7�;��͟�i���i�������8e�����SE�L�ȉH�G�a1JΆ5JX�I���+�Eu��v>[����ܠ�����i(lF�Y)�I8:"+����|^*l�F���o��{FW���qg��ʉ4����5`*��L�f�L�	���'�3�w�v��}G�h��s޷f���37ie���`!�K�2�4V�1����M$��Bs������uq�D��f�"-��G�i12>����LHE�+k��k�#W�����,��[�-���N(M�amе��z���a�/=�Rb�����ɀ�8�	�$z����*�w1Ov8�b� xK�	+���_��{�!W���`�a�3�ό�.�s�6h���V�|�_��SE�RJ���F*�m��OX:�r�\�q�;�'Qvf]�yn��b#�C8A����sN�z"fT'd�3i�L;�4ʹ�����D8��G��������u֯-�>����x�]w3�-`�sO�Ͻ̕&!a�:~��S��)��,���[�}�yz�)���y�u�Υ�ި�LC|��՗��q�@��>�N����(��I)�,2�VB��9�}������z�'k�Lo��I� �p֧���#���U����O��*~CR��A7l����
����ݧ��~�σ�f��������H��F����H�T�¹�kI,ǽ�!���Y�G�R=�mc�rM��^��&r�1�?�v� ������g����c�Y��럆,�^����o�ǈ���s���&�q�+��L�[��_�[f"����?�G��4t��@�'���~�xi��#�(eѦ��讁�{�"�Y�b֯����Z(�{bDC����R��9teaS+j�U����¼�/���wg݇���]�r��5��^)���!�*�	��|j�\pI:��~Y�Iu���y�x�X/
�m�j��5X��U�oK�ԇ�;?���͑}�/�Vx��	sY���]�T�d��]�Yg������[G�F+�K}SJ]�� �����]G��Ыj4��[�]v����)f2p��X����B��{��fU¬��v�q�qq��s��m�x���)le�՜�V���y��_��w���SR8��"�8��,�H�r>q5�S���W����*�[�;�F!��\9�&��i�}Q�L
=rO7�,f�$U.y��ܒW��?�wD�}�si X�g�g�u�O�LF��C6���и>���w�r��	q57��IrvZ��a�vFJQ_�Ey��t5nu�)v֪���d�r���:)��ep����f�N�<0�X`��4�P*�@��}L(P*��ޑ����'��tV��Gd�4U:BtYn�(q.V�BA�g'�NY�kg�N��T�}5��t+��N
M Z9`?�kZ	Đ
ii����䥅PD�q�J�[�AH_��:�zPPD�KB���@{�\�Hۘ';i�f��L*2�q�9H�*+j՘^Wn�#w�"���
�CI�8
g�
ݭ؞Qn��nL�
Vf���X�ugy�}������������~�Z$CT���4�B��^R�Os�;�P0}v_�b��6��ʱ�B��%�U������p|Q��z���e�`	����|.��Н�KA��J�tk?_W΂J@�޲�e�4������n��9��9��}����QZ���P?xŉ�x3��a�ZS܆^�� wSrKE�C��qA��[(Qݺ!�b5^��!s��K�dEm� �8�K�b+�%���(9�3fa�'E�Jɹ9�҄�޲�f�'�ⷻ��4G�/a��)i�]5����Dzߑ<������
11?�b��вq��Q0]�FK��A誠Q}�ܭ����n �K�Yª��bO˛�3����svl�|�K5R���J7ju�g�F�X^rn[�:^S�e�ӄ]ح��XNi�k�>ɢ�˗��O<ҫ��ZJ�/I���f��_8�9r� ��)>�z�f��%8�i��O�F�A��������Rۣ����x*�R�ʃ�po�h��{�XXu���l\R��[�he5�#��5A���x�<����\ac��� �:N 3H�����K����w-|J�P���up9h~s�%	���0��1B�P���o�� �� �G���yA��I�C�$��ǭ(:6�<��yO�4֋89f8�C��7��
���_���Q��k����LNyMz��B�����"Mp@��j���.�����꺮��0?��It)�ʓݲ��$��5�ًK�����9n
����u����9�ɷ
W+�4w��:��r �g{��o �V�(Q*�8��������2��G����`�1w	�E����s}%(Q��J���
� �@� 3)�I+*�+0�oJ٢�j�G�4�8��LeA��
X�2��6}�7s�2}�Xm��3ZIpJ\����f����يr��w������	3�����^��%��=�i�F5uq�(3p��Ҭo��h�;g�Ԙ=�ݺ�>�������d���b� RZM�a�6�#^�0������Ő�ƾȟ���0���	_�RiiS�9M�"W�d�Ġ]��ej�����'|���x�X֙�����p���w�4;B#2��4�	{��&	�.�5��_�~����~#�ů3R4�/�)]�^id_	�];�.q<��Zv,�K'��ڣ���x��l-0C�<�R�D|����-���Ջ�k8�GN�?]��,� �k�����avB������`�7��>��i�
�������m�@�&t�j<���1dBu�G9�C��,� F�?am�DVcR�hM\eR�g�S��FB4���H��\|�y�i-��xp���pG?�����u���tH>���*�&N��{`�[�ǚ���N��xJT�0;]�Wjiӌ���H������vy�wv��g�:�C� 
��@�f�@r�u]�"0�B�*�5�2���m�|�V��g����d�t��z�;�j|�gu�>4����5����nL�){���z�>�Y�?�4b�aKG���{�-�f"g�*Ӏ�G({�}I�@�����L���i�"�3<0$a����򚫪:[9W��l�?��(S�Ѣ�%�H�u�ڼ�˼��%�0[A�5o��*H�<�Wi��U����I�1E�%�{�in���
y!�H{{=��扼Q�L���H�a��b��a40�������}�V����p��$R�r��_�O�l+����&9oM���CM
�{����j��@��k���mw?Ag4�P"	�na��J���⸧IsU�%��k8����Y_|�:�h� ���
v���wφXdf�G����R:�:���6�/�\Gŝ�ȉR9`=�����BU(
��M ܅)4�G��<x�Ν.����o�|ˇ��Q`j`/�/_�mj��Do�ls�0ߋ=ؒ�g��qJ!s#���:����,])�-�"+�ȥ���w
�����%���诬�t�;Q����K��W���˰�C7=z�d�p\e���\,vE�t6CR3MX���ԟ"%+g���A\����m���%�a�o�'4�˸���r�ހ���?#��K�"�_�2h���ea�C�8^k�_$���\F'�O�,<��=ӟVWbc�p�W}��t�`#�A�6B+d�C�������x��C��t����eJ�*��U���6<��d�N��`�JF=	�5��@y%X$�&�%�2��p2�Fm��@��v���b��u�?W��b��zz�N���_�5������'8"����:!u�۝��������r<���Tu���=1tz�9�]C���Ѐ�Z��
$�G�,ͤp�.Q�Ż:Sh��L+)�X�� ��Z�be��p}��l�+Bh��K��"�Z{}�<v��[�AR�`��RIh�8���4,�%�p�o�tNi��<ٯ�",����3a8���Q�=�1k(>mP}/���Bi���Y=]�5E2x�}�׃y�[\q�"�h����J֕��W�|�ä�.��
'@�e0� F�
p����z��*,��1�:�� H<_���F��~
�f>i�<��8���L���m�eZr�Nr[8p���-PO%�:�k=���9�M+]}��*z�u:_rr$]ED�N� o8������I���Y�6��Č����fJe@�q1nr��In�eF�	V��^+o�"�h�31AP��RE��v���rnw��<8�9[��쑦�p�?/Ҳ�џ/��}��j�*��,������"��������(9���������$֚e��{6.[�\x�K�0>�2�m0��r����M	��Dу��@s��=NT�e��jCM�#f7�G��#(Z�V3EG�1~J�@� ݞm�A�X���}{��u_�����]&����˦ޱ�3/�?�&�Ղ׌�I[���j���lV*��{M�0�  ���3������{�B���|˻��=�6�B7u{�o[ko�i �	���RP�Yi������g,V�S*��J���,���n����y�OP�`�\�����eY�o�h��Y킹�k\�N�	���`-��m��xjH"��|�.��[��,�b����9��(3F��t#���	O-�2]"ʵ�&��f�����%Z�b*}�+��l#��U.��+��$Բ�.��I!��Y���/�)DĠN��Mu�$c��Qk�m� t����FVЌ�|'&�������}��+�k�x����d� Mj�j|Z��3|C��� ̅Ұ��C��-|[�����H6�<*�1�L��t ��]�r4�K�f8dc��&ƙMD�i~��W� �o�EM��g��H�6$[W '1j5��a��ͤ�@Dd�k�:库T?`�i�~z�8��/�ըz[Z@�e�GeJf��b���eѷ��ڊsy�(ȿ˂@�b�ʷc}�D8��m��x���<NB]�k���\T�903u�-Cկ��U�9M���u�?j��7�j�dЙhyU^4(ډ-���s�Za����~����E��L��D-��@=��#G!?��b�#��)D�Z�.�Vh������xO�o(�F�Ts����ӁBQL|&�{��t@N�E�Н�K���$h��]�.���e0�;��80Y���� ��>��>���Q";�s����0�O9ʻ��)(���,�t��Jj��j���!���*[�p|��]����c�fu�j��E���^�"�P ��}�'�]���+-�1�Ӿ��b�?N�hP���3�u�~���\�^���-��.���e�6��/+�7bl/u�4^g�m�12�h�����m����
��A�s�B_w��D��[��Pv��Z�����p�c��!��䈣w�2�DB	���s�C��һ2���@���l��ìBS �`X�#�\���������:Sy�r�L��ĕ�u���w��:�hoU�ˡ�V�^wɸJO4	W�Ys�v3U裂!��u�kY5��s�Iɥ/U�x����Dy�Gy8mVwi>�!S���S��wuyX����(<n����s�����^_v ���5��M	����^�6 }��[�T�����v
q4v��ro�I)��Ȅ^=�;���{.�>�h�S�r�y�Ѡ�Y��v��,0a���HYu�c�	�;�"P؝TT���1T�}A��Y�	��~	4m�������2BL����5ƀڤM���.�B=�u!b��^b���#����~�_I�jw)Ky�*�g%O�&�i��A�I����s�g�7�G�Ђ���9�����Ui�������R		�N� ¶ٞ��t�����y}�؍e c?8��0�u���4
ܻ탡����rSo�@95&8��Hܕ�҃��MqkZ-���x����J&S��C.!lğ��C��N���:�Ҡ k���Td�z7�;�ծG�FJ 3�y��.��R�?4[�6MY=Mk��z�ơ&WYʋ^��];�a甶A�i��Z���eg��D�!���[�!����l���״!�|�?�6353�W���K����x�`:!���#��;qz~����X��ԣ�ĪX�JQ �NFb3���q�6�h��^��[�B�j{r��i��~����	�gu�S�?T��L�:"���3�_��һ�J���P����q��?ן`n�?�<�e���/������1K�5��Ax���ts:��Q+փ�՛`��/CM0w�k� ��[��p�_��ᎄz�����lɴ��@�r:*S�C�1^��.h#�,{5#��\Ȅ�P�� �g�v����KD}���^/�AA}���F�2R���}�'�8���ෝH?��t���r�P�,1�Zw��_c&�1y����ĵ���'>`��s���㾨�Ҋٝ�X�����7������^��C�����(=c����#�)Ճ����V���J�0�� �+����T[��.�,�^�]�pfO�?8��uz32�Q鲧�,.v�pq�� �>���h9��ml��V/k#��W0��h��K9�]�ӳ?��^��G�n^����禑����8?(h����X�k�[�Sc�5h�X#�Ф��qX��Dp�_��$�&������/�HT�S�1f� 3ƣ8��E5q�v�)����rE�_n˵���#�� ڟ&�����C���@賯�P|�4����>��c ������6�<�l~�8��������C����n{��Q4:KcT�ŝ"��W�6)61�J
>y=ݹ�0U�����Д	}ܵ��PS�UP���Ȇ=V)�)�{HFrHK�l�)��p*F�pp�~E�2;������<��J�Y�H;4���p�3[WT���?t�#���G�c�B��	����x*mNu� �G�e1�a�9�� ��J�do�R(�_��T#-���Q؛|)�6�W�Ͽ||��H�!�4��4�Ϙ6���za�iy�,��Htgn�F�,�-K����%O�(wc���>!��c���߮[�w+:˼�����i1�J��H���v�n�r6(H���Z�m�s��͞��0�#���B3�
 ���z|mtdɂ�F6l�P?r[������X��]����4o��$�^�0����`����7�:� p�����f��_A�� �ۅ~N{S1qy7�q��I�{uV���i3���5�im�ǯy��jb�[>r������FRb�5�m������{��h���LX�ё��[сK�IR.�{NM<�$V��Q���ٝ���@K��Ɍ�1��S�?-W��;�Ъ[�(�'Q�s��rx�z2������N���<�]2+1���Q~"d�	� S�f�yܐ�<X�V�8�v���2��Sw1|�� ��i��5Oi6
��c�=𒯤�>�w��Q?�y6vq���rA\A�纋K���<��x�j��C�t���܃@{Gb��7x8p�.}x*��H� <ęOl�e�O���N@󈳌hM.މ9T�*P��Q"�IwPc5=��1�e�i���nδ�f��B�%i����6���I�M�M�-��V���>�L�&��v)�7��c�3q�ƭ��㱏�U ��w���$���W3
��^��=�&0�EE#	�yz�&�@�g�L���:���9r��~7�!�H�@Z�`{��^����Zby t���7 ��BIv��ń��
����	�����B+��i�Xu��ܱ�B�}�?]�躜j#W@�|�?A�e�3����}J�'w��o�7�Ѱ�S�8�dJ�C;�3��&��=V�y��� Ƙ��k��R�*�14�����d�����
����z.E��c��dE��/���PN�������A��ɨ�����Q���?.� ��pf��N7��v�
�B�<��G�E�������<�}CN�=��W��R��׆-$ �8FN�r!��B�V���rO��&���j=�s�%w
�Q	|Hl:l���l�hAE��y�bw�g_��O�a�6Пw$k7�̨����i�o`kN��z�Iq��
�2x;�$˼u_��j�:�R����'��.\o��|���r�yB@����'a4�&���^Y����{Y��{��/\&��/蟪2���r�9���f泫�'>ƃ���E=�R�P����+
�x���r����M�ʪm�#��[rI@"l�,vf��}$�B�˯0���$�c(��1�_�_�Q�x_R�F��O�z�[6�v.ԟ 	<���9�'i�Փ���`I��^}�Ш&�3��V��"3RP�OY6x�I,w���O�� �h���o�$:H3X�'�ǵ�Y�ֺ�~t�TP���!�b�y�:n@`��T��:���r�;���tL�Vv�K6���Vi~V��|�!jG�V�d�I���{ʆ3ҍ��>�h� �Jz�*G�%�{�\o����ðo�b, ���p�m�F�6wgs�7O�n=7?R@g�2��l��;[�7��Mڡ������vDS��r���Se1����n�Ҙ����,�@94�Pu+B������ۙ��.:$���`�v��b�Rc6QC�� +����ʖ��jm�C� ��	
�I�b��й~�+]�"�j|�^����Z�Q���܈����ӞX wq����6�'��v>�Ș�l��#Vб����ڑX���P��,�3��U���@�^w	jn?�Gd���D1�<eI�������i���p��Sy��?�،R��L��\O
s��O�d�+�z�P>@V5������ZTU&뤝�h�0���U��A�U�[�㔇��(�*�2����	2��ٹ�b�B�@m�3f�á4�����E�9k�'*賯�Y|.G�1�AD�c� �B���$���
e�/{���+�ދ�uR�_u?�sL	���o���
s*r{�L�����Zp�ۙV��Ќp��iZ����^I5��t����0>>��]Q ɪ�S�	�Υ��X�4V+�M��@�@�H lJ0,���\o���v� ?ǖ���0_��6�C�4��&���D��N���
-�P%��b����kf �a]����^�woD�����a�ޱ�9*AT?�K���n���9gQ�Ϸ�`��U�֞���ɧ];�8����u�?��g`��C���0��2��$���r��Ʒv�"��}�(���p�Z{r]	z��WP�3	��1O����&gn�1��	�)��"Y7i�������C��,w�,�	��}uG=��ȭh��*�q�Zߵ�Q��@�K�`t� �t�%��y�f���ύLg��;V�Vy��+�su
g׈H,����0Y�s_9n�Ѯ�Z�ܠHH 3�$1�zرN�a42��?W\`/�h�T�G$�leԚw>�6RĈ�ZE�~v��2��#{�nO1���Yam�psD�Q_�u��4�;sR���  h׳��	��POǩ(�B�7qm�،mS"�	���MS��K�&�L�jz�js���H�_�����q���_<���V�6b���X��N/�h'�r!3'��#0�m��'N��1���	��!PQn�n]���d��?�x�u���T������!������n�]��7,���(j������8����rەgI��6��H�00r�!P��D?�?��h@4b��.���bzx㇫���d}%����C��qd�M?��d�n���(D�H��^=���4o��,��7m﮳��A=s�����&�g��"TX��]OS|�Pɗ��2YZ�'�V������Vh��l���?e<��5�ʮ����oѤ�O�:Y�r.���-R�¿t��R!p�鯈����eՅ��!j�:��9�6+'��5�늚��_pq�<�#V�S���\O/�J0&=O�&�u����.�Ne�e��?�<���X��~���sh!��$PV1����<Yy��G2�,{ߐ���˓��?d��P��E��x�t}��{sWq*�D���y�4Ƈ���W����N�Ҳ�n��'�Yu�Mޚ]�w����D�?C��!8��(*��P����n)���� }��i���)�2��U�Q6�WMc��"�u �_gQ���Z�����u{C+�Z+)1�"�@�X���2��.��<W���(l����E��I��cӭKq��f�o_�c���x)?N�=D�8w���y]ܚe����!�]&[y�z� v�d�w*y�����Tt���T]�8I�u-V��ԙ��)e�ye�<X�/Fy���/N�2w`��o@م��Z��p�U3}M젒�݇�ުAW-�
cYٷ��{��Z��n�Z(�ugj��7�f��E�jx	�,)�ooʥ� N���v���4l��4������G�S�!�#�����U�-�SH��`V'��Vdi�B��n=&�I����ax�����;�b����k$Pn�e�k�����ՂВ3�J��CZ�Kd\ֹJ����T�S� ���ؽ�S^�Rt�}��*��jE�ŃmƣX ������!Iޖ&���w�e��+Z����,�S�K�+t�z�7[^΀�4�F����bu+�Q�=\Z��b�C�5�B ���1z�{)*�0���{�1�&��/�j��0��ϡ w�L[+�{�,"\1��nN\J�24���<�A]�,�롍����a�����$���.��W�C�F$7n����F'? iIu�Ńi��9��P�p~�����#�\�f�l����k�$�๴�W9;��b�LAY���o1@6A�$�1p �nc親i�Ȣ��P�-�$h��+0����c�����;3H�i��K�]H*�{�g�N��ۤ~0�;\�O��/���빃.Y)��h<�
8	�ڢ�.����⪮����i����6� ��݋��YvL�����d�zT!͜rY��1<u�gX�M��3E��;�R�V���"Հ�P����y
�ǄC/L�M�������P���o�´ɍ��'���l�����2�e��Jk�Y����I��g�	osD���v���8����o*V �]�>n@N�,j7�h�p�\SK&m�{����4Đ�o̵C<G��o ���{�L�9��� ��:�*��H��}��0eԶ �X���'������2'�J3��(,[))A�J�e�$����]14�����vL;/��'W�֮�as#6�;�^�@����e��[�XPK_,J���e�f诖���_���!�8}Mq=K��� ��)w��Ck�^"ӼA��r�x	7��K͚/��U�D7}�Ο\�G��Ry?#����
��}h�ЖC�'��Dg9�Ne����� ���
��|��%iB�
w	w��L���D�{�-�����|N�ȟG49���{\��L=�u�Mɾ�y�nFC����wN���}�N��U� b[�1lT0)��k�d2�"��.�r���˞�:���H�.馅�n�
^���Lg�N
�Nbl�5`��3q\��z'
�"�C͙j����oL��1��n�9�)z�l��/�6
P�`�\�I�	�;�=k�m�j��--�5.U+TB��ؚ�E���@��%xbb�Yܐ���
Y�iiL(��1ϧ�e,W�,����h��(2��]�L��sq���kɑB���W�#�gI�����]�2�rh ���p����sU��v"Xh����)��n��N8mxr�O|A�Ҳ��Jn/C������jḭi;0]�����R�qd�,t���<�ק��G��y���uQ�����9Ģ�ސ9pI�d�p�9bpvrBF�b�Ɵd;n|&(%�[���";W�BH�����jub��a��Uoל�S��Y�.�!zK_*b���s��&!���d�4ݹS!�#�֛\'��&:���*��C���0���p
�I�еO�7ƵwS�n���}�'��pJ$NC�U����5�.QXr�x����>���J�������1�z�����׀��"g�������ܳd�[����\�nT(f�
�T�)<H��Ӕ&z͕܋��_�X���'�^w%�0���&�]@�"�k"Du������W�x�b�7!5��SO��ïk���6�|{6��{�xlX�]�rZ�����F7�;����V�#s��F�\?Sn�7̝���z>�vgF��,���l��=��zp�J�hؐ(l��_k�E�iնfK_���pl{{5��	�q�?q�ne��e���F�K��H�7~����`yc
��|K�4ڠ��+��Ϗ'��,j�5��|\�Y/�F��Z��3yX[�v���ꖬSG+����b� Ԓ�A���S�녉�ENo�-ƿ��WB������IC��e��l�<wӜ���7x�Rv�Ñ"�F�t(�}���fy���>�y��8�:��.��	��r|�T�*=8�]�c���'��/�p���UY�D�I�
¸Bo&a��v�Y�菞�-�т�p7? ۘD���=�_� Y�4t����&Ib��\��nԾױ ؞������ht��v�pW�W���YSؾ3t�8l�e*w{)3c���]��l��>-���o�z4 �F���Ȳ������eXL<q���5�1��6��b0�z��t̂,<�R`�c��P�y�a���G�7�����&H�Y�-\�{v~T	\�/�`�M&,Z���DQ��. ���F�l��9�W��L�ɞ<����c͒���1<�AT�y���kf*P/uEM��]9�����d4�=L�$4d�f��#�{q]�P�K1�:�=�ʳ�߿��R�3ݚ�dw��P<�T��K���!:A���܆I�!t��c�<��ЁD[ΌHW��>Ѓ	60�䛄��<K����DnADm��hK#S�$�*a��O���.|˚Kΰ÷f��/'ޮ�,M�$����Ņ�k9�j{9����ypϢ�;���$�PkUI�~&i��A�M �QiyB��M~���ݵ��GR+����/������s��џAjy1�	V� ����8��Ļ�?ZuBAʵ�fH�Z2g� ��^�mx��To�|4uC5���0J�x��]p���-W+BWB�����v���݄7 ,�G�ҏ��<��A�����uk�p�����l��Gp�
B
�%���o�<�:څ4��v���y]�e�n���{YB���Z+��w���5�@�-xꈢS�ބ~�x���j��'F_%@�+��(M����k�!���И�:�d�v��M��޺��#�~���vF�k�u��bB�l���筝��8}��A�������:
VY�H�Vq4-�H��D02q�|Z��Uƙֿ1���A�m�:�������g ����g�:�+�&m���.焳�^j���/�@��E�ZQd����#)�����郧�}�?��:�Ϡ�MRy#��;[�$��Oр3U�t��t�y�ڒ�_�)w�WW#�B���׻	5�T�W�~�\F����r�A��dh��[��٬�N�����=�p�19�C�g~�!xm�0"�!����I5�i�4�n)�E��ڰ�8d����d<��Q��S����U_Q�cwZ������j�Pe�gv��o8y?���O|�7��?˷����vo����󘜼G��\?�z�!R��NZZ��
�'[�ե9��r3Z�CG96W���xp'5�K�30�4}�$H�Z��9���J2���b���B;S fC漩�=5�� ����0h�U�9 ,�'��v�`D�^\�&.�����������L���`D��/�5�A�3��zb"jf�hB�R��'���4��P�����E��j��0��OX�H��+~%���]�lw��׏:h�㲉�<~U�ӿ̔,dx��X��b>�U�q���`ODa�a�A��jlZnq�X����&����w�M6��9@�$Q\-�]���"�q�X�R俍��p�d�<���6���n%�r�_��W�7V���h�AP���V�Ť+������EH&(fǋ�y�Ǫ2`����ITm6�m������x��a��کN�)LJ����f�;�#�װ�M7�B���q(xh�-z�G��B�����	x��&䆋�T%��`�:O�K�\�=��=ߜ��!�:UX��f?T�XAmJ�_i��4׽��,�s�^yc�R?Ҥ�>BmI��;����:��3&�<p/��"��x�;�$rShT��blMRb9�����fy�����7�����PY«���ř鶳��$|� ���^W�4^ �U���6��v��b)�F�����w%*E��4�:y��u��s����f�1��I �����ʩ�u("���r���Q>u�Z�Q ��vXjk��6��_�=�{�F�~��~=q0�)#OS���S!I����O4��fD��8�l<x�Z��I`��%!����1�&6nR��b͌�?9��]G����SqK� j?��;�py���*ʇ�L^�T��pghL�8@��Y�w5Y��k_�dn�����s��H��qY_�k�pM�t���`�{���"����8#W�%���  ��`fn�$�`=��_]УwS�{��TU���{�����ҹ�������Ǹ}�D���-.�������R捠�'(b�OQ���l���?�J��9�J��:�C�D���]�N��aZLgx���0�j�.��Ɓ �Q������m��J��r�,���t��H��'v�2����~������Xx>ӳ����V�H�Y�`$���ژ8��:�ԚĞ
C��j�Cm���w�������W�l{��q��W��&qLX.��ȣ�7�Vr�Y����K����ڔN��/�Ѻ�8��*2l�^���1yV+
�����ZVc�k���l�T��W^�S�8x���5�l��sv�(II���x��v+���%I�v4��G�ĳ"Я��-���;Y�u� �6&ύV� ܩ�����ŔjȽ�|{^��RHR(f+��\���I������]��]�L8)Ӑ��G������s~Ce�O�Y�n3K���q ���u��:�\�*}�z��'-���w�z� $��#����V�� ��)\S�q�\8@�B߼��v#�'����@�!X�?ホ:=�ꍭ��QP��C�y�	�P�^ױ5:5��)�~@��>�B?�¤�A���L�a��#��p ���v��]� ���|�/�â৚�o���6�C7Ap��ɮ�A���'�E�ͨ�3����%Fԅ(>�u�E��o�BN�}��#�sn�`��Z:hk���B�bԞ˭JL��*��T�Mp�OjNwr$,OW����6��U�?�!yh�T�Y��nw<q��y�8��w�va�9�tdk�z��<����y\�E&c�d�	�TY��8fA������JN�^o���j�ؼ/3��U�wmhl�w�K����x��x5�lz�϶Y���%ܷ��U�*2B����:>�3�S��r-�)ZX4X1�xp>����D��-���]���6\�9C���1����C �ei�[�̓���^�P������Ҍ	��d��+���;k�9����ڠ���l򂥴��&d:6IY<��Vw��d&B� 0�\��.f?�E�[����ӗ4���@nc�����r�58�>�)�W��%��~�N=ji��������󉆪�ƺ�M2W
��B���/��
��|��[׍-i0â���m���h��W�Z+�PR��#��f�!�D����b¬o����?�AX�c#�bX`��{��k_��p-�"��]��@�9�}Q"�1�Km;5��(�Q,ܩ]�9\����N���.tf�l���v���<OҊ*(�*���.����鹧a�ay��#>�wF�~N�i����\�Y�l�i��Y�N�.O;�m>�g���4�(���Ǖ�	%\�$~��@"Ov Yd�7���x��R��Zk�8?.�'g7��Q���n~qqM��(6&Y���4$��kl�]��\˲_Vw0�L���"�:��X�`��V]� ��b��?����hI�E�U^h��b)\~�����%��nV-����8E����1潳���5��#�5�N�+����ӅX�D�a����E�O/D��6"��+��A�mtR0�G�Nv��t�܄o�x�3�"��`�2��o��@Y_WBp]O����S�%X���Za�2ٰ'�TS�d��D�ؒ��b�(_K�"�X��j�]=���;x�v99��,�5�����$�(>�� ��ݪ���H�Rpb@�K����?u�Y���H�݆�'���
Y�WҼ��צ�6W�eS�>z�z4����*�cI�9n�4z�<S6���ա�TvBFX�xʮ����i��Bd�SR{��`ϵ��e�z@�Z��Ȕ��S0�О9�w>����C��r*�
$�ȳ�3��?#*bCq>x�,�.�l\&�%��K��H�e?{2�Y&���慵����-\��^T2�H �2-��Q�>��_�ZD�$oUIw�\rD�aS�j�$�W�V�4���L��[X�/�{)@�H�Z���ѵ���M��O�f:��U�AL�M���{��v�RV=�}lE�@��}hA��i��4�]���W$z �3$D�6޹�~���8�Ҿ
m^T��b�	�Q�t޾�ކ�#�������⬽����T�����\5 Ŏ���.�S�%F,�l�ot޷��.b�)ڻ}�bG/�=[<�<#J��X������*(�͜)l��y/[CP2l��7�ą�oj�w�^16K�����:|��1(�?����7�E����e�!��ǉޯ����W���S`�d?'��ځ6wБS�sR�K��(\
{S�GŹ��0M�D �D=����n���t�2��K.s'Y��;�`���o{��KK���W(ǐ��G� �o8%M�쯌���+���{���z�һ��Q�p�%ζ�Wrk���1�!m�ҍh�?b8�q�
6'O:Ϟ��@LN�[݌�?=�I�G�rU�+�����S�K1L�K�|��	���F�sN�s�^�=k��3�Zp��}kj�Lp Ozi,��?�s	���X>��_ ��pe�^���O�q�h����Hī�V�y8z�h´�6��#yǉ̝;(ަA�����\��2�):�mJ�5'{�����Pn~��6Y��0kX  ꭂ�ya�c�G�w(4mb�1=M�z�r.B$�r�qwj�A�Q��!y߁���m��R/ыY�d�����r;�����2e!�~�J�X��e��R
B�g��&e�a�SFe��/5O�|��q�GW�*Q��E̬x��s�4e�l�#�w]�q�z@��hm�>���k'֒���Pg�|�r�~w�*Rq<
O����"��w>����v�e�\���]�nu��[i��Ǒ��[`w��>gN<ۣ%�=E7�������s��':":�ֶ�����&VY���<���]]�KI�s�m�cbÝec�S�1�W�����d�"Gs�j1v��x>@��J��1��8�#���B%H-�!���*���&�s����x�սmr$]�}�@誷U��¢ۘ��-�L
o��� �^���Rʗn���u�Pr�z�7;&��]����=^�I�#�p%���?HAa�@Qk;Gh��#��W���v�є�wD#`y��n!X�X��=JXmoJ�F<pxz�w��"�9��u�Vb	���L�%�&��X�_.S��[y�)T}D��/-2M����ѥ�ͭ��:
�[v��D�J������G� ��ȗ�w^�H�����\��6&�E~���W��Y�v��؜���XG�_�� [\��/8@�鈪�g��')4:0�l��j9��6���+�8�Q% ���*v��'s��|�A��?��b�4O� ��\r�7�3b�������?ͺz�¦_�Z���"5����j]������+�Ձ��m��7̊�l(8��͐�S4ӳ5Ǥ�O<�T#��u���b�v�Mp?��*Fxi���=�]���v�g���M-޲*��Ѕ��<S$�C�1�m��ڮ&FR'N���}�~	=��&�&�qO}�n�R��rI�,��aPBDEh�F;�;Jv�9�Q�F_��1əP��sm���%���a�EaTm�������0'�[�s�VwQ�2lü�����h)<��h�3�b��ϱ��������9휻���8�-�W����nN����^�D�����q��zb�{rJ��m15S�)�9ޘ�(�3���U�aHM~�S��
�ZVR?��1A JX*�9pB��7_5=�SK�P5�j�<�$�� ��c���S�\���zβ�O�~;��+ s�ZX@��E�*y��`����KP�-0،PY-H���Yc��ۍ�$�����y���;*�bY�m�A\/?���C~���e�\��7vV���<.�\o���9�ï��vY��E�rB7\��y���t8�$�.]唬@x�Mt�=��'k��	04ˇ�߃A&X�"�>Cs;�Q�IS,#�^w
b�gۈ�p(μ1��Y��u`�*��y����o��N,nӘ�ǈ�m�u�#Y��T͚!�".��y���o&\Г.�O��k'��� �cT;��Dc�rB}�Fm*mq�X�٭��FX`���s�%�Fi�T32%�!�Ŵ��m�lF �%�R��`�oGδܝ��*�����5�4n��2�G.?����+o�A꬛c��WWֱO�1���n{�}�!�1{�y�~N����KI�.�t��T�
�&τ
� �*��:5��e
'3o�>o������`*�J�`�$jY���ݛm	b��ӻ��F�;�i�L���z|mC{����L��;Hg�ah^RM��1��8� OZ��~�L�Y�����n�<	:ɛUU]�i ����2re�V�Ή3>�챧p7�� ��)��6v�"��t<�8L��P�q��~�eju=h�`d|x�'^B��Z1�Xs�L����n�5�x�U>7���צ��t2˟��������S�Vy:Ϊ������L��C,{+�&V����]f~��hb����r6���?�������kܧ[�X����Y�����a.tT�n��XQ�� K8ަ�����oԷ���x�dq��epE�5�{j���B9�hG}Y���?�"�H����C-���R>F��C�d_r5��7��s����� �DZa25b����w����P�{,T��y'�|>s�[[_$�{�c5U�ZRI�5r�Ѯ~B$IY&A���*(5�V�6Hq}���1�ucAΗ`��sl�QՄ�<���8�x~HC��c|�9�Й���� �=��^��Y3���6?U�%Zm���0I�Vc����\��ap�4-�"��o]�{S���$�Ĩv��g��T���~���|<��~)���c�O�E��$�f]�a��u����Yق�1}v����4 N�r@�l�}��RN�N:�bEb@�>����� �\&{��<��I )�Gש��;#Ʃj8��[�7}#�r]c3w"�����w�����9s6�ʆ���Ո@��Phֻ�Z��6��h<S|����"����ٳ��F\��bJ���_� �Ѫ��'�7 ��Ӝ�~��������(���6{��g��<w��D�:zS�;�[Y��uf��I5����� �lkԦBw�<�I�q�;���z!�/�< 5������t�'a��,��T��S� �p��̷��m=A��LӘ��%^���i	t	H�L���UR��b}.����'�K��Ѵ�_�T�[�m�j��F��Y��&��N0u�5�w�������w�:I3<(ujjh�6H�>�#�*�/my�M�[�̢�D���� M�dY�Gii�]�k�1���A������m���3Kv��4ľY�lM�{�MM���"�׫�̖~)7c� kқ(��9@��?���.����=���^�1�j���	a^�V+��?-��c�� ���>���V�#<��cff �7F.���qA��1
?�S3)���ׅ[�a�Pv�Wvv��$�`�Z؄�3��1�g4�n?k���F���h��<�]��Q�P�rL!�C�zC���(R�pY�1!��0�%Z��������o���a6F�p�Tc!�#c��_����T��r�������QK��F�e@v�y�v^b��e�V�áZ�cQ��=ڒAB�R�篇&�%��l`�.��D��(h8���c���(%��.p!%�]������´i7�!6��s���%�G�a�;�P�6�ӳ���3�5�oK8�]�P�<���m�1�����1y�/9�;{�.��fFBA|�h5@�����nxg/�n����1|`#�H�o�!�~���#U�,��"Ilk�s�e�O�`�S}�j�q7�1��ը��RGPn?i>I�;N�`x�`8�G��m����^t{&,ګ��Y,�Ddb#�d,.�y&���4��g���q�z��/ok�s@I�d�?��mş�<m����t�'��"a	l�!������-t��T��cˀ8�%�1�,�*Z���̺�Č)0�¦G��;0�霌(�
:a����˸��c\����0yhq�}�Q�Y(��u�#+N7����0��A>�X�/��֫�>c�!��UK�bc�`B�o��z��ʙ�r��z��
%����K8�����uV��v7x�m�K��P��"�TͿ������aA4��w��GXm�dk"�|���m�`�5�����Z�D9��z��,
�&�Q<��8�jbb�"�ܦ&�3�� ;9K|+y�V�|d��
ͷ|�ֽk�s����,@;��t�%aL�oup��K������j/�xb��q�F�̴��jaI��0iM�| jt��u"����G	��SH�ڎ�"����t j�� Ҙe/�I���Y��Q��o�4����o�$�cuC����7��՜�f��T�D�
�Y��8��4X�'�=龇��ҒZ�K�,���L�5i�&�jf�o�0�x<��B#�2x)Q�{:K��:e{�s+�.���b)l��7PhK�ͱ�X�)pEH�AK�J&�5��������Pw׵gg�#=~���X�(��t[�L�y����5V�P0��W���Y��9v���4Y���1�u
K�QM�4�FA��4yP�u��\�Nui_�砙�~�S��t��y+*���NӲx��1|�Y���ݫnE�_��u�r{q{���s�����(�������nE��g�� 3�(�#�mn�#�o��̈ATu-*�~�4��0dti7����o~ݒ!��5ƫ�8c���I����S��*��n��L���_w��{�^4�"��g��;������Sq�i$%Ҵ�+0�����a�U�RX��!���q����8�)4u�ą�������$	ѶB�30�^��d��/7�q��.��J��@���"�X<+<�H=F�Q�vA��1V�v����L��R�#x����8U�ۡ��6�����F��D������DeI��Μ�M�s�^�Y�8�r$��G��n�N�
�g���p#
�~���ޱ6I�D[/%@'q���\�q����X=K@e&�<�U���`lI�8;���i��L��w�#�����fk����b�T��<���&N���&6j���NZaGK� �a/e<������i�71`؛�~�q�Bi��� �YRڧ�M[�	�ɻWbG�ˤQa���+�%�9Wk-��dj2͓������>D�
��<Y{kC#����eE���k��poC�按@8�������쾗�_�I(�q�{L;����.Q��T��7,�r����~�#:&����G:�@tW���
���
]��Khj(��U���wl�	!�_ʘ	��ώ������o�u����iK���%����U��
�vo:v�u�_�ڷ��؊2q���u�)��0[|Q��ئ�}ŕt ��N��y:� ����>M����,�f��D ��V��ܾ!��{F$�JI`��Hhn��L{�T@p]���r��e�N��s����PY ���\���&Oz{i~O�����gP���ڸ�T�#2��ӛVzG�^�ӆy������"��eQNƸK���4L 3�ED���9����Ax�T���Y�����<�&�^S~X�@2|۶�w���21�%6"�{E�Ⱥ��X{Gve"����jJ��|k��\ʆ��s�n�1i=�יO	Ҝ��;"Q����MG��n��ڀ�ݿ6��b7M&iX1�P��8@�����B�$99&!������LM-�>�����0R%�k2��%�q�I��� ����~��f��-Xgb����ٌ��i��`B��:ޕPY̛�T�ügz�s�d"��GX��Uc�jH�����4��< �`U�NumMUjY��$p�>Mq��]�G�]�=�Rט��q�L'[)�bЌ q��%��|��+�3����
�z��DZ%@�ru�n�0��Hj�Zj9��z�fwC�r+���YA�"Qj�<�����J�E�s-��`��YE��k�����_�w3kj�M�u���5֨e�Gq��p}������<�)��Qx�}�k�'��V8�({|��\�˯�\��ԛX�t,�M�1�,7N� w��D�^��&5e��%��צc�8���č	�F�aN�h���0�W'w���j�X����Nf���_ͬ�`9aߩ���<y��c��2I���d�{�=�^�)PÐ�~6��P@��6���b�n� �#Y���ȑEFR��Co֞0��o%��ER;Je+��eq�HuC���"���ՏK��"#}6�Q�e��L�WI$�_�-�b��eͪV���d�.�um��V���걞Be٢���}ڡ`��E27t�L��M_�ɽG��<�C�4��s�]�<Gq�"���@5'��εXN�W�y~Zo<��GI�� �����#��ώjՓ�[�q�95�Uo嶜FOcO��]H^�y����;M^�l?��M����ϝ ��)�s=���QyZ��)��
j��8�k\�܂V&�
�c�/���]5F�c���+ɰ1 �u�uMB�S1y���29&8DxL�5���M��&U{���6�p���gpS4��H�]��ɋ<�c�}�Y���@<�� B��ET��	;�wûNs�.��R���gk~�������wr�_��g�60��3ó�"r���#Y�y���f��vӏ����b�M_�2Ʀ���2'���Zl~�*�#��]�_ kP��yFR�|h�4>�s���\�ы����-jH���K$lW'W�t&�ׁ���H��}23���q���ń����Y���up�s�&B���.i���h�%�����z� k`rG�A�(�
��	+�|��2�>�A��`s��th�N�z�#�������4�6
p�oiB�����}x\N�'
[5��B�E9�co�z�[=D2�{;���ـ���&��e���PTyJ%���6��ŭ>[С~��'+��@�Ca��w��"�6C�dkR�6��p:K)�:�-�$�Kp
5��jZ��ýU���K俆�v�7��e�D@y���d�:�7%���Tz����}����"P:ߜe�ܓk0�Z>{��E�纀4{l�c̽V9�2$?w�-3�Pm�.,c�^=�b?������pBx�&�,'���\���&M���I&� �%�e���.ML�������~�] �f�l���G.D�Ա���S��l5�,�qLc&#B���� W��}S�P���Z��_Q#�j�V ��j�,л���x�@Z*FΜ����	c�+v��pH�/'~��hTiy0W6eT�Z��n��7�t;2^��G>��;ԚL����~L��9V4�ro��"��)`��6wp[clD����p+�h�v6y�1����~i��Ph�i8�tqƨ�U"�|t�fl���a�*��̺�s��$�J�:><K�����?�%���8��q��o;�GW�	5Y��6G�+�B����;��D�i�I?��h��/�������i�*�?~��Y�x0i�6�/����ỗ`!{���>�C)�9� y���He/���~��:�Nԁ�:��꾸\��&��ޑ)� �{Cf��~��"�}bP@\TuUϮߊظ��^[��"$-x�0�&����c_]!O�c7�!� �\}ۍX��}e0�VI�'�?o:V�R����Ȉ�rh����\E�[��G�/��!e-���<��"�>ا�B3�=�+�.p=���`�����&�l�n�B>�,d��#3>ag�U/G��%�����D#���w]�n�C��AObK!J�������:������S2x�g>�+�?��̚l2vĺ����/4�c�e2Ǽ���%Mm�[xV��κ�Aa�2��j��^O���ρ��z���}n���\�A�a�G5y��s>AR��+��7��8a��J�����j.\h��H��Ʀ��W$C���Q���4��y�4�����'�"zR�,�
�@��h��Fk�Ta�l��o)�3��goX���4s�Q�� �d���,ūfY~w ��*��e�*��^�n>vS��@����>��^]�4Ѥ�́�G�>��<`K~ʺ����rr`3[��0ܚQ���RA�Ljd��5]��(+�p�\N�o�xǈv>�B����;OJy'��*�rA����t��+�����L��++0m�%V{b��.�l'pA��X����e8C���|?��K�]�뻻�����E����>SD���!1O�A�!SR����}w�����%����0p��%NVD��c��p���ҔpQ�G�h� ���F�%��"bW91E {����K���|e`g����e;Q=�E{{�N�*�f"����~ƺ��A�=��T4a�t�Ǔ>�3��9=3��d��w�@�� XG�7$܊d�!E\3#��y� ®�0w����]ar�JQ��>(#���l���^.�`�"8wezf��aY�*Nr�uA[K{��u��|Mh�9��\� n]PI��򤟏~�~�=�R5�-7����.�2<���;�u7S�]��"���I��̰<�u</{�V�`�+�����%�
"D�>ur ��*�]>2��#���|��q#r�a��K�E�ݧ�$�E�Ga:��{B��I��3;�@C�?�~$�,���2�w)6�xhUU��U���Sw�5IaFzd"�/Y7n�>$`e�H�s9�F��2���@�@��9�}"�������F�[������8M�F��,Ԫݽ���y:�������nB�+h�	���wFd��ҙ�\����M���ѯ��wzx���oR%�`*1jX��"�q@��Aa]V�_�W ���u�D�F����H���aj(����_(�FՏ�y�"~ז��c��ʸ�)J�2��rG$���_c�a/�v���uGD�j�2MT�ξ�G[#t��o��6� X1x*6<�2`��*�J0e���lXp9{��|-��%��1eHO�0���6���Bv�Gƕ�~bD�T-�P�#��Vؿ>��U��3�J�+ߒ�u:ipN���Gh"Rė�^D�I�./ :��o��Nz�H��O"B���ݧ��$
��Y�� Ro��B��s������\䣂��[�R�m�<p�[�n��J��Q����x��C��87-����w����'��߭�C������M�+��i뢁;2~�7�RX���"-GgI�X�Q6g�� ��D<LqEM�
�o�c����e�&^@�Ru���]���5%�S:���IΞ�C���P�DM�S��G�N�E�nV>�G�WW��g"x��d@ڱ�e4\%�Y��⋖�f8gO~���P��X��[5s$�m��i�?zJ2R��z���|Po�36M��[�Xҏ��..E���B]+nk/4i� |-�����'�n1�+����z�i��x���	%����y��7fu�� _q�~�Ɩ$_��޽�<rei�S_j�?�M ��ъ0�bs���q�/'q�_�JaAs��+�SI\D!�7h��}%FV���ch3�G���̫�E[+[�����D4~@j�����g|j��ۨ�6���
�Q�+��,�-�F3�}1:hL/���M�Z7�)��cϰ�nQ]��f LO�st��Dw��9 ���pP~/�A)��s�-{Ƴ�
eя��'T�v<ET4
��`������J{1��0���Y�N������W]���N*�T�=׶�ܜ��tB�-�T�M���\���c�^чPǜ `.T�]u�o��*S��>����$ڡ\aJ�����[��r��,�D&=�צ�5
26?d6��1r�b�hs�f�`���_��8u/��T@����i��`�EI�͑��w����Y���}��ɐ�;9��F�����[5#.
;Ԕ��\��H5/�����s��Mw���7L/�'���`^�l��*��
�3��<s��$0��w���#)��\\9ٽ�0���o�Ę���㓓��Ő�@4�~%�����viYX�xH7�gK��~��D|�����K�L��-`������@]u��[#)�w@zK����3B������/��0�,M��W�s����� ��6_������wrOٕ[��F�r�|uB��� }4��b'u����kgv]wSVS��5U�b��d.����a?�"�+_�8��F������gy3���'��GE��N��)'�_��]���n����rw��ɭ8q�!fԭv��ҠZGV?��0/!9쐦z���WR��P=
MɱA�|9��E���ZϜmT4� 5V�3H��%��>�{Q5��G:@0wR,(�h��$J�H@�PD\�`k�$8^/'k�ݻ��V�$�Q�B���`]�5�S��fR�e�`=M��72��U������k��6>������!9��g���.�0��hG$=#���<�(
.p%C�����7�����y�=	#�9D�9�q���@���op���t�wX�հh��p�=f X(U6͂D��0����"� z�R;�=�2�v��!�:|6MV�Uy� (���XwB32�ξ�璷��J�o�<��V=�ug�f���r�lU�f��K@�_��r*���un���/Co�'�e�v�8`�{���#|/D 7��+2`z>��+��e�R#z	Bzۓ�����4�b��ǂ멧�5��{.Fap���?��.t���q^PQ&Q'y�<��ǋ��z��������Ϥ��eu}��C4�h:,�$#.��]�!���p6�'>$ �0-������	NΊ=Y䟬q���^P�q�ѥ����c��3����@�ᅏ����Ӹ;t>2�CR|��a��n��>���n~����a5廞��)���+�y�e,�9�elX�g㡴�?�m=�[���x����B�-���n�>��h$c��ISo���;K������X׼rj��ǀ���W����;����^٭�� _�y:�k�Cu'�2��U|��t��P�;e^=��b{Uf�]�������g;(�7ۧ��Cg�!`k\ui���k�/P���l�8��=�<{K�>2��w��ܑd�%s^&ΐ@���n�i��H_��֡���T�8���|$ߙU�|�d7͎S3�=����7
��@�|2�ӗ��<��#,�
r^�'��:܁z8���c��!�52��6���Ak��шGE���f���N�X���vOh)��H��� F4nb����*?���rxlO!z�Ix���ݱ? .̀�h��R��f\�L�� ��٨>�4|D���cmyL�
c@ "D־��j�h�F�Y�X6"x��m��x���Y2��v�2�������������p� yZ����"6g!���[��o�l+{�*����oK�j'�|�&c\��=&�{�Ƚg� ,�\Y���[���ie ������3����,���q�i�cD1`>
����u,�U�sE�a�G����+��0���k\	[j�XMR�[��U�@��$Y3( �E4�Π7�52W��2-�x2�=��}��#���P؅unM���r��ɒ^���%[����p��84�0���[e��q�	n��� �<r�����4%= ���p_<�G�&P'FQ/��}��+ʁ��(1��/���"�\ ^�.?)$SDK���YN����aZt�����Q�7)c&d	��asA8
CE7[�ؘ;L����涫;�:pxk.���A��%�4W��/M�q8^�Bmk��K�_A�W���݈��o.;y�"���ɱԚ��EA�z�Äf���j%�'1[9j�@�D���_VDeBU�-߭��P�0!�q����ڻi.�U
�Nm�W��=Y	f�J	�B����ۆ8r��[%���W-�&Eo9|N�J����uJi�~a�E0�m��� ���hj�K"�=��uȫ��E�+s�����+�N��x�&� �ύ��g$j�@��H��ԋ�C�d�5�~���'���������<b��õ��Nrh܁�1��8Rb�
�fm�GE����##	X����Z=�l�3b��LdT�mz&�`Q-B.������t�����z=�e浒M�a�ؙ6`n���If��F��O�l�����ϑ@��D�;=���H�v�jc���0�ƭz���q۪��|ޖ�Dn6\��T�ʬ��x��Tz�'�|����@��2'>ܨ3�L���+���We�H�P
(r��of��+�zHQ63Z�(��)^��-@
�N����z*W$B�O���#�ۼ !+���2��n����$�/
rT���Ѕt���:���Wli*���,�߅���͝`�I@ ���-��=^��Hq���/�V���*R�Ý�i�9=���FL ���4�?��Tk����WT��C���HP�����jh�?t��u0�X��iX\��90�?���,�Z��?�:$�nɯ1%IՁ�5�*W�]ԌW����k�,���L�ҋ�-�^,���%g����H��	��!��l�e�P�ޖp=�5�g�zn�IWLեaGlp��Whզ��M�f�1ML谲��0����0H?G�����������vs�?�8H�Nڰ�ki6��2!�E�/51&�Я�L�P�la�%�+[ p�|S�skڍ�&��^B��`���iyS���%��	7��`�>���G[�Q/��,���J�L"�$~�T>
W�p�BEq�r���ዿ��$�h�¶����w]b�%�xG�l���g����V��I�Ⲱ�Q�|MO���،��ިq-i�w���{�J`��6wj�Q��_�0���mW�C�w�ך�`�P����g�繠O/�x�=-�?��8�]+���_�k�i���/�u�j\OS��ݡ<j������
��ib�T�{�Nr�3�)乪��,�ԑ[0�������b��=V6�(�ly�=�V�(RH���˞Т�,W"	�6�S��0�VS��W�1�	q����1|?��\[m��Fc���M��X���� �:�
�>^ �mZ�Y����0����"���v�=����觘Y�:>�3�P���� I)����,�p�a2q�B�A?�Iw��
���4�2����M�Z��Ђc��/L��(D!��Oe#�����n��P/&�_4�3Y=�UPRQЦ\»o}�\c�i��U�������|��o@$���. ��C��HAN2<�����#i��x���I���� -z�s����=���KV��zz,Qb��saĄWʞ�0�Z��/. ��6�~.�4c'�Y}_XH���O"�J$9�8���5�M��昝�a �Ү����c����!�~ ��J�#�іB�^0Kt$-,�9�O��*�N�p��66�1�s���ۦ,�Q:z�y�\^�j�gԨ�⭱_k�������I�x��ǯ�?�i=�4V	]O��ki	Qh��2DҴ��T!�*��T��27p�B┐�Âд~��It#��_]�
�"�tsW�+��|d8a���b]��*�H�tX�Eʋ���m% e�Q*��I�d�p�Њ��e��ʔ��C�uZ�o��/
�V�'���b�����j�B�v��0l��4��Pb�I��26�F!�>�!��� #��2�S�7g%<b*Wd>�� �z����������p�JwHmF��j�D\���,��l19�	���C�C�R���?r�u�x�%T$��S&�,����D05��x+J�?��%�ࢀe�����۝�	M�F}�Q�3�VU��LQ� 4���ÎA|:oQ� {�/i�v��AJ��	�f�� ����.x&�ʡ&�Ӧ�r��( ��Y�OD%Q�B?�f�7M��z	��);����0�J�(/��T��yO��7Ź_������!�I�F��D�����E���zn/��J��VFE/��A�u�GZ銩O��Қ�Q��A��I����T�  ��0F��Lv_�q����E?@����Jl��~Q�_�o���u�zhT���t.)������n�C$���&���z\�Z�	��B�k͔D{_��n�9����xX[�c�5�^LJ$,������Nn+�J� �_�S �4X�8|��x��=���8D4�����w3�nr,�6:�0��N[n�(��Ÿ���=�o�nG�k<j.b;X�Ӫ��tJ���"8Zc�{���y-l;�m���	a�<Ѱ�h��2�@��-�H��{��;ې7w�.�Jm���[��ۖ}Q}\��=�h�+��'��F 2������"���l��J��А'q<R)���y
iƱ����MCa��o9,]�G�f�\4�ح.b��5Ln�,g!���(��F:4!��Ne]Mu��P��������W'݁��;�����z��1�m5p��5��N���T�cY�X�sa�	W-HL��G���ݥ�<=a��U��ƅ�SE�
ǅߺ��Xa�7PB�� �w�T�A킳�Z�|�!xOX#�:ܗ2�:�f,��J���(:������FE��)�M�^����6$7����ϼ֨�~�ڭ�!u��ԁG'��"�����0D��H$��	���r�I0@��.�k���w�0㒁���b#���
;Q�޿�j���ԝ�_։�]�̴y#�nA�vl�4%Ma�`��]yKAS��=�oأ��B:tG�Sa�`�շܲ�����ꁫ'�X�a�H����
F�BH|���;.p���ܩ�Kh�S�|6¥���_B�R*��������b��� ǳ�qt��4CѾ!
[�w���C�D88>O��K���3k jnI����z��7̀��n�c�����7C�z�>'P�J'�FRcNɒ�6i�����?�qCVNF����r���=�}���3�a�r<M�m��*�eF���E"]��86�;4����X_q˕9�t��sg�)<�������L�U�@ �)��t�E2!�B�}���ͩj�c� ��{l�_H��w�����R,A���{)���׋~yhKɍ�f IZ�]�?{@~^�	ҩ� ��/����k�R@B���
\��,
�S#�:hѩM8��Z��W݀�)`| � �T|*��A��ڲ�];�O��C8�B�i�s)���r��Y��u�s�Q�^3�*?p��_;w��Ї����=^vg/9p�Z���+^٪����H��j�/��aT(��,:�~eW4);P1�Fh�e���!�gk�գ�5VF'W7����_�w���[ytc6�>m�t����*�qE�n���E?xIszEf8���n�MT���[!0ev>��wl;d{�o�)�D�����ѐ�wP�Ί�o���3��6�e4*�R�E{	�kٓ�7םU��'�_D��E��k"-�o��tb�u�M���}p6��@Θ�q�&�/& �s��F=�f�( c.�kerp� z=̲:�S+���_ԾTJ0vXz�3* ���S�r���6B��!u�������;��dPЃ�<�j2$�$�B#'���� ��&PM+��z0C��Wv�ϲ}??-X�>z�U��$�r��n��;Gk1���i�n�..���;$�O��xOG�W�/�����ol� ���x��rl�1q���QV���PX�w{#��lv��NN4�����Pu��h?`�?�)�!z4j�8��z�ؐ�}���S}_�C  q,U����C�
���_k��u�����d��NsN��:;?,Q�m9��хKKc�����_N���` ]� I돉�D6U8a��<���Ł��;nK�P
���j��ǓpQ.j4-�އg���]~H�KY �V᱄�qdYꛌ��Ci���ټ�8�U�1��1ɒ����4z�)��#:��v1V�CT��ʈ��zV)�<�fyt`���l_��l��	�����/7�G�}:pj����' *���(��=\���jZ��沥we��[§�=ɽo���o��ϳE�ї���|�IUN��Si]�=�eI�������K`Ί�^�pq�¤�2��ܸ�mC>�z8���9�Q���a`=��W5������"E����0nW-���1�F,wM\�0{���Xw��S"`�v��@g.;[�)�:L`)Q ��@�"��ds��ΆPŪn1c��/vsG����P��X���+��L�5���*���.�G~����I��H���S
�JտEfA��n�\^���fˆ���a��/�DXO�m~r�a`���v�RiY���8��`X�C�D��y�YO'��H�a�5S�&O��[_�D�n�%�ҥ2��L�N*�\�<�����~y^�I�U��BߥY��:tҍv�T�����Pi�#Hݳ�m�G ���,�H|g���E	K~m�ʖ�� �Ue�&�@�<SVq=�K���A�h\Bo(h�G0���R}���y2u�!��aUĽrmX����Ǭ]{��Qtω38���|��X=��7|�(�]�K�K/b>��	�};W����rn���wGI拟On�.x�"�M�"�gF�p�(t�$�$��Oz�cz�
�e���PvP ���Cѵ���^�=�U�B�B/���&U�v���*k�HR��ܷ����xf}k	�������[��C�@�f ^��<@�߿b@���>>�y���hU?��v�"tM[���>�J?�ea{�r\H����O@ޜ�(>c��Ο}j~hvO��1������O��Ug����GC�QR�X����Y�v[��=����n\���`�Ɣ̿'��oyˡ��#���N�#e�.׫�9vQ�>�-Ǆy�ED.�}���7�,CY&����[+��U��%��`������I}Zg�K�X���'@�:����0�G?��X�6ïG�.q{���*��M�˃�y
@��~O2�?ۇx�X ��y�U7�|�����p����t�����hFHI_*S�&�)�J���"��7;�W���f�}�����ɾ9R�'��7E;	i �^2{}��L��SDwC�w-�vE��>�~��P���*J���d}%��wǫZD���4سrl*x�mk�shŠI3
J�St�0������ɿ�^��T�#�@�����R�Gv�`
@5��j`�י=S�����ſ�������"Q` ��ڔ�T]{�eZ�O���.|���=��ゝ�Gl ��	��}3MH>aFk�R0;���w��l�IDD��ڌ(�"pw��2�{��:���C��Z�4y� ��%�1�S��e<�A��!��m���I)��O��G�Ҋ>�i�5�[�T�|x<>�[-�>����iq�uc�<i]���#n.h4Z���j?�����2��uc��Q������ �7�ڥ$�$W�Ϣ��m��9?�e\�#�A2%u��e�6�b´�^C���h�P��=k�雑(��
��\��eń�$dF�l��h�g�[Q�O�߻ހ�D3A���@4��X����`Z�]�}�|�W>Kʮv�F�gp6��8,�,�mj�t��}�&�ǒD�e�ʅ��Na�y��f�s�I��l�,{_�y:&a���$؄?C�k��3������݂ӐG3g��)��1z�e���PR3�r�\�~��!&�XO�T�Md}�:��0����ҢN��4�=գ�'��X�x|����lR�л~�}1V3=i�8&-�G¤_�����Kn��mB�O��<�0�0��<xSuN�lI�H+�q�f�gfY�����s�d��k���UP���.G��̘X��U��&/�c�;*7�C�ɑ|��P?1����1��䳮:J
�F�]2��,�,m��B���X���p��%��d��xC�ROg$yNU��p�lկ�P�n�i�s6�/s�>h�����GN�32�]�ڰa�R�8�&%��/}��>*¨$t��U\�*�>�����Wa�%���v\UL�G�����M�G�>ۿ�'E�
��(/9[�X��W����L����*����� z��6�mҸ� �fQz-�`�$�0�U��}���QX�	%Ϡ��y��ʞd��3 ��<���E�{�W
�3L�>J��y�Y���MX���M�����Zb �Z%=ǅ�o5G�
U14x�v*��x�2c���_.�$aI�p�Eg@؇e��N2�����Z��}����.�D;݋�2��>��-~�! ~��Z�M�޲���m����)��٫��}JR���T���~� ��֥!	��7T�t�]%	������
n6�Cu4�]��T��������3)o|$rz^��<^fOQ4,����e[}.����k��KWȰS�L��MD�'r���h�E`��}�
ޗ��m��eP�j)������6Tmɾ�V�ViU��2���({m��m>0.X^r'�y���n�	D����vJ�]�+��iYe�qB��d� <>}�|�h��P_C���\�X~l��B��br}Y2�T$+�y/N��ŲC��Xn����Ldޣ`e��,���v�:���c, Ӄ<��L���q��5�N�� ?,�A�WR�%w-�:��W3����k�Y�t�ާ�|����|���?e|cY�x��xzT�8������ύ.+����=��1Ա��T��$�6��6j���F����KΨ�m��1�7�ޛlL���`y��χ.�֣;Ԝ��j2Ňf�[ٰ�N���'1�Pϓ�8�7���Q4pם�==�f�^�:P�4zEp�0�_tڱ�#��z��Ę���bӆsF�j`����LkȬg���qP�  \���/m���:�I ]37� ��X #U����qN�8��˔�S(={�?�3�^Y'�� ��](��\���6�&��h�R��ń #_w�V�ۇ.�+m�����>�K����a	qg��2���lࡈ��2��۹��+r,�d��X�uz��}�N��x4M"�-ױ�����5�1���N�O"�	���me(���4�:�2͚kMx~���^����]�ߣ�1&ZHW�J��P����%
�⑾�y+�Wjw.-����-ϣ�ψsOW� �����b8���l�g+�̋z��ڑ��o�C���=��:�΀\��mBk�Ư.�u���X���	4�=��*&�M2a|J����h
������擗��O����-*r1�e[q*��;��X�?���4�����,8RՅ��X�����o��q���u"�@��UK�������jdW�������ÁRN�\��T�6�m|��7�;Zp��!g��1�9l��>-[Ws*��zs���F^�s��QX�r�G�%3�0JÜڢ�`��:�C�i�0j�ѷ�#����2���<-�aη@�J&^kK�1�305ޔx/���'w�����V$8I��8ϥ����ԕ��n |t>�����Z��ÓV皫^�Z%�L%�� �'�tX�^�dܿZ6�!�A��O�T���
��P����ڏ�6t��C~I�O�����W�������	������*�?J(���g���|��t&�`f \s \�ÿ�
�{����:c�%!������p�;�O�����Um��qp��+#Q����7*;��Sŧ�2�
[p�D	{RVFD�N�x�ǵ�WF��µ�>�������Y�Z��h��4��oR�O�y[3�&��@A$c ��h��e�@7C6%�N1���`�(2k�Ye�1���5��_js�4��Z�]5{F͛���A�ŕ*x����>LX��p	^��Yu���Oj���Ãc�oA�Ƹt�^�QG׈�|���yܒ;]�_�`�\�9a���v̋*%���oc&�F�;��q��Կ�:��|�'�W��#���'ub��>1J��e��Ya ?y�%�n�H��ă�X��;x�{Œt��:���������!;>����&�������^A�ߘ�w��hF��c�]�<Y�<5��Ÿ��v$m�S�����Y�
���4U�\��#l�_c���i���
�����9vLB�%-�5T{��*5vL����ۗ�?:� N��)�E���ko	�F6)�AYp�W^rq��BK��xQ�%���z
�螝;�50c���h�GKƆ�#�c�V�  �_�Ȝ�c��P2)����mC�^��q��^�4�	�*�����3��eJ�����&��e�t!���ѳ'b�싨��edr�B+o/gC\Z�I܏7��UjU�S��nh3!��h5}j� Bq���N�j�c�eQ%��)2�/@��=LA9P[��j�Fٖ���JZ�y�Zo2<��ݽ�h���Ɋ�`Iw�^2_�j�L�#¶j�ƹ�j_��׮u#9����{�����f�:�Py�F\χ�1)����Qw729rg���w���
������\�u|�������ƫ��)E�GV	���f's_���\�q��7p�"��4R1�ӫYqiF���u������-|a'���+{�}`�#,��T�sm�*�8���0b���	8��'@QV,���<*�,��K��|(�~�e�Ԏq�H�o��r�'�O�Z01p:���B��Q��Υw*���U�i4I�A����X���<�Ţ��W���|�NBI�j:~L��Ph�!"VC-���eO7>��诀�:~4>�U�3Ui޴
6�W �y񪛟M��K&i���f�O�6¬��t����iۼ�t����8�~	�^Yy��\+
r��i��"`Nĳ�m�ϰQ�,h�8�vբ�ʞ纫�_��?%e����`���^�N���
�� �[�����2DZ���CΎ�d��buE)���<;���	斣���H`����|bya�}>�şT��F�sH ���%��[V����c�������1����&�e�9��98dkQ��`S!?����K�F��Z=��w_ϟ�M�����;��-0	�*�9}�˧$/�8H<��=(v=u->-��d�^F����sU(yG&--���($W��@��m}�6�H�"O���"-yy����X��J�/���(�ik�6x����[�°�7iX*���a�زiˊ��`���찀b9��5���vt@�d⬽l���O�0t���3;)���,�U I(B�C?mg�8V��>���t�����X4
H��_#3���^M��l�QP����jӉ�Z��n8��T����l��P�(|Ea8b�r?�-Y��.`�_X��L{�O��	C��ٕ���Z��)k$�g�r�گ=�7�Yو��D�FJlg:�%�찖yr;����eO]�9�������-Ƭ�KEK57���|�B��1ݗE��;��#�E�u�|��^s�]C�d�X!�2}�XBTޟ�G&�Ā���<&)FM����Ԥb1n�?���Vj�稜;���B6��z�\�ǅ~<W��m��O�$�$��v"�EӢ�II���j2���~<�(�O���@��)ɪ�D.\�Yy�S}����1��<��iڰ�RC^�̸������@��9�l�SG�76���)=<� ϓ�q�@{:�t�b�+j���Z1�n~A: ��ASU��fm��c� ���/���u�$z�Z�͚��5������'Y"q���ْA�0#<W����I�4ɲ����ż�x�TB7�!��`�FY\=�&�;���a��E>�6���ݺ��ճ��ҊAw���%�*A[�nM��TZ�F���@b�H��O��z�x�N�N��ə��b;0Nę�pm2c�����nX	��/bOD}��t�����ȇ���Q��yº�J�W
,����?���Te���:��m�)Yf���q��YA��r�2 �>��8k�{ן'a��m�yͺD�k�b�E�eۺdB$��s mF��@��c�z3�J]�������{@Bp/�_[b7�Tr.��Y.�[��9�D���XӞ��-�ZakШ����6o�[8R���U(����`�N�
 �����j`;b�I�;��Ro��8j�Iz0A����?��H�̎�"���[�b`�� "L���(�ի�D,����7���M�S1��Q��S��-�F���`x�1��}�� �`�~�r��=V�&��`48�^<�Բ�Vt�2�'妗�>T�7Ӭ��ډ��O�qba5-��/�X04�5_�������q�u�Z�A �!ßL�}49��͙-a�'��N)�:WVo�����]�
���`}Y`m��;�A��&}+o����~��ˮx������7�4��.t8q��#�*B�B[����}����s���t�H�K�y��%��V�\��f�V�������W2fK��fs� ��%�R��ݶ_v�r�w]Xr)��g�J`�֙��u�xС�ec�z��1��ʡ`��ˍF	K�π�C'���!�ap��\��
�Q�)!x�ksG@"mEa�r��7��[�i�-��z��t�Y긚vЃ+���G�A�YҮ0�_���Ƀw�S����ik�G��GP��r��q��c��Fl.Q�[���-��jP��'Ԉ�|c��M�TE��c��p������T>j�[�=�W=���B!ߤ?+��ď�	ʲ)�����XViA���X���`��*��D��H�I��M��*�**��}8�չ�8��)�O��rЮ�)�g@U���d�?�X>:9(�y����>u�/�>p9wA%��u#9ר!����(dfu���.��U��#?㢫�]i�٢��Ժq�<����`1B"���o:��YW9�\�y��YQu%��/t�{q���Jm�T���R)H왶�����g�`[����u݅�p���^) �?NF�*�|�45*r�W����㗈�|{�P�zƶ����z�=��v�!ݟ�ưϗ�7>瞢�v��:Lt*m/�sK\��C�_�*
�����Cn{�V���"���*��mf5R��٥�4�O�^��*�|��s�B��H�LK�f��i$�K�*V�u���	XG�6�_�鋳/����qN�����GZ)̎KaLb^]�>O�.�/B�")̭^�\�)�s�H<	��R�,K\5���f2hC�\��n݌�W�Bs_��y�B�Cݒ"�I��Xu��f��Οk年��Z�8�d����|����rg�~7�>��[+��yJ��I׫m�zt�X�-���:{�����-�/��t�"�z�0�P�F�p)�����q}�yy_�T� �	iHb��=zb����� l��7D�Kf��0�����@���A������*�<D�c�{������/Y�=-�����n5{��_`i-���]�����z=_�����vժ�����P7v��c
���6��ҹ�V��`u�m�=�\�4���C�gg)�ۆ*���"��`�����ֽ9�_ɧ���$��0�`%� ��ZF�_A��E'��0�xQƮ��tf�j��]6r��s'��'�FGӂ�v�4��\xie��\�璦���_� Z��WxFM�l�cq\�����D!�7���a)�H,�kǁ�[�J��8�
� 5��vi.�e��K.��bH����e��Β
�3w�L�:-�%O��t��x��/˙o�/�a*��*s�j��g�c���/�%���Z'�K�$| ���ۨ:)(ZT�@*4�K+�Ʀw ]�5|�꺴�%t�=�^��U=t^ś=�a�'��\Uf�Ҭ��e«D
* �{�=5����X�!S�2��K�L:��4q֟,_���飗6qhT��f¢Q�N{��`�����s*B�;��=��~��15Vb���w�i��n�x��d�{ "�=l�1蹇M��� ØǺ#���*mw�0�u�D����y�DۃQ���J�岰1�x���T�Ҁm�Eyx����q��Jj���?����<�To�<B~��K��=�<��A>0�'�czcQ��i��f��w��LW@��b�@��S��i���[�A�k�H<�P|
I!&����.W�{\��?���(��-��u�X�\u�%0��GЃ�:uÙ˦Ʋ+<�����_z4�����L���HV&�� �(Oa;B�yL���Áp-�8�̇ښ���B4S��XQ� 	���:�DJ��2��T<�[�a�O/�ItxB>!��ط	4� ��]�F�K*�h<	����ld�ʝ�%:��o��ʶd�RŦ�(����"��y�M���}����@mA��K�̏0����I3����QM��Q��G�(MVT�,���<�-}���K��6��<����-N��8H�fL2���oljq��H?5a����}�~R�W�`��c3��[[iټE�$��
j��n�b](�v��/o�NRN�.3]{���ԫ���?_����[\~��l�ܬ�'��	������n�e�ݍ�%���P�ܶ��0TcMKg�g�,0a��ȋ7�L�\(c�m���QՕ��Q��D����.ݸK�x~V�g�G�LB�;&��咮~��ѣh��C�@D�
�|L����v2��72��d�w��%62Dei;��>U\MK������ ��Qϭ"��#KSq7�k��=�����a�ٱ~T"g�g�o�gď�1:a��B�����t��v���ǂ����Q;(ã@��}u��n���#�A\�{
�Gz�XWU�h����YY��ɀ8���\�r��C-�j��a#���-G(Ǥ3r���p*�f#}>_��/�,W���ċT�H��K�M�
���~2{Ui�B�>	? �|�kO��2)�cQ�f��P!G��u5�g�±/*��ț��m�(%��j��j5k^K��[��5����G"u��͹@����;Lc�)zNr50H �?ͦr��*Ccj�x�z��񾺺�
t.7+7nNT���y������4��޲�{�����1Ѥ���.�����7�phV­�
�Q����G��5�T9�zŰ�!��[-͉��6�u��!�za�N�k���-IP������F��0�\н��ײ���}6�I��Ӷ!�;�������a�=���\�n]�\�ќ��И��Q�x�x��خ�*N_ja۬����>s*��L/�R.�r�z z���ۋ#��;�o�<:��mv�\:m�4%�{p�u�U5B����s�Μn�)�9�y`��)���&Ձ��]��/�#�w���������Tn��7T'4����ieB���"�ދ�U�jS���bYI����G4����ȝ84�`��O7�K-I�6��Ĵo�Ep���%��%
x���/�y<I�*]�;:II��YC�Z�!R��Rl��
������qg���j�%i�Fu.�Xf�9�0i�i����Tx� �:빶ҹP��.*1�4/�
G�L3Č!�Mڤ<&��A�*�����Ց`wcLY_��J��Â����tQ��1�����5��@&T��t����άH+��/��~�hM��A9���� o)OY�P7skIH}e���oXR d�k��'�����ⓛ|>��l$��/*6-:��v3���F���q�6$�Ze��.����4�u�-K���t��[n�u��~�����ɘ4�B����Z52hb#�1/�TDJ4�01Q�z7���O��̷܁u�{���NDl��CŹ3�)5M�hS���e�(�D������Ӄ��m���1�^���]EЉJ�7ġk~��8SVG#m�Y��f[Y[��0< �9Hf�;��$����8����g,�z^,sF����Ч�q������T��T���p��"���>�LL�T�Sg�,U�*]tr�sJ���pw*0/A��^�b��isƺji�@(�R\
�9��I30!��`�3�U-�s
9���j�mqr����V<d_s�b_L ݹXG���m�[Н��mݕ]~�I���V/�N:�ۆޘT�nj\�8ߕ��5n=�D��E��w�Q8�7˻+�XA?�=B�ؑ��%b��7�Q��z��8A c7�֨@m@����:��&���~�8��;��O,�|��������P�Ť4+�yD��R,�t,��o=�!��!���M��@�r q���`�L%�Պ�z�-�ܙ����ϓ�t��F����y���ǽ�;�K������&Y��wFIV-Ģ6Q���PU�t�Q�����NV=�+��W!��_W"t� .����~}�Ii�^�>���\?P^�A�4YV�Z�QF�5!E|����x�V�?��ŋ����hI%͔�,M^��R��(�/��1U�
�s���1�����U�=|�=��K!N��d�:��<L��0�s ���Xo�'������v��Hf?��t��l:��+�^�(�q��ȫ+.l�_�n�wM'�nr��]9��Ix��]�����c�φ���|w2��ZrD��=�, ZɌ0��y�!��!l�Z�4����|ͧH���L�)��W��1�k�c
�}�]Q�	��l�pF&Y$�X�D���=T�#3;���v�6E��._�J����CL�Y�
uA_�Y��n��;��	G��:8�u��������y!NWj�~��v0� �]�\�����)�`	:+�n�u:��:�f�>*-?wx�N9�"(�R�*G���)��� �=�����$fG̾�\ً4��W��
D�}�ǟ���PQ��䌵��"!�]k�kO�{�Y�& Ůǭx�f@�b��2x�~r�6���텽�(�3*Ø�2b�
� �Ѵ��ls��^%���ZP3��xO!G�fS#�\;q%���PRg���Vv�Of���O�}��$�	5���Lۭ>ǻ;�Rk��%�ȁ�b�N'����c��tW�g�2��W�O�g�K#��st��E�!�,d�C����j֘����Y��C}:m�5$��pHF����K !��#�U>�U�_��j��En`�l�(?��t�I9�(�h�e��:CU{��Xj6N��dOЅ">������t�x�	ERWD�B
X�p�y�+N���(���[ax�G/�S���ׄ� �v�4�]��U�*���(<���0������� X�����+c�C���
�A��z�,��Ė�k��m�J�VWƂ�]�a�����:?��jw�%tоltq8��se���1(��	W���A�lT�K!�Ѣd�D)Ze��U�����z��(�EC����
�r��Qa��B+�.�2 ^�+_�Ql�&�u�����n��>���_�����U5�A�����Ʌh��I�/���U�K���-Bُj�Zx�&c����H�����w|C�k�1H�^`����=�&���H��N���n-9����]�C�[������pD�P�|Þ��u��"ŕ�T�"�Ep�ѯ`K�j����ɒ�.�`R���4�h���ゃ�)�9��" �y�@O1ZȎ�~�U6�U ���nl��G���M)�+.œ�pa�ɥ/D�8�H���q˭g��ݭ.��Ĉ��|�B�k/;�a�.k^��D�}Y�`ge��\곢t���)+�w9��z����<&色���_O���[l�N�Wi���6�����[c��w�^O���g�ܦ��VY���S��s��G�O��Q79����`�	�g�b��$4�5���	�C8Y�!U;�,���.���s���p�p�/GoѮ��22�-�4��-�k`���(4aXFl؍��Դ��w��V�i*�Bn���5��v%!)���Ǫz���(d���Juۂ�2��>����VLs=�`I���ALW�oG@���:��B�\�x���gf�Ț����5;����j�[���B_���E�7�AjB�/���HS�HfI��\l]�\��.���k���qrX��Y��u��o����PĐr�-F�Ud�_��>�O���q�?�M��X��T��[�}��Q�#�������J�9Eo_Wk�٪A5���]E)�g��aS�#RY6=&��ġ�N�HE܀i(r���3ت�b���B�O aX~�^�߼���0�W�M�*���&��l2`��(�|�_.8;-$	���G��o�^��
�.w���9�h�c���������$��ĸ;��E �%e���"I��[Z'�te�@���|����Z�&�`S]���
��!�I���߀���b���/)��m�>����ȓ��o�g�z@�^��?���,X�N��; x���4�o���J��-z��;�a1�5�j���"p���#'.�0�θ��;1�����$rH�\����ל��Ep\3�^�T"&w*84z�	���VY.L��%��4�*�E8�9����*�8%Д�̕�`������M	�PHО�e�������|ϖSw��Ԅ�<�7Md;�;�ƞƚȰe�Nt��$�{\��nC���煺ԑP�B���z���Qw4;貀Z��<��u�ݴ���W�o�|�6����8����b9��>@y�1���0Q������	U���4I��)>r�P�#��J3\�QuDֵ��R/��	�:0T\E�l�zk��M�=����51�粁��
���P��I2s}q�,6��pц��K0A�S�R�z���c	���Ҹj�CqK�0�P� �r�!8���m���(3�V�j�^���dN��Uiߟĵe���K�?�FT
Պs�K,D��1�at.�R��[�����G��%����#ܠ�]Bv_@�&�BO����"����f��$��_���k�t[�ú2����EBڜ�N��Iۉ��������[#�牄ꌬE��W9��:g�����~��[m�X��
��{�k��G��Z� {g&�D���,����&x���]y��|��c����W�y�ǠŞ#XC
���"�?|2�tk�:9�l�ͷQ:������=���_meDT��t�0��Z�������wSVu�r����$;�9��H���D7�m�"4�l`�W�LpT�L�:�\lW�~4I�:��:�L���G�D�k��{�<��T�����N=1�E.�МI�k����M� �K&�LL�x�����^L�Ĭ��}����H����ڄ]� Y>�+v��B�56���f�gЊ8��`���y �t}���v�,{V�,Ȝ�ɚA�,��֤��N&�݃D/(3iv�ԝk$�����~���Z��|�:	�8�����GP�V������t���ԍy���P��z��>S�}ME!7�l4��W�r���|��?���[�xh��+����,��b2k�0SL��]�SF�]�?G>�R��_�/�^����0!�t�����,��1W�6Z���oh
�7?���ﲊ�Su#X݁��~_��ˊ��]�I~��M�'�r��2�&�U1��<�0�����3Ȓ΢Y_w�{ܹ���q:�ok� [��T�����R�!�j�eқi��cՎ��d��]��rq�����42�9�y�~׵n�2Ⱦ�u6�^�{}��9-w� H-��$�n�~��KÒ��8	��I�YK$�U��s�\�ױ�.snØ|�d�F&��ے��S�k-�O9���H�"�a��({���$�]�@C��lM�:��	|Uɠ�����;B}s����;�y��yB$�h8�~ߐ�΂U�>ƑC���E�3%�z����"��2�jK(�T#	n~�)�Z���#f�0���q�]��Wt�:+tA+KxܑV��ߟn��^��;�I�I0�'�������0���>�zj5?��&&6UE�mҧ�����]P ��̿���[����-7�ꜩ�49O�'����E���+���N�j�U�%��4IV1�@����E��-�ȷ	�c|\������7��\@%K=��Uмǣ�j��T�!���dyR9��0E�u��#L��/�7�
��=Hf�9g{o���e�����F_���$NR4���Ŝq)�s�H >�U[/�U��T�^��A<ŵL�ȶ�u
���g���[�.s����G6�ªI�1
U��䎪���� ��~��H�(g���7t��4���o�VG���%�L�Z����� d���ǋ�x('bu�T��>�^C���<<�ݴ.l�wk�f�ã�0e�߳����a@��K�W6��щ�G�c��)	�I������)�hz�#x>��i�1�9����?%&PoEz��$]�Y"T��w����	��eۭ��ڵ�
Rn����s���K㱝;6�Vsb�%�W�����-��Ue�8R>73E2�e�_*_�o�^^�Y�AR"�6	+3CXf�o��L'e�C�P�@R�@?y1�>�ò����ЮH�l����ǌ������O{����8�cF5��x�����D�y8��5�SN�? ��O��嬌�?��Ѭ��TNq��p��"w#�agO�EFW�%�$	V|��֘['�^Z�U��=i��?�L+?����_��'�`
%�� ��_���S��x%���[�V,{�RZ@��+bW�=�A��>V4E#�Aڎ�9�^�/JHS֗�)�_�\�߳hR����71� �|�oH�Y�NMǷ2��/קi?f�^8�i��N۩<(��x5�Uc��4�)���K͚E�r�)�y-1t�2Hs�;>��O�1���6������'��^� W5��]خ�4����$�<ឧ��{�ɟ����w��[�۾ ��]}����S���Bc_@ �c����m����Aϭ�)�}�z�"�/���5?�M#����v�{����p��څ_�?Z>9�#T���p��֟�F<�U�c2�5U4�0�j�mxz)�T�<}!ʽ;���1қ��$��t �	0Z�XC���xT������#�L�Ӣ�8\�[��"�UsL�{y[\������1gj|����,�h��M���hG�x�2=���N�󁯅fI��¥M��҈��v�O���A<�A�p��Q��3g��{�����ȧ�oPr��)�ˮ9j5fЪ�iZ��л��D~�ħ�f{3���P��U���9B�8���	�%�Te�<�M; ������:+!�����?G0�"�3�n  Nh])񹭤O������X�q���G_4sO�6�1^��D�,O�(�G��k,�\$l��%#��H��hh:�]��)|ñ����Cy]�����ʒ�,K��*%��������a�nk��l����]s�rQ�v��.�F�;��mSuR-����oa���*_��gڹS����B&�����,<(;�����`������h��\���R�GnJ:M��I�4
i�1F8w9�*���.û�F��N�Y�ˆ�i��=�C�	M�*��է�N��;�~��1�`���	�t 3��%��-4Es�~1Ӯ���X �5e�pUI]��y|�*O�+�~m%LU�z�n��a,J����RC�O�l���\s������|���׫�S��~!�lAb�!XQ+]�}`��v^h�	G�m��[ ���FM]���[5	�FW������ΩE����5�k�}�Qu��Et3�ى�AmAi
@H��Jh!P��� �}�U��J����90����g�"up��|��iC�ÏH��x���ʤn��M'Q?�@u���'t�>S���!��g;�.n�J�K��o_`���@g�����/2�2�2�vǲ��B���p�|�̛�96P��ת�ڑ�U��G)/2�w�OI�/Ю�[J84���8WͷK=f�]e����k&"�k�uo�#}o����Օ����ȅ��i��ۮ����!���>v��YhV�GI��U��^ K�5�YV6N$aE�KYxC��_�11R�f9�0�aO?x�N����M��22��&��7�xO�S�#�����9}ɸ���H�� ;Ά�85�0!�,Ơ	���^\5�K����4����Km8`��^��H����<��e�nK�
�֏���?B[�qdw�P�H4<A�������\� ��VD�N\��i�>��5��va�I�&�#���Rp��Y�&8=%��Au񰳕7Җ�럗�VJ��-�S�Z���cJ��5\��K��d	�2[�*0K�vU��MTҚ	J8ܗ�q8(RG&�wO}'��b��/f|�zs%ҷ�ϗ*c0���0��"~y퉡Pj�6瑠�Ge�/*�_\M��V��)����x���ƱB�.Ā�ȝG�F��l9�y�p�^Y��дSS�v����٩F.|E��H�S��P�����\NA���,��DAIN��U���� ����(��T��c	�|<X.��������F�p@?Z�i��j�0�lE���ԉ©W�ս�f�^	�c�~a1Aip��;�"�'c��
t���>��V��[6^���Q�\+�3�L�N�¹���2��s�W�2bL�;k�JG5/�E�&��eE����hB+oW��r�G��Z:���������{=Ci�^fÿBn�a-`��Ff���śj�6��V������>����f�X�����?��yd���� ;"���Ս00�\깘܄�)��|���ij���J���y?���ୃ�s���c���l˽䂤3%V�IK �ҥ���@�BзϽ��?�9�[�4��3{-�8`2C���-hj�r�x��>�30�����2Y���|k���3�τv1�㲧X ���HZO��+�� �&9~����3��>�n�M1%F�ʡmNv>��͖.{�1)������f�rL�֫��|����<$e�C G�Nn?�dhd6�X��r�%�k��oOf�C�[5Jr���J�oGa"��q��q҄���8��k���Ě����/8e;�i?�{
SO g���`��tR�i�A�G���oT���Q����eH���<Mm����0��O7������:�+�1�����wx�^6���D]���3F�$rF�^��݋����/S8p�S�˪T��ϿZ�ҽg*�}h5A�#S�+A�L*��{, = ��6�"'��C�D�zMG�u��tΝWy���g���\�'a&E��9W��Ͱ{`n;��Qt�̌ۈA��Lh�O8k��t\�[T��S�^~)(�Tw�g@}��*��O��i���P�BY�}D����&�'���+!X��=�ѷ(0a��xtL��;���������Z�;,*y�b���M���=�Z��d��ߏ����eK�!���5M�$Y��a^R������ F5�FD�6M	;|�G�]�*��n�[�?'��K�Ѩ��!Q>�A�M ��;�v�e������D�Ʉ�om�Ģ�흘�/�h�RL2�'kQw��=\�+fpB�D=0D(93�Gqp"w���1^r��M�"�NS��=1b���SN����֦b���~���$ћ�"�~��עY��
��C��Q!� ��z��>	����*9�I�|�����^?[��4c;���#�5���]�n�J4#H��$\4���:`s�v����^���wg�~B!�@���z����]�v��������d�:�y^,鋭���*�*���Ѵ��8��`zn�6"�CC�+��(��?��i������# ��[<f7���H����3�E@K?yT����1�Ӊ��^�͏2Pì�Л2���.��ccYB��Q[��7��m�q�D�eKJ%\�!���n{�ƗuQ9m�=���xk�hr�Q j=P���!O{� F�T�}7B pUR4�	����#�ɸ�S�9��&od>
��8XRE~��I&t���ʮ�К�eY�Sjz)�;`��*a���jݑ�Ý�f��������dȼ/���j�H3^7$���Gb��)I���kIΧ��ا)�k�gˑ<"k?�O�^�2\���Ry��g�DMy3 6�0R�&o��9��z�o�i�gtM#վ��KEڏ6(]�?�UL�4�yrz��vl(�;�"?{�3&:����f�e��H��Ʈ|0���!4/� ��
�
􉼝�cYv�ɔ9�4��0�\��RP.�[����%RB&̽�a�,�a_>�cWlQ��M�lY]��P
;mT��,F��̧���R'9�(Ŀ����7�n�B�y[R�mf���������,G�_��Pt�Ք�>N�W��l����P�������,Rr��ۦ�z�;%��j=�Q�z⁗U���S�-��j`�k懢����);�ż�_��3�#�)cq�]��sg4n�DNG�����-,�ΰ��T�XroК�X�Se/ii�"`-� �`��H�J���?Y��$n;*h9�5�h����J�6Q�(��X���e�8��N��WM�* t{"�����N�����Zjy�o؛�8�}PNp�BJK^UA3
�ٿ�1lF�7�KLR&�Uܲ��N��*��	�j0�pϯ����0J	��+�j��;o��zt��g�x���Y[��Q���G�L;���b�6O���FY���xK�Љ���u�8,l�Ƭ��6y<�C�Iq5\`��鼙�m��(��I�+��,���)�V0,aQ1b~. *}C�����I&�Ӽ4��k7��!~g	���_���,a�zW?+�*׌�]��۩��F�l�\�{���*�bT�T�k�ҹ}�TM�GFi�B�*��X:�w�����!�;�B2�H�ţ%�����X83�Y����?V跟���E��e����3�Gr���z4��ՑB�s�Yu�t�v��~���ź�!�2�:��R��!�m.�~FU�q"�7��s��Vtk&��\[]Gy&�5qX(m�.���v^��������w�)��X��D���A��AE�E�����6ZG/eC���ˑ�9����?L �$�d��[�xA�qӖΜu�l� �^��J�>�%���I���1���P��+[���?B���q�
��?�施�M����#��k7�|q�n�B��\Cq�������L!k�_]x�*�0� ��<\2L���V��;��?��tr'F��l����\�0]����}=d�w�
ɔ[��{����j�2k�a�(�tlV�@���W�w�����b�1������r�u����jX��4���y��e�d���
��V;�QB�Q�j��T��$v��;H\�C�\6�~��7��;�g��g��+T!+n�x�Q�K��d�,�*���HG	1E,�ԫb�}�����-�+I�3���b<��~ ��:W��-p����&Ε�%!׆���/������*҈��$����RyV2���,G$�ղw��h�؇o3��i+�NH6!��r��C	eD�e?B��fo�O��p��h�z����n��k�?w.b�c���8������4�ύ��k��ʻl���
�e$W��1���3\��C�OLG���\7;��egyG��$΅��5Է��yvwp��i�&�M	t�E��ہ�m�vL��t9����Oa	YC��)�J#�Z�!��GG�Q��4(�������!� � zzg�h*>�x�<�.y!z�ܒ�C^'�˴>|�M�r|h�n���j�Yއ�ڶ�E��ۯOs��07���S-о��h� E6!o��m����y��u�9�������$G]�h�Q�>�G;�L�5k �]�غ���R���2��N-��y{W�e3^�$C�4����Օ�0s�@A����I�	3.\��1(�]Nv�.N��6mw%�w�KP����3v���!��q��0V�����a���� �~�j�K����+��f�J�e Y���"g�BN8�>?a�E��2]NE�iH�I�&
��3a���z�-Lm@���:�ˣ��4"S����{:��%�V��˜�V�/縳@��)vֽM�_��>5�p����)P� ]ҡ�ME��G>�ɐ��0������_��� �Z1� Fizq�����_�,�^kP��]s�ju�gŲ.�DL�?K�x�.~��� Rh�@�����H�T�� ���(�*�����ܓ�m��������y֯�<F�5�����D T�\�M*�Ef�ׁ���B�1ΐ���o���~Є8m��.���k����K2߂��Ep�n'�*�|T��|�v��i�{/5B&�C���8��Ĵ��Uk�	*U]���1	k|�8�#��J*u�0�����Xr)�Io���e~�Bq,ߍI�.��`�8$�0B+()��'�M�k�<ޤ��ſ><�/4�}�V?��7�N�qYY�%� j�b} ��1���F���*AT��ZV���8Z��6"�=��J�,�T����k��=Mp9�j�4Aq��|��	�4Ө1 (��F?#��L���CY�(kU��]�S}��E�K�t���j��6n��/t��W�ј��V55����QF���dm�@����
f<<�Lh	�g�F'cܳ
c��`3qX���+�����a`*�''�8N4ٻ?�{���jf������j����\����r���[.tuQ %��)�?çCSp�����G���վ��!�����@�)VO	d�1�7E'�@0��f%�������^9� 2<�\�秓�P�{W/��v8f�A�����N�e��?4���`K���!<�v)P�`&�ÁQ9����?wH���������9f�_�U�: �Ua>�>���&�Q����U��!2x	�U��p�RH��gy+��s؜��8j���:saQ!\Kg��c=H	k&��ٶ��a9���RF��Po�	@FaX�մ��D�� gh��~��@�
�u���}D��B�h��6C�l;���v@�vi����M]���dNkO��fW� ^2�9���Em؉���,�|��)�'v��HnG>Ш-��������uF���y��@m�j׮�����t�<H�) �̬7
�e�2�
�~���V��~#>��Y����,�� csXc78�ș�uɳn��2aY�������M��09,,JA���0Wj��_y��3�v��eV��ij&� ��\�&i��	z�1~����l]��M��I����٪OS�U�G@S�*�i��~�a
~v��4���>�w��&Q8�A-�*���пl��/9�=�X����g�zc��R
8�3Ԅ�B	s�3�CR)���g����]�}��p�ƢvM���E��.�߹��b�&�%/���w�5����i�A_�{��&��VNk2��~-����*�J��r���ᯏ��F�!Ƕ#���!�����{cw�ktiC�U�|�'���^����;VI�ˀ�avw�>�4�c`T7:s�P�CF�u�ӝH��	f���?�͚+K��p�E^���֣���i���|��L���)��8�;����	7Ry���"���!oa�B��^/!��˩Y���ϳ�]�2֋vs1:S��3���s���Q��t�܃�*�������&�ˌ����
���`�
N���w�U54�"r.��2��v�2�ԣ/i�"\+�p�H9ZJF�,<^��XF���]/ �X��1���I��唬);���%/���z��潒ծѹ��e����/yM=u~٦�$�#y��˹;z++���x��D|B{�)��`3�f����z	�hg1U:���q��ܼ%o	��z>�f��'��N&���kj�q2�}�t�2Q������7}��9gӾh�b�!�zo/���c3R�L�m�fǝQ��\N0�nG.�T���g�p�����"�y�����;\R`���d��,�&gq�0�r0#����!2��f��K /�8�k�F���w����V�Y����������%B�cT��Gn���i�&�	dN�o��M`S��8�hkD2�ui�P�������bӺ�N���;hU����c�Ç�^��}��?p03/4㵕�? ��(0�|zں��{�ID��fl�����F�o~n�E��q�t�.�U�����{pK6��,�Ɣ�i�N�����l����3��u�փgqL(r�]�g�#`q�Du�S�<�Ԍ���N��6�?��
!�Ka���F�"��T��{��>:����O�W"~��]��34W�HW���]/��!p#��anu r�k+��u�o��?1%�f~��������KU]~jH �6�E
e���|"�X�w�'\���}�QBt��#�Wo�E�$�С|e�s�F�fd��..��/����L@��+N$	�X*�����1�o�G��x���t*��1������G��i��`�a��(2i?M�_�o�[Pe?{fi6�{һ��s�'>,W;�'N/�e��+h�gg���_R�O
Q�?i�V}W�ދ���,g^���E�u����qːdC@Sk�h7)�����'@N3����é?�o�o�{����Hc��z�A��m�=pS�#[V��e`�?[*?h,�:M��f��n�g��KuW�jj-�s�ud��iT
�Y�$�t8=r���W�uM��6WOТo-��)����j*t{��ڈ+��Ι��&MBGZ �@;b��2�U�� ��1O`��$�u��Ž����s�oO�cA�.�j��K�}6�T�O8q�:�e^��'H7%�G����~6�	eC/�6(��g���$��`��ɈB]l��@��Κ)2Q���|�!!���0���֣.��T@�"q�/�ܩB�s�
�xJ��d�_$�R7_�|��DO��g�/}�-8'��s�h}9�mP�/��6��@���-,@�ecAw����B��U��#In�kտv��H�޲�a۹p.8	ũ��p�E��Y��e��!�Б�b�Q6��������@ڃk�G�Sr/0
����_(c�smІ����qI�y�}{'����&�,��ؗ������8�0�;y3�_l�9��t�~���e���
�c��&jwS�DZq[Y`����F/j�� E�������@�����!�3n�WW�͵,����ڭb��ycX+Y�-�:�=��qc3��ДG���2;�p:����H�zH �P�6B�� �lu�v��Em�	 ����[���m�Tr�boE.���_�[/�*Ֆ��\�Ve�������y�5�"S��]�=��KnM�����|i�um֦��'�C�ads�S3�Ok&�~���8��%��w9Ɩ} ��Z��=������`��֑%���`3���Z'+�����p����n�Ȭ��Z��f��e�z���u+��^��`��� H�� #C�`o��D�Z�W>��^�]�ʴ�������@��B|���>]��`���f��ۈ���R���?i;&ߑ�� � �7�S��yyOP�j8�p�qָF�V~�UMF+�5�|h+H�$=k��<�t���^�Qq�-P���J�"ۆ�Z4Ds~S��<>)�}���kEbEVdxl���Q�~-%��"�t�%	[�Ɓ[b�6n��`�h���U�^a�jr�@��5Eo�q�����&���S�u���E\h����t����ۇ��]���M\��?�
F�i���Q����>�1���+۞	E�r6��5C��Gߒ�./�����'ɐҵ����ɛK?tp{�q��2���L��3
>��y�A遑�b��b%Y��~09��-��Jp�z1�����o�����3����8	�I)�R�W��ϵ_�Ou�iO���(�y����^u�&P"������M
��Uc�)Y�O8�\(���lY�`�2�)Ѹ_~�<���5!,O���:�@O2�6(a�3>a�R�V܃qv����p��Ί0�D�\7yG�U?͋�z�/d��Z�WR�I�W֍�i��8��g��ؤ�W:t'�y\C89v��j�?�e��2{�D������;�(1�	�Fa�^�7Z2&�g��֝��F���#�H�p���Bn�����f@g��hR��R�B���ϳ�u���E�Z+�t7��,p+��-��H�����H�_�i�)[v�RZK����N\���f�yV`�j�<Wno�a_���/��
\�����E�{��:��4�����S7f���z1�<䊄\�N�j��^��t�;��rȦ�����b�g����V��c����{F4Q��̄��^'F+_�l�$� LR(������i L�[IE�:�@��^��:��5�&ן��\%�qc��������Rm�W�\����6�e���,����s���~5_, ٖ����%�ղ��K�.���F!��b��$�ċ�"��a�����Z�Vb��;B�U�Ɯ�4�?��Ӊc�4��=PȁT�� ��8����=�o!�j���Zj6�^^t�p4�(�y��[Y#�5v�EC�M���҄%[���\������B� ?�~鬝D���9�uኬe._2H\j|���6;��m^�W��t������Q�?y�q@����Ėt��{e��j됞xg�өs�Uſ�Ϥ�C�y����keǈKU��8��7���ٯ�p�?��}�Ȟ�5jU�1]�<��p�+����"�q~��hR� F�����*p�k��M��K�[�̊�^�U�熍��b����;m�A�O�JCY��!}�$�-���7�Yh��6YQ��g�ؑ���^��aA���îarJge ���]]|0S=T'z~�b�YQH�� p:\���U���I�ʗ�[�?p�����튑U��bazj0��f�q���\1��"T ����<?���ݠUK��,����vp{.�.�5�֗��� ��d<�u<yy�?-�C��r����P��HS�RbJAO����|��:�^t~C5j���xUp��71�թyǨM�[B��^������Q��'��c�D�woD�"q'>�C,2$b�T�_��r����c�ع��9��Mi�sD���!5KY0�~����C:A �t�>g<{Qz�v� �(~�s�y�j�$fׅ0�pY��(nD��547�R���q��)��k�
� �L
;>i�vS/œ� ţbUg�a�r.[b���
C/���R��N��&.�צ��<0{͎(
�1�u޲iR�1����-�,i���FG��0 ?-��Z�0=�����_4]�z!���K�֪2�(B(�휭���U[� ���=T�r}3��<�0�&n��F��7�2�ப,�'���p�^NŞ�-,�HϨ�ŏK�%@��є����Rn�斡�y61"k�k �G�������� v�f������
(Q��j6�3�Ś�.DrB3$���L�x��iT����c���O��$���wx���ݒ�}ݏ�?]�V%�D^�4+�G`+lO��+I? s�0�.��Ɍ.�
tA�gs,���x��#���3P�Ζ����.�y���Rw���Q�Ț����m���}u��T]O��{D�zg ���W��͔9ߐS{pqsNI�eI!��E��)\�=���ݸ�i�WO� ܥ�<�0Ըc*j4��NE���2K6� 5�Jp���h)T�z"=x�z@Z�����۴B>�m�J��';�\5����%���0 �0�ךּϰ�᠉pI72P`7��?����_6I��K���-j
���T  �s�wk*���Z]�2��_ͽ�yGA��w�G��;| ��ܪ��T|�{H�+~�`����5fO�8b{���BXU� Fkt�<�a��#Vg��gu;�Z���fx#��R���6����Ovy��(��;&���vvOt`�hY5����ǼC����G����u'����x��p���W�x3N��KXBp�+�aM�@7�U1^j]���U�R/�� ����z��=9�~�%��~b�Q�bG8F5���k��h�<FZ�qa[U��T�)v�r��	R�����P�Q���Gk=q��'�A��Z�eBD�i��Osf�"�V����cN��.�=V���Ѹ���*� T0�6Pn��U$>��J�G��ڰ��L�3塙KW �I�m���&I��|��F� ��U�S��<��)k��m�MqnH怴 �N��y,3���4�teye���Xl�=�j���B��D�X���J�W���;�^=��Ă�x�d�<w��d@v�p�m�\�В�R�p�����]���Rm�����M�*`h"�"�"��|����͟W�%���H�����ԙ4���� �Z�A�<EI�T7�73P�Bu��Q��+��q�/}'o2]����3����a���39z4����g�6�ݣSn	������WA
�b�z�1��<�eD��jS5 ��!�/^�tl5 �r��ϴo7�T� ��߀@N��4xS���s�Ѭ��Z?�6}��PJ�K4<`�PK	�$�B���iڹ�8����q�U{�fo[L�����7��B��7t��u�d�+�U�A=�C@��,f Ժ�}�
�I{�i����-���ԗ��3���/r�zd=hbI���x9�8�"�6�W:D,�^o�{_0��џ뷂�%�����nx��wyDm��P��3>d@Q9��G�u$h���r��	I����@*"���O����o�W~0rTN9��v0���B^�؃d8M�q|ki׺=��\�HP7�Ej@�䁿��T��R�º�o� ���!`º��$j��8�4�jld�ߟ=,�¤5AUgn!ՅӾR���=c	-T����'$��R�G����Ⱦ�:�#��_���m9J3���ύ��Ũ���'���H��*�i��Y�:��W�.T2k��i���K��T�hЉ�:���GGl}���E֝w���-M=�z��-����>����/G�������)%�b�a����'?��x�4�鼥�B�)�ɤ��O�/'{[�Z&���og�\��2�6�b���g���6t���|/ȟy�&4I�'5�B��W����*�����/#g00�6�4N�-�4ޮUh\BΎCT�LP��
�#>��P!v�@��A�b����w���i����š��N�����j�l�0�?�Ú���r�� f����!�{�B4�Is�p�0��GS�{c��.;q�<�&�
6��|W�+>����R�����v��Ws|�G%aIPJJ��BaQ(���H{�m��K*v<�q�B�ʻr���;���GOڛY�,�ك�'�FO����Y���k?݃���aQH�$]�x��u(���3m%U��`��������)�÷�TUl��QI�ҟ+��Y��U��D����y��kz�7�"��>�J���$E�ƹ����몽����뻮D�	�5�օ�����y�1yt��%8�3��v�D���������.䗠R�F�.�kT���LM�|eevD���*s��v3?!\���]��$���3` �Q�j�zĬ�>u�>���c��u�5r�;��N`����9���kc*?�R�����4!��En�nI_(���z����{���s�����6�����>B���$Q1?��
�P]�sS)��>���8��x4h�V��ؽ]i`R�u���ƿϜ��3�,'H%���D���Y���H��cB0_�W��Җ͗�-����S�J�Bա �\�.�/�����YË�}2�����aa�j<tڌ�'�U�_2��(��"5��jc�;}�*-Ҟf%���x��,Za�D�0��Nl	���uY3�"'��T��r6�#i�HT�����(��?e'�kR�Yo�^1tA*�+!_�7 ��`ͧ]b5�Z��pe}3
�QqfF���b�uN��*o��KK��8$��O(K��Ţ�^4U �wqe�/�Na��Y��p�m
�GL?��J����\ ��ĭ(p����U0��*�J�҆���*�b���µ�	��hԙ�D�H�X���~t��벞qP�w�(\����qpk7�u�KV�ި4�-�Ÿ��A0��I=]� nG�7�j��O����Rk/�7^&s���4��V���_�k�S՚]r3�)��9�$���$؆'����I�U�;P�}m�7<�9�2�-Հ�spk� tH���6_[%4�&'k8�\[e��<�i�R�LO:��̦i��dY[� ��mz��6vl�K�8��$��h��u�%��H|U�VI��$~���]�b�a�?f� L��X����u;�"߸%Sb"j���b�>����Np|��S�X�L�{�}��*D�_�H�����̆��8�����i���A���8��Bz��R'��^�AA!Ta��E҇ ��In�
2�!�V���0�OX~�:~g�9jA�,S����)?������&~�Z��%wnҌ-9Jb?��S�G9��Aۭ��Y�7� P��TX9�~�¦'O�E�1��yQ�� N�*���'~<���=�������N��	)��Y!��#ϧ�ͳ�;����I��yR��[*�����\�bE�u�OPS{�Gq�'�<bW�p?x,C0�ԭ��N�䄺O�$J��U����sd#�'�\�G��Z���F�0�h^feE�B�M�U�od��� .��z�Av~��F|P��H47,#,��'[k<ԬV���޿7�oH8��,c����%ɷ_�F�=�,�������K1�����ĕ"qhiΪ$W:�o�=�2BK�k���������O���3��F|y:��q��`h�JD�~��g6��rzTj�[z`bCw9цpdf��J�Ͷ�頀�Ƞ�uu޴�H8,~	U�=�Hs�s�W:�`𷶴�p���s���M�h�-`����|���)�Dƅ�j/�D�N����n��?��_���>�����M��ڗ���.hq��`&^��(�o�@��m����m4����D�9�����x��B����:��^X	�_̧NZ�Q�Y*y�r-Ī7�o��_�Zu������@Z�r�&m/.kO�s�y�7��Ŷ������'R�,��7b����!wȌ-�|5w��HkW(C22��'�X7K��1�@����C��YM禄i��d8���-,!�B��8����ͱ>�:�;���P�4��A,c^�#�X�	�V�+�P�ӽ��,n}T�(}Ɉ�G-��P����4�ղ��o]�L�p�o&'C
�{"��$���;���'	V ��6x��XTz�e%���d����0�;�}V�eMΟR���Q��&�0+fm�qd�����fj2���i��pz�w�A�0�ð�Pd8�]W�B����ܟ�ǲ�Ibd�7}��-�@>��ƹ֤��W,�"��@X���D:&t$&q����VyW@l;è�nw)�k�b�8hz����Nm,�#x쎛�'�ڨ^w�7�E(��ޚ��޾���R�G^�45v��45�ۑ;��.�m�IA-=U����P�5k�uKyP��"��%Z�N�U�U<�-<b7W���i���C�q<�Ļ�j��ұ;��u�.�@����N<�?k���>x��o�ri� ?͉���K�>@2;j�P:��n���m]3!G�B�e7o3�9P'�{���w���������xQ�6Hi��ɟe8��1|�#�z��1薁`6w۟n�jڦ�Y�+�z���o�0��y�A�<��	G���7z�>ކG&�+K���~_F�p�E��%����||���7j�f�$Q���c��zo�2W��>/"(D?g�Ѷ��5#��)Ҁ��a.q�H˸c�G�ImWs�DU��O0�bX�^��	���@�"��[�?H��I��Wo�K�Q�8fj�ܽ�����tuh/72�%���%�����r,�;#�+0���������*�[��4I:��1��w}$1�7R�����B��,�X�X��[�qaM(����tk�8��hQdQ��%��+F�e��\�H�{H�ׅ&ģ��M)�oG��_�H��Pu:u�`�q���
Ԅ�
w�� �78�����&ہg̃��?f]l���4b�~Ơq:ަ��e���P&7������'�]O�M�{��`69p6Jf��$Ti��y�R���u���t)��
f�	Zhb���l0�"��Lxb�՘��|�׺���1mq�X����!�05�s�נÏ��!����Z��]�[Ѹ�-?�����s��<��V�F7ܨn��������*q�%�;��ͅ��r��|���Z ������̥O\l�z��Ⱗ\if�lW�Q ��4��B�����[$�@_,S�Q��J�ǥ'��Y#��A���@-i��$��X���ʣAr��
���?����O���S2�� ]z��Hp�'�M%�q������<E�� ,`x���&��y>��G��(?\lФ�2,ߊ�WJUz��1c!e���(�I+E_Kh�K7�Y+�k960���].�f��#��A�}(n�B*[�屄��7@.������(Ş;�4{�N�I��3+����B�_t��p�#�HF���>�[���U�r��P��9�6gPͦ�<��Y_v������L���Y4����<��F>پ��Zɯ��J��X�'_���2��Q����<%Y�z[�bo���z���V��j_Y��� ��0��,�dV�����;�S����}tSҜ�S���o�&��OX�G����U��� u^A��y���_�#!ɜ���X�Fw�n��XWҸ=C%�x����!	=�#���\�'��՘,��@s��v���ڶ:_��q3�E�V���V���=���Fg��\���<��F1¸�c�jpP�b;ܬ�T�-
HWЅE�w��F�� �֘v���J�n0ӁM=��6�$ͮ��a�g�H��"��e:f��R ���V�D��T���v��4��
O#���
�BM��&�����l�Dd�L��X�TZA~&�� 1�Ȁ�p`���?Z֙��ڡ2nDF�sr�N$���O����CF���d殷3��?)���u� �r/r�d���w@�mH	m����U�L�&�yRC��($�)@�b%mO$*a�1�y�1�*ốˑ��M5���k	y-5��.ؼƔ�Z+s�ۋ@ 7����I�7���n����}�~�˱��d]�٩�#0�/��8�,З���� A�W�+�u�k�&y����{����'\B�		����N���f�/��{���!���AoN�������1�x6O���ȇG�a��`��}_�?�5d!>�9<�r*�8;�� �}�D*�0�}��xU��Ye���Yz�"��턺[��6����$��U�>)���d�x��I����&�Tx�������R�Yz� r�u�:�����&.�Ya�� Q��*l<B�4����x�H�����E:7z�q������]k�
�{���S��!vrnǨ��3^�c%k�t��p|hj�����*�_��z�ߴ�0A ~/��_}!e�?�?3�
��`��mȝ[������3��^z��4�ޅ]�g��Y��i1�c�)n��&����"���"��B_(��|�CG�������������s�FE���w����VId�����m�b!�����'�����/�G��jz���B��m�N�8kX%r����W�\@�Å�n�#�ӈ�x[���GQʿ�7�����
���n��%F��?�{dȢ�����loS�M�D���S�m󫹭�'�1y�>�^sV�\��e����5�$%C�M��l����j�H�ɶ��$��)a����Eff�2� '=	�n��\��Ȕ��R#-�wb����<����A�gB�`��G`���G�#�9&�Y�[�=܏4���.��k���z�̻�Gk��p��<r�g��v_����`��w�K ���3A�@�B��L��|��
v�i
Q�(`���AO]�|�j�jl�ClNx]��#��9f����N �@A.h�[�NJ�	�f؂��PAfC�Ѣڝ��H(��"��\F���њD��}(��Ή�:�L�`-ZւC�|��O��O@p��V���d�\������!M�n&��p�D�51��� ���N��Pc��ٰG�j�Lf6P�I���E�d���_g��C���"�v���>�\�4 �jw���ʸ���'cn�<CLП�r���D\�D�p�O���#.���A :�OEx|�*XP~ƳV���C��/���5��g�{��LV���5KX�(,��, �!A6Mϡz����n(W.����溺�nG�����;�=��	�������H݌1	X�#�uR�u ﻯ��b���(9���]U�{K����c� �j�L�;p�9D�����g���3�7ø������q�����GO����4!����:��w���n�?b�y�R��e4�|�wOgq��G>��R�7�������p*❜-e9� ˫�4
��g���òj/v&y�P?Dπ�Oa�0��U����! p�+	��1�Ĺ!4&_�8��&��~^��֣����9�(��e��՘Q�nia�eӸ���6�H�?�f��r�;��OAu�Ī����:�Yt7�W륲�����a�k�[_�n�u�^b�	D���u��!9�P����	��̇���8!�i��G�o0�nQ�����h~���s�h4]�Ѡ2��4��V|�:��U��#���b��m�Q�9Δj�A;��Yi��*��Hw�x��*d�W�Ѽ^?jю�0P�s��y!�Z&^
+"Bu�I��ޛ��I��k?����VP�o�"{v��!�z��B�5N)�4�Bt��4�.�(�o��T������3��F���.�q�CL����j�.��#6�9Շ޾���YM���������je5h��\���`�SaW�M���t=��G��\��b���3H2�DoD"�?�@qL9��6�EN��E��RyfM.vv�v��gH'�I ��9�5u�	����P2Z�0�5�|	S}���%���L����f�[�k$]"0o�_�����%�X��;\�З�!2g"���tA#yY�움�ק�o�R�0Y�I�9��fw�b�a�6�Hxe�H��\���Lk[r��J*C���/�4�uZff�6��KVS�0��;�Jg��5�s��ɠ��2د�`�˕�Á)3~�ŉj�}��O,���"�ֿ���u��\"6�����>8!+yTŲ|��2I�ԭ�8�!,�ω6Ntw�߳ƄF�c)��y�`�k ػa\�ߺ�*1� ��H�T�Y�1�o�����H�%���<���_�$@N�Bv2%��BY_#�����/����7�	x�u��v�W�%��ԓ�Y�ڧ00�Z*��,��@��>���7�"�w���L��Q�R�H(�^�Ϫ�p1��:��Y������lq$�{9��tr݁����j��Z�vCǪQ�I��AHh��Q�'��C���o�,�`�Xc��(rl�m��/0~�2=��|^�ޣ͵hx�Q�"�
�)�B1!v����a�<����,jV�W�s��EE�T�ғ����]X�ܑ���;P���r�C�Zf��	��A�ɚ���d���XĻ�Vd��3Q�G ��W����
=���z֪	n�ŌF�J�3���MX����"���E��e�����6�Bb	G��a�l��jzRN����L��T��.�5���;ٿЪ���m3�i����w����KZ���j��s3�� ^������A����Zm�ߥ��BtKŒ y�KR8�����%"�� V�~z�5��c�/�(7�m��dI<�ݏ��J�@v����q�gC�]�\��P������xL����������� �a��dP�&����Ül��ˍ�b�n� �r�����jy�c��;B)n	Q�$��^:ȲF��ů_�Fp]@7�߀�X�(�lsAC�K'E�q��\�or�=�a<��-�ߐz�-�A���S/��cQ�Hg��A�@P
���J���k7	� �I��>0�CE������'�r�'��\jtbF�`10>k��y%���&�	i�1����!�z7�3x�8�h8�$�
ml�EI5��'�t����O�������s�������'.D%kSj��3E����n���e&ur�Y�gX�Bī.�D�r�~��V�¿/����]�o�윥�{:o��`>zy���Pom�Da�⊎$V�.އDR ��ݥ$rK�D�nĞ�Ж�dT�9稖ܧ�rޥ&z��aޜ8_4�/,y.��W�?�p�-6��8��Y�q� ��<r	X�W�{c�6�)�͛���L]���C0+[!�Fb_�o!R���=�*���|����@��0����)�ݞu�+�"ܨ�0��
��N�[K̀��`��,Y�+�׎������ۖI[�-l�Pz�C���jQ�r�����23W�r�a��qk)�S]�-vĹC�.��D�g�^���U��
 ���Zi���r�q��3����m��;d�w�	$��yp#�L� �.m�=	��&^Ж��4�Je���5gNS�g��g���d:LA��k[��7Ǔ1&�Ơ���:���[j���E��i���YBW3<c�Gͳv7 o����;5�<ys]�
j<��*��z��8�zV$pq �-����0b��;�:o�QY`�ڐ�
�ɽc8�"�U`F^":3QM��:$3Ʊ��5& �\�ۛ�|j�h���#��Cb+��U���w�!&)�W��[�Ʒ�VBF7,��}��q(����	TJ'���]�;Ʀ��r���h	�tB�m���ݣr�~�~\��b���Eo��uq���<A�?>4�ڙg$^A𪫿��n �9�s0�)ɜTNn�t���Ƈ���фx��hW� S��25��yAЦw·?�|�{��EDȂC�	��mww�Pq­XA{�ӊ����(<��q+�x�[�:�Q��s� d���.Ձ)�Q��}���p�_!>h��&*��>�(�7Һ�$IlK��d|�h���i}{���H�ZK�����>0������ Z	�ꜣ�|V�� �9 �,G*+����v�ߨq��w.a��~�DE����F#�/=ѩ�nCVJm��N�r(�[VC�y�H �����������t�ұv��S]V�+̕R:�ʋ�ڍ�D��C���l��{�h;|S��\��+������^w6<�{@糚�CN�,kq��~o"�6�Z�3��T�G!Z
��ǐ�� ���̧gV|��� �c.��q/L�h��ʸ�Y��������:
Ca 3iS����5��`A���<�,dn��t�jq��2慠����v���{���C��đ�#�TÍS0�gH6����O���̴�c��<0�3��c�b\}�LK�@XQ��A�<���:nm�E�p�:<%���K"������ c��g�I�pF���(�b��N�`�zB��ٚ�m����c�T�D=�#���
 W����{�0������t�;�R�;CJ�|�uĴ��w9ݸ�=j��֮��V�V*�f��x«���$9�r�Qs�:x���X0.�ܬ��K����꠴�B30{.l�6@N+u+�W�(�O/���U�w�-�����L1E��,�˧�.�Ķ=��z�x���Z٘�zRݻ�nv+��3Y�b������G=���u���]6�߫����śU���2���`<����bo�h�6Z�r��<M�y���M�!��³��e�
�v{ŋ��JX7��,~��dB:�}6��|D�I �08{=����cD-�m܊�G����C��E	��Y��lh�adAJ�k�~�F�����������������H��`�7%�pU���,*狎���I_���R&�����	�m/c�/lW�E�u���Qf�ū;I�#�	C�ʷ�����E�7�	��6.���}y��3����ڃb��՞r�����a�7����@=�e@Y������R\�i�#\.����'sɥ�-��va�k��	xʭ�q`�D���M��!F���haT��Jl���&<{g<�'�Q�i(���w
j���Z�������b��v�k�������X6wx'�p8)��:�	���5�;.5��r�](��>�^RI���[B��.�w��j>ށ�hi�|�0t��<���H,I��<�����ꄬF�Y�ID߁�*����L4�~�B��JT�μXR�l��B�mґ#c����U��x��Y\�)X�#O��b�8���Z�c�D��r�p(��\���?�/+;���j	Mu8�ɕ���v�����l�J-���J9ЇU�GjU_Oޭ�y\V�n8�H�$�Mi�����Nğߡ��L�2�$���bnA�Z�	����1��^2VֈL�39:PDh�3l����v���m㗩k��� S'�Y�}A\�V��������WJfy�N�zH���9S�
}��w5�T~Tru&o,��)�%4�@�x���t��|E����1t4��Ik���J���ݙt�5t�d�����5��7�Ӎ�̥��� I�!�וÚ�������	�^d3�lFn� �R���pEC~�17W*i3sk)����_ǶyC%�
�Qƛq���f�2c��cdU����3�6�?1챙:��݋��v��|>�[È�3�Z�W�	����&��2���~jEѹDV#S��I�����i��^{�+����R�\��Ms��w��Y�<r�~t�Q�+�b�OY��b����Q�7��EW(Gr��l��]B@T��jчb:-��-X㫉j/E�>�������l��gȸ�G�BQ��Ig�}Ģ8*��#�E����MS��	����<N���ğ	�?V�FT%���M�#μM����ǵ����i�6k8)��F�j(����[��N��&��y���Diߑ�gB�/���
k�i��h6����a�����mW��0@��$�mȝD������AQ*��idь9�e��� ���[����-q2�"�~{���h��	xQ�K8Љ[�n�H�ćŜUt�vo'�T���A�{��xv����ݎ����w<��
 �`]ӪR��:o����3����Ҡ�
�>Q��~�f;��d�M�P!��M�d��0m��Х�g8�n�_(�b�����N��4��+6m1���S�X4^����
�X�v�}.�U� ��w�D<������}5�L�~���#\���XI�ŗ��|d�*4����Y��.'r��F ~�-�#`�2@���*X-���~v�2r��Q�Wꌏ�x�Z��%|rr�FR��u�=���� �&��ڍUJ L�O��q�6X��nٙ��I�ܶ��av0t���c���VP�򘽗�ƴ�&Ռ��P
���(��l�,A2��K�a�m��ӉC���_��'���yԵ_K��У��p�p��؂b`�\��h���v�g����O�I�S�N�(�E�M�o���{��1.0=�\�#�1�����[p�o-4{�1
��+���E��%ĭ��0ήI��zdfu�W��*��Y��ױ ����(�ε�!��c�ܝJ�\QwR��$�H�9�C�<H _�u"��O*�%c�U����K�O��j�G�̆N��բ���K%�+�*��Fx���|{��|U�;Z:	,���x�up�q� ��+8'�c��'�V�
�Mmkuk;M�{ �_8D��uzyN�R[ۢN�%f��Y\}���!Ӕ (Tc�k�����;,]����N���i�#l}G�1�j��}�U��闧�]�b"\�&�����u@��ͮ��.o�n���O|�1�X��|�ٗ-T&s�����.��fv7���G ��x]�5�M��_����+X3�#�x��ᤦ��L�Ŕ�#���O� L�!N]�j�5n��	��0��]��#���?,���GW_Vtrd�Q�c���PM���d)BtO�T�K���&o��,��kN7ozE����¥L��4�Z����S5*���4[d�atwk�v� �.�*�9U����YVJ�z��;_�8���Yv�X�[p��A6prߔ���X��4�9Z�ě@d}��_cr|tR�1�6|gUǚF�ͭq����̑�n�ӏ�ծ��B/���#k��T�����G��W��9���H��;�q��
#�J[l�a݈�r�9?�@K�pk�(�xLV���M�įA�����c�N}<�t�M�+P�2zmB�`�O6��bj8C�!�D�֡��j����bؤ�_�Ң�7~��Շ�!�Lc��)b�^�)8�?�	HC=�@L�	�*@k����#kB���*:��?	�s�|D�VHC[5'{SUD"\��� ��D��U�q�;�����e��a������@n�s�"X�P"޾��w8�侾����þ�.����J�0�� yV�jXo�k�6�t�3�%1�ρ�3������ft��x� B����ERd9Ց_��@T45��
kI?P�4L�pvو�N��� ��*mŵ.(y�����-����Z�n�8�tpP�Ѱ��p���qr�;y���.#���(���Wl�����l>a�j@շ�{�I@z.�˦'��=�/$�&�R΋aG�<.��*���Hŀu?H̔� ȀSW����Z�y�3��-��5l>�e��x�����&��3���t�.ϳ����DMղ��*<p�5܂:��)�O�����^���)bV(�n��cHg8D�i"bG���?��%֍�\`���ns�1����|��ړ�nl��mo�)<p��ri}i���-�(�-����)�{��뗑
��[�V�����O�
W�A�+j�P�U2=<������#�]N_�Pل���U�TĞ�*�8f�Ѕ%`�䁻�-�]}m�鶞n�{�� @j>8�M[D��F[�̏�"��N��\��vL��ձ��W��PW�Cp.P���0{d�|��[?�s�#a�{#@S�K@7�aK��:l`{���g��	�f+�L��&�{��7ܵ�@tg�d3!MS��c!��l>xdk��M��b0�;����7Úf��5����m��B�&�-�ƭzM�3�(�N�j� E$Q�Yx�{	N>Ƽ:�Ѝ�}積�D�`�7:��/y2)R�#���1,��a��x�;��A���>tL�H�y�'�;9&_~H
s8D��GN�0ɵ�O�M��ҥS��N �a(����~����:�N���Sk��R{��z妩4�@�<�j�׆�vhn��d�"H�Ժ���}����-��@ |�g�;G�$e%�5��&>2�wtJv�K��MG���i��\���^$�����m���D,��U�l����k髧"��wn�=��� �W�7�����2��X�.0[m9��њt��S�(@V���Σhё���PILO�2���s]�O(P����`��~q����%!����*x)J�,H��uzZ����M#��<�>e�ო�[k��s�\̋!��F-À��DS�F-�)_���J9���ݷ�L����$������+� ]�����t�ý��wHX���i�-���5"�B��<?M�:t�7� ��8!�D��
B��{c7��@��d��6u�ƛ'���I�F���S�z��Ux�}0o*_ї�r���+�5E���@���Ӿ���EA��Kwv�oL����2�Z�֙��e��'�NR&d��+�i������0���d���w*����~��.��z&�M�,e7�p��lLʙ;��(��F�h��"�jE�i�����S�'��J���=���x3�87��ş2J@@���sA��e�l��I��Qr]�J�6��l���NE��C;��~��\�]9��^ɷ�Eҩ�hԄ˃u�j0:�Ye%k�*u�a�ց����X�yN�\u�!U�}}�]���FX	�H�6���Ӧ9C��v�����ut�Uh]�2gda*2M��?7�v-ٝ�� [Y�y�X��|�/��vY�ީ�A�����]oF�Ӱ�E���lr4X��HΣ2������{�<���nu�g�)Ą���n.zx��@o�@�pyy�f~N�=i)X�
�u^m�w�kT�!��s�.3Y;�E�3�opE�m��RW�%J�.R�#.�:q�;c�Wa5�[诏Fu��3�.�G��
<?���uV:���hp� ���/��v��]ȟqb*Β�)_�
���%Ϛ��[���Ĩ��i�@���
20:�40W0Mk/Ι���=�@ۇp���[�#}�t/ܽ�W���i>MU8(6)��9��hg� �(�cxø���jʧ��Hr��>����^�#Ю��ZQ�����W��ͭ/�uw�~cx^7 ��l�7�KCEi:�����P-I��F�\�X�K#�< �׽��%�*���HM=���wgPL�E⦎/�*�~oHz̳9��J�&���-Ţ��s��}�̞W���B�6���6�K�r)!�IT,E[I���S_6�	QJ�!�3l\��s�?�T�GE���B�̀W]=-�W��2�Y��K3������##I[�EKX���+���Y����{�ު����&��`��7ͽ!���|�"�̐��P��rȾ����;ǫ!��xU��4?�7�VK�A�rX���H��EԹ��=��k�}`�N�Y�~;g�;��w���H*��`%�'����-�y|�E(Jics��+Q-B^K�>��Ĭ�פ�	�s+7J�{���E<��{\Sgd�,-=�f1�N��2DA��Nc;��iI�'(�]Q�YKG'@��������NI}��j�O���5�<�;=�w�OW:\4RS�D��'95À�������
7��c,���f��)h���5ѭ�Ju�k�/��5�#�d�[^eS:U2�mp�n�$�[�N��&Q/sRf��E�#n��ug	�{=Ч� �G�����vͨ�WF�����`���VCݏ�a�R����&�:­6�x���0H_�²r,�8�����
�`4���>L��^mu�{6���3�5N�$�'s.]?���N��d���X۳�Q��%qU+r|��"`���rL��p�7��e{�.�p�sxY��G@!���*��%E��6q���	�����8�G+J��c{%��`B5k�������N��w9����-�X���u"�,ޞ���͟��.2��CWP�%}(KӳO[/�X���]������O�Ls�߳�@����C�G�9�}Y�]��&�ǃ�,���FK�j��������
*�5����C�L�R	���6J��.$�M���DmTE�y�3�2���k@hv������1��<&J�(�m���>�{�Gk?�a��q��EOL[I.�F�VP�� C-����T����Vp��m�����:�y�kɏ_n2F96�煠�c� ��{�����f����3'$��� �{r�:����5�갍Cvi�l�e�h�_c�Cr��M����E���r,
�њ��p��H��y�Ry����+OE�(O�Jʢ��^�����+:M�uV����d}A��>��y�_� �1IduU^7�cG� [�Tm�$�q�ei0�����[�m՞d]ܵ��w���d�+
ʎzTmu�1�u����C��P@o\g������풿���g�6����a�*^���%d�"�=>�Seա�fm(���=rq+X������I�@�E�bIˀ���C�Ւ����y:�o�x_��=#�h�>Pc�� 7;Ԫ1�mkh,9'D ��c��[���S��(+\��9h��6Ls�z�{E�V=��߅Nr	���NӅN����7�MH�^��^r-+f���f�67\���>G�n����mc����ۗ�7x��e0�n�~�h	>躣ݮ�4���_%{��#��r5&�c9EICo�ׯ�����cS��;�����@ucFUY�]�!�y�(YFT�B��t�dg���D���ۆ�iYU�V�Di��P[p�G���_O3⏡��X�	\�3��^�$�w�XE���?T*t�q��J��V�%05���RB���*	qV@�,0���䵲B_��5ZY�)YQ���)t�8qj�J�d��>�*�LTV�B����an�-}U�x>��i���ɥ.{7.��W͖����eN![p@��I��D�����BP뜗�FR���6��RG<�m�9�����#U�M�b��0������e�e�Q��#PH%���Խ�S�f����[��n����zB�����_g<���&)\�>�3����QS`�J���Yb�{�5�BkW�S�HB�����-��|h��������
��:=!���Yy�|���v68N��t��šJ��k�jS�L+�>�	�Z��C��ׅ��7�.�����Z���2\B���k6�G��Dy��	���Vc�f���{��){c�}�_c��y�!(͌ d�ט�o��q5�(�N��ʳ�	*y���G�%tj�x���$e��G��j��2O�h'Y1��NԻO:���.�E�)�@��[$��A_�Q�fun�[+�ݿs}FW�!��N�S��&�0�h*/�ԝ�v8T�)!~L'��Bm�7�V��f)�ݛ��>x�<h �T���UѤ9J�\7I�]T�FEr���_�r�v�}|۱�W�u_�+n>-3ޝ��ק��QI%s��+���ˍ�~��L��N�-9�0�����p�8��E�2k`��R����Q$�E��4a��1b�!������"�I,���J'�t�ҁ0�ᏎC�n )���^���C�H`�=i<��k{� �t*���GxB9(�4*��|O(������@�t8k�1G�b^XZ�:e�����U�zB�jI����[��������q�\��K�ѱ1�y��<�ə���u�qS���h��TƕH߿%��9X��1�˹c(LK�<�jA>ߙ)����p~@+�L�YӮF\W65���?���^��?kW�YCSHʰ-4�� $9��R\��u�����n���`�tp�+h�}�`��>�2m��m�-M�x��*��F�}v�r��گx�IG�'Bj�����<�EM[^x0��XX,�:����{��(e�AY��{�=w7T�/I|Ե�7@��*�<h�= J'J�^2����6� �Oi"q����z�.Ǉ-����H>�{�BHdH(e���*#i�R����=�Kd����3l�Y[��Tf�٬/{�@�@�_��ޣrzd�;�q�0�a63������D���xJ�,�tu�nzOj%�фH���@qvv���
��pА�2&�&�Y/�E�Ù��?1�� ��S���gB��ƨ��"���ګ�Շ�5�oֆ�~'��jW����E��&��4}l�v� ���i�H��}굼������ua�Q"�4�m���������tB��3Nf�%�;���? 8l��<�eb�囃u�y$�7�=V�RY�<Xk$v�j�_�ѥ��/~�pae����ei�Ks�L�)&�%t*����ڗ�2;.�G|�󪚵Ә�Ȟ����<��
�ҳ	�$�t���gC�e1�S%�fo�<D�5��*M��8&g�����{�i\��.5�UB����s�0�J���;	dV�,0~��QBS���Mj
����Z�n�mf�^�1���+�i�-��k����ܰ��.���	�_˽ٶ��`�����E.�7�P<�KM�;�<�����Wi��+6�'یT{6�c��^G�j��S��;�{ �X��9&�/$�ـ�δ{�T'Uh꽑�cI��K
�
Sk�g�&�Kys��-
��7����K�@����Z%H�ZB4�����+�mC����QZ�q�oH�v�q���3�ia�]�M`  �o����s��Q��U�t�>@��"}h$?Z�i�����cX�@��/���~"G�p���sv� ��3��=yм�k�~cNBqBs���noZ� t��b6|Ew]�I�>K�$g�2�a�u�}�R��^v3j�Ɣ�����v���u�?����}{vY���j����⃏DB�C�Z����� �b�]�x�X��������}�#��6���h�A�����)����yaxڮyʀ%�$�40(����="��wDÌ��,��g:�3�+"�������	�<����k$�+�z�ʎS�R5���P،�Z&90cd؎����Еyx��ӭ��Y�K�e������=��R�q����26�N�X�P��(xuC[3b��Ea�˖�K�o��%W��������򿂆��?6:h+l!k
2�(
~�� qխ�^O��bʐ:i=�<"�J��ObY=�5f�ql*�J>ri�"������n����f�@�4�\�����]��_9=6��w6e>g��C�>���>O �	�� J����qdV��y¸��lH����-|I
K16{�˧�m��7t����4?��5��}?0�L2@��)#��xN�H,���P�'��"��LpGC�����]��L��hoBS�q�(@��t0�y��I���H���ڮ��b���n�=��
PXy�C#��پ�C��^�xT[I�"rF�6�\
�&^���Y�N�\[	h���0�{f>�P=3���t@�>�Z9iI��r҅w�\Dp��c�'�"3����z���G��L�6l_s6���lL�k���0q�0�j՟�8֠�SJ�����U�n����i�Q?x��r/�<� B���y��f��L�T.��4%���kB�b?{�L(ݖۦ�2�(�8�5����gY��}�N��@ĝ=4��X�����͵���nIn����&.�,Ez���t���i}`��3D�j�տ,_q�@��he���<as"*��jC�XLu��RO���R�8���h@���J��tl��3��9�:��؞��v���TL�n�x߰r��b����㥉�k��[W��� �eJ�������6V��gH���p���i�=��NA�s�2��霔\���=#TB�܊=ݜ�7@_�_#SVs`M��F,;p�zQ"|�9����09ц��4�ZowI��r�3�p�������	���y:S��c��l@�ȕ�'R�t�^�pu���1j' �~~ނSo8��c�W�`��B�&Bʪ�.��Ԃ$?z|���b�?',���h�e�O��[��=W}w���H��f�*�G������K:h�Xi���u�P�p�Y)�P-�>�3���ڜ�E�H�n�����V�<�Tt�E���Y����b������vn��?�qD>�顩RMRi?v�։e�
���|�r�!#A�؈肶o6T�k᯿���U��н3R<m�H�)��U!e!E���נk�0ڱȊ�#pw��a��T�q'>m���o������ �.�)'�6,���&�
i�����r�h}ⱉ6u�]�A�W/�{?�U�>x�8>�m�������.!�6��8����%)K)�.T(��7�>~���MB0�}���lv�W� L�~䜛�N��)zΚ%?̞:�wv�`ݶ�8�姠�鵧���,팎�gbHM���Q�Z*�;?e;J��<3��N�|�r ��IS҂A� ���,�ˌBe�&k^m�C*)3�##�.Qե���w�]�?�Z1� B�
u��
n���44���v����u���ߵ���cb/z����~�E��0{�0��a f�V�M����g��M�~���yυ�P	�/�Ǿ,�}L�3k�v���_+Q�h�;�bEH	�iu��F����k��PA�\�}y���Y�����@f�F�D���1F����?l �����#K^!�:W�А�p ��ؤ9.�)�H�aĘzYଅg;�bB$#���5�okU�;�_��O�N����?V�R���)4��]����R1E�˝��FoX8#�]�B����B��yҠa򇃤�֔
�&M���o�r�N��!��Β�7�7�`;�M�����:�ַtg3'�A�7J&�7�v�WI����1C���P�X.V��5��D���p{o̩0f�{@Ʈ�%�9��mG�Nu�]�=>�H�݀
���k+�p�	��fz�w��&�#�]oL����8g�c��I�2,��.��j �a����Ї����t����(���:����_t<�eWb4�d�3u�`p�Hy#L�3���O��*�L�ˈ��#�&�vL�v�Q@��y����~]�v���c+R�yh˞���+G5L����
~Ah^~��)��.�%����ρ��&�~Bz���r+fg�
w,�����w�x�׀\%+az ��L����0N�ӥ�#h�-�.<6��@�3������b��*]N�05e�E��R�>�*HWbe��5��l���+[��=c:]k)��5�b22~u+�f7C������u�B������=�I��B���P�//�0�[i�T��V��rۗ�_&�r.䵍]5�9o�zw
K8/���!Ze�L}�e�uG�K$t��ɟjUE�v T��G�gҊt�JF�Qcx����᱾�U}D�E����{��w+�ץK��	�_%�A�_SӲ�f+��_�R�<e~ .ׄ�BP-��"�rNs����^%i��1��S�ɞ[߉���3e_ k���m�;�Ѥ)U_�Ӣr���j j�̙a���^��V�.rи�R�1��wtXX��'뀑%�=b�#���j���܈(5K��	#��\���9��޷	��}B�Dd�ꖆ˃�cW��N ��p�|���)b�~�[R�Q�M�^L�� �_��Ǆ����Ծ�N`n��Pҁ��J��$f��;�L��h�M��	��E���SB�jj�(7d����z��"��hE ^FH�!�83��m£�Z�׆<�.<v���&�p�[�p����R����º1^KQ�腃�qw��n�(���A��r��SE5�,��٣���3p�m��`:��Dmu�uJ������Q0��2����!���>�s��m��q���nc�����Tv��4΍zW&L�'KP$���qO*��mzlɍm����d {����M ҟ��?U��F�"�]ڈ�:��@w�?Ӳm�j�4N6��e�~Y�E{k���GX�zj��XL˴�y}�!���G��5P��n���Z���Gq�|�eg��v�cp��_-��M5�����
IG�u�Q�@Α\��ws81�6�@��'7�Lg����Gi�B�R^�5�퀭�6��P�6p�ͱ ��b6+�E��D� i��S������-q��o%9�5�dTeZ�J冖?�r�:�� Vb(�sr.�s���)��Ot�,�'��|0�u�y?�JNX���7w�h��K�TM�k/g��_qD��'�h�)T�&�ƷE��Z�3o��õ	��$�<�U�	��Q�f�z2���3^�f/}��\�ܙ~-ު��mq[�'"�F�ʍnu����W�p~���q�{M�[g߫��&aI�'IB���`3�.���f������bS��ѬS�i|;{��k��PN$\1f�@0�x��C>äN�]Sc�׌��w)@�&��V�V*C�����Į��g�՟'��E"U[��E�۟[����p�6nP����qA��b��ӈ}���9w��DY�v�x� ����G�9���h�a�Vj�f�*g���^)��>m��Z!�1�3ԙ�ǻLd*;{TP2�=���E�O/��ʻ�7<ţ������H|3�as�ؔ�����1Ɲ5~�Ub���-��ish���9V]���7�(b�f2��q�ɖ��!œ������C�8�����Fhm��'}k���6��Z�[s7�����w�m��_u8�:�"N��״hVY��G�h8�	h��qĊs6�d�&J���5�|l�9Q��˻�?(HU1i�'���}�k��mݼ
͐uo�Z�)��b��xغ%tDl�f]���_�����}r�r���sF�Y����i�9T��!�7��xQ@��>�F�4Y��~�����P�7��WV5�<%������e^_yA�,ͬlH�K=�x��@��� ��M8����\��F{F$��pu��0VE���Y����lu�xWd�v�w���.���K���E4_���>3�`���	���'��F� ;$�WX/�3�U��>��5	�`�
��-D��7H�xٍ�U|�k�����J�}�����N>x�{*يf_'�B��\J<��m~l�N�q5
�֮V0c�p=g뜇�V�Y�Z��y�9#�9#� ���}�#�����e*���<0h{�A�3r~_�5Y����7�5켺�~1�FZ]��9X�	+�;:Ǻ<�k������c��s�g2�s%�)�/����a���Y���b۲JH�Xgݩ���l���@�f��wU�<M������6�c��nȭP��<5��r�PtZ�p.�݅�:����M���͜���qG�E�%ѓ�Ꞝ۔w�S�����n\�ܫ\����d��m��S���jh�0���Z��0�eb����>{�!�I�M�rY���e#E<��}k0ieҽC����q��Z
C���#Ťh�L&̺R�M
5�Pcw�r�$�T��5��GÓ�M�Q�o��Vo����y!5o�7���j�-�O�\q/]�J��tѶ����%,c\�!R�dG*����$���[�A�����n��X���b������^&|n;冺�'̬iŻ;]��� �X�V�8�y�R�Ah��$���e=!�j�3�r�F%���j��Mc�SWK��k��;����cN�bI��;ejZ�8�'�]]Ꮊ�T�q�ۡ�:ڼ���P�
�x������#v�x������0�f��۱-ET���EQ=�۾�7a��d��4�d����u�֢�ѼF8�$!�NUu��ML�z<eh���{	�+�q]�(�����~����V��{.|�CJ5n�T0�a.�?���l,&�2�O���H������,׺�>Um�Mrn��f�jf�Z��s�D~L*����f��͵�p���0�[\ę���ן4�C{��<�ΌG��P�)�R�T3#��J.��7Iq�kt/FS�蒸������[�ɸ�b�:������+h]�xW������|Í���� 'X�͙ӧ?G��(�L��zC5m��H�!��ɵ��/�ψ�_+�T]$Tʫ���X�Awoj/(~=��$�/r^�u�q��_�bR�5O�.�O�ߕ����Y�7����]���w� ��ZZ1F<_욲A�ey�����w�,�$�+�'Kk���{#�=8�������ⱺü��d!�|r��r|��N�j�7¥�"㕂6);�I���WHA��@SҾȈ60������"{�pL%�P� ��=øR���b9P���Ֆ̬�}�{�8j-v���Nz[]��9g��,�}��k��,�� _�xv���ҭSq�h�Ek�I�ۓ���G�~+ˡ ��&�d�O�����FP� ��ߦl��+���\�@M�%��DW��k<���#���u�,ϟщ��.��DF���
@؛˪��ܼ9~FƲ�J	�����'�=�[2��Z���@0[�JlIB��x�S�;�qV��<�c/&O9>��7��`V��wIȃ+	)ę���l�<!M�2XO)��5����}�z}�VQfU��!�@u��^_u��2D��s=�˽1�a"���CVx:h�(V�:,��3��i�E��!���E**�r,�)����x�_� W���ư/ҡ3̲��� �Z��	��+/�}*���ad�z'�%M˗Z��.��FfL
7��7�<�pa�Ձ��̄��0�O-�����\|'���HTW�WO�|�[�ۅ t2�N�w���@��.c�>�g4�83���}
�e11��D�ɴ�v�V+��#�3��l?�	����!�E|a�e�IT�T��:z����څ��ǃ������%S�&��kQ]����	�#\U.��{���@+���ea�$up"�1��f��/l���{�:�fC> ��%��^U�8)ɴၚ���W��Y�(s�h˹ʫ��jՌޟNE_�e+_5��V��Y�8��+U���G�'e�J���^�8_3>Ć�f�žn�D�̄T]78����Ǟ,�T$�L-鮍�G#(* WL�u��5V�4���m�/NW{HtDjt�^���H���������0���ğeHSy��gffg�N��� �$ �uMh���D���]zZ\C��YT;ŏH�S�ANv�X�hƵ_uz	�4Kئ�B	ȅ��@��#=H_��P�+.���1�Ǫi걥F.*�|����Q�"�"_�z�?�f����p�HK��S����'q5�Fj
��a\������9�-#�d��V6�)j�M��Y��g-�&՚ڜ]��$��ѕ��M�Y�����I��$�囁�+ʿ[ݰ�m=Ւ�Zs���T���g��e4+Y��i}���6�fMط�Y뺕	��uku��i��x�"��'ٿW�7#	E�z�֠��ϦFH���M5t�#��� �S����"��d�[�X��bJ71l(ѷ	C�ϴ3�gw%��S�&$��kkn	�J�c�Լ�;����wC.k��� �R,��5İ�h��i-a����_% >� %ǐe%_�C���\��E������(��&Q!u����bBܻ�\gRQ҅�_�O�J��`�%���\)�!�r�R����&��(�>�Z�^�Dq��{�������v_@�Z�X�9�I-����Eh!"gD�R�� ��x㦙�o��}�2���h�dk+��[.��^+޸
>��`W�N�|
r/J�tѼ#�0�+'���3ۃ�|؂�"A�j�1~S=�lcU�r������(�x��[??�:����R���� �g����T,h��OESW�~{��*hG	~��W�L6���T0n���Õ��,��o۹��@:��I*]%a�j����&V;ESP9KtLI��:�����jRC����ϫމX���*��$�`����g-S�K�6 �.��:S���	_�O*��M��ξ/�{�-��E�Ij~5w�6PjNm�t�������f�E9һ7�f?K�������}z鄴pEN`��d���M���x���g觴h�˂h}7̶���'����x,�j��F�)	 �Ƽ�g^X�\��{g���� ��j��y�:H�{v��K�E�6�XPV�yZ��^Hj֪�e�y$s>��ր��ծZ	B��Y��ŏ�[���m����]�c���$�!Ɍ�W�;S��*A��1����n1�p�kW#�?ьӷ�4���� ��2�);'QJT����{]0t
1��^�P����ᐗ�|ך�ܼ����B��KTI��N�_�~� �C�Ɏ�j�;K㠮��(5
�n� ϙ��{�4+I�u򹉡��6�1�IQb�`��I�R�a4�[��S�aVɺ�>	3�˛�`�av�u�͓ܼ��|�G�ۀ�Cc�cG�m��p����fL��`�2�w�L(U�|��DY�4�HJ}=j��,�Z�z��
�|)`X�!�>(&�):���O��J���[z�E�]���s���)�\��������br�����P�%X�M=lJR@�J�T��=�Պ�p�@��n��gʄc�X�v$\'�i�52z�:�p���$�Z����>��`�/�'>��ɬW�f#��_����X�WC�5#� ���I��v[s�E��yC�te�R��+�o��yg�K���vz��-w#y��]YC�N�f�0Ěu�彙��Q!�.�������8�)�f��qu��@o&X� �Ʈd'}ʤ]D����K ߙ���ժM4Hcb#��yȕZH������s��:��K�Q�^<��HD�\2��3.{)��!� �s�⩉i�܍@��	��5h{�Q഑R�zJ�?d���'^��s7VgJ�i��eF����)p��Q�>R�U0�d\r�G�!b��/R$�U��FȌC�RǤEk<ǑX�&A��.���s?5gFՖVG�k�����$-|._�lBP%�y��H�����|x���p���1���$��;/!�=� �����j4 2Y���ʾ�G�I��) ��H��9��iAś
N�������\���yj��礕�M�0�S!���(�5�K:�o�,ښ9�;lb�
I�Q�U��;����r]ƭ>3��:��{|F���q�������6ȏ�T�+|��P���	�A!�8Y�K��tA|v�� _K�l�z
n>#A�a<G�|��b�����^���2��i�R#0�~Ϫb��<�4��{�f:b�8|$rP"G&t����%K>U�8�>�l=)4�j^��[@�xdG���W���2�Dvຕ�I��������"�M�	�����..���E����M�2J�tҢ�>U�4�)�Wl����-鳍��n�X
�D$-�4P��B.��D����M�V�d�~c�k	�a2�i>�Z>�Xy��%N�hlY�&�A��,�F�g>K@�KH��ѣ��Vw�h�"sZ&h|2y�j��	�sC���G�0d��� pW�6��O��h���^���ܻϥ�5C��Kwi�C8���6�>��2�{δ������l��雨�o'a�05�ѩԀ���B(� xT'�ۤ:"�^�� �>e^�{ � ���n�&�k�S��!`S�=���HY9"��,3H&K1��i���uͯ�6�pi��p�<�{�a����Hc�D�l�����kR���Z��d�x�CnA5N��=�~�fO��/��S}ٌ� �����讗k�z�8�}F
�� ��#�-�pL�m͒dut&4����D�����9w`�����V/�c�0�q��P�U�D>Zޙ�"����oJ		������.�e�\+嶥��҉����ʶ�,�Y��UصHs���^�7MS׿fR�II���KFFv��Tg�>A����1���}e�/�4��$bf�����ۚk1#�*i���έL ���Z������帿)��w�:�����pJ�ih]:l#�O�S{Ny*)*Kխ�+W�It�&�����N����Q�?�`9�� �"� ����W���Uu9jȯ��٣�L�Է���*e�U�CDB�)�	�F3s-4����w��_��/%kR1y��,��ߗ��,�6h��'���9�Oō������RR5{R���蕗�qw}��~�ޕݍ|�z�W7�v{&��~�[�F����m�߱���V�+�i��W��`~���!*�긲��J���'Gzg2�"v�6�_4l�x��Z�l�D�܀����^�
ΈB,���7v]:���I��㷨��b�q�l ��[S��AǪ2�S�_a���1�9���!u-c��>�A
����[_A�	��F_�柠��!tG&��0�xdFLk���G:<G)���_4{�w;��	�/`'�47J�O��]� �2��6a-P~�*1M�S��n2�[�$����W��gb].l3G�&�7�E~�B��0�=��/����c��B���`n#�� �J y�_���m1���)�	ׅ�8&��:�9ШE��~�x��z
��?��;�0�����ZS��$d��Tr�	��>�#�M13II;���g68X��QI��M���M�95iqK��c�M�h`%t�I/K0 �#�9��]`�GB �p��:RM:e���oR���a�<����H�26�����o���� ni̔�����2�~���Qwؾ��вiq���L2+���Q���*�����0ttbW��Ae���ŕj��⍛J��ǰ���	��PF���l��{��:c�O$�����FG���� S!k��3��F�享>��h�2a��9� {}�3���RΞ���6<i6�ʂ�I�e�u�q� A��O9����<׮4���WL�HLe�Fp����I�]:�Ӳk;>�b�~���� +T�hϗ�#��"f���Si�J���@����R����7 ݾf.�ڿzL�U�Q��E�jj`Zv	�xZ]��h��z������w��}��l���#9�$��eD"��u���] �U9A*Y����
��ǭ�>���S��L@���ޮ��2��3y;p#�W�̞ck�I(����ؕ�4[��}`�rҵ�~����YZ*%���q5��&���������^��lW�z&��xf�4�=��j��Z�)Z��MOBJ����KcT�_M\q%�����!��
O,�e����T���яt	���K�p��:�ͼ�ᇫ���/�D�QR�q��L���Ͳ�2���0�(�q�����+�@K�d|�ö�����B�����(��%��gR5�J��Jd�/�`��ܞfM-�?I����Q�����\k���H�U����p�̽�� AQ0�.T�.�� Zkj���l&0`�ɠK���|���o���G2ns���*�f�ͺ<����e-��(A��e#���ߥ	�
�04�����kV۸�V��5E�[���$����-��b^J���x9p}�@7J�w
z�����_q�	��A�^lu�����������OY)y��Ƞ!n.�ET��iM������sBl���4��4d����ZB�IӾE�w5Ï{L)e}V!J�|����)O)/��-�e:|�4n�� �c
�����^����_��	f�����ٛ[)B��y~kvd.FY$/mr�\�����	�bf:a�L�]N[ gG0�Bx��\����LP��m���4�(\zC�ֲ흮�J,(����۰{k!��CN��t�#���-�r�cU�"�B�w�q0�Kf�Ta"���9`����?�e:���N�%�{UӀ�F�mª;w�w+PӟЃ�K:77��e��O�|ݣ�B*?��V[y{�P�hcȂ�����8���H�vW��N�V�<$�ލ����=�PU��n?g|�d��f�l$kD�.��E��m	G���P��Vim��T�>�r�6���3_�J<�G����}�F���ᅄm0�\��?g(�c�����w�f_;A��7�Io�T��%É���I����&~q(�*������iG�l���i%���/��袈����
C\��yR/���>�/>!m6�>�sȣf�a�Y���Q�gua�1��P��!��������o�ar&��p�kW����v��pz�h#>x[�x���%?V�zr*��/x�o/LA��ƈ�*��kL�L&��#!����@�_F[���L��k�I���`�#�?}:�T��#|��]c��:�ץr|����KA���c��j��LF��� J,��K1JmT}gJh���:��t�%Ǫ��Ҝ�?	>~J'S�,
�?u�{$Z��[�]�K�\?�_uY���i�i5��L�@Y��)�U��/PY;yŨ<:�]E�m,���r�7��_]��6W���k:>Oϗ�����Cc�Ψ��w�c���w��U�^&�Q�N�7-$�k���I>P��^TH�a�HB���zE�t�땾%�{a$�[���W֛��zY��YҹzAc�b'2b�P*rq�yk	ӓ��Gs��HOQ_荨��t"��_#�㦩+P��T�N�K������JC�;�/d��U�=��;�r��T`���$~W�[�m3��	���-ZA�/܏dS��6'X\� �� :�U�W�;rlYM�����ɽ�Dw��L�!���{�$�Ąo��Z+�h	
S�d�1�w�5������ �2����q�i��W��w5�٢ڪ�	�k�}����l{f3!�;�#�9�Љ�50�j"���ˢ�{��c�Z���'J)�4�M'�;�H#��i%t���Vn��|`)5��
h]}���:���z0^2����U>e&�k��o5�<�	Cв�E8��<�)M��h��@z�5˹�ӣ��$7�O}�N(��?��D�� o�ź�5;"5�Q���H��0��L!��.�}�}Qɶ9jK]_	h(�gV��"Zs��<�~�_Y�-�@�
1~��~�e{�z������U`��v���x�m��?���o�/(Y��fԀO7Q��k Ι��beN1�r���ĝMF17b2�
@��T_�zD f*��z?�K�����[Er���8U�E����>^��IF�n�.�d���U���q�ȸVz�K�9�zQK���u�{yc�H��,���V|c����N�B��_�T����U��K1� ��~d:�:�	��~~!Z~�
O	>�Ũ��3�|�u@YtA��3�ߑr�B)��>8ɈH؏�H��pzh1������n�;��d=���.��0©���I�(9��E.*�leG���D����]���,q���2uߚ���s�g��Ȅj@�=<���?+�dwo5�k�sn�F����T6��5�P�|}8.�X�#o _��_k���u�B����e�א&�y�?N�Mɴ�Z.��9�o�x�*�|���*Kj|;�ԋ7��o٭��E�*g�$T�ʔ�Jf�b8�&�N�'_�N�����̪{�L�;�+�Z5�	��`�˗>n#��z�{��l~�U�8B�sd�� �Esy���0J ��L���Y|��W§c8G�4~|zm�ӄ*q���֢�8�\So���ML2	a	ʧ*D�,�[�3a��}��ٌ�c����ca�PX'��3 4�b{������bg'w�}�}hR6�^D>�r��5�.}L����U���t��r��F����"H*j�Z*� �;���)��_�BH'Un$�z�6�uO��!=�����--azw��7n�ߘ"���Xєp������?E�I,�ᐡ����Kt��Q�F��i��q�+��\�D�� Aӟ�IzGr�Y�����=�6����cu�]����Ю��~t��������!��	�&�X��!hM����B!
����6��CG�n���byM�'(�CLX��#�k��Q��q���+	��-)�ht�O�ӗ�賊�/!����ˎ���L" �e>G��ԧD�͆]Cy����뎪#�[�o�X�;���у�R��zc�1=�m��洌���d�oka�Q��J��Ҿ�%Y��>ZK������݇៝��PQq$M��|�7���0L�p�&i�V}B.��Mo@�B�g�)A��zg|�}�	/sx�#���]o�8�:3�����I�������Dn��(��u�@"�&��j�&� �UB.Z�.:��{��^�
3[m���b��@xo�K���������|�^wx���py��1�kl'p�Q	�;m��b������^|��F�,�iO~�8�#z(���e��r:(�D �4���1?���i�v� �?��ܔТQfl��T��Φ"��Q[i/4jO�]�4q�cY��i�&��f�������́�7��J
� �l�*2P���R1�KW��[w��xJ~\LL���=w(�ԅ���9���J?D�vBS��3 U�e
ټ����2�7����8���Ob���t��Llb�kމG���C!�`	���Ks_�a�ᱺt�:�.�+��gY���ƈff�q����K��� vMԽQ	�%鬔36X��Հ�=ˎ�������L����K�z��i-L�78܉8�u�Lp8N�����Q�2��j�:^O,9�����NjR�a�8�'X�N�������j��G�c>)� \�e�������J���G���.�/��`.'C�� ��)��J���(�B��24����[��X���f'?�}�i���c��?�L�
��+#�?�*n�b.�O�X�
��Ap{�=�Pg�uC������٦G��[��=�N��#�#�pLet�c���I���c���a� ��v�es�=UrO������ �ޖF�a폕���$�0���[K|��%������Rةq��6WZ���0�=f�AkH�)��j�e�Y�A�.}i�I��:�%+��@��m3�F?�㉬��z�����Ӗ�$�R�>���������(�>��!��T�d��'].� -�p�^�`6�O2)j��u�^�P���νA��&�;	�dȼD���b+|�LDLI���M�[�>��Fb��o`�x�[�m�aG%���y��Sj�bK���`
c��A�h�����s����y�G4�����7��@�5FC$�����Ɂ2o�p}��Bt^��F�5��G�Ub�Ƅ�o_�ܩާ���5�Gi<<L��V֬�����
g�n ��[�@%- ��<r�)刄Μ4'�K]�UN~��	�%$n<�Z��SzG�<�K+"�;�h]FM}��m�&g�7PG����_!
�V����� A�o�9Q�Ȏz&�`�u���7{��[m��b:��f{2$7ǭ���k�������(Z���p9�3� +0�ASw��`�|���kz�&��j���
����hÔ&��O  횋�o4z!�/M-���!��:��/vz���g#;.a�~J�>o��?��$��e��T؏����Q�}�%K��b�y+=�Nfӑ��=&�:h's��sLЙ����
���<�D���ZR:Put�ס�]�� ���}C�՞]��&���u\b�}�=����_Ň��Ə��Lo��@�Vz8~?�Ŗ�I�E�B��sP��X��2@"��v
CW%�6-��̭j�����ݪ�`�ω�#!�4}�8}���_*�:_ʪE�1f�2w;g�\ͬ�@�U�O.RI~e�17j_a(�`�hŧ��-���'�8?�J��%q�[ԟ�����m��TJ-�>�&��m���[�ˈ%+3E���>�I$�y�F��s��\~4Ғ��/
:Bth�^l)��z�C��vW:'!ϛ���[뱠�X�x�KT��8DjO>@���U��3e���Ө�b0>ΓC���~w�&)Ur$�l38Tf�?y���=�z�
��Q:��wGT�8��ᖥ>���E�R��-�4tS�LrI�Ba���VKC�kqf�F���i�T&�=��
����|ZY}���ݍ�r��Qi2J�'1/V��[��!�s(��
a��@	�g]^�3J(7�����:ˌg�	|ʑ��B��8(C��U@7Ѳ���r����UE�1����⼣��F�\%մOP��z<2j��屳�in`/?.F��zl�#G3t?�;H(R��=Ѯ��v�I��ZOqu��H��b��G>Y�Y��y��h��(|��y4����l)&M�l�����rT�D���F�����beakE#j�A�&��&��z��RԒ����K���*Hi�3��E$�l��=(ę���8ܾ
��n�v<6����ң��嗳_�u
�a!�?�:�9k���A?w���snR]Q�Q�X)k�����_i��>�vk��6���2�UW�rbaȼ�D8����;��7J���B�EZ�e|��'�S��7��#¬B㾺NY
C��Ԕ����s��7����&-�� ����+s��YKȯ�) �3��G(p �S�����^�z�Y%"�
���D����̡a��c���.6 E��PAY����_�U�3ą��T�7��sC����k�6
���suZ�NH�uV��.�׫r��؃��>IO�N�z%/����1w�A��c�t����'�����ۺ���cVJ20��S���^M�+��~sXF8�2q퐒��4x��"g���pz�{)�N]h3H��^�y�FCh�[��k݄�����iƏy�Ο��į%�$��z(�+Zu`��F{]��$��-�j�{�u�D� �b����m�k/G��v�Th!kI�iZDԂF��fI��Ic��᫠��y|�x���[�=�+P�/�� M@���#٬��Ǡ_%_�!?���^�*�$�l��@�L�w��2┶+0�CI����$�0�d6�[���bŗ�g��ƣ��U��b��odk[��S�~���j�Q��4~�=���w�ScU�a��T����ga�!n7�Mr��_�L��
�'懪�G종�k�����>à���.1��f��a"���9�>Z�"��_��l�f�hYK��p�n��$��/��x���[z�6��^��a�r��-0Q�ĪB�1�F�rJ�d=�C��f�a��F%o���_�Fh�:j�Gw~%,������O�䑧�.��nx���O��_ǺX��HO�ˁ�QB��}�ꤞ�����c��hj��Ѯ�ؽ� �������dWf��laE����7�G�|�OX�M<�9y��QdY��H��*��'�Jދ�)��V\ڏ%c�ZO��v����uXٲ�?|�h���<a���1�(#��w�%_V���-��P�e�' �t�p�(���V�O� �'�_��,R)}z_�����n!ZE�rl!�_E"�Ǧ;'��1��eDB���w�R�S8[�6r��ݳٷ2���W�S^�
��.���`Q�}��c2���t���V��4t���LX0{�=�ynH�Ħ�H���4�E��S�zW3ĉVt�ś�oPB�N���ke�k����H�ԇ�Y��Oʚ)������ b��-�CN����B���ȼW� ŕ����`���'�R>��0Z����˹��н?�|��|[���1Wr��F�T��J����q�}�B��_��.8Jx׮S\F�&^�G���{���u��*�.��Py�ԥV��L�ƶ�=ƖՓ?f�sG�컯q/ą
/��q��Yf�,ܕ�&ݕhLC~Lɧ��N1`�cI�	M!�m.RL��O��+����ٺ��l)��1�n# �_Km2@���B�����(��MCű��%�픜�3�v1�h�g�Ĉ���>k�Rb�N��j��-�)E:/��G���H]� �����4߬��Wj<j�����a���F����b���?y�#�+qH��݌(���dF0fN�o?N�;j��1v:��S4A�1����q�11,%"��-�)<̎*�D/�����:��{d�	q�^w�N"�J�CBT�a�͜c� ����0�O���<�0��4@�����l�mӊR|���x�,6t���B��C�Ɩ�y5)#���*���=i_?�	u5\xM��U�� )<�~b�J��W1���l=�Z��A��*���`��G�G����dC�����f=�#R����dۙ�Mg��?/I@oj�ʘ�c����6疜���A�
٫E��V	F�ڑ$�F��ROaߎ�:x�K��틴�VT4g�N)��,��v�ɑ��zH}~d��1[��d2�Z�k��[R�[�Ԗ:l�[�*��9�PM�����U�%���Ͷ�8��8L����W糤� ��l,'��B-��G��R�P>ç-Kc��ei#�Ē$
M�8�mDK"Pz"��a8�޶u�c>Ʋ���r���
]b䜞"��v\�ڜ��5 ��2_���;���|BP�Cr����<ػ�ks��l[��OD&��ZW�h���X)1�!f���d����aa�8G��t7A/6mu�bD���ce�6*{?n�[	�I�Pg�1�j��T�+>�k�z������?�>r�i�����5/Kc���RQG����27~���8�u�=[<3	ӻ��n�7� �A0���G��#����Mb��``c�`��0���*i���i$�{ĹIt�����P1:u���˔M�_�`��?(C��9�,Y�x�`�s&m��w�i��n|�C:��.��i���'tzڒ���"f~�?#�`��I[�����86_�*�az�����09έ�7?Q��T���hW�3��K}����Ď/�~g��z��'ӭ����^���x���n��k��Ĺf�aѬ��5��D��}3��x?C/I�N���&L���L���ɏ�s������eg�4,��r��z��(f̛4Y��3�?>M/C�91�Pgy�%��u��XRlu|w �)���c��Q����r"Ƌ���	��K1>�F[j7��٘݇d��`$RL0����(�ak�	3����N''�%��TGꆬ�kjj<#�κvг���@*����>+�@�P�j��e�����i�a���pQ��$3��$��������Rc?E��I	X���}�����
�ȢĪ���B*�D�!zjJ���9�@,S6$�7�Ж����pW3���w^���x_��_��w��SJ��ߙӽr+������n9���pQ.�nK�Ò�4�� =Kn�6���F��w�ѪN�[ôep����d�eA�p��p(݋ �'y�r}�[-M�`�R0l���t��e�����I�z j�X�i�����Z��� �\��5��7�ӹ�㨎�SYQEmI��~&����G��NA�+�P��n $�!v.���@�o�����6�I��%+b�^�x�+�4����m�
#C�F���T��Aݪ�r�%帱|ƃ�7�h����3�md�����8���7;�}elB�	aQ~[�=������R��f�4��-,��fT��7���`C�	v��~/q��9�r�zYW��kɢ�7YӃQ{z���?��ҽ�>�.���k��zKS^<10���޾k-6�_��cdX���ynoK.�۱1`%� ,���a~�
!�����!tAX����=v��r�
����u)皔c甎J�m��i2����I)��!W���f�9��Z�ѵ1N���1�ę�B�Or/�Z��)\�j��pZ��6�lD���������K��&���;�,�#��ƻ�A�\��]�hCx�}�R<0F�b��Z��/�k=q��[�9Z���*�gA^���o�xenޛ�=�)�����H��f]����}��Jc Ao(�<��.�NY�W�߸��dݻr����ޙ�4��k:h02�v�qm7�'�B(�\�����3��Mi(w��
��Vg�b��rP�~���-y?����m�ik��
��9�gW���q���W �		��L*!��
����Z���;��C-e�����¶��CP�{ٳc�oX0�0�z��Oٻ]�<d�3x�W�7NL�0W�u	}���B�[�Ξ=���8��&�U�<�ӓ�u������xl��G����rMj��(Z���H>d3��N��뤆�c�O�`��K.�m3�4����n\kOs�J1U�����:W��z�-��-����_����O����V��a�]IM��@�����h�$^�e�J�`�{t��Ϙ!	2�4�Q�2� c�@n�73S_�T�_Y}�<�:��O�e�3+�6�2G�s���X���[K�q%����0��ϴ=�J0��@*�~`eX��+�J�H'י���cUC��)΂P����4�
]>*��6Y�HO�L��	x:3 ���U�0��=����8\	I,�G.]n�ž�d�;�tz���,57X�Wq��K=�0K
j厝��6��_#��� �^��;�F�Զ�l!���}$�^T4!ܯ��)Q�H��{�}	f�����-�9"����8�9�9K���/����}�H�Z��8P�:�%��iw o1�CMU�J'�;sy�>�j�Y` �wH+�4�*ד���7%q�6��<D@V����K�Etĭ�Sj��+2�#�v�]Z�ן�z�tH��!|5�_ن�c�@�{�������3�*�EՃ0�������)S~����.��s����L�B�O���EB1��xn�|����0�d2��3����s��|� �|�����^�ZU�J4A���{Ge���k��]5�oFo����(@���R@rJ��;�agi�����G���%�͜�n�����[�j���Y���8������UI�غj�c�o���V4�8���o6����߼�|�á����WPG� &A.~��|{��+�ܸ��o�sc�(�V�B����
�r��SCy�Q/��G�,Ly�{I���N5"�FS��Co�1'NA�Ԋ)}-׃0�L��5�C�{�/b����h�Ғ�Y^�~�!z�z�;ACݚ��؏�u�� �3?�a��f���o<x�%�I^2��W�z�F*���K-s�5��������8c��Lۑ���34Ov���f��+w}n�Zr.�,mT �奫�C.��k�,G��r�>;��I>B4�ŋ�eG�u��s���v�OgP�����iI�ć�z�{�s|P@
5�k0�~��8 �Lx�|����h�i%��p���nR��uƔ�:�-s�W�x��pD:	�.���\#e+7�Q��9Uc���P�w��K��[������d#�);gVEe�����A�2�ޜ��0�g�;P���e�-�JAr���c��E�E>Y�X���j�lߋ��!tˮ��?>�h�զ�>O��ˌW���gY��P�RF��[KR�m'm�WL��RFA���kQ^���������p�hr�
��	��t�N����{�L<W38��ۊ*-|ؤzR�
@̣D;��&��yұ6�v�F�;N8�}U���.B��~��E�@+��f"�w5�z�C�NE5��\e�B�_����*�,�:��>T�MJ���h O��'Z�Zw.'8X���Q�����i�GnC���33Fk� p�������yJ=zN;h��B1�*ݣ� ���=�0��;�k�B���/PHEC��i���~��vM�h(��Lx��E���k{z��r���k3�KCX,ˣ��bO�u�o��.��u4j?y�@�6�~%��'<Կ���nU�1-�P"�����L+��ߐ��	_+P���p�cy�Ǉy����������m��g���HwNoA�o��μ��{�4օ���`tDS�6���mE��ߋ���0�$�wLQ�R: ��.����p�|֩�~W���,����J`���aa;�i��<o>�{�S6�[���ݕ@�¸H�"���H�c�AJll�x��Y|%��"�\����;6w�T�ZdW�X�=6�B�%F�I~���kqi�!L�$r��q��A6��>��H��@1'�XC�4̑D���cF�:PG]5���&�ܭu�5hs�R�5��++�)f����FU,a���'�����[�k����2eb��vg����7ʎ
[�x����x/F�į�Ἇ����f��"��ݷ>��خ�!^K|����]�hRr�Ѫ�ay�֌\x䦕�%�;���;��ϯZ/���w0����d���x�������]�}��9���T0>�8#� ������~��2���Y�C�i&L��U��.��;�c�^ȼ�s��q�d�%m��r��n���&@m�ѐ�\$x�FLJ�}q���ʆ�?�5�]��Z�S_�L�� �#'���&��2��u�4p���ĲIY:6](��9fw�[_���N��k�H=��^�Q�s3��1&WIn%�i�P;�9F5�+/{��7��UC�J>��mK�1/H`���S�7���%8�� �Ѱ��u(1�*�E!��P����g�G//1"Z�	N����m�]"��J+��%�����RٹNy �`v��b7�M��A�^^6N=��Y}�l��ۅ�;���ʎ���#�V�n�h��>t�%�e� 4X�����[v��dX�W�I��|��z���K�J�K�U�3�s>J��<�u:���@w�+;�8���<�w>P�l��a�N~�&�]���|�<�\���[i��� %�>Ʉ-��#+�P{��qxhȺ�IL� ��d�\-�E��d�����V�ZgPmj����v��pUw��p�8D��DDu�1!���3�]��i-�[]x]t�t��l�7�#F�C3���5���#nb!B]��m�RPa�h��znrN���Jt�]��3�����E����CS�	A$݌��e~��AVAm�2'4�5#�J/�:���+�C1�/��7޴�,����锣�#�1yz,�ͫR$�[4�e�nl��ʧ/���.؇��A��]�d�@q��Yg��jЦV5).�,��cO���8}�4X%]	;�&�q�N�t ̵��w;n��]<�*�ޛk�A�F��>Wj��D�	_����͝�L{*�LmQR��ɃVY�A�z��@:���9�)`���K3̒�� �CJeZJ��>>%�=c��B��%��̐t%L^�M���*W�F �����J�1,���μ2�\o�~�BM���d�c"���}�� �A�p��������b�>�1�by�������yǌ����&SpsF���0qS"�R�a�3㚐�k��;p��e܎�������Aeʆ>vw�Ƒ�m�g��)�`0�0v�Ɩ�
�~5�E���e������ ���\��0��k�'��܏b����~z*L�!;�7,R�t<©�V���nJ@�:��n�K�!=2(X��(�_D�gV�;si��Pw�骶�xĢq{�tu*�m��F!����]���	A������A���0ǜ��y���Gb枥!���O��#R�S�i��M�(+�ӡ6LY���������>��a�
��6��q_�!��Td���|����J��� E�j��Ё�+ψm�Գ}_��ƞM�!�L�"��Q90l�D[ȣZ�d:��@cz<���St�1O)��߼��0��k�E2(ZdG!�g;:���K8�þ��y:�=�(K�){B������|����+�#��]�LXpX����뒛�`ch�%�����!	���׸GUiTk�~t y�D`]�CZ_�`�v!�NIV7#-��?Vp7;E���$"5Mu�S1�sܓ�8�Jz7+g�?pe�h_��.�4����&���HL�@���$h1�^��������S0�<;����U��o>F�B�֪'�-����W�a�kuG�5�A��N�?.�A����6��KYF�#W�&�%���h.��U��y&i�����P��b�� �'����ܕQ�W�@k���K�?U�m��q,cɼ;Wz�u���"��%��ʼv#�n�na<z#� �UhI���ԵѠ�1�
�,8��A[�g�������ZIKΈ���p��t1���ڃ�h#���{;��x�Qk���xk '���2^���
�Y O^���-&p��������a�E��b$z�1�) �7@Y����B����R�6�A�9*O���0?��Z�{jŵ�g�-�������)���`���d����q�����J�ի��'���k��61��|h���X�w�9��b�Z��q�p�$������8X	Q�XJ}����TltIa*8�)u��0Ł��<����1�s�N|_?��3wڮ�mx�ay������`r����sd���O��1|vZ���J�'���&K�����W�rr"�djkl�Z���Lv�u�&�eb��Q�\�N����>C��5��:�I�D�u��^��Y�j{�W[��݄��)ޙ#�Z�{xE8�ć!{Fd��X_k�:�A,:i����zt��h��X�i��(S��713�������CH<	�h�:�^j	`i#^V*\.Li�+�v5?���a�	��aYm�Բ&٫nTӴhcS2��M��`��8���in�?l�V˴t/=N�|��3EjF+���E�TsF7xv�ʕ4h}��ZK�E�w�wt��q'�!>o?��G�y���=)�����8tӍb���-5�$���s��_+����{�ߪ��Z�j�#T.f7=�m�~������3YÛ�@����3??Qֶ�Ĝ` `��A��]�ұ��ɉ�����������M��� $�nxm��oP���W0�����eY*��eU3�������������lV��7��|+�wA�J溇)P���v��%�}�f�I�cμ(�b�1#����h;]u�7�?Ƚ*�����K�3e�~�B�<v�'��ل��|�ٕp�~��F�v������%�4�e�v9��ЛA��j\�����}(�����6Vu�x�_:�P���������JԲ���+�a>�%.|�.ϥ��f�!.�GC���$61�5:� yΑG�b���������D֑���o�!Nx�.l��I�JT��� ��$��[O7�=3��������;�rD]G�:3���@Up����~�S&����}%�O�>�	��Nq���
���#r�JT�����ˋz�n�bV?+�_�i����h�=}���ׯ�%�)���9>��#puׯ?RW��E)	id�v�����W����[��#W��Q.�n�2'����\G�����
,�$JY��AQ=2��!B��l��G� �%���"u��*���6�N��]^d��ȱ�ߣ;��ҙ/�p�Q����)ݐ�	{щ�8�gr)R��aܸ�ڇ���3�-�b(,��V���n��Aa��{>�TQ�-Sϓ�i67�#|��+*SL��ׅ���iA� i�����U�u�7{7�צ�DA���\�u���M��0�q�oJQ�e�	�A4���� ��ø8a;?�x��,5ⓜ~�Rf��p��$5�	���ʘL�����F�����xm5�K��x�T�`���dc��X,[+ƌ��f��c�Cg_�s�Lp��[7d��D+��w�]3e�؃w�d�����}�o?��Ѐ�Z&�;���1n�v�)��*�L���<�H�$����"s����'t8���@�@��y�i��¤x�"չ���a�T��9�?�3P�&Of!�ۚ҈)�n�P���d��,�I L�=2C�v��S�kuȒG�)�e����%��<��N��;�dk�˿���w��;��� I��mQ���J)*ŐF���-�Rg��q��PJ:��
����ю�_Q+W�����}	�������Y��	����"jZJ�+�~���	쓆p�Jyn�������!2Ϝ��m\N�F�r �Wsm�F�.a0��s^3x懈Kp�k[�m�h�!@2�1s,�%L�Љ9xK`��� m_q;���J� f��N����b	���[^f�q*�W�`�B�b������ycɰ��ru�����dpP�%�mt� �t*����zt�tN�m`u�=�Z��Ws=�M�,Jg�}[�L����������z��6������²ͱ���E���@,���xn�)�x7�}̑)] p ԧkp~B��FݶO"L_
��=DsxC0�x�a2D.����7����7b>&En��8�sHP�'{dy���)PC��mk􋡠JC���򊍋g$<sj�K��$ӹr煼P���`�"S5�й>_4.G?�d��ex@k����xޖ`��!�:q�L�k;~�%ِ�:�; 1����Ý�MT���L&��sjE�ǝh�?���]p� �-c
�&yCɪe,�p���TR��a*��=���D���;�g�<�,�-��Yu�5�:P�Y�S����0}Q���fw�H�b�f�l�/�	aY� kE��'��7������])�r�٧ t�R��[�L>؊�տR�Y`��a�Ƿ/7w�!_΋S��V��M�k���@Oм_�	M��w2b�}�Gi��� E���ƾ�]%��l��~�oy��2�7��%H��щ0�H1�cVP|ℾ+fl�=z�R��wv�]��$R���BM��'S��#��%��E�	��"0.8�X�6v��.�m qD0^5K�%��-%e5�J�wk�Wi�C#o w~�rg�>j�̝m�b�?�V�Q@"̒������[M�����@l2gJ��vn�$��(arN?}2h���0���A�օF�gF��K����e_�P������SѺ�]��� ^��4����5V����9�x2S�f��Ik|��z�ɵV�e}>W� �lj��p�b#�L� ���\�$-yJ�����׊��}�"��uU�H&7�J�d@.ZQU]uV���S�Ӆ!f�-H�\�T{�:'r����`�E�
%�W	2��"H�׈�Q@��R,(n9w�H�Lەb�C�Gb1Bpv�-.��-M	ܰ,�A(�D�'���n8����"���X
'��M���gw�A��,�K��blE��b�$SZ+�-���jZ.�B��n]-+D�^q�;��`���S���\�r�;k��B�ꀪ0V��߾OI���>�|y��N���1Of_��"q�1˙���m\�T]�܇��E�D�WX�K���ܶ�2��dV�B�҅y�lcy���8�Oz���P�j�]~�A�FYf��ķ���)&wǇUU�[��N_�}M_����~�L��������a^�Jj7V=�씝!����𢩻P��]�yD�$<:\����9�i�eQ(��oѥbZ��2\o�bu�	� n�"0�юs:���EEw�f�;�ҹ�]�kL�=���O�Q:nC�m<K��  ����i3G��
�����H�Ezn��;���ֵW_"�+�٤q��g�|�e��5L2��ѧ0g�1�4����s���
$����C�!��H�GK���v�H�J�Γ���f��j��̏K�`�q0� �,'8^��Y)k��a�=�@zd��~J�\�m�C�g�d�1��b��R=�����6���=D`̸f�K/�<G���#4��xE�{g�s�0�Lu	�[��Q��Ye��#�up߈V��AaSgi�y�7�����o�Cc���.Ĕ������E�du���a#@>?)�c����k�*�� 8�7����T�p�KH�X��p��oC�i_�[�<������$�p1Á��q �%鹵	�0fȹ�������1?�|�����N�a��:+�����EG,�Zش���H���˔����qT���E���]�6�K)�i�Φ��^��oD`fR�L��3�P�����&�=�B��s3v~%��쭮�9�_�B�}F�A�f�O��/1^eх��wqLn�P�S�5M[br����l5;+
�p�Ֆ���]�ݩ�������,�hi$s6�*�P�1Z��]�[6�[lE�1m�|3F|j�~����tHx��y��ǰ�v�	,C弈��S[?>��@��T�k��UGT7���`�b��h���\���_26q�5����5�YV��=�\E|������;<喌�ؐ�ۚK�����:T>3@��_1G�\�T,���*+'3,q���:�vx�NY�:7�{r�<Ыy�����(�aa���j[n����G��yl���jta`�������Ր��V�	j'?�m�_E٘�I6Y?��m���~�'�N��$s�$F��tp�t"F�9�(,�XT�%�&�Uq:�����FB��l�gGv���@�Y�t��Y��u
����s�,���|6-����5Y��&C���pey���.O�w%g:�1a���O���	��y�q�i�-BϠq�7��OT�x`EС�+׏�Ѧ��C�D�΅�S��]� �lC ������1j)}\ExP�S�	��Nkn�N�q��jՄf�c��&�a�c,���-�7}�1C���I�FqaMCT���Zr���Ak�kxϟS�C��Ji��"��#�ֽx`�e�A�_z�<��6b@��9������n�:򡹼��� �BŢ��<�g&��9R�dۢh���a�W����4�+����UsPq���N�R0ѻ8�l�m��QƼ6y<mUn2C�GԞE ��\�ǘ��}�;�zn�a�
f�_Q�}8vP�)����R�7�ȴ�VRֵ���1hGc�4"uF��4�9^���j򐅭�F��w�����Wz{��O���O�S��S���W[�ڥd�P?e����Ļ#"��]g�b�&'oY $��.�C#7�hX_1�x$U ����^�'.:���L<�ڽ��:�vFe&t�y aL�+͋���m�̟�$?8j|���]�_U��\m��I{P�Q��7�s�?��[�S���$a."d?@z���d}ʚ$�\v�Q��K��0v���ntP�L�Y�΄r��>ul�)\i��"��p�5��W���n�S��xý�`�	f`$��ЧX��X((�e�������E��}F�	�z�/T���}�6 �H��Y�R�KP�;�,�*��X���عzO����I�e=���X^�F��$�)_S�����՝xz���o2��-�㣯�.�⣉����r�i���6���D��Pr�u�na[\.U>��)&/Q�^-�&t��Y[T�J�&bD3���!�p�)�q������	��(���{�JL��O%n�Yx'�3MՐ�"�"�Ii:������U�v� A�c��l)�	����y4��Q�_HY��C/�+}�����N6�=?h�x:r�3�gNH#:���{@U-�X�ύEC����b]a�DC��;zar�:�C2G�-W�z���]c��9&tu`g~!��0����ϴ����1M�%�x?'L�۰��6}�@��6+��09\��pj�h�b*t��"�?1෠�T�����{����5e�����*z�S�ڞ�Y�`�]���Ҏ �� �����I������Y�3Y����j�<��-��L|�nK����rbv�&�ĸL�[�Q{T�����I�N@�c~�j�T��mk>�=_�����G�"q����! ���Tꂺ�"�j�$W����XuMZ�zVE
�@��=��m-h�k�v���^G�k6���Is���¼k���~}ř&^9Ӡ�#2���<re������aͫf'Mf�}�i0�A�sR�+ŧ��ۗ�z�*�ݜ����tr�]1 �I-�7)��M��}�Nl\�)���#������}-�O\�ٙ>��9�_Q�V*,�����-����B�}6ұ��hJ%B�8�����W��D��7�ޢD��;B���6���1���A	"��*l���'�%,e�֦d61��_gl���3�۶�(Z
�m� j�z�����H3�di��Xi�~A�Q�sҺU$����iD5��h'd<zt�>]R�oɯS�J�� ��|�x�~�ے�
^�:���$*��zd�.\V�y�X���ycw��ɂR{?Ds�iQ�C��,���I48����d�8���H4�7�Z��	�Տ}.�^��<x�����d1C�HE{Y��8��m!B�~�T�� E�iC�?���ݘ�S{� ��r�",_f��^��a�C������X ��"���-�,�d6ݓe��g�o����'i��?�G���)��%�s1�zdyRV[�̽$��h�{�?,#Z��_��Iy+�©��T}�����ߪV6|fl�:�\EԃR���ط$\!�����	h��i�4,�����l1�7��>�Ƈ�y�X8�]����Ri�8��ȿ�Hm�-�@K�Oﵖ,1���RY�(���g+��1z�G�~�a_��R6�\l��qt�F�\��[��U�$�\g�a����m�],��ʻF��7/�Z]���
0�(���Ev������ɹ�A���W�2{�]�e��\�2,[�уF�=��2��������9��wgB��?w�6BX'�OP��^M��DF_@]ˋ�*��UL5`k9�lfh�H{T^���Ni�|UǸ�e,ƥדs��h%��>���8N7k�W"���8�u�V�(��+�B���9��V�,�x�.��,����$��Y�X��f]�n�Z]j]p|�d�;V�7����Y���ID��7���i�;�q����74u�]&��<�Y[����UCX��8�CH���~f'�Ou�mK���n&�N�@�ƌ>Tu����*��0��?���q���,%��ڠm2(4���'�{�i�D�d��(p�_!�>��7����e��g0h�#S��%ۯt�����n�d�ʽ|�,��Hj�s
�y��H�lWw��(SGt�C"yy���/-�*��D �^���b��pY�x�z�G�qEV�6؀Z|z��DZv+̯���
%���N�**�u�R��C�!�!��<��%}!�a�.oT�!���i����J1��=\��Ƿ� �[�.皢{�yx��s�F�ۤ}��aJVя��I�/��ųu&XA���-��ձ�`�8$��2O��2�~J����ozLo�R�y���I���A�y�ĨS���[W���	,�W�>�-��S����2½��uGɿ����FKH��uWr�f��3��Yc)�;�=�2ӌL�X �`�d,�)�j�#Uc�k�w^�ǡf��OǺ�I��QRa �<��zwU���o�J�l����e���TRL�\�g��e>"����� �& �s�6U���NtY����O��/��j���l�ʐ����� �s��(+=s]����}���������s6�7d6���L|^�F�����T�,�&s����W������n�]�^��q4��7��r9C�R�%���ꩭ[�`&?!*5���ͣ5�\�v;�-�j�Wr֖H?8�b�_���ݚO��o�Ůy�\|��u^�œy�z�&�k�7L_��#	�M��l[�H��@��Ʉd!C8,dJ���ˍ���'[��@�����/�� �ػI9�#Q/�=���!77	s��ʏ�c��C��������	�~��r�air�i��^t����T�Ӹ �B�K�5��9�n>����]9%�����䋽�<�	U=#�r��F�m:!	(�|j��Չ��3)���W�_o�u�Ӎ�M=N��y��-iwa����m��C����$;�L \��Z��U0b�w�#?��V��e�A�XI煆�z�DO�NDA�XG�ZOy�U󛖐�G�C��C��>0�R���1;$�Y��;�x��S�
����nt��!.t��I����\��û>�l�ܷȉO��5��簠C"�������j
��MF��}Y_�x�^J^�z�B=P��<��BOU������ܵ
O��,����+F�[�x�C�C��r.Q��e�4H�+@1"=�Ǳ�����gE�������g	�ʐ �Q���Z>g�Pj��W�g��)c'j�.+��K,�>��]��D�w��e�M1j��|�hG2X�
���B$"��*9a�)I���Ï�x�4�������:o*qч�Bvn^�7��	9a�۸H�SR�6�h0_��%�|�j�dg��D^DGr��.G3s���|	.V��$"��/ɔ����w!h��a��{�^e����	q����WG�E�jAņ�Us;Y>z���]�C��O�LN,���LfK�z�w��z}3���(q�e�y�08�`��.����8o�n��b����D��9��@��-�1����pR���b�KG$e��C�F�!Zq(�C+|'�΍��뛺vR��[��Cg��a��A����ʸ�\�c^3`^�9l_``��ח��� ]�WT��Tz;��|HzZ7�jZ)hŹb(��8�QE