��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.hP�r~Jzܣ�JK��`�ɼ�d@2���a5�m�1�*�i�)���LD���p<��s,� ����+�a�,�e�U�2?R��ӄM�Uc�{
,5p����nT�DV�N�v���9�ҟJ����zi.��|>�-F�� �tse=����0�bI�F�Fu7l�r���M0��n�kb�B�~KV�h>��4�H������{#��C 
dm[㘷���Ic�-Z�(�9/���u���w�v�f�z���)���X��&R���$&�~y�u[>�͡n�>�uC.{-@��� ���_E� �$�#���#�"[P��7�����k��;��}.ke�F�M��	����|tm�2�,,ig�IkQ�/�b��zxݫ��H"^&ZP��y�w�~��9�3H�����1D����I�%p�at���;w�����DH,�cT�D�P�;����k�D���:��_�tP�� Xhv�v��Iv��2��dv�S��I��'p��
�7_���4�ee�@�s_r�x$�������r����-� �^k#_d��Asܫf�W%doJ�*����> �"8�������G��k���"���G���fQ(�<$k��w.
�����y�5�΂-ԉ��?������"�T��h�!�P���ګ��ʫO$����D��L�pjJ������m�+ձ��|z����g�nYU�a�=�;JT섟 @�N�N=��؝��v��>�S2��pa�(�i����Rؚ"�;b(�$)��]H-w�i�%�-f˦ltIk.�+��HcW�-'��9�@y�Dv�1�X��I%�6�`�X>��?�r#�ڹM���P*��N��/�;bC�A�B򎜷����)XՈ	�;5��%'�$�[�C��Fz<�3��K�ߐ}C��e#�V|p�%��L4��[g�e�����Q��2D���8�Z��>_R����������p�dw���`p��i,(���;�a�����?��(�2K,�#��=�0lݘ�W�?��:�G�=W��L�!���,%a�]�0�5��L�/[.�_�%/&G e@,Cۖ�_Q�m_�s�RNXyH��d��+(܋�`���]gy��AD��,av���<�}��nO����T��+��%G��E��9��S�B�A��r�H����c��]�L�3�&���W��w��"��c0�g���-�l���~�W0�5L�3�=Ca�/��� ���P����6??���uۭ��!�Yw�/���2[�b$�Q����Y�e�t�?wo�1�Y����X,����S�yGЎ��h�2�����&�P@ѝ�B�哛Q�K���Td��)������~��z����r7	��"GJ"�9ϓq�Vbٶ���I�_]�rґ����D���z�s:�簷����*Մ��0�Lt������1=�#��g�6�
Ҏ����*�{��Wd:��+� �2�Z�PEĵ���(�%�e6��/d�hU�x}�ɮ���DcN��p{����!\��v�%��܏GGz���C`��e��"�Y7�T�$��%}��,$�\���c<,R� ˎ��r��E�.�:��Qپ��#�`�D]��mN��cB�?�)Q��~��`�����P�i$ ��&�&�(�U=4lIO���x}xW�S�CjT/?A��*�_t,�J�f�`�D��;,�*�j��q�BF>�d�m� y^9O,US�>K|�PL��LC�\�U�1q3Lwތ��舧�(.ۮD�,T�6X�}=@.��?c�(O_�ߕ�NVkR�A8�|��"u!Һ��;#�]���]�P�NIa���� li�H)�b5���85�AE���$�I%��cZ���/��cXq5���u����s�fk�7��a+krZH�dZS��2��t�"�\L�Y�0�nb�0����G1ءb	2�Ư[��kO:��ɘ��j���.�N��Vdc�Vu� �9\��ч4����yr����Z�~��2]�3�Cow�c�g�Bj��4^�s~�qF��Dw组z�P[-�B7�Y���uw9]��E�S�-*'L�:����TOs�P%�B{1>�>��y��Deu� ^*��9X�4W/�cJ{*�aF�'/�G���R�yµG'&6��ā�n?j������A��>-_�Ё���U����y������J�L� `Uć:�;�T�-J���T��O�czF�~��=M�, :�T�}��m��L�_0�yK�3��劋�dˠPwJ�'Lm���Bo��xl2E�TY0_ظ�]Eb�7ZƤ|߃�!m��􁈂��$/�hO��ਖ਼���%����w��k-�9Z�C��5N8�m��p��N�$��K�s���\���;ؤ�̬b��0���MW�ʡMĕ�S{V�¿?�4��� ��/U靖��yB�G��H�= ǟl(Qs�G�G����'�h8�nv,�&O3b�sul��o좿
}b���j��Cy﷦���$��U�T��Ŵ1�sG��Y�|���LQi|���F��>ׇ��&限ퟝ����?|WnN�q���2,@Ȝ6_����9���5��A�T�$JG���OzLv�_�;�ƨ����T7�1�#U5  �<N�@ḓ��;�ޘ��T�׫[�A��-�uC(�Y�F����jFA��BN����R �ҏ�Q��iq�>:;��*��$�!�b�|�.۽bˬ_1��sJ��!�a\~�C�'j�`���s����}SI5���[U�NƷږ�u��� �`x\�Q��d?���/����eL}L@��f�o*I�]����yB��H4�Fޒ�����OM�U�9�؍�Bc�ĈC�;=���_{���&FNF���u%�3�Gs�x�@�&�X��qJ ���)���>�pd���~n�?k6!U����	?#�TϷ��/�L��c��v���ϭ)���Kg%	 ,Y?�.��ӓ��&��F�Fb��g"���tb���>��J=�$1��!б��XI��� �PC]?�6?�9��d���X�XJTءj�ĸ(ic�]t��\��⌸{�	2)<�Y׎>N8=!i��5�A�ӭ7�\�c�0,��P�P��/.�ދ�̾�L��Px '�އGL��=�j�Jc)��#s��]�0F;h;�����k�y3��Ŝ��?����2�p���1B/��!,m� oS�";^���h��1�Z_En�+΂-:w��S�и�b����.�]�詙��5ԮIrݟ�?�/�
F�N��&�oS�D��V.L�?��ۺ�Z26x(��*\�yt�:�*ڢ���t��e�BUAP��<�j+J����M�K�<z��V]���*��h#&�m5<o�dF?�
^�ey783�Q@�H�~g��HN��  ���"���ŵ���
�d7
 ���0Z?�6$��Yy�Wn�M�=�^7�.lDӓ�#���3z)�9�����:N�x@~��O/�mE[?�h���ف�<��r�LSK򜝕����V7�Z�2�+����R��5	]���֐G��F��@ټE��վ�b�4YX�����l�K���W0?�8���4G�G��%���=�U3�|G���@��B��޺��x�@�q4v��Q�<�{�H&�q��"h�[�0��?bг�E�;�,�#�{V���)�gL�6�"��H��q*UC��rB�Up����A!��w�B2�BK� >�~�2Z�m�My�1���̂�V;@�%yj�AN��fR���!\7�DJ u�v/�b~�	���8$+�M�Zx<#k�$�L4]�B⬍����e��� x��ޞ�'Ha�Yq��&��H ��}k.��A�$��:?���#�p��aZ�`��Uw�+��uh�(��2�%�\\��Xw���o=�H��dI� h�$�OI���õu�b��������*ۊh����%��ׅ<��w��M�fN���.�(�}�3�Q�8 yl��V3ۅ����,H%�LTb��X�UR?���ӂg^߇��s��Y����rYXW;+v��Ǿj�J��̨�|���?�ي:(����>ӕH+��G�+�$/x�g��\XwfU���B[���D:p0�iÈ7��4���חB��u�b.�A'E�LD���TVOq��nƼ��y���	�n���$�XO��������\3!E�t�CǗ�C���t/-2�xgxs��S=4�z#�ZW���K�rX�,B/�cØ�C8�K��O�6��������jXL)�����@�i^F��!�6UM)�s��x2ϥ
y�p���w{/��<[uH�R1ifU�����լ]�����Bd��Ϗ�5*f
 r+�
sM�[�q���N	�Ǿ4�5j�Gf:v�KkmV����v&aC��R��U��{+h� ��.o�Uj�����`2�`�-C���6�%C��UE���M�{_�P=ى�%|�d���?����yE7~��1i����)c���f�(�@���t6�G8U��"�b���m���� t����m��:h��CU���Æ��0c��,��6����IVV��o��M�n�/��k��q�y�����R�ˉ3b]X�����!���J���F����﫪�%4�:5J��$I��I`�ҏ��5�T�9���ʹ�u���ᘽ{�۵��\Z�������BƠJ��Ŋ��!�h�'q)�a?8�F����IYٕ�LuC�L�P � FU�d��T��X�/�P�j��c��V���K�x_��JЪ9��![X} 7���(�G��X{@r��LV}j+�&J��Ņe4�1v�2����Tfy�,W����p�5��]s���/�H��M���}2�q'
��"��ωy�9�T��*�7)N��>ꆪ����	��'���j#ɔQK!���cLOz'�딖���:ˌn/J�*t��$=����`��k�5un��)-����+�k?��x
3>O������ۇ�K�V��Zv+i��Т���mTx&G���(8���n��K��ȯc��I��#���Ǹ 7��zm��2�P�R
��}*\|Ԋ�՟�!{"E�{��Dm}I�3�,�±���]�M�|��C/�l��"f���6��I1�9���k�O�fp���ޒ/�={D#C�ؓn�5�-�u#�*��.�e&� �;�]�E�dW�L<>yq��K��E�8�,y���'��Qh�*�G���~��i�i��R���҂iOL.�)
��f�ӂ�!@2;V�*� �m�0��ܮ0��V4��I�H'푁�du��ވ�Tg��-?ş�8G=dv�(���c�<.iF��:H=�D���G:�Pj�Z�5hΉ}��6`@���g�\+����Q0�,jn03�Кs�i�yzz�Z��'���*O{�r�M0G��]e<fX눕�|^;E��n��&y��VԨ�#���Cm�C��Q����-�F[7��j�y�y��0���!�� zb��t�puAԽ��`lR|��]��V�+��dA8�B�����2�u���&��&C��)U,�tP~�z�!��&��b�(�,W�P����$70�q¾?��9�b�ɶ���x ���}S��5�І���{���[5�.�u�Jj�ƬSj�5�W2BQ��}�v*<��<�`��M�U�,�&�:�H[�Py���b�o?ˌSH��F�}��؛,�1+Ȑ~c�.a[��(�@G��iJ��FV#��lH��C�s�v'i:m>��?����>�¡�%�������]��p��#�����C�<j�Ѩ+��L��<�g���������,q#̒:����^� d��XX	qTM�{�]���C�#Rx���k&�j������2�}�T��GyI2��U�v���yy�Cb%�f�(��#Ө�!/���(w�}����U��!�Ѕ��fg���#8��Y�I����m@,��Pb�J��h���
4����Z�\��^��x���ߏ)�$y��A�4�>3ĎQ!8oM]�Jf������ 1���`&�k�C#����2�Uͅ�%�=$�wŘg�:�[��(����_�v��u����r�b�|}LaU{��Qc{ˡ�K¤�g��%��`�j}�_:`� �=IT ���v��2�����QU̮�֩�1�g�sb�FbVU�x���Mfx�0���J���p@&�(��|��_�?���B�x��L��˕'�qT)�s�Y������FS�$A��1T�k�&�[f���>����T��n-��W�7Z��������2���s�a?�Gk]�����$��*�B]L]�nog̙�?4iL�~�N�U�����jv%_��A�;XQfh��Bك+�77� �='땸�_%Φ�>�y!L�V1�d���H!��D'�����o'����^��Gن��ږ��<Y�*����X� ��R�{�HB��A|�g�io�����.9a\# ��[�8��e���	�*V��=�J)���{f����3�ߌ�̠>���h�6Q�p�ۧDG�9���IU^��>OX�ƣ-�
�ٔ{��$ڥ�Ȭ)���|��yR,�`Ȓ�C����}�Y�ua��"�*���H�ϧ��:D���Eξ��߼Q[=I��;lK����o^r��<���Y4��ǃ{�1��W��a
$�'�"�������㘥]ˍOo�Gf:��d0