��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�g�s���nGФ�y�$7��J;�a����d�x7JA��9*����|�Vb��`�F-�D�/��nB8��ʾ(Bv^o�����Ū7���w%�8
&����g�;��F/�k�ShPd	�����r2�"pk�Ñ���
H���ݿ$u�,+��G$$,����ǔш搓�Yk�^�|��)?�\]���1�ϡ��t�	������.�[!�a�M*�������c;3��ȓ2�k#�2�`��wC<�;��������i��C�UIgf�E@��E�y�J�F"o�(�_�'���+*�[zM��jH�u̼
!y>�N�
p�)Er�J�A�s
�`q��B��d���;����'X�g�d��+}gS]�-1�ou�mHm/��L�L�8si�VM���|���Iף���tr���~ �V	��n�Ғ�E	a�;�^���� �f����kW5Č�ۧ��.�8e�P[ZVr��M+���))U};� &�F@��4�4n�	�����v�3��F�VE$�yޫ���J��G����z����j���*�A��=�[^���{�b����"9��ja	�&���7=�q�A�t@-�bE�f	�<>M�ŷ5q�)|ݰ���2WS�� ��7ϯ2��Ak]~y`Ni��n�s���>��b��e�V.4D'ב[��L�����.�	�X���Ly7�Z�BQ��P���-�6E���/ÿ8�?(}o����FF`0�?�lj���fG�����ʍ�"� ��hv؃��TF�f:��{Ns�s���[;�������|y.���
�T���g���M�r�	���g�HZ�PM=��I/�1�r8����y�ZP�R�����!0�3K�b��R����i`�ҸG/�QN��w�C�-e������.��%�%�M"!�%W��1��$�\IX(��C�|���FZ�;�K
C�A�0�K6�8.��,&[2�J�Za�&�b���F�{󳫆�3/�m�����o�0IO��J��ne��P�?��&k�-r�������S���^80���1Q�ေ�����+G���%��IN暁`J��+�� �N�a��F��E]��8n����YU�#�_��.�0�6��uWvþ��+��ydԓ'���H{Y�A�� y�b
Kv�H]��}W�!k2vë2��6{�PXX�Qbb��2�V)����FB�q	��0p�����o�njt0�¼n�x4p�.Z�T����e,���<�Bw7��6}��L�!]�fi�\~�G��aȗ�4��$ѻ�����~����~�VD����[�Dﻸ*x8�!2���>ʪ���WGދ�v�����%Y1�yT���5��'#��$\3���E���Q(�6�?X\��PTO�i�����1�%�� �q/k�a���MA�롸��`�y�b_U�3�~��.im{���&q�إoMw��'���ݿ�O���Yg��p�,�+�F��IdٛNyF��ЇH���wj��-�8{��q
����;�~�ͱ��@����I� �OM�o{C�i����h½�}�m�3�<  ���r����!q2������'��6BWd D��d������/��!���|�D�r���(x����V������_�^Jҹ�ԉ�x�s��чǿ���)��?0b�|��?/O?�H}[<�)Kl�.v{^Hʱl��J��7߰�:�C���Z-���u~�����~q�:q�w���k��.�ǳY����C>�]�FQ`� Ks��ῷ��tl�n�Ҕd��8�;�G��DlJQ3��Jw����a4�PJk�n,�RR3N�SU]3��˨�e�2T�ׄ_��&ᄟ����J�	�s��m��d&P�*D�p:�& W�V|� ?�����Sq����X�K�J��*1>�k��x.��<b*+�\��D��1�NԞ7"�,�^���[J�l��Ӛ�TlP2���9���u�~F��#�T1��>P��a:�؅�Ŝ��-!Xh�5nU�t4�,m�YA�mۤZ��)_����Ǐ�d���x�wLg�XV_Ty��Nт��&�Y�e��@͘���5ꉐ�h��n��sɑ�%m�4��hgb���d_|�c�!{�r�c]��V�<��E��D��_i��RՕ�G����L��U�
1����|_��˜��ݛK0�k&,�����N��3N!'�|���*�?'�I3��M����(�ݩB���	a���5~�����eI��;�Y;@pJ����"z�P��~Ȥ�[�F�L
3�	�wHU�2��@J��/$��Y4�ڔ���٬P�#���z�c�m��4j�:��26�9.�-�Cv�y�Aݹ��o�7�*U1ɳ�t�,�2p��д��G�'Q��BJ% ����^u��;Z�i,e���O�����>�K��!�*�S�	V�����U\���­3Ca�M��\ꠖ��-t�V�m��?�e>;�Kg]���7H��р+񷉶�p��y��`䳠��J�Ċ��j|%��i
B���.��U� eUZB�� ?��Ԗ�^˞ё�w�o��[:n#˼l���8>�zjz�T� Xg�%{����M��L �K����F���SJ�]�Yj��m�\0#�L'�m��H�r�e���-<�}�)��oR���{�0k�w��AvA	�s����"BT)n��
~:����rV�OS]O��N**��s0�|e�j]�}��q{1�Pe1���E>�!Ic�V7��qY�#\[�0��oAx�Ľ[u�����(�<
���� ��r����]���݀��[A�X� �����,��;���.�o{(N�GJ�ΒO���}� �$i�2~˅_���Pj��'�e����͙�T_G�|mު��.��c���/��@0�~*߸���h6�ߐ����?���S�y�DȒ�%�%3<��H�HS6_�tE�$ᡥG�
��_T�1C�����C�Ai?�	��ф�O`4�(�b��f��'�!a?D�>Q5"k~2�٬O._�?km�[Zz��9�גK��v���lh}J����Q^�D=ǋ����+�a������!�%�~夕��^rHy44򙝩Y�-�'t� �6m���*̻���̓��L/_�����LZMY*�8�Q���'��>��J��u$�v�K���3��'>p���o�r��3��~���8� ^���n�sh��p��l=����F�%1�L����ڮ��8b"Ytl_.��>�@�S*	p�=Z�XD6��]�k�a��6��'�Q��o�Gnv���HK�,��ź�T�w���LP��}*x�l��������%6��Vns �f�:d'�8,��W�
�69k�w9�H�Oo��\�i�j� 0��0[Y�W?���8%/R�_sQªXG^���gp��5&y����Չ���ۇY#� #���߶��u�H�;32v��[����8���)�X,�K��� kd���0O��e��pI�e�o�������|�i���$˗�Qv 	;Zj�EdÑ䫧�+�����b4�]j�O���Ed�m2\�w�/5� Y�������4g�3f���~l�#Q�5*���6�	�Ii��aB�����D�4��w���!ܒ�x�}��pM<ˁ�Lj�r&�^�Y����b�4�O���9�aC��d5�n��)�͉�-��ogWJ�%��Oq�oj��fʭ����՗w�n?>�KY$i�Bs+��M�{�q���f�c����&�s�C�����Y��\��Nx!�1'�PK5�����!��0�5uw!���H�s��_�f`�_*��J� �|��G�߉D=��>\J�𶉄#����j��?��s��7
H��i��
�^��A�P7J�P��!��{���]�@��A�4r6&o������~��ǖ�5��EJ��zM)�[=s��{rV[��4o�h�H�7X�T��lٿ�Fs��&�&�.R$0�*��U��fy����Q�.����3#}����E��^�������μk-~�J��}8kZ�*	ݏ۳��4 �؋��=������'Z2�#!�On�(��pb:7h'�����1ЩE�`��+�^9#<�S�q��)̊�_'�}Eu����X!<�3&����5�B��6�����W���~%F���/�q���%����sA�o�wR�ł����y�dԂ�ҩ�Q�@!�K�éA��TD�0��c�gZ3eH�o��*�h3���'dN�i��6�I��p;��/�h�H��C^j�9@��<�啥��ѳ,�0h��Yo�ު�Z��1E>�|�6���9�-ar~=�g(m����!b��L
����jM9�a�ˣ1~��(���1[A�G�wh�y@����+���o����y7C><�9XeFr�8!�'J"T]������m��	TgO��*k�����YS��Z����|ge~����D��,� v&��B��
�p���<�i��ծ39Q3h{[&2�L��]�ǧ��� ���oR�_�%����a�}�Ě�n3��A�.uV�7f|�,zC#�Q�p���;/�&���l��
X�A�;:N���?��PH�E�n��
IBV����vN��Ai��J�^r���[&�kRl�W�����U�m�5���1k�4�u,3k���&�0a��2����F��er)
h�x�䋆Z/��J��;�?��%�ts�����D�c�s���M���|��!�
�<eq�n/���Bdr�莍�7�Nj���^-~x��s�8��?"J��:�oS�K�.-7]>#9{*ag��E��5�/�S5�?�%�!��M{F�D_~�����@>��~���-sK�w\���t�s�0I�k�=:^�2p��k�/>k�_�]-����!�{�����/��_�[�EM��������v������
�|�k�t�4Y��W��o�YA�j�z��\��ʸ5Ijq�9S00
7�f;�̸�"G��RH�lI��ӗu��
������<q�QPü�p![�u����Q
�U��$Z�1t��&s7 Y��p�� �\�~H~�TY�Y���{4���3.��:����G*h�����(�&�b��P���e��YU�y�h&a�V�; c���Q��l\K;Di�T������
<��j����EC�e
�I�N��@"[���	�{	ʳn�x��w�ґ@��ObY��L��^JЬ���b1��k/�^Z"{����q���ߓ5�뜆 _Y�ϓ�չ�wi�75'
#Th<��)˲��[�c���=,d���,��|��
K�wg��9 ,���8�p�V.����ꄏ#�Q�T�fφ[���F��-�W�d�f�3H�htT����N��e��_������.CšB�y����g94�������.����vv,�=%Fqw~1'�F��3n�1ٵ��_|`���<C�[2��絋t�:�sd�KP�ՙըSx>���KD����ѝ��P!�}P��H�j��˓L�P� /�$�O�G(��[�,G��r�#�"�>��^q*\f��H�������KMhvp� �9�;��E[P����?��'�����u�Y��o��J�b;�*h�*��#���f�B�:;ϲ�+�u�I��U�z��	�(?���o�!�x�ɵG��j%������3]d�0�&%��RY@pA�	��Jz��g��Ym�d�R'')�f��%���;)��_|�M#w��-��I]J2�0�5JKKF?Y���O'�%\�R3ϜJ�tdrT�5���>�,�Yn����4bj�N�hs=�����>� +帣�LF�&,��L�>�qX9<3-�;��=>J�0M���`xc���[~
��H(]�=��|�E�����̋P
��<��*Y҉N�C��V#�[B�I vϷ��I��$5�`�*l���	0/i��1a��.�"kQw�vD
H����ݤo��U�k����3��h�����Ӧ0 ���J��DL?�i�g;,���Ἆ��8�o��1��'A�䢚�{�Ud�^�t&���ܨ]4/������=r¼�,!-	��l?#�*�z���<�T|Iͩ�9�6)m��{.�K��<��`b�r<�������:�t<�� cI.����ٗҫŷ�EiEZO�iЬ B9U�-R���L	��)�D! 5l�n_9��L.a�C���3Y�;_�ԗ�ý���4�l�� +�tVH67M/dJ7P�Ӵ}IK������l�~�=Q���Wn&�����b��İ�ĉH������Ӿ��t7��Ս�FL#�NWx����`�X9).J�]6�h
K�  �2��u�F!�盎���i���� �?�������I����
jna*��%v�y�3cBʬ��-�B/H���Ê�8,`٤�<#�^evcw�jz�����w�8�� �	�L���/* ���_�`t���Z��?��;��H���O�ŅHR����31B��Dx	=��?b���`��4�L'�@5"��-��ꞈV��[�v�f5���Q����~�8-�����Q岓͐�&���p��ܟ�J�E�v��B4��p
�Ҋ�B�%>�^�K5��ݨ�%���R��Zh/��3�R?��\���Y��?���U�����*p���WE��WOR�c%���]��f@�^�@� ���uT,��c6���I���J�z��	�@�����6�Y��܀/�ʑ����Ñ��(�0˵MM]܅*N�'��eo�JR8��u�}��/��q�2�o��C��c<d��I�T���
+������K�K����ԫ�"*t�טi>�-�@�vo��Y�~��<�FNg�G�����<o���~�/}P�Aӣ�� �=Zb���r"��I˫E=��f���x��;MR�iGH�U���N���E��X�\��_R�������[Ö[�ĩ�0��#��;�Q! p0['�Ӹm3GM'e�g�=x�ꮯ�$C��2o�U��b�.�w����\��E� SܾCY��(c�lȳ5�ڃ8H�`��p��]�����/;%ڰr�T�,(0ڴ%X��ד*�ǰ���L��k�S37�
��7�r7�В�L��p!6����^Ua-��V&�zp�����nș��*��)F���aZT�o�<�pW�����f��p�-�����rZ�����h��D�!m*��:���-aJ1�_ A�ܟ�2�	ϙπέ$�`�
�_�E=0@r�LX��wP�P��ߔ�����TI�%��S+�O���2��xB[O0��i�:��k�ot\���\�m�I��6�ץ�7;Mh� ԫjk��7�y��CX���O �zK������R��.�?�Ӱ.V v�6����ޔ^_E2|#�E�6������Է�t�<�F�^�?i�mh2�"�΄���tv��V͡����k�u�k0�g��65���0�&1>����p��̌y�]��d�6�p�onߞg�7�?bX�IKP\��QT�;�(�3my |���S�+�/�i�T-*�M�T�ڼ��gy�ihH�)���s7(EZK�����=`ýG��6�x�O��!��a�LFe�P ��%|��t����bV����!Di��� D�88_}k��Z��#��kWi���ޓ�I}�"�$��� ���ϑ9�Q���tH�����B��<;��Ќ4�[�Z����"C�HKu��8e� �˶���`�R���Їe�g3��Hw�	��6��Y�-"���9H%��gh�ʁ˳���e�`�������f�
����شCn�7ۼ�9W�|^y���N���#��T�~�a$ne���Խ�q��'�V�l����`��X��/z��xn�l����i���@�&P�
��{�m�R������v��*���9��pxhA>� kKʥ���KQ���L1�����X�L��Q�mj�XN�{��>E h&��s�܍;y��wDȟ��{�h�GjU��)�'��|&j��W{�Iy��M4�P�g2m�??�2�dg(����bz��9��c�%g�I�>�o��