-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nX2C2vB+Wo4BYw1lscTYeG/4qveBht/NvZo0AUE8I+QfKlejSIA6zEeR/LHgZqtK6G4Qpim03YKh
YioTNihS2X9FIp0uU1mX8IGa2+UERngvuA/f7B0wxiXJMsqHLcq1egQwFzgEmwFlAj0+suBumP1x
hj3nYZfFIUMH7BSLbD4ITv63RXfnzEZccM0o+xyX45rXkvFTIRxxgIA8iKvJqQfPGV4lvtBG7HTx
JP/g25sLELNwWeMZ9nJ89g6dtXgSJErATAe5l4ze8LVKdtKlO7DJ5lHRza8RvTuMYKJgovpjiKA3
GSXCBJDYiWYpNJmXEoqV3aX2WYnc+I0ok77Y6w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
0wfky3Zt0Ztg8K8+4wQITKOdyeMV+bdPjsegMKUhMcmWH2ATZa4VWj/YA+QFXiXQ8717u/QliTSd
STcjJKzjn0LdnI+R+3B9Nm0m2JSF+z3ok6IZvRuulqGbHUfLYdx5lACReWd3d6SBoR40AOHQOSHw
MZYdmYb4U3U02s/wz8X7fCqwimkYSsMTWGiSkwOnxcxc6cpyv9uz8Xag8uIhucxTA6dHVgK6ns9w
YNe3JnBeyqCC8CD0haXQQ4BfdhkxAGNakO6YTgiIUb7F0HQlhqqyY0OnrjeecwpM/tHnVjl+yMRo
mjcMeRV3UYU1Y5Ccq/TV6wQyQaH7GZ/svbNtdtQXVC2n3RF49tOPlEpOnRnCtHhFghowAZXbzRUg
EvvreFTcFeq6OqNAgN3CLl4dipyRBL76Ch8pfvwwRHf6IxGnpdF+pcJcYPS02zUNbThRbXGAwSkF
OaLPTj2MHXaftVcfvQ2YN/tbdNEoGhKqLTwGmpJdoIW7l+gHEA6j2RrhXm/aMgEaDswqMS53mZdZ
Q7zDkbN+Xt2VpEgF/s5b6tGR7ASs2tmRDBFEcyHDcvZNtpNT3M6p0M7RvobjFC7bJMFZy3+fEUhV
uGLr/q+3+BWhYTUwAo/TRZCniXUNMVqjP4Yd9cFXZePHcpggNcFClxKtSpHdIbLyhQ5a5s42L8l3
tqc3i5s37nCJxT5K2HbUVffS+MLupbUE3l05o4fxlrRftmk+99+lRtttpdgUOh7S1HutIZ0vjvRn
qWz3dSJ3S/vRtrFpSv8ndi45kpEQTk15Kqq3rRS/RyMIA2Sw+Ih8b03M1gK1O7EB/XeUpDJkigGM
D9JjgRfPOseWTGdCVqByDsYhagzV0SGadXGMt45P0FUUlrHzlFgMenOrveH+yymE8CkW675fT9Hh
8FrGbpf2OcYZ4Me8jpEpTpVHmIQbW+1dhxkhvP6KTBMnNaycRF1Q10YrGPjfPking20ESNRGsdkv
jBM3+BhQCmHnBu9/jZciWqsYk7Eou/hZCxDWX2L05cQl1FxkQwPIAUVTrZAeHaNI1qPqaDjFluMT
1yeWyXKwqK0OkxMJv48cWcj0iGTnBdoaxV2Rs9ODFu3qlIFFP/gYDd1/NnbW2+vaXKVR8VeB+E69
K9AYElhUlTNAaKfbAvcrLw/ykJTeLPQdc4+BWSXO7npauU+HM1qCW9FxRXuonOwAtOPZYM+MvJDT
EqWBoEFYvtuVHcQJF85C8kzKZ4oMIxFDl38XRY5Bd0MgqyM4Rdhsw36cNSLpshC4LLaxnGFuKeVu
OzdlsBF1sj0MKNs7J4Yhy1Ypbvvj/GNIaFn6+KNHJo7y0yra1oGroFwfM/Srz8OFCEjftQfVw+b8
LvGvYXNjus6TtP8dRegREdZKHbJzixcdq5n8KC/58+QfRhybc6gTy+oyUv9QhVZCHzuxMf73EBmS
t230BdzfaqUqrdvFCC/H1ufXI447yGDv3T2eFGOC05EQnOjVn9hEGSNmggJOcVb8nGv58EEqkxxF
NsQ0iXMj2e5uLjU3N1sEpNwLAjw5dJTP0MCtmC1yetj0C7qK38sbYhKhLZQlqCXJEcJNbC4O/ZzK
SBo9GUf6v/l9/VBJXDwjt1rnHL0hPNWm+BD/vzS04vXMMyCkzu6bEzX4z/1O8yVUmkoKhBhuvsMy
H7w3v4AdYi+W0wSzmapn+7Wnzzi92l3ktw6Z2qdoa3TtuCajaCV4o7aSs6U2p9gdWAnyJqzjyFdM
dJFeiOQmUT5Ltk+pg812iK6YVGCjF53q8xPn80B5AcgxsIG93Y4x1pwoceO9oXQTcVzVU+8eXDRG
pSFJGhEYQikIhu9kIK80J17jgw8Kt/i31CAP1e8h/XQbCQA5zZ3B7sQJXt/VaovEJMaBwF6k+1gs
cmZp634Uf+ezopAFIveDygBWPWXxPXtLGY4XcEeTfCJBOFj6Tn6+l2Z9Yr2GEGwsF9De1lmW3qE1
j2bmVjbbgpeSutzfjBrNPRp+mJJpLB91wffeU1vdAm0y4MQgBAboGcpfHG0LRwJHVSlk9dzBEEgw
8Bgop4lwB6Fxp2aZxRgN6sx8VuSLlHbRy+KbV0tlmuhb8JCgB+1dAL54rfj5yz6FUfHiaKY4TvHN
swFhhP149u8llkoBhJG2xgpkUPprmdKcMQ3hKjr9lYxzLCOdt2KufkyDXJQhS2/YiQF/fawyWrAN
mPKIKU80NXUbnFEY2yxuz/pa2F/w2ZP4rCweHFB+gXUmcKTqeqs/FkbQY4L8fuP+v3KzFxwfeUho
0ErL58SBjxUMIazYVur7nKoeMGjKKStxgQbzbJC8igVXXpzElvWJ0a42NIOZGceNWT9+1n7Uinlv
pmMbR1ejLpUFfmCt3ezUf4wTQRtWLzZa9i3spuB0vEMIrXZtD84mORZE3IMEQrdr/pbilvQeCzma
RCIOB++dXXKNpLdwdTE5ixLZHs63CjCErCUDvCbcArq37pkxHpoN3HsIurMTzLbNL/hA/TFsMUeB
1kdbo3xIIBw/bGKLTyYGseVppLNQknKeqRVPGY8PyaXvw+/cU/VpLlGlL3xus3P7OQcjPGTqIVVZ
/nANLcgcOaJtSECiKQxEq4RmfcMpGVcJXCifvO/OrBam8ffG6aEObdCKgg4oqMoPDkwShdCqTV/C
MbpPPGdK6eqLnHhDQCLq4WvGsEtw0nEif1EB2jtA97FZZBgsQyU83WapbqDSQOCiwW9wNqkJdSEX
+yyPvLozl4jTMz6y4wSq/jlXOH1ZaiFZpWS8tVv57lF4LmZGDCZ4c4JoT/ATzXEVkaFc7blkvqug
GIcWZCp92pGh35hFh2Wp00Sgaywfs86s6OMuCFmqY+LNYHfaRee6t4SZFCxstLWdz6aDhb6D7Tz5
vgwNITTXNJk/v/rzeBWna3LesYwLf8v125o/763hiTAa1yIu8l94BEupGuub43wA9PFf+Az586vk
hjX7bMEDOfuHP5F2E9XVreTD9VQpbt7PZyq+NgnbrkFZ6UhxwZnEOtsbANjGwQtYy4mgArdrwaD7
kGhov8ltn4il04k50lesyqAaFdiN1oIQoHvJ0ZZPAtD9jG0nzgDh0LoLlAqtRzR5itF3/gvsHoXx
w1jDI9QMcp7gHQqH6j7fBEe9KKJ1Zvu193OlD/ZNZyIJPeTmkfvK2/nJhwtNUXE5FOKwmY+3RUNA
Lve00Ie0pEj5/GOsND6oJ8K2z5yPV81ouoG3cAwWD0qv08buyxy9r8H35lLPurkHKsGIrXitTH7h
qgoxWG+FU9QV7Azhsm7/5qBYVtCAgpMwS0QQV/ARYd97gLDJ2PogvBSWptLiveyklsp1JPIeimT6
wB+0kJThjKEWfi5P/UBeAkJw648E/iD5YHwSfe4FRI3kXw9R5dGUqnYg2CRnEaPHM0BlSOmBktvn
0BIKafGNFz5gdEeO4i79RxOcf7pxI+rOGtWYI/48eMXBupgz2w09qS6zH5NCXoQpRFflWbNkhBsT
PN7Jn3lBCA7HDmqhBw9xF4AwwThtO9nDm7ROEjCaolIVHjTt8lMit6hDuZHyYSHJfbB3rTewCc+A
Scm+5W/TMSI7XEgqQHOHCdYa5Fm/y6vK+Jf7Oi6vO7WE/9IS39GR5OWy4/0/KRx64XNDQ83GNxgA
/2XWHnb/XZ5z24d2/vBWdUq+Eca5Ib8pyE8WOlLJRQ9y1oaIldi/T1JaKDCCz3gj6awvTPdSS9eK
QInsg/JT9wZYKJ8ta9Zg+8WAsxAcSHkpjMELixsqE3fduPl7HwSIqFAJ4iSX74NsqM5eWpfXYVj3
Pl0SICnmYHMyjAQ+9ejJhd/nyzpiZWcq8kMk0KwdjdudLGxC8rcLQDmu/vENjeUiOif2LRHcIeN/
iYfebELm254Csk8034C92CsPNRg2UCihHsYP/626VW9HD/W6uYCb1g5lGwPXRRg1YL+Bkbnuroae
T03bOds5WFNRqq8GVa7QCtkYhT92aCMqhcuSwHz2dGPTeAhrVkLQIenl54kDwEEGfSMtpdDIHv7w
5VRI1AsfeT6bVeHuQqwLk7Baiwckd5K+DEX1iakYVPhSVtu08hEaRW4JOXua9u+ZSzKpiK0wN3iv
Tr66WXSiI5UJZLvFVzw4lE0ZS6xr3UkrcHwBynbu2TDARr9jpPdHCP6Ro6/Fc/HTf0MhXxLCWnhu
25ebuCdwn2c/zrWrCKge5Gs7qYrePYAfvmCTsopS4AzPe5WiFpDrz01fdpy+Q2oXSgr5qU0SmyJe
cGAYKSX8BLEwNwNBS+fWxvCRNG3vDRjAVrQx91XBEbh95SU5DWT2mR/PWZ510ztq2ui4ZJO+q9Ew
3LaHl2xN5+e7kgnmQ7zg1Fp8wXvtXrUi7Y7NRy61PhxxHOovijuhC9UJRZK8Pwvkdk4puSP7/ATB
sJcItRvJPTpmrme66EOci30Rd6p4YWScklS3USyya2G9m2qQSnI8BU4pSv3l8OlIz2skQDdoF283
RbaxDMJNOUQr8hJ7oEFtnsubL28Uv8DsnuK3Uu5YF2VYsC/MZRURktftmEGTKxKa2YBDr+neYIRz
MSijyvGC7V7tRr8/Urj7GHtZ+PfEILgZ8Rssr9zjYVGP2xPWw8jxkdah4I7g1V1OTjvHz9BTo5/t
3p6r3d6x4Gt5UFDrWAA5sgaGEFw5u2REPSTpHY/Z18MC0m3QhhEKtJ4KV0FHDHWru4P1VDU2HcZ0
0+B6KMMM4IvSJ1TXIj5zN5BxY2q7w1Of5BT8uGAGCZooZ0lq3h8EcyaD34oFhrnPCeERvkfenwDV
3yUNGhUjRRKMxRt+Xkaj60hwxw77nEJ9G3uxBhsWcumFYTmH+ACImJC5+7EBA84YLuEUGigK2k6J
UxV1e8Qz9dCmGK9isF/dB3/lDVz1TIFyLi6wq0iFAzDH1HBDNH4zlXimTlQSZDbp5mriZgNKnwHr
V27z6rKXLZfGNxeoY9Nxw70X5eiWEFhWAod6Oh5gjEFKMNLeSWsEtvBagH6uJrBuNud2QJ98iH74
oVw0vYDgrEQMbjubBTIwF2PfSXK4n04iCgl6vPBkHFsJau0deoTYUTVpXKkVOs6NdDosGgIbss/W
eod83ZiV9Fp+kIg/RulvpRjaGH7g7T7vZ+fDt9TicbjUXMe6D7e1mWD+gShNnBq9Yz1BRpqxftUA
8H3cjAq1z2AcfM9ENX/VBFCR1bXLLZzjMMw7dDL8VSZ2ON1OkGjpnwgnp+OWKZsiNRwwJX/+duVw
wE20ij6eX5E53HyCQsTISlTaAY1B2hH6m/IxwLpACmG1Apdtq6roHXo5WbWNHQnQ0IYhNbb5kNPf
dpA8ZvcHY0fV8K24mm783B/Uiq3RgKuCKV9YUJe3ZuLEbOj1wwXnAhAxwM5pwGjhAOPTUJIwuZTv
F7vLuDZxCBek8Qe2wN8StNHKdSpmVQq0rthxgplIJ8NICI6iuLRDRb1Avfg2GVuxRJvdSNHYJA2K
BT1eujbKs4wm4UmNgy2AaQfQWK1nbmdgBZNn8s/wpC//bk7amGLnY2e04y84OLGiBdUBy/pHrivR
xXhHCd4NV/NnhgT5Z/W6ezpGUzSjcAxkjm5LoKXN90mtc/y5SIGOGvQIMKZce2kPg/MlH6KtfNBf
hF7E7L1kfsRaRytckzMLy7fjxQlg2bOOXs7Ya9nND9P8XAKtvoHU6/pxiwwJCSVrdSgS+8SCng6c
uiX4NC3tCjVL627x+M93/KLXD/HkL4LRJ/uf0e72+Itzt3U2KXKnYyC/Xpnweoxo8Sd4NZm7j7S9
15zJ2mPT4BN7LBTFhd7bZBhIGVtigz4PGTZHlRj/ZYqKpzVMKMsgS79wubDPQ3MKcVDh0vmX63HB
5Yjgaws75RpNPaThE7JJUVs/Bd/BDVrbiS18wMBNFtkVsx+unxmSIP1VeCLdaS3F0bfjXz39W9wO
bJ5B059Ifftlg01rVQsbhxaibUEe9KMcptKX2o/82dYlUu9zBXC4EwXHCPSoDJEbnrFFTHtgDUAc
99P2V2fTx4GLpRb+5JKYO/nITZkdN4ZH87vSbYAs2dKHCzaGGzmNQo8qoDZX4DWV+H3ap1SwMbnx
vfSkIg7hQmEoyIp8vWcHmZwkK0oOSMekBfnaHrhYq+3MSggNs5xtvv9C3ZO+lPiMKilThhS9GnSc
qmvulvKwK4ZtcRwJ85jzqlFkvf1GX9vjwmpeRB7oh7rTtRvOBl7/Q4Rk6oU8ubwpe+s1go5YJMl3
PZr4Mt0wboBlNd0ujiu33957tvrqjhTBEW8YRHX0cNkJnBJIfNEdCKhcL4PGYZSVXIUtiJTpboRX
SzgxtUt9lru4jozNigf7wlvWkjRqIHqhGZjaqrJDulnh2tAzci8iKcBZ2zClVK44hJqmMASl7FPW
sTpk3pHEjyR9tgy7yNQI+/MJeV0CYNWX7tdSEjog/s+iVu2ybUVe/A2GLm1h6PqI/G4QW1KNYwyZ
xzs9U4wAb3bSOwb7s+zZKItvy1swvAg2kNXGTSTdqTWb6N1IopJwlRMy7FXRKwIFV4fmnkpxfpnX
71dcOW6PUGbG13awheI3vaNT5P45Mu1yKJRvx4vjqdgnguRjKKNOEiLicUjG8ktDtpAk0q0OgOK6
fYBmo03UWf26+Kw8KliXe9V5OEm4sqjisvMEVTHKdmG9KT6ZQqIhdAU3R1C7YvFDeN35kTBgc+Eb
SVsgABcR+blD4WdkKb4lNrLTCw2QJ31gAAoizIQ1n19PajCxlu6xH2Z+AQh7MN7HejDnlUNeUtxV
ciOQ2y36sdszbIof73HRFi2o4Sho0RjABu3dt/vHvpgX0mHorIWs0q8QGArk1iwQrGvHAlNZVY4u
YSbIGB8EwIU2lsVst4TFpa1V+5RlmAiio0AzQAFfEEOkHWg/q7sd2J8444XXZXCbu+DXQUQl1mw5
+QHrBVJMeXjTR7y8KUiM76DNdRC8RBvmw6HjNI+H1P/P1ImFDAL4fKJcoSN0/Lahl4Do96vN71LL
OO5R5iiUO9AwPJ0ixqH+Ng2HtDhUL7CJ+OBwUEU7Zdc+/cuUX8I0e3BGXbAZnuZckltQxOUh1j4T
0su0IQ+1VcdC5rTgHGudnFvq2WE6e1DZNKgfUHwoBpVOsT19TpLE1smT9aGUz75tuZLsG/yEQp8z
WfyzJul34F9E2IQKwD8xrjwHAQwBifgA+zhHe8EcDC/vN4tMdK+1EX6ssWv1k78x0wkI77YZlUKw
6OWuGvqR3kCC3B45/KOsGZ2nOwMdL3ZPGAEgOyzted9GgiBtRCQD4FcuHjgzmmvCQ40JAnUlb3UV
JhwpuXo47tvoXwEkuxYIEooP31OUZXiJNjvOL9NS+QJdQ6a9GUI+G6UkgKc4pRX0y55z0tc3TZ1P
qnMkXvpLC5xuyo2Y4akyoiirLCky/iuvEdtVeDq7ysm5P/9lrOfVwpruXrAIj5GpMpegoGX9ORcz
o3O/3ZBcyLpjWG1tATa1ocMEQLgG0Y1S+cflXEO8i5KX4eDkmbDBvWGS5FdIBbAiImFHdb36rVxC
TRFSyFj54839Oj9s+hGltWzoWXYmhpVUOMvn67pxR5VCAdDwa3aA+jMOSMae4O6ga9LrIWXOBotb
WZWkWP5VLQ9ZYz2ZW+Q5gDxx/TUsuTWENCtyaRa/RJ5Juck6oYcnVqJT/nxbcihg5GGUfHuGHtb9
KQ61hCjs+miJK8bhgU6T2frhIJn7daxuOOInT0aRTlN5CoB7HCfl9q2LkJbIbGyt7JNa5YJzovor
WmglwKF56swjAGdmas+geQU5f5LdkBm0SIAT+v7oCcuqJ3RgSPNBGSp5ToineARlZxeNwJEFaaeK
vt9vOTvQoL2+BSeDcRjqF2f7XwOgnZGqfIi95MFeagSgA5tcU/6a1a2u/YZYeDi/9HPpl0OBtqjF
l12Bi4nSYr8ragE9aQsIs/9bAoEH5cpqKI8wVz8zdo1qt4Pn5VRH6DBwXhrwe9OtM52/TIvixi0v
ShuBEnfhFUlh1YYh41ZtPxAD0zK53WJRU4bhX+8mQvvfuT9YhytSzhrhSNJsClklm3Xr2uVWnDTM
YJxEFrDIAq+qPt7o0hVWKPPnhs5LO8HM4+zZ4aEjHjAxNgeCfQmC5TV6RcCVzQlvPkTdoHad2UCS
POAe52SA3g9ut92MmCnQ3bObQS3pxE8l6OykOAgTgrzleuyT+2tqJLi7m8ukLIYI+Bt3SRhP1FaI
TCV5CkFPl1IBZwGf0qMnk9JM+jMyoF5dAD4yTbfvgHctqfQvtpZHfut23a/oARl9q7T0yYO9Cilj
yW80vry0GVccrhFNXXE7o4fs1s2cfMqLlMBQL45bko1MaOZAIp35pMSdRaznMThXKlQugYekMR5w
C4zIMXqQfNPZ+tahF3YgztEw4MsgaP1JH4MXo10oqEzbKcQt+PImwGzJklhf6SuI1jfzmWH28J6j
RRtnkoyTjn2DYj4/QzOjBHmmjsr4oc3Uo+4YG5Fqn5EzSV0J4+neJhiQEFwTls5stzFrg8H00rgP
eKvuA3pJUkOx1IsJi1nER519cu/O+mYp1zuAs8K3WduByP2hkIwQ8OYy0IoMDXMtwMjSIg5bh8Tn
BoTCdn/pmlEQxADKhbqXbkH36Yz1UvU93zTEd/+zzTANL08Cup9RFBa/12/AuLnMD7bAe1bZ+ZFr
TGNmSp3QjjbDFw5bcgrNsgXCspkHMvN2MLmw4h59L9XTTWuztFWoefrW/YHwScDpfPryd8P33VG7
dQyiIbo8X4Q9dl/lWKC1kkunFVCrICv7if4ewDhbGfKTeYmkbTsTL4cc6zo50QhmI0IreRLfP7LN
tljZ1NX+tpZRBQgzMK1/En0HMFcML48/HRto0N6drMeZz4rnm9mG/zrMQwqLYjSh2/6j1J/1Qigo
8YmffUEsRVfb9yo1x5pmn0NIuUeYlMpmqTIbwaIt+SYlp0yOVu9Ocyk8xc+imNgjWO6oFjqMAoy1
pzBb2Skqiu0FPUO/n1XKYTUwBHWr10FuJvimGWvzyqwk2G7Evr7T4q97Sl91eYWLXNxesnIMC/1O
wXhJvjw/BrqPASWiGFyF94ffUnucIOOFuUZshPeGW8+HlYY9akgOaE/i621IDZ4W68idyah51mRl
1Yrxx4BA49tUHwpZi7SSXARzpHUPhOoNX69CKFroIFHlXaqXWhUjwKUkvzqBPgrrR8kksKPqACTi
/1uCcqZ53qjfedowySCqynq89TAofx3GSHFC3lbutIShSNbvbL07udQh+0dKbaCQS3vrbzcGfYdn
6M4KheDxjOV+/V6gKyCVeOZBClpvoqNw3M/DCZMvoKTaVylWKHsg4jk4IGexpzwhGa79c6bsRlNX
US1Pbl8LmvM9Id0q1juUh3nBMr6Pu5mve+0orRoNnEPTwf7AJDJRCk81+rblnLMf3Ki4LLS5ssFv
FlpvQ0tKEamHNK4GvoFjLrY9p9XvWxtobOtza4Z3p1CMEaiTZSpVBqc3w4BlbhJHX1mdmgZd0T5b
CZGvrQseh4wqDt5o+PXHDUNtsfkmIMrpPO521zR9Vdexqj2FWKwNnT1l91W4rvVQCuqEjKiKsQeu
osY5SpbNiKSdml6zrk1NToEoj0sHMig20GFjDOWL5TB6XcH8FO7HvxK+yiBesCLY7eVcj0uyD23M
NCMZfyNoU2ZA8gqTuHsJwmGJLzGCuKxt3AeMivknjQTqAVPETr667nOUcAalmw8BDFVYpYDT0cGV
dOU6RmbeYp+rHYBg57Kj5+HghmAyeHGvxeTFwYzBAVt+5mEJxVnDrZVSm7dlrhj1SWRUVjcXHxlB
tum61RqSkJcPD1eKmkIZYp5ok5a2pJmD307bGYeaQbW8rQp5xmus9N7COBjz/y7PjG/7hhQREE6v
AyW0c0FGKoX70hSQt9hdXtmUfYeKpaTKS/zm+Lw1EcutzRz/yWs1Lj6nixfB6sRNqcnHdNwJDVUX
HOOe8ByJxu7+p7yMQtvKhpgQBRHBRUqqUjgAzDIvq6hfeTEeE63/4M7/yXq7v1FSiHacPS2SVgIe
rylBr3mwqHlCJxGwJ0NdC31n+T4lD8fLUhROGrJ5o+/m0o2nYDfia/faKwJzGC8JEN64L+3Gkikt
J7ajX2fucuxR3ImYydmMKRIDE+KrIOoFmksz/RlVuQcmVkTRft4Soq3G/dofPIexa9/zDfbkBd3q
xE53vGLgOd6gAv8UsRxLfbqsEEW38zvEFg2h2+MJNWXh+2a3cOWKBBlCC3D9/lBx30CMrjcbeiMI
ZpYuOfxovSTQXKtt+ngH6MSERuff5bR8UFxh3hPO8BvK6BAJT6X+jp/NlSaW3VIETEcG1NXp9Ya+
URFn70InWPBp//7aryNeb5zEHmLB9IfDnR3Q5Daet+b094pxGKnFnTz1y3+4+wtVkJ27kqjJfFq0
DsTXWCBPeTWwZvoUP1IV0dS3584bsLwJwx5SYadrh6LpN1i8+01esInHmqpiqQTZ/RhRbJw2BFP3
wyRGb15zTlIOpvHdh9lgf5sfFZQBGzKw3QmZ/K04DRBReDI+CGJO7M/4rqy2uBx/1ofPVW1MbGJz
pk9WVJhgUv0w1eukUGd5hVEli8zoZ4oWptEwXxIEDOzk9nQ4VTK8nLxxVd9STGrWLLuX8E7JI5py
QgQa6r0wUJZy7PQs7MAlvDHsochSFDAsAde1BnH2QgLXhNzy59FZSGbPs+Mpho4PWjNM8KnYP7U9
QN1j8nn0u5lLqC0g95QoWNmEP2DRWJ5QdsUvhvyEeKF1EL0TFmrYZLrL75DTqs7mC7+RQ+tDhLFL
toWzbwsC+9Z70ktW2OBb4sD9KneMAIozGE0TBWCahuy+QBmrALMNVb9yqDcVHij9yYxNfGE7INJg
s8BZfG10DxNwBBrF8aWf5eoEyx+wiKxjqWuR3hSRaAeRFSDGN65DdVF6t6Cx83/CUrzIrRLkbWfA
IHDUgInVIsirUu/SLwV0zR+7MHNVFfm0pLt+mui2Mt9pd9IAj3wjSbL5x3/BJ2jwo0xlP041BZKc
znPYY7PEkoOexOc/ib8ls9Y0n8NTdRjKeNQFarxTc/szkaxBu+4hSLv9f7syjc8lV2HhMMbxLsEI
vHDZAmcRue70zq8pUuW1wuUrnHbLZkMWPA+ygKoCIoPd3MzhrSiUz0cgaoivzg/htgB2e8+UemSV
gy3YeiyrMqtzjkNTOr9DCH6nvLil8sRRWBdLd67O2GZ4OuisAHDAftGljvGjual8c5mrppI1j80B
UPZKIkPxV1i1BtmAb963ocR+re7+1m6c8gs/amorzuuHcN6P/Mnr42UH5b2eXed1Jbkoggm9yj/1
CTYcsLp9fcfwDFXrW2ERZZaH1NWRCIz5GCHSC5ZX+/SSpkGrdvxkpTi7viWiGWbdyDK1CCk2EZUf
qNPPzhZhoy5+1E7Xe0zAczAbSFW/AONZG1Xly61WIGxPZEEtm+2axIdSJI6nOfssuItYpXvc3R3q
CJGaXNN2b8Q2EUpxc/6ou+xo2tnXuYXVNIG4ffzkPd9nBumv4VwFGTy8SXY15neyOWWyLfK2P3Vw
OAZZCX8691QXXU6YxNvIuwkJB5gPlDDdxgV7Qlw+r6weYcDkShOoxyBjuet9VFzQHBRBzGS0kt/f
nfwmE3lwe8ieMEch8wFJg9VAzqf/9qZzfNkizKiWOMVjVWgnSmfB3Iu2bZJ/5Ht9FhOzvFtpkhkK
4SFffcY93IYEeW/wRcWQIY1X4vz4SYd/krx2j7hlBGp1O6vfWqNyjyvObExNDhoor6cdVxU3YgOw
yUxxwP799EY+dA/uu+7FiyzGAHPNTkWWvw7q3KWGaMavvysQ6/agW5Km5Zd3eUF+dz/dHtf6SUu6
vFRcKvvOYPPtV4Wp8Go0df3YNmpqh8Mz3gGUEq29xVvVDTOb7BdJOUtQgZn0/ItqIUmBdj7ByYr8
1WudqCAhD2daNiYKRobqmlv5dW6qn4eg2PAVYi9DdCC3PfdYqqxkyIc9Nmto/VX+hjkdeVDVcLYN
1nRc8zSwhtt8TlnKlBOMmdQB3XCuww5x6+TYRJj5SNgQwtEaak4G8VAstJgHcsRi/6CJ9RFpIUJJ
50qdnN7PkNUZXt57Ub/aXhfjgHesH41SIc50m+eF2TwahGlMI8CfsV2oRYAXI1uEBD9K+UQnBLBT
fsgYPQi0yYwCRbLdWXBu1LMtAWt9Gjbt8cem8CfZdiTaFeSmpF+jZ2WZkkTWs/37MYSzw7vCQsxx
7tIyqvCD83jkjTvlY6D3bdD/kOSCr4GXO2VRceZgvoRHsMCA/lxoEvStvyCQYwrnCrkcbmbV46Qf
INXVLMF/lNoq2xt+wGCXiv6f4f0a23ZwCz4JiftKQdnSmGCCxOAFYITmLMGFdcTf2VYqIdrfxPBF
GnA5PZiLWaSeIAgkWyOTT6qh6xCxLBzNj7p1105vV6esdIMadlC0Lb2JLlodcLr6pBZUVN98jJzX
RXz19EiDqXTe/sBw7ww0q9LG5JpdaM/L3TEpwZtyFMImUv2nG2HvofgjX5VZBNQzxOjNqclstmc+
jF+nxHdsXrUXCUXMR71piOymJtjUQsaUmH9XuhiHS6a06B7iGEEhaSlvBQSZ9kVzabjBQJM6gSZC
Be/EXF9XQGBHNHMinxmhVwW1q7brhSYI7G+k9jrkAgvniQVc0OhRZaMybKDBO9NEwjzD8pcXMErB
JuLh8mL3IDv4PESV9nzW/1ki4d9HKS4nJmi9ziXa78ddeMqqCEmBZ8brf8B/gussrrIv0V2kO6Z8
jubTOUcSjeM0xgIRw7Cg09UU2dCnVDILF4t/zPB7f7Nm1fPH020dnGi53ca4RKCZWc1PvEZkZSJS
fVMH2Ll3iPjbaaXE/qW7XNyMPMTa6QevfnJNXHlnso9rtnP+0QVAjKel9CKpe9gFQM0h3UlhE0Hp
kLm4cbZsuWC1fZ5PXbmiCnVR3U3uzWQt/nxsTeTkRqfkJISUrWvJgzi2enSu5IKEjBxUkt1Ez5wA
tHpizKYLz1A9AO9+g+u9YJFZDQmB0K1lnzlRbynrx0Da697vzW0Yt7l4XVaoDA5b+4m+u3QDhbmI
upii0TQhPCG6VQ2fPDUCdCzIZsEeq1H0Mz8Lnm7iRRGJMySm32lFjOmWJTPOGPcIymlGuThHKqhH
VsnmsEvNPhTFfSMhhZOEDKQ1i7+EgxeIe3AB+KHAuRWTvOhBf+IIwmoQm4E+X0p2li0LJnvC4IeG
rwNDfHJ3UmgW+efP29gtuoVbovyU03OsQ1DZmoZRB+t8jdrgHt3Fu8VSzryEWx4qw3L3TwOiXoXE
QFEkQu7N/+niNXSlXrldbLNBAGK33lFuNxTp0DlxS938x4uCB6HZKh0d4RtmPseYdB6TnTyYoyVK
JziM0xvOIbb2PGPmcZCjr+/YJpUCZ9F7L+aI+jEMF6M6bD+DVNMIXG16gN4mA1hciYVTMJ47b27t
uHoaN0s3u5tXW49VxcAQe4th+rUp226SM/CTkra0Fiyx2t4r6ysj3nqONJCRLcziIjLp2sKEGgyq
w5obC6Wn2l60SJEW2xJNUeCMVjOXROHlJAjUCy3O9Mscs7vcdoI0DM+EZ6s42Fu400z0/UDaOa5K
GAlB89AknndngS8O/GQHuLL2oC96GLyFMjwDzVuCwM+2YUruELId0e/e7VSBy5QZnlBwo9dlBajf
FssKrCyRsxjSOgYWAYON52T9HNta3O8h4kr5mejClk4eYCDB7V0HKcWDi9Y9CvX1L3c7hQS7Ksi7
cJVSIi8Zh3UtPG6R3kXwHiTodAcCU+z4TAen2MYQyAdI2YIXYrZgaxDIPeGxVBESHyrWOvpK3y+s
aX439EthVzvTUP8K7C79DvYc0tqwfe1FJU7J/aDZaL1nSzzfEibg3k/RZXmOJd/cAnuge+UlYOAR
slZhkA0skveSkQLQvLqTWuLWYqR1Cf6lVC7VWSD4dg0cExo+MRU52vs8iz9YpMBGaynvnI8gFy/Q
QOzNIKmtoaKjTW/quWhEtcYBH7ptrLb812egeBXI+q4UUMAAR8ESgoHa+o/W6m6Id6zMeBp+2Oo6
OIRhWjMNIMo9CP3aNUF0xaFXg+kambLE47wvYeWsytlVMiITROGjBB02MCH5+DLixrocQ9Md1qeW
7enX5JUcZ1hc8eOfk0UfEPjDxxo34jA8jABaQV20kcmBXnItCa2JFd2D+cS/1BltD6HLcei3mSiN
G9NZ6MLPSjBL3fKPg+mU2UNpYd7KIwDcpgLDi62CjUofawnWvSMMUyqJVG9xynE5hAhi4awkGRVY
EhALlU6OSvkjFCEpiVkHh+VGlTXVc00O5yBCelE9M69xcA8BAI5tDlG/0ybf/Nc79QsTpX5YQ67c
HyD+j3ZhR7GT5Prw+HQj99FzjDVqp9HDOS81IqNcJLKwhBjZW0JREv6brvfGTB9W0C/wVo9j5Yei
iGNbvID/nwuSlERIHDADnfR8QaXwIGjqlMM8BI9I4L4ytRa+va5r2WAhzgtcfJZgTXPwcwvh+6pv
wocIIQlx6oOS8yTU6esl56xCv3wpWsMWD5g9+ldik7QSZoubYRqTYZgwuCv1B4X8ggrArVJLmon1
p1YETnbgjwmmUjVtM1w38inNnkwixZZGeWzJ7U9XaV2JimWz6eevWwdR73jA84tSE1/GJwbXGfqT
qzAG0jaOaWFQl/TwVw+qbYV4ceuxj1ZFkWoGB9d5Nr8V4Ele7m22m38OrZlxR1Y9ks/MUCH1SE05
+xw/c9UX5CXIjkWptakDda4FwRzq7o1RisCOuHdtMaYcHdCN+86GibV7OjbtNWrLOjRFVIdkn1ib
mMlWCWejwya+rQFG8WmO4fJpm1Lv8st9pdw8QlmFeR8bHjHsrookBQrByi7T+aSvQN8hDQYMs2fH
MjEbOvecA4VUVxFkcEuBbpXf1qiq6OeQ20JZR8jtDpl4pZVg5zTd//jTLZjYtFCYAO0f/wj/CZmW
n+ZyeCFtT8z3uUnLZm9zTkLv7RGsyk9dSdRTn3fI2BpRyHyWuGIAqFtCrRWaX8O4zqII09FlNLer
I9ZipWfaxC1g6N4rK5El+E8p/doVHyiBpnuhxjlUrFbWC+8ug2lC7vZVpwi7UQAusCkt7MneIsR2
beZg0qrQ5c7uH4YRq9lQ0DrTD5taY9riHkzx05eFaE39tMz6569EQ6FTFdbwNpcySYDmWiXv8yN8
MoMIh5T5CqqeJIQz+pezGZJ9dHAvAlUrgEWuTIRLmBD34+C0XQZG07mwBSmRlMNcngX0A56XzqQJ
AUyAx9k8T107MeXYa3U/PmZJI+LAdXWUIDlkO8bDRfe8jD6FvCYnbXtnND/2A/J9wHizNUrQMLcu
/YIutt7902bgIx/BeYQJLwNZyYtIYB7EpCVZt5WZZP6/nNJ/MT11516+DVEx3GwsY1FV4aDX92m9
OgYfnpZsRSPryhfJOkMcD4IgG4t5EumTe0s2lcHnFqXqCgdvc85QNFlvoqGEfhGfCOo9ZWS83vzk
lQ/94Xtv1Jp9RzDI43O1qVGnWG2qI7w5Gpy2C57jPyxD5fgC+6Tk7VMHAfyVRlW4bcSf1Vj6jB5e
HAFT6IaGeRYthkOUgM6mUAYFUrBa8bml7nCQI6yABvQaMx+Nwp+6+vSUhVPTOOIApV1MaGnVBpCf
Uf6PNchMuLcRGKT4jn/HSM/cLnFfaoBIWpax2kEiTGmjh/DVt3hKL/H+t+L/K5nv8mg4gD1Yt1o0
og9SC5h/tBzgWuRi6tXWNHfZvcdDDPZ+bgfI/os3M0kB3ebXeQHaFUnCs9llcVhyFXnJsf676vTe
p+Q3/ZUlydWIcsanxlDiwet54c9urvLyGGq/dhDYnmeiOs2iaSW6LCk0G+9xPnVgGLViuITCjCT9
/hki8GQqF/aYtJGH4b0aaVp8JP+qJQqzdRkuknjDEu/gF7t+c1q0ys/X/B2+XNFZpPN/3TELkuyd
Cg8kb1E9m2SVvK/mw+G2nM3sSlTlHLw5gWvm4TeqwI142qmLsvge4dC+MKxeqmuYx/Za4SUcSZF4
NVCu+t7EVkrHUuqlPfSD4NMP57M6oL08WY5nYHdSmtfNQsh9wisFYFHJRmKY6uwMoRGNLctNaN+J
20omxzBkho1IdgHmAyMak8hFKo+MiNvCzyx+bD0uE2Zi3suB4J7VaMoQL8GobW+u8sBTIJMfpmVK
t5xQxMFH9lNDIIpaHLZu4t80HHz7XoCdmn+5eB2IqYHyYPx7GRLRbWpRSX4cx3n1+jsct7FqdeQM
QEftHGci/I5a5CXYVYAVntgZ9s15XT0tSDlewqFR2AUU/mdxOvABmQEOJ6vBpWKOgQTlB+hP0HeY
eD484cbpI/qmpOl87/NBdjeqogXtQgYqedeyG4LyI0dgUsMmOxp6jSeBPB/vlPA6VIKcRaQzP70i
DONzINlQMvyjZv3OYwk+6nfIpVWJ9mOyohrD7NRJ0Kw9uy47WJNIdZ2hZnFg6q7HHS+wCjUOPY5F
jUmEh2OinPezuIZ5CLKmzJariUwLuTnDY0iICPlxiq5zIKbvlw/WUsodyoQbLroJbP9DUpji0n2M
7wSewPAkTtpiI8RWeWjG1QRGuiFODPRJmPFZcKU8q5oV+EQwPe9hs1pCyWP8Jl6kmzvvGc8l5TJ7
xV7ACYWXzk6fWzjbdocpA+4ZRdN3HnwRm4mjRsOUGZlpG6xWdbrSVFrJd43N2B0gRwPJa7PtWSdP
kXCWAIDsJFL8dwNu7SMNgu9jn5ZLEIOS+TD5v+lurNkbKb9tvfXkvjSV0KPLdtTUN/8xYhj/wc5I
oUtedPLIFjenSE4mO6Kpepd0M6UA4HEpmm36GSeIrIXiV1fZ8zrrHGqzjfryIYzd/AhJ8G1sy2Yo
j9WyblP0cfmk2mieAY8ULfkDLbKmoPZFSZZBQRsAFSx5nXwlR6cqOvZVGxtiejduknvLDx+nwLkr
/JjwwmXBL2hZNqhae5jgZNvbIQytx6kniHSeXefH0g6TPFZTu0ub/8TkCKeHLVe2qfPc8snse0qE
h8PXKA2NeJEoKZC785y2ayn9fapmilKCya5KBfrXGYjcvqy9Vjg5XJSAOjRQeR1nK2rlfY9g8pAX
Vx0G620lC+2vt1aOpBC49G+fMcVAgHw=
`protect end_protected
