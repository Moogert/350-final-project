��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h6>�����W.�b�]��ɣ�L'��f���JT�2n'6�Z�= �.(� ��n���V��cی9qT/�	�VZj]�(�ͨ��Z���A���F�|�bԢ���fF��[C���:�CۈH)q�1k�{o�!��%�q>�d��>@8f��[��V10>��k-�_�s8�']�> 8��8%`!�tOD��x��lmS�(�V�oݙ�Y���zP~�8�e���R�cn�]�� ��u�=N��Ǣ�s�+�n�ˬ��p�t�pW(��J��tQ�-y�)Դ��?�
�u9��-d�8��亠�FU28�{�]0#�d��	� k.6��k="=���������x�ͼ���8�%0�r�Q�6��H�!%GH�:�QvYTa^�kiVZ�	`P�4@�kh�r�iYZ��e2��[�Jū�=\����&\e����	_5Q~�)wG��?�g�8���[�w��?����-3��N���x-O(xuƳ*�l*�T�(���WB�ĉ)�/h�e�]N]߰���BS���nO������so5W��XZ?��پ�B���'�oxͼ����~.�x����#e3�F:�~M���$)�w8��9���:jK/�49)�VҦs<ѵϺ��1XØ���^�e�NN��#�f�������Bm�G͕L��/|������f	MHS����R)�H��"%��ĥ���œX��S�ZM^��������a�!�`c	*:�75?7S41���`�c+X�O�(�]�i�Ũ靰����je����9?��Z�����uҰ)���U��` p�1���y��3�~ƾ��61��C	����L��f�ĭ�X�r�y���icZP[���Z�}a�bONuė��c�K|��w�n̖XW���Z���[Y��\Ч�Ԃ�3)k��w@��w���4j�C��'��6�7�N�	� �s��ȿ�REh��������҉��:�] Bk��G,V��֓
o>�J�ûfd�>��b� ��~�u�a*ń�a�e�my���ʹ�ů&�D�0����?XC�j0�����\U�5��F�&�����n|�&'�b��������gA	-4�~����/r�8���D	B�*^}b�%�tX4���Qoz}�~$=���^U#M�n
�p&Ht��*]����6�m�Z��V��0�M+�H�������>l�O~Oa�Zή.vf� ��.�����U�<�o�n�F���ATf���@[���7·��FM��|����?-����G|R�b!��2rl�B��Γ�rB`�JVvf`g��->�<�~6��,��hΔ��������>�a���\M+���|k�~Uk�~�	V=�&"�_�?��������Q��84_�'{�L�,-�;,w��$�=��0[=�2݉o���A����5�#^8��e��b�����h����6�x�(WA\7m�P��SG�7��4���첿,��ZN�4�4�=3��P�ζ�)�t�Ul�vҤx�[@Z����Za`�zEa9�K����0�3q�fT�ʬ�H�q���8 �;��'�Rh�]�&�a�9.?��1����M���4}����F~B�����2rd����y����`p�,���k3�;�I��𚉷��bKs�G��]��>5���&*{�
����4��^#f� �˴H�D�Ux8bg��(lP�*�]��,#�~r��X�3�E�9/��#:vKd)G%5��B��Mǋ��CN; �7��X��uKEAG2����`qRֻ��d�t��{�}��q�*-�ЃE�˓�-��I��I�#�)7��7vHԤ������r���������Fk�-LH/�,s�g}㷞�֨x�-�!�3a�zl��`��%^��0¬\��������ٸ[���6�Ŀg~��s�a�uȃӾ��z��cJ��4&��MjT�q���0�R1h�6Wa�;�-�tR�6�H�ָ�-�I�z��ǧ��+�7Dd��D�̕�rXe�4�=����!���oY�[�{t$����ϱ�Q
���7_��[����6�Rx�՟�ۆ�ϴ�͎t
J�ɢ�޳}�����/|�@�ޣ�Ԁ|��Ll4�?�����;��Ff_�?����n4"��bi��d!�+��Y���q�nF���
��*\�J��A��C>��&���xL�o
lp,|>��Bp�����=���Qy����/m����cDl�(�����t������u�'g�x�弢0�X}Ҍ!*�1����b�r�P�c���jgN�=�K/�$7�&�1�J��L��W����՝�2o'��hC�n+F�,���@(��Ǵ��������Q�̘wl����bu`w�7��/{�=f�4~/^q �*r��'��z�<����#�J�籑#�z�#�� z^�\}�C Q!����
)��s�W�`;N��˶�A��v7�d�/%n%�m�b]��D��w��G�Y	�Z��ӯ羅�q���)i�8��׾k������j���?�8�C`�4����Ym"l�
W�2պ��qM�qi
>(�b��N4�gz⡡~����%���@~09h%�v3wl��ߞB0�Ĉ���,����$&C)Y����p��G��)�\ #e��]{����	��^����4�^Gd=9�Q-�CbZ���j}�����'�Y�O��b���zho��� 밪"���RM
��_�V"�Z8,����e$��H���L�Q��-�i�׳�Q�� ���va)�r}�����2^��&7�;�H��n�K]Y�%�{�oyL�)4����S� �4y-Ka�iײx����C��+��� ��B9�P��3`��(V������u�9���huս[ w�����\�s��I7��3�z.�«�@�ןa��Fs'�I���jN��&4>+��j�L�QD���Vu�nH7��x%����hS���-6�3'X����qL�p_6�$`ڨ7Y�� ��;�"��	ٵs���j�$;c�>�Hz�W�{)��`ŉC����wo.wIL�j�7��3dW�#n{����"�U���
!�H��z1��鯂�Ks�̊rsO�=w�p::������mE��&tQw