-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1xnFhLvWvRkm035PwXMaB4uNNktZ3D9tfrTJcgUu7viYnhps2uXfJz4i+p5p/k7vqYFV+2cmoAJw
LGoLR4VBF23Ha+ROOYhRNQ+S7DhFUGltyvOl51uRqTaDmTG7k96CenVZW/X7Zg76B6yc2qIdk4ly
2zzEvyErig5EXOKe2NJx1XcZ8dnf6ETffx8598QV2NPJGocBB2P9k8V5NWb383Js6TaE0ce6b81J
fin5hl8/3XyNnTd4sVr+VUE14i7pYvfBw0Iv6WfH7xR1OKh+DLVjhJXTi7gNkLl3eyfkXsax38JT
W3bCAmp+gOI9KmIk3kHgxJB3WuCMhgioC/KVkg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
m12EjMHxZ4vYknbMZh3iUL3H3aJpM0jMtftoO0NIpidyY2eZI6dyI9xf7uWRHM1Bzu9wVuluWGvO
Yj9jxkDbaADxyX3O3qUuA6mY/AMTzt2tI1I4SPmRASiP6uTtPacMhZHXNZs++pkfrzEXZvoX8Kfk
ovxsPPUD0BoRC5Ii1FANpUdKW/bC41yCf224Xo3gyU5mLtsMJtlaAZk/6AQp/2sJlSTB7LSNM8aI
pKPPoxRxYvyroCieTMyjAqDJBmnellNtVbdp3zObKkLaBj7iYkIThlKr4F/5nx2LWf/7jGwy8FAL
CF5CZvWrMXZcIh2Ywt2uyt/1aCVotiXloQaEhFQDAM38i34C9KTRrZWX2/pFWnl7WWn0zxsIBaju
cr/9sMZB4N/do77kFD7Gb2sZnr1RzTqATMFgYrrY8E/nea5drFv79nrXxE2V84IZeMXIuqz3c05f
b6J1pwVxqGarmb9Tv0+YDGRBb0DOrFRvp64g/AerYIofQL6jvuvuZS+hctg0/dSv09w5+NgRvjxI
dniV6dH/RRMXBlXnf22F+AdfvaHUFYe9Cmf5+O4sJ1a1T7YSRu5hNyDjOb5JkdSaOyG4k+bsOLyu
nQdqfunet2unbBl3RM8G8xlbPF/k9GDrgU2pQnfb+rmIRAuzXO5MLYLvHq/uZbzfKLgYpDQ7kNYj
MUD8yvIbHBcrhI8S/qGQ8nWmift3P9N5rpNN7Du3z2oxGqR9Z9JZho6mfE5d2g2+6nShwJtISJhH
uHSkRD3NR1AKsPST2EYkIL+wiB02Zy9O/7/N2dgbjU0R+6aJGdshO+bkhKCyWnwYKs/YTPUnL46j
F6JS1MucQ+CA/bmk1xzbpAaszLxU0uYgdjJJcPuNYDaxh7tYwdbVU1lZ4h+bOAdVS4LoHC9prKbS
2qV+zE7xsorxqKpndsYxf2nUqhiEHrxBpAbWyekZwcavRflZnsfITpYeZMBVX9WOY7/nGSWng4c2
kMG779O8bXyfJtn7W/FELaWRxbMaS1BC1q7+dWWz5B96MnZBozJa9lLBqD6eRujJivV0KmjgwtH/
nB1oXEHp26K5ldtO3et8P7tcRbbl/0PrbdB08BIorJIpIpJHQzy8vt2dV1rblEMe3PgwkVHdpz8M
f0r/IWgU9waaJGVzQlacK58B5ogWW4bP/1NU6Ix0+tgEQOF6yyEqaiWM+m/fxlPzD10580QUH/+C
OxJhle9KLeEFo7udPM8rkhAz7lPqxy8R0STtM5uKpr7dy6Xv7yDU+3c00esuq6B5tMeqqq4dvs0W
2YI5ZvMQDQzdZd5DKKgWgZdwqaCIGix93dT0obxzjZBJd3QJjy4ihu0dYwKX5seu/AyK2H8FyFQB
pz1HCk6XOTQarMMdEqsBW/oi7RMhCeJToV3gI9vsoOk5uLyjG5UVqqeRgfFDnmkppUaH/V6pSYfg
rZ1uADtP6MROSmdWuHVIv/vcP/J6l4C3pAFEy50XGiPtgexR5dpGRznN6BQ5SiXttyL1pg6Mz40n
+lErqErKxjNg2H9zayHG7srzScp9b9bkPFUhj6VnKZINq7LbofFWyE5unnMNiIxJiD/8pnxZ+lau
1dC+Zq/d8OUdKC7/h5li9qrmX4n8Siyw/PyXhOh4eOPRfNiklhy6GB9Hs/PPRX4nSHTJLlgcu626
V6GafwvyIljeho6mbhQ72z5Yvd7s8gPLPWGIjncupVbYzUx1lboE+9Aa+OAsU2vpEVMah06bX7Z4
u1LNpUOp84SNxT5e39zveezPcbSJlDFO3Rotx9fw3HoZb93DDOO3toreHROjUaBQgY9ljLlUez24
OrtUkawcDrts5lRWkiR9L4S1yRZST6dce4vF/6f+wIY+iw4blrU97Crum1g2UXpg/734tDGAngwH
g2HmMAkwAc371Q6mQN4QmHb9a7OEn9C6v18Jxrpxjsrir6l3KML1UqX8T5dJCREN/bXrFyGH9IoN
J8vPMXsF9AhRyPoyTNe+bw9jR7+fe+YI1NRERGLLE75Amm9qIp1/JH8jvWgegHP3lLqFjJkMrB1q
Ef87kzH23H5XcYtQ4RnPSQgZ96YueEsDyE0D02UfFCq+fUx2OoZryPoisquydwmNhiNXWgxsMfOj
64KlLJrYaN3eP2wdgBLEcUTr+Kt/Zfchg8keyN6wFfto45f8zI9qCwuugD3kejvX05kvQTmZvK35
X8rL6tp3IGfOXDcuFciiNh/T/nL/KmZ7KQkm6YNVRlKyFyjRn0RHzzU9wzr8pIfEUDKZU7Wvgi5e
z15K76WCm3RrBv8Q0Jn5F+o/e0rWEPPN1iHMNpLY/LvuiI4WBCUEg/A7TG3rfEWSeFa4b17K44Vr
4oWgOMrcfhcFgacxVaQd92wy0ICrP/9W1GgDL5Ywq1Dv4TGp1GYcJPdzJACL5TYBEyfMNlkeYQz9
vC11NCHATvnVhn8FLal/xnBJA5kFNnA3UPlh9SHw5JnWX7dK62IQfg9jE08VFcvWlYgujY8yKOPv
RrMI3JFS50QZxss+tlZGWGy0+tZ1lEe5BhVVgxipP6xSLTsRTjJ49YDw1YDhVZpy3gs9S9pcVOn3
XGKU/uID52GB8te2rp55fGFX0+t7g1b464H+seAIKtkVc4SbiwiitM9vK80UFBouGxYR425DN7Op
i9QtZjX//Qt6fcTHc1MneOlByaanukvbSqrxiuhU1oLUAvq2jVsMj5T98XIq62bLwE7bM4kzIANZ
TMMg7RlM8xCkNEa3IC8AuN0iPodSSWpaICWt9BljXy0yrAMjduVmphXk3kvkOvaSmxvvpuvzOKAN
ylNTnzNkb2K0MqTtz1WiJbcvOmb/F7WF44mPv0sqdtryLxy1MHYp3rPqFBKPjdRmbWDE5EaXTWye
nKOXZ7PKrGG91LVk2s6Z0BVFpYIgva4eREI9uhEZ/ew9IeZo3ypkCs6srfwXnMBxMHGOOf1nDXSX
P1Mj4liuPjSwectY6NTodlCW4n3ayHbqkHZqFwda2H+3DCaFRjhjQBIjSrauHQQPs/D5Ve7ugGnw
BI5U84e3EpaI2imj+WlUW/BPDgBtAjakEFA32ov2QNdi6JUlmdJDQJn9CDXyPJk19mRTlgqz1crF
yUWIc3D5INH17+eOPnxQ/51TjQxIIxePC1BtHRomA7sPAuWsjMYqIMRNM4OjYcbufQkGoMn04zIx
nt4NqMSETHt+ALw275R291rNlJPY6brmxWb62qnoz9Ra8c9bPRwc2upCLrtL+U75i5ZxoTuthYSH
JLfOvX4RBtWtidhV2hmAOeujmTdDT6rmO06Cqc5HqxumCRWsH4zTr9IkHzAcrMsPiEz4Pg9EnNcu
/NIoyoLu5zFuCxgjUFXgMSAEI9kcWFdIFXn0TUcMqJZAH9s1pEj+27nvUif2zrj2LjsuUxSpqLUK
dstbV62Qe6H5aKyuV9weOdLHyKBMH0JSlEhNqiGGkjymzXd+zIdpA+b2KuVaDG9cznRHDWC9JKzb
U6AdiW2uYR4d7LYvFvhiZVLCNC9DjERyOV/6g1MVmcI8aTQAs2z6tgD8ypacv1nI+xjV9UKUifkp
uSucsSqFYrCcunkeima93mEPN/T29rHW+StO5kG2aJx/pWKoSv0n1aA+jEjEuM67s4bXrw2+e24O
kXOkp/ucj8HEvw2SMEpFhqh3a7dtySahGDHKqs1PDviM8M27BPZpyFD5OmY6bKYGVcu6qonccokg
/C8JgvaaQQoC9kNtc/2pMomSbUwdXJjzRHyFHilPPCEKA67jXHUegK6W3ixnrWgrJPXKAyUcmYO/
mE/tP7TFatA8qlSTdB8RrDfaask5RwpthskLTe7CHpPIIL+uslYFlb8ZgAPnJQS0NQwp25WFQw7u
K3EtYSsCsN6SDskfsmZhOA2N539puCamef4P3HoMidAn0YhihzGWcIKdp/lWDHLUMS6Y/UO/AShx
xjtYYPHuY+X8hsEOG8VUS7gbNLsxRBC0F8J2dYFYFWXltBaNSDV6xfGslD8on1s815qruo7QEhTU
/FZpMwTxTbTodubs1M3yBS/3yERZaVFWDZ5kiQWeful9GJ836IeKk+31qfBvOPisgTyT68yghBXE
s89PpE8OQo9ONfrVmfDYq+Q9lg/AmtRRM3ciliqB8VMJWOY20aTyPzXNf1y3W1uLGxihnOuC6eng
c+KjjHhX0/yHiKmaiOXySp8dQUwML+CrTlOwfw83u7aN86rhVaUr7TrTCRbPZpOm58qebdv11V+B
1OunCJZBKJttAJwoo4Ke32iC/cSTknZGDvw0Z5rc8YHQHQmy2mhpmnueaG8wj03C9EIRhkhLkQIi
OMC/BnaLYCUaS8KF/kUEkwDCFXPwhf3qMKeMSQOzPrcqjgqpkf6GTwRlaEyUt0B+SH0Pwu/wLPg5
SQ5sc/qNYfztJ4gFc1N9/ZwUor03sr63vWWNKXYAy+NfdJZUwvJuYOpi2NkjOL51z/DHNGPEP2zH
7Jd4H989EzCxCg0/XuVmQRG2lZjZBkB/fFBfUA2c+Gf1osEbvQifYGqSBB/EXooTvBKPBkrjXTdE
q++QMT/DcDbh/EwbbAZisvrluonfsXvhAk9/giXUVsuwEslD8jTupD2COtsk2mebQbSyAiLbwWSV
DOJ5tgDJO0m2qyvAujmDZ7qZJopuYJx0Ot2AWGNIx1TcADXEsdVug6tP6Ct9MBpchnwJFwy7Rxz1
ITwzNiUJoL//P2R7uRnY+qKL2+pdFu/udMzPhaGP3bUeOpqaxLV/OhU2Qn9oO/wx9ZmfRxVhLRM7
9yQIIZ5R5zkL5IljiNYKzTak2sClnjLj7J5kfIfgb3rzm+fP6fOKj3SdH28dUDAn5DXuzp6gUA7h
koHsaZ0P+dH+PRmphU4w+01FEffQEiIc054PEdpEnQV87lnBzZY4SjGM22kuBDMhJo992iocSrdH
r7UEkCwizp74NE0m1Tf7kviEoiWvG8nZ64yNE8h/ZCO2VBTdYhCzaZwEEmwaW035H/RW39iTGjuJ
DH3x3n+bqphgyOaq+c387XnhVWJwfF6OicvhaHHjLy39jJIF0g6MmvQakuduvqgjW/sqBsGy0Bm0
BprIsU8PBvO3HFzcqEBtAqn+dDAtv/oAJu+XLUmWeNXqOgySFkE5kK2SKrosbY/tmP2PkRpgslVQ
A7Og6L3TLyMqlD7vTt8/xpFgFJmVlA/vOpy+Dr4VEh4gezpuJh5YTAkV4WGsQLCaflc1ZmrxN8o+
taioMPQxICiuyN21nWOiZny7PqbJ1rp+OCtJkV9B/eJqgG2mRp9V/Y/wOKRbjjTLb4/ddRPaRT6A
ZXAY+g2DDtkdOpharzPU94SSP03ZW/9oM72vX4BmGZ+5wMvKXVxIzs7QwODpNnbpguOneWPxEZFd
pdfbDu3LaeOrmuHAEjC0PpqEw5O//TpjKnV6GotR0uDKYgUaqfkrBh1AWRjNR24s//CZemg7Nyxt
H34UOjMUhJ0CF1qelA+pEDkRlQ/5o4mptMftmFuYuKEmlD52KGjoluzfcEbaFSMkRouIUmvl3k5T
vgq2mP0dI7SDrtP7xznQajMt4Z07wXPory62yOdE2N15NQ/xzuDGTXN6wqY0xCwu/zRIDqzvy7a+
rwBuYv22yHugBdeGQSrgzKxk+/zUNFRnYRcB8MAEOXQlDu7St4kX6oQ6VpWWk7UI+NcXHiIh5GjA
591/TUtXIksG0jXTBx1n24+0wZiHtznG8xXbxJaZ3oJTn8BY33s00Y3lZz7/u3sl8K+kqJoSJird
Q2eV70jqlalBn3wQx1l1vabqZNf3OYSkYFp/9udwP+V6tsEwX5+0EKsPJgW0QrsuPdMeAbBhY8uC
F9Yi3eD+PCzApnU3ZWOAhU+O9P2WFooFxAdMUqUr7PtR0cExdSH++6zAT7uCz0JAhXxpuPsQ6OLW
2fhVfMmb13mEbs3DHGUPhBzlHYI119Fq131cElUw1eksB8IY2vyj42y14dRMTCS6bsWO9cspUPmo
m4zt1iCp+qN2eKeRBvX10jsyV1EzyXmdLQ/YiwPnnVOLHQGzjGwrGvDgYU2KfM6YGfxtwZYzmubd
1INkP0FxI7YB1YmNSbUJ2wsQKKzf/+Zumr2SisAhn+iOZVyuZAQ5WVDAmennW5KKcfcbvH4tZ5Xf
tqqG/8D18t9fc6Y9lGb1+6MHZ+wNxTqzUsy5NXu2f/ybkAyv8ehFqCKbV19oRHbh3hktJLhs5ccO
irWMkuv5SD9P6E6nKFRkqs4c6WiEjXAVVdg0qjmj43UeaPs+xEaZsCBULCXm2puHZ/rSj/DXsPfp
t8gcuC/1lD3NDw7sFVwTMNeOZFyQgkM/Agpq5DxoknlGrc7bJRZD3k1AJCPB7rQ4HoPjDsO+llho
6WxNRYqPtFE2hKxiq28SSaxDlRWT1HQ7ECK5tgPhFiwiZGvUntNZFWetZx5GEqwYxGk190tV4tcu
U8Xu3cZwhF5XR++eVgipLhhHeESy7BJT4Fe4Dyt2Hb7lsmZKk3xZKY9RN4jT/UDkZPVj+DvcwL/K
UJHJez2R9MFZfg6mz/NkCZnrNNaaazHQo+TTiX76K/3aHAyPh+atCuJwrbyUzybPDDJZ71zhSfOy
w1LHMThY7wxgeEy2E1iXR4etBs/6Yierd9gwCrQsIMaFI5/X1BYLWh65y5kR21ABnj2Eh9G++0lr
DHP/6qHL4NxDjEUWG2e+vGm9NZTMPYlzARuZCA735hao/RC1wxyNVKxuDwhEOOS8mn3huX8hQN/I
9pi1aUPXw+9E6+9d1pRAIJmVwFm/iL6vgs9bx5fXFLYCBCNgISE5eHSf9ARgY1ChHszwsz2Yx+Ca
K16+rgAcVpS8jSqi3s81NH/dXmdFJFfTp3QnangJYP6xwljkhAjC1Zd341cq6AM56zMFFBnFFvdZ
xVMHeqILl49IwQJXxi7MH7er+gsybRM+qVcB5pFd0iTCCtQye9RLTlIUH2G8OsX1m3AUMMbMmgAX
W2D53lTZHx7SLJX+msoy7wHOPYk96GA+5NGrx1zO+4bMRVBCuLZkv5W2IK4MLrEThz9PiRA2FrQA
LvI2qGcSRmgniTkXM7sog49Kmb6FaL2E/WRCB5bp+iB93WXFY3ZyxnNQVYBZCuY87dQf4JMArQbk
MQ9NFsBlljEQAWrhUBe06HJIFPtzsGcQYqFf6q0tm8mie5lX/iiD32G98/JUfw0Ebja5KosRuAAi
LnqRWLNMh0sVybGIkJvFueQ3GTl8Np97eEgPuV881zp5CXaCqus+s/UVI7uYkpfiwEpbI/szdCU+
evUeeDaK0sKhJ9CA/KSkNhygl4sMMLvNryWE43fH7uLzdFeYW5uax0u1GXTkZm0h41KtT09QFuB/
CSYFPjzfq/pBrx2qyF9IR/+pOXnHBQraCcXvFwqWx36yHlmbbXoHMADSPd5XS2UGnQuD+KPyS9lT
KoQCJ2hkn1GbXOM00O7c9tJ1vlXrEw2Wxzxt2K0daT6wRidCz0AUdRWsD2wMtIOQGSjc3kZs5aAL
CE5pX99ls58O1KpcjCtLETdaobhUkKTfVTVOPFJ1bP30wzN9ECEmD/szu917lCh1/0+gCx7CnFEC
s0Nm/HW064yyZ5Jo2k8ojRLcu0iE7aZq2h1ZSLNYvNog3aZOHUkFEU4p3daFhlCNxHj9MQ8jBxuz
I11gczbmOgdgtZV1ahQygLJf5Zw+VSDhoDJe2zNhMi/w8wSbOGUajWuCzyNusiWl6EQYGmzvZ6jw
tebsXIlwqc6+xTCruhMdwA7ZVtROpvh2/fGLrYi+oigIpVpVKNz24NWydkmcqBp+rweSQdS3cbwT
XU0pofI1EB0SURuHTgyAFmd5h5/QiUrMVbWgthKAqP2VO38KuhdlmSP1l+ncKac0gneAb24PNeAE
Ue33pY4LXEpiF63XTxqHJuP9iHqIxOt2VDA8WZZUOaeO7AA1T95ANZLjpsup1Oq+13YFc7VH21qn
1oVYWLU0vTctw55p8kpEoinHaveMBsHp+0wi+dF9y7gtcHJ5cIsnJc1O6dAKFiQqyZ+QgGoqNdNU
yIQKjOiRWYySQrrlIQm4OGrRdtKnQpYfXUoIlsfbeXiqAPfERXJ6INkbwnt/2VNL6ZSqHDivW3ZH
603fwJ5rWNgFiBt9ybY+a6Po2ZD8kJe3kp/FV/xk3XlCgF/YKkZVXuHoy9kFjb6dAC8oWim/cA7E
jgkGpglr0By0rfHrNp1KSW3xeOb5xV5doMhjbLblGY950VEeWaqPlbdEXr5D5GAYkrKDWQ==
`protect end_protected
