-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lraae/VZH6J0yMXrlrFYsblnoyAgPohHWdjuuoAF/YigEDxiZoNdG4sEY0yG+mteLb5TU8/fFi/M
vWBOtCAWrMlyjm9iKQ7vvZYI+9+BemR6uSvTwi7YAPhWQ2LzpWQf+zvi93rsgeTQsO3ohDJPwbX2
9nAv9IZLagA6UKcAiT/rCTUBs388VD97X3R6suXbBoWpXujJflhTOZgQc3vlhWWUqKYvCdIkd1x+
//cdgejm2Uw4IjQTT0C6APTSvTI3slOriibtVXoZIl6VSrvHxcqCbmCdaBLqdZ5a9WDF0Zg7glqq
VjDoLpEmmDhWy38wkl8MY9gTDR4hxHnNYOPeQw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
LRtUFvAMTOxKxmt3kT3YNdRdW1NEL39nQ2nHNw2YtH33bdSsmEunr+JW/ssY07Jvpigpd4P0gilB
3mmEwM7yqLYc1XIulKeGmL+kbehwSHd8Lie/VJuDa4SM04mcaZ8/qHCK3ZtiZbelZr2R2BDY0oaY
NaJmjHsKdWr+MZkC8bBirZXjS7okTOwt/efQgNR02VVQQNM2/UVkxll9egTHak5tP1GhTssxgCjx
b79YWdndRRh/vx5kSJEL9lDCldVpXncRJSPrzgs10jhkEgkMhz+r83Htrae4BJT6FnM5Cjc1td3t
+5MEUJ20Q3HozIyTDtq/XBiKOCUcXgQC5Z7nl2CC36jtLHFYN6Xlg/nzmaqq5KiJnWRD2vQReWYv
dp+357e5vGKFBZXlN5f41T2K2EkOn6Ga6E+RWon8r6/KWNlW9i/GzqwGt2rahmCBWCZrE5FRMlhs
Gn00ktCjCNm22dNDEdtJ10oF69dX+vwatcRZmtDBGYE3vkANhdyLgwQFl/y2LQLq9K6zxR96pTeF
29DTk7r1yOSkT9CDgvigs/IN2k9djwp8RwOmulB6LJTSARY9zPyY8sDm8zmw6HzVmCYiM2X3/MAR
gKACDxYuGteXkyJzhdo5LTmYeCyvkJVH56kfH7d+WxCN4He1KM6PflnOHhOIL6FX1XF6TqbMxKQA
atkIbOO/Zpc7sk6VywYuyeP6H+7Yi6t8QfEYkQs4XzoWJ8KcSwNe1Hom1wCkszOJFps9WndK6RGu
WVr1bjfSXsjZd+YnQZeylxb714LuS8c95fpVI9tXjRRv7e3ehTK0TK4KWCR3xWvBtrWvhKJXUcH5
R68hJAy9jbEJ8cEj2ii0YLmJTKo7Zb88ClAv1j/xMnM3OPHgtD5omf9KXq1V2eD2v7qMDuBOuvHd
53f7srximZ50uvGSmgeJx5HZzMf31lH5mwZUhqvyx8/xcOc9NGzJF31onmqIyQJh9FpT/C8iUD/j
wB0K/T/9bnHdR5sSO0UJqn7NTDNDKgt++cwGeGr3fUu6vgeXK7Deh+bLjJW3xHAVs7oBpOhGXaWM
uNmZxHPM+lyzbGNIxAUhtn685YnOEflgKBGzce7CW8elxq8YaSKitDjIyE9SBiqhp0qQ1MFZXP1c
r7EQecw7ZLAGJqGc8blMPbedAeqTX5ETmFqKZEwuLA9ib1rabCkZBfeJQAe7fkniJu4IPj1f9dVM
bI72gnXj6K48Kxa/sSk5IAYATIRhfDGh3zCaqCfUX817AlZBEQjUDr+FxFCCAcUe/SWuGymIIkU0
RumwFd4JSSMDy+OjZi5OiSpidrq8Ss1bGFqzai4IXU2eriWleTHmfJVJsuB7C12/Txi+m+vQoVbb
Wwc7HWUBFIqRfOr+QE9QrVUQKF2ITHcL6WgFKZlowem2RU/sbrzl98zCgFH4sB/6GMebwx4pbLvK
/4xY+3OyFOZvuXQx+Sox8jTSOzcTeRFeCBd4GxnwuIBpd17rZW9Qwoy7Z6GrIDKGI+tOfdD24jC9
dZHwQVKRofLIMVxpMHNmDwY/aa4gN32Ym0tFfwjPeUQ9dJuVYTFq4AiDUxPuU+1TykTPqMF1tmfI
EQtJMuIaHtV44PARg3FKaCmRXHnyK/P7Fu9SlaEa3LApR0Rd8FlJP0NB2L2f85w6gkd/jzmXj++G
cfWIEklVg9KM0LGL3uMg2NsqAZxRA5c05VJNfA3f3c0kDs9WxsKGG2x4vXGf/ddYB0idlQuqBA1Q
Zss+HRM9xpgKS0E+f5F0yvDIdKdfAbTOZ4gzZ+Rh+jF8hQRqUjPPFmDflHZEOwEwMppvIFnqTmqd
AsQ58BX7oPY33CDqQWtm+cCcdOKQv8ywnMMzc0KPGw9V+67ZoBJfxWDGkmEGFxUKLW23qv49PAMN
VzZ4ClwUcp/eDkAON6IVYW/4wp7neumioviKC8tj0W4iRQxNP2rVRfWlcGRTRcluxDQ0LqCv494M
JXEnLzdy2AF62loRmotUHHrzB+b7q//WrhBUZSqUZhD2u3wl2XcWNZv8AYZrIPk71NPyVeFj+0qP
vvkK60MpBpxFINyxSrs40hvugLPVOKguCyMsTL/K+83gYe17YJ1Shg4/3nGZsP6d5sKS72m7UPNW
+ZqnXA2rv1zSj+zjW3Q/MXPRafyd9406+NSrk1EabSy0lGj4IR+hCyJ/pbsR6NvPuc8XU6AcpqnP
Ye8npaW6jYM3Zk8q9sealFl1EGVnxdWv9Lbko0kwSQdiahwCP6w85ZVT0Lq2RSyGhFJ2XNv/7Tqf
nKmE11O/xHzBppTcDUvVa0zuV0ZDDyp53aLzV6z5it7xskpOIRTa9HRNCEzFiLVGcjcJmO88sobh
zrekiJPX8u0hxYJ6CAJu1i/1b24Gj22Hny3xO0/6JNpj/FJE86sjgscmd6pWi2SOtT+JN9paYkiB
V41vsCLSlaxWiFTNpWueO2olzEF8bJJR3QvAqEP1fCYZ4uSt4aRUXFsaIWtJ0wvnqtS0X7f4b1hJ
BX377ftLncltfI7rBIU6a3klM6vkxR9ZiVTUwVZTvb+d8cj3nSv1sJ75I1DNyBsF+1bJLiqdLEaa
d4mxfw3L6qRdlu89B4MAPNSuCwwDBfyxYZZXdTGnHQ3Z9hVLH435fxCWZnPEVPncVcGX5jcVye/g
0IQ2GPR8n13SvYast9YhlxyhK/Pz/gKAY9amzKncqgC86eWBLCnSWYpCWJEslz1o9M79Cj1KAyCy
deOKE9s3MOIVnmx2B78U+GHFbaqc2PwY6dCGzovpBDEYka5o70vXbslEpwTlDrblx7p9HlaE4TgZ
W4HEcWsXHHSNnuFLU+D9sGHW5FEusSwyGcJ2rnN2nZps01sFcJKNyLXUOdeGH8Ccs33iHXCIljdU
N5rqmWKYRZvkBGnBUi+skmqou+XwEqexrp1Ydcrbi542qLqlXcIbCjz80ZqmvSy+H2lzSY5Sng70
5WT/IhSwhqbLHkEX5/V/3pf52xZ/ABK/rgbOOKbUXm1gjxz+6nW8vOhIf7gRhpWKD4A+OVgxpizb
9OrggyI0XMDDsMbXPrV0mCiY/mzTTAa95zUIdVDdMZFQcGf97eRuGroEs7SmHjnm/tOPKjpQ1UQP
5eHpue9ZE6Hcd12xXFE5thPlSnaGUhOHwG7UTPFh3TVBEtGhvR9XWh1qqMpKI4U3HzBhcMQsnNhO
i4OlhtEKb3KXj1oZhljusvmDE1aZ+C5odWr0Y7c+biPqO5/Zn1G2ci5jwcSru0dNx9Pt0+3lFiBh
JR4dg1DxiOdOVzEefuFTPImvJochcmTerogvPqlU+VL+C4u1vtNkEsfU7xr92JiJAiQWXNk8SqUK
fkb+5fA8UFjcMnx64JLnMoMQKeBxUrdgS7cmEm3CMyg/VMRnPoib4LX8hsuVvFraYJPQtOWPi9vI
nUL2fPdVqxGPc9cGE+LFFP/o7I0UBKvYULrwsKnQ4vB91yXJdUe4fQQm0TVWLl9d/AxCD2nUrAIh
N6IHNRtFYCTESibwfb/FBwHJG3UDeZVCRU8F0MgKACltbqHKpFRWRUrLGCJvIqZbjWGkElkws7o6
hr9z/HgH7EigwWV3Zd/lgYvmGrRd9oA1/pIMyqeK5mqN3n+BzoDMPwZYDKX/lgXpdR3U4XnJutLE
tLhSj2W/mqOd8w/tiQGlrpF7b1r8o7jCOBHDcV114Ma6Nr6WY6IoSTWFevhd8bzE2yJulH6xtNyw
PLIC09Q6635FESZL2yUFUv9hatvL3xURGA7o3dLAeMNPmXhwNz/ThjNnQORH8akhesMLf1iWcdHB
s4qb2CFXQwuYfD6+8vC9teYN+LbsD/JGWWo3DodnAM9FEmDymfurogN/Tqq6zYiEtfAjEoi1HRHT
MSkV77xhXJwNOBztUTbnozfcXPirykSudvXK/DPC2uMzUbhL2M7lRQyiWw6aH8axzWTHPW/LKvDN
VgR4r9unmrRApozGdj7pjTdpS8DrP9+g2YDP0l4u4wuHEbC5GB4+KyZs5dacs8O8XmsWz8cEXw8c
kzo/Zup2x/fE8aLZJm2K6yisFmvVkz98f3Q8vH3D9JiiGXS83ZongWMxX/F7ih9fugDRkGZXimis
NO6FX3M8u5t0X6dR2tG9msj4vf/WgDxYJfT2+HCEgb+v20CJDw+CVx+yATyE7RcskzsUZCip195b
NDSqkv4ddVEOqel+0MDdJsg3wnwVYuDlASw2irDet9qUR2OsVuz57++6HhI77Db8tteokScJfflh
YLSxI7Aui3gzqt+FPyszrBC/OEjculNsAwNiQgwr61FdUVPGgxIJLmKaRIZ8VAf6CTx2ogREtpd2
StwKOVj+BFsji4KpEJ0ErxL8j8eJVHwzqT6FDAdslOHCfAvldwxDmf4GM5uV2HwcL6gfA9VVzaAb
cmJNO1kZbXnAIWpxhG95lqKWEzcrps6vWE+oMH4UDzwa8OcSQ6zxVr0P43th3BzHjfUfxK6r3cdV
oNJfIE2PK2cRYSGi7cFgh06b0utfQXQA0nq7ncwu8Z1OubnQvwokcjxYCWgM27W2p3xfXKvZjMQ5
N7yQsJId/P+j3KtTLo9h7k66oxhqUw6bii3ehKMAWdGwdVL7JoJ20p7NqTZDsb+MCOgmpC0beUIw
yXLf471W/Tk1CQAeJr9UjnmHysl1VU65wroE3njlxzBscfZft9uXeqceNTsS53a7jFysZLuZETuY
nN7ATDy1wg5gS69wlfomIyzmhZgIES8wRptClF3QmFMO5kRLx9882miKYTpCKzro3t5USowv+4yo
rFRO5bbmN6t2qjgsrzWnNv5XO4XwZqUs4/2/ztiAx6Rab2FY0HjwaPoBNXnv7oSn0s8/AxPBJVX2
uk5itaHE2FvWVvsMamNXWyXZ4M/9HoGXlkKF2goq+pKsIMTQNK7OtAGr3DVBA4rYk/SZ04gQLEig
aqqMUx5NxnZ751ZtCtLb4kfjdXBDiTWod5y/bbX49gQDM0bG6TtcL9HXQDWUBNhf+wKEBwQ9gFK8
AdMJJlFNa9Ylf/tnXkvuk0+PB8kn3jlVXkn2RMLj5f4/9AQzo2JW2KfVU+5rKmzwmapjZV4dXK8U
vOX6MIw/kQWxqg4JQmIyNwCaLtswyzZT79FdRPMfCW5EEW7vWllKS2uX7LbL1ayT9tgBNVXR2TL1
YDiMaGIINwnhwQD7lb47m2tdy2vs5IJ3C6kf/AwiYPtAKw66yypXeae9U2uRtQ3VMrDgS6W9C6YQ
BKXsWbdNWKITqH0UAB2JqKGvHy+gyHG1/S4+wWj+LFgLNkAZL4rBydRzscJbaCpGUXaRpCKsNI5N
wO4IySezzz7+0oZWfV9l5qPU3vVRzhLHP+9O/6EhF+CmEuAUEZ0fyRIEVtlm+kpriCV4o7agsaBv
5qPrA1/XHZYAcCyPfdyKPQ9zpmrF/nEDEwhKQk7X0U2L1KfEBn+xPuU4v0+PQouDZSV0V/v0dxv6
Jmj80zFqBoCnnFbjIySk0R9cDiY2zAuDoztwe3S71XbzPNWhGituqlzk47Us1ekBXonDAi+UMFl2
YOXYh1CuHNxFLDTq4QMngO6LRsbxisRRba8JHyyZt5/gq1Uty4fUUio5OyKPv8S6cyoyPAW8XogS
RClBIGzNaTe2gSIamfB/T1EPDn9WrzPd8/xOVUgKl9yJ0Jm++fuv9p/mAUbdII/jDLrO1tWxAwwo
UkCSggoxQPE4h8PVO/hyPAJEJc9anFNabMUpa2w7UPS2fS0fGM+YZ8sAdoOfXdihkTFtBeu2B0xe
kp9C/RTKYx2wDb4wUWK+xqqeKfRLVuww7hZw4Gr4d6Z4p7n49OAesb2vvOW2XRHkizuuMjs8XxsB
KU8S0ZJ40kmcuTDbJ/3byMXH++Wu8syz7idJx9wCb8uyOXqUZat+ySbZf9I5027UY/gRu8tFygz5
chr0T/Mbm3aHkyeQlpF6RjkTIqH/B+LwoFFM6Piak95cbC6Nd+YlBlKHFjUVup01wnwpniZqPwTZ
yo6CZSFFf8+Ef2E5NTC8jd0aj69/ntJ+ekgudAzVFyY79GSQzLMoUiu1UrkdSltVVd4VAvkWUqy9
WArtIFATvVf2GxggnWUw61i711mPY1n3kctY570X0uA5AHh/CdDQ/twQoB3sR+vLusl/E8FOX+M6
tU2rz8JkAC6CYXI/jb9lJ2K6SPg692L8WoRYFzNIaD9BhmQBEWbc/4wWl5dvVO06puSXL+iQE0+j
VNm92FRq/PU3Ng3x8J8UkHQAvhNWZVjwPcPQEoXyfilq7zbD2gTV1UH1VdJbDMuN6Z7/bvgLiHa6
TpxiH10UlRNQpNjTjTKoDaZvHOz5YQ+8wPzO8lh6hdiCEqFcWGP/DAQeAcGb2w64lRItUDPWvcbu
NIYxyO9U8t6JTneikdl2klRRrJMLtf2IEPazL29riAREEyYbGMRy1P1H+ZXpkxUQrJMg+hTWpcbq
0ffv640ufSfKLJeS86//A/hECEtT7RX1pmw/L/31PC6OgENOXO53kCk7xA9hi82bYMKV7VtVBBpv
qn3JglYE7lFZEw6ofIlFtUQUB46VAkuqz3JZqQrLEQBLxKCSRzxeLmA2kf/U6lAqjOz/CKAriMy1
DmuhHhRcW8QkI3HdwGRYVFqTgl0KBsqNZirjNQxhdXCKXBKVYJMU3e0rM1G7ghIh9cLQ3/CEfURk
7dOHL3vc49NfaNpp7ot3Cwl2Rx0NElg3A6B1M/AbaOx5V3ClkwGytrYUy3fK+jzGCHEdaTE/l1DB
N6h+5WmfBivLwgF1dOLlqD97GLW6qxRMR2pfsn44ZCh/MobVU4N1WjSNuYYnX9Prq5omw3GYz+ky
EiTSvdrzUBge8Za2FiAu+x/OP4BWTQJaMnc18xbeWKnabTTa1rt1txRuB/dtEKqJmQLJJ6KeGwOc
YIDmKOvravYlpi0t9HuSgSi5t/JGSAYIpfpn2fShEKwzZzZLUVJHA5fLaiftxkwkEso7rnGNQosl
8Yos86+ixhZYUtM2lV/LX2SREwooza67Zqycv6SjGokvG/sT
`protect end_protected
