-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RwWYxOfJQno6DKVwZVBcyfbfkx1yrpmtyss9yKO57i3reU9d3N5JXqgmMGkMMNc39TEQu2Au9bmN
tcweCEcM257soCuXvGjY0o+A7PSeKWV2gk8I7+eW641TZ04YJ0qcqstqc1vCs7hbZ/kMP1h+aeg6
dwdVtLTtEs6GPhi6WW7HCVXyuWXLf48cagSi9Ede/sEQT/1VrASRxxeXH9lmCL5igK70WzOlXIBq
rwXK04wDGQMXP0Is3tQ0QhjFbg38DmCjg11rBn5GBawRUBB2bJb8BJ453Z1Az9aN1isq8b0T1SSa
oEbmcKPBjiLMGdhV0ZRZGo5ZHsol2YPjAE/qZQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9488)
`protect data_block
y2JB/oStkbhXTEFGJ1ZsXcVa3grjLzV5M9GOTFVHvGmxnbBPE6m3a++DCxH9cNi52cRzMl0vFFil
AZElUovhNXOGU4lZbn884BoXmAbnbr/d8Cwt1x6II1Xq9XF+BKVoWN1mieoe8k0c2QJQZVB3XbN+
uKf91Xf2IASBuQqxW8OS4tX2mQWDyzsas3tTTyUIsEVQ+gzuX3opHu/syKRPcWP7XUBioyJHyi4/
bKi3kMvwTH493QjJwb7ai2Hz6ndRWspY0eBb/ch0yDyC6RguPgFtSk76MQvS6ucHBmEMnr6r5lG4
TWzePsMGm93Ny6BxbZ+9tZuuJnDw+mXEP+Qgi4jkWDXcwZriFhDFD6tU4u0Q67z+M+Us9N5azJ6n
YElB9ku5RibdlTYYTj8mhKcVxy7WfSbnomp8AE0p1Xh63EJy7PGtSmIRvgFUjmV8ECUpNj5dMm6d
7PK8ddgg4Zlxo5NRYPwNs44HOr9rDIbJQJSzlbaG78/QE/6AutrcViWq31vKZrLCozbLD3YMvkU5
yFcXQA8aR5S9YIr8hqVqsUrbbgpglk3EDPSeP3bg46irrbYMQ0tYQE3BLadlrtSQ8MFBAJC+iiDd
sIe2Jkwpy845Pa0Nke27F9nm5l1rKM9k4Mn+H3xXzffzKfM6s0SSQDJ1lVmUi0J+Nebz81gwDjEQ
m514nhkdbcFA34K0xXn32oc/+4eTkZmOKVT0uQAPaLr5q4/Z5/XGBkIs2/c/8LUh7dFtpc+bJLah
+5PKcOmJzN0FsVh4KbkEmj/NgfJa9SnPmdD0G5BcVIPC4g1cCKmNXS1L3xE9fu8PcVXmE3XS/5cg
O3QYLt8uP/fEiKzU+fddDiCTy5wgHtZJN46sePevCaJyV8cKK0juIr4bbNZG0LgFDZ6YiN40u01N
w/QtHt0oYThMSwKLGMGzx7yx3lDLPUVj5l8nd21v7Dhhq79xY4jbiZmtQ5gBMpfj9gQUugieZ4aa
fOiNHAjJ6v0Hyzvk2CT09ftB3eNE68oIhWXXz+F3IBAIyP89HKiXhlnqNa8dP/jK8+RERpKN2w+N
u07fGHpYGAokOdfhYGqrsqrVib73SeELOPoJ397NrbyH6kKy/R0rgwkmSTluExpEQ5P3FDd59prx
lFwdFC/75mspxoIoo0odAgEzQ5B7J/C5v1nXHZRCo0l4QnCMeEwnCbVk1+JqH7F3v3gXEBygQszB
zdgaUsjkdylDLmc4iMzDN8wqh4xlbYKn62rWB7Sx0uLfP+dqYHkudz0Fz5VsP1vULo6aft3ub+eE
hDa02uoci2IkQll2Ccz+5rd9JBxqyUQw1+/j5hojOj233OYwkuMrbDWb+GPzEhgI7/TjoOsfCnnc
DwumzwGi2EZCbE+BnX+EU8yysBPrLfTDj6F1fb8YMVLb+Sqcpvo6MwFeV3uKJiY4NROMPAImqPVu
1UOPaMGq+fqOwxKHRTKUboO1Gitm6v4e41F8hh6Bot9uoQngJAA/MV7H2hocO5MNJsZoJxh2z44+
IM5RdXQvUg7kx/A58NSiFtSgyIjtC7DTUf6sefdzr7DBRcS+Ip7vV1XgEICU8fhii4VDe4aN3TVy
FQR74pyFjeofNJi5NblnvmAR2VlbmpoeZzqm8nfGL9SRKpjkhiD9vY1xemz4F8ELhtRBzlh+Zt2r
NjgFztjZ8rpvKL0VL76hgbjbEj41HnwSmqHtfhcYWxq9u0Oa4aNJiq4rt/Tn5m5jqvUU+xbyKMih
SxcRRKqZNR0Y8dxVFzXxDXIImzNt4ybcTp/qbL6hQu67K4a6oiU2H/G9WUWk46LTTIHQuiNsus0g
B0Una8kSCa0yznMIixBf08VFXYqz6YCwO1jg53jhZweLwaxruaPd0m3cT0YhGmFp2ASTxFm2tC+h
6PoUnX26PeWygtcm2pCBWIGM2lPoSg9sGFMPRYrUM7SAxbJ8OiG76LEaVxVPZEH+zTK6IdDlEmkZ
mpK0V99RdurA4GbyD3T6hrX3lbdur2LwrvKV5SB7BLzozvX68PBOZAaDDUykZBjMiqqeRJJPxMOY
j0TTD4mG9mtZobIgRpOzOE8ybhQmt3PO43QeU7GIL0V4oEgnjHAjZSnWwv5Ctb7Wb4KEpqzp7ejS
i9ZPh7WUWM+VSS51+k4LtC+MkTsVGTQUqq1KBKVts3cxD+t2mVp8wr4myuF7sri1m9jmZgAQRBGL
T1nQKM8w5OOHAn89NCWCuUFR6Sl+NoGPEPGqgqMNgY8uMKlBu72adXHxEaJHxkZowT64tWm1nLas
3Sd/UEV6/y7c4yQKj+fE4fWPyOOj/MqXErN5TGLWlVQltLKq45CwxVdF69C+f1j/e/zbbQ+xfMCC
sQ77W8gTSAT1oXDqJAXnfChL8nE+Xfp3FUkhMe4G23vVw1tGLLhayfoKaOnx/umzWIL4GW9W/1m4
zQ0JYtdD46Exe1h2W2J6Lj9EE3mUXwLlTNUacTiD3WWBplJLehFt4R+EvQEJLe4C2uwL6SMorxQN
ZdhctKpuVetFDNfIIpwruC/hEFPF+0HRrrQ6sJOrcec/X624uTTuFWwW4EtPlWb8xbddlkg6/O8N
A6/OO3hk1IF8LeaD67lX92WfJQp63T/Ct6BK/tjrhHqf3YE+5WmGThq263LTZR02/m1unpSkhypT
Kl4tDlVhCJTIgqoV9r+1EkDM6+KXAHT0TKOIffnnvKHoClQgsFXEqAZ/vGJJvXtEKCcjO1YBtpMY
g3jox3q3cHoSAfsKGLKWS5E/0+Kp/WeZaLt/RTB8xss2Ae6cKHNcLklBLRn3vzis/R0usXDWW8Ng
s/QqilZCc77kpQ4Vx/fcUuuF4CaSrtnewgQIzvztqM8vQtVobYBwqdehOkMYegHfcJdE79E66CFp
CBBjoKctj8pgAnDEcWLR/EmEXpLSQt2tCv6pP2dIntaCsNTDGlfhXy8Xsy++VE2D5shByprWoFar
VZ9ZoXX5A4BiFVTgdOHVuy+iyOy6S+9busRPUQ62lBJ8SkJyFWwzAhITqgFJo2nJNzxoeNh7xLMO
3RLteTzV444hvyNl3FjMEI5T7xQMavEPQx+jhmnvTEZ4Bd9DfSZINZ4Vhk+bg8mCFk4ydQx2Y35S
GrRo/X6eSIietc35K8WApEIWsIMI7LN3FAAmWuJMx3p8YtjIfHgs/o9hZkI3ko0R31wxbdB0nnsm
bcQhw/Z1iS7JDCI8Ri46feHpdKEoA4iErMr+aYlMnBiij5mBnvDWCyI3gaNeZdPfL3rhkBhQ+5Ex
r6Nfm/yeqHB8Pb4ngDS1kMhDs/WstlGuERBqt1YHnPVZM5JpQDv2Ch2xNfph7ccgdOrPD4afiB53
m+FvaBpZjJ7nVhna4ABP2b/EirZCZc3/VHev2fsZ67HxTeBva23fbNwFMWXadkNp88ruPZUaWIaG
swYHOGWSyJlMlhkZOiXwev5D/j5nL0EVXLygIDT9pldm2rFBJo/AGZE6Tzy2JTVEK7cWJvN4imf3
0YcbVpQRdbfVkwaAJYzOCtO+bjx/AaxXaYW1eENg0p6WsxKu5Y5gSNY+aGBXMVlQXvPDEvNHmE1y
ckGR8Z/A7o4yzyOwVu5mwWVZHMNki4HkqxCcVYriaMWoDDthZ7WeAwBJ9BRm07KF2jMtWxA29rUO
Qjc44Dh9jZfHPyNNkFQtix+VCIl+8XX06sN01tJDI6UggOPl3FSeGoaOOU/ck9pMt3Z48k43m1G/
GdUCnQvgakgUDeSGO033eQmi7kqHVJTegrxEU+/1qSMyRJF18x84YZD11SwyinG9mqQa42WHlqED
DNKgpNNSkpDEhKrP7/ES6qyKIArFhPFBZbSatnm+KHVfMDWcvNwiN+zWXYCAZG28RIUMpaONk9Bq
2U28gUq8WBZLP6xug4uExk/8X4+tBznTzsn6neK1WrBtF8MBcyLYBxz+dwOQiJlTYTeJTkHZ61mj
vf6GDmiP4UgAS0MlyAQAFu8eunjA5Oh8pAQLgCgCpX4APR9wTfT47M8f58dMkvkJ4b7/A11qnvqN
2l8hAJ4D9UKhJT2LPmsZbew8fmNKaeiMFTbGI/MrYR7TAvvmBvNw7KKhMXQQgX7RXh77vXRK++vD
Ml1vCr0fV0SO/Kx4dnIgUdoLTzuR3k20PX4Mh9y+9gTbHal4F+xUJZxYpgCeci8LLkcX1aZwGchX
cY+c3nzZ7vKNTbDivOnYlSQ4wKNy+vylpbeLZ73jcC5CMLHZ9/p6tIJaIRttvE8a03vMo14Rr6+d
OYIjoMP0u+E17XFXCFMwFeXtGavqQhGm6ya9EPg9u+DuehpPyC0f9hO3li/LL/+LGB2m3xEvs/dv
oNhTcrtLe0OHM+AthiwAonp84Br9x6luyOigwIAKjTNwbQ7PjxsK85rc2A8aDGkm7/PJaUjvSeaF
sQM0dB/NCTl6954WLTR4G5+BWMrO9yKCizc1moV/Qz9hY7EqL2FKhhxPa/IVOUlntrTU7ZIQCV51
YoWR5y94Up/uz8nYifsTOODEuqsPSj+4oUkg+3iNB/ONiB3M6qaQc1rqnrs5YF/6cRbcNPkKgDjS
kDJexI1hO0PDvzqBrACYQSW5snnfBnid3j11K2nlapInTuEaDc4UAzyweQo/ttChZxGFACc0yg3p
BIsDxGzE7LqKrVRvdMMYaqAhW4il2+5YAdbkzKEBeQ09Nx8NN4toZXTh2tZIgv6mzGrnOY6BX95w
QxSMbNFjiT1QmWgHDxBRfeL1lB7pwf1e7OtmyPcNlU9uDaLX4xEB9cJkZ/XWaqPvyyNTAGV/aD5y
QhU3AJRGbWU78wvWB5cjwxD9X9fdT8AIZ0H2I8VcPHpaxl88MCZXJkapmFS2tKW4ozTYDJDIIRPd
+C2myrGJrISvju3OfCcOFuHjsAZsL9ATg//FWQX0sJ5OQDkcxiT4Ki2upfHcOjsKBmDmVbjISLI2
v1AvRY/q879/gmo7TSI1yQfgbfK2vaLDSxOu+GdGmw1xP98fo4FNGUptuKrW+f06WtLI7rGl/jV2
lZdJ0DlFcfjL0DX+Sqr7TWicoWQ3ZI9QBz+3yF0moqryx0rbTcchpKyfGW5YoeO+T3a+jW+avSsr
fVr/WLoCRWe7ydy2HeEwwPoShdotimuVnmB/TEdSj07o7OicANzpeVx2MU6g7JAXgs9CthdMbLpt
WKP/fVZDNiirTOMtjU1RPIGJ+LTWGstY4EICpRqLIovv2U6ZUSutGkEbv926iEk7OTOGqu+BLwEI
kGqDRMOg0zYLCjMbsAZdRwYmqY1V1q6Uzsc4yQms5PgZhub2G6Ktb9HPXrwB5fMxjd8IECpGJbtl
ErPJzSlnMLH6A+gWMS7bzKF4oK3LUwSf1jpydg4aOMbg8BYk1Y8QqMrO5PkjT/L2ShBiBYfcpvJI
7XoX/GW9sxBYa410Eea55K9AqXjJ3ghygimtnIZHIPnoKlbxFx07lzE5TSmuEEGXefSxxVjFegVT
GtzChGRQ1QVXI5yjuseQ1QgwKtNHGWpPQB3ttkbytDuzUrflBjMS9vQ+6yckk12N8ktDCj87A4Q0
2d6ARvmqoMVvuHZO8v8puALH5vI/qsqEDcquvZHZzCh0nDH1dlqMTUAClbrs97G63Xr+5SVWv0VO
xh4Azpz1SCaae2IeC1CItmvUaAFZdb8Dk7xiA22+Tx4g0cRLmjXPbVEcw2mzmnCO0fhjFqt9L4BX
QeT4MNUF+rZslHuTp5gMsUVlnjq57lHeq1vmwwTQFI0Qpb3PFoBsGc4YZO8MC3qT8I2KDv1/3Tit
fj9BGq3/eLf5D3Z1D1WzMfyVBRqUD+cUUmdT01gdCdB6xqgna8Z3Gn07gBuPaxtxHNDNZazSrJ8/
aFDIPcLmBFbsZ+eys91Sy9397V64lYtao8U0oAOgQK2n9CHOMtYRLbFHJQN9pk8P5ahBBm3NycAi
M6YFuLFi/NuwtAW3AgDJahVidGjJxM94WcvK7a/RqRajINzLGwirOJR+FwMerI4suuUa97zilnap
LME5s0UPtu7aBXZ3NXbgich+VogC1fDpOyJ49FFfbphONXoeaewetRCmKZQhkeJyVmBTbwWlko0f
mg6Z1mbSc1NfspVyA5kEG341I3sAhK7aESCMKrh+ry1U1eDNAmcqhi9i7V0io1HFYOo6lVZ+RfCE
k85GWRCmX2wkEz/NVrhNoktLal5QUCFdKu9TLrwt5ZYrWYXfbSTU9tcuym2wHYWXLOnwWBvgBXZM
BxieD3RFfzeRDaFnS+eNIWHY38tvPT4nYxMd5sfXkwMwaXwEY2YrJBhEpM1T96FqO+3DrEPIhDsj
7tcIVFrHAMzKMrFbNh3XQQUQOnEp+jOhSi6ulZ5HEO2Oi69ImrakVaeM045hAyDMqdz/+RO8h48V
a3i8/sJyc5CgPAAsPwyUoZulH5wuK+cs8i1ZYE/eWDHW7BR1GXRNroe69ujsjzjZfVjKHCq5jDDm
00yusmCPqzF3DtIQICIZYaAFpIaXbG3jeziQeYCiQqtpcst9l+9DZVdVOdXrELQzC+G6Sph1flrf
Y2do+p6o9AykOozz74QfI73UTq4Q0p2YNy9SNGc8wIGrkXHXXGDA5BBiHOetyWcZwMzQzyP34SIM
gc27k3s4JXhX7h5TmHztKDmjzPpZK9+NsCeWyrSkMwegKMq29XYPEFWUXYyO83UZZXZ67C8KPIon
wCtj5QgaZkUCX5pEPRjoQKdcyHlt0n90MbB2W/lerT0Dub4TXGwPe2zqQswS1VwWtJNCuKDryY6V
uodnHZxh4KQ3JP3V83b5FLBIeDesdenspuKmyArtHPWxIN7Q6QHY/ab7c+BCE0T2ph/7wDBySG1h
lqdn/EXo+l0ewSGdyAHcvYFB4655NjqJg8MpyOXyM5CBCsh9tYO1IK2KH9LJqHudAjXzRA3J1hn/
oIPulg5DXRfaZoIUfMfiYNe4Hze7PiqLKAnxBmMrSLLLIBCdb1OfULsldMlsSCG5FTrMwaggjnjC
dghW82vR+wmoGXo4rBNryk7L+CXFQQ5TZlHgswGNCwSwfrw91OO+HUU6iQCY1IQm60DpPy9bmxX0
uPFfadCfzYK+lsFyJgP6qIy8EANbjU1//JBpbAS31Jc5i+xKzvrYiMpoN20t+V04pTEMg3ezTOaE
ZGNBVwjXwi7VRpriw5RkzhwBTwe9MgRkRfBAPDji8JWehLGA4M+zuDQBEU8KHiQiwg3wX//b9W91
87NO5aQgNpl5uHCjEmGrWuMpSn7pSXHWWlpKtV22izm8xMDgfIqRwZFkl8zea7GKLJyR44PSu1Ke
5Nztg+4/lsC47O8wx1vqcDVCtZRp/L6yZjkvxfyk99FQ/5/SmGR4KxXZAiZ+ezT0sLdtWUVo/0TL
7l5X439JUrzMxQhRpsRAFzM41UuQVRC0DB68OpYsDea6k+F928QKMAxQ3qiKseGL+4wGWB6o7t06
wE1yfCZKPPmKxGIBBprr4twpeXUYHoMHnbLgE+8YXytJAJD7zDS+Og9tObotUu77Bvo8QnMP9eJN
dkEHWtTQXABgPaGEGg9fIG+CqgVIR6KewO2E4pLjWqqslxXDDvPCErTsU1CS8H3tAVsxEr2wuHK7
X10Gu5/FfOno0OaG5fGYvGuO2luEzpQiGCPHMsCL8Ghp/fB+0qZnko4tfnn1/joVFWqnWGJtOOPA
Xrq1UAaadbAwgZ9y/gCxAuq9x8/PzDaYYIL0ioKCQQhBDCF4bQky/hV1m3/lecTPmrFir2UfnvjI
ubrtegQWJxVLi8cTgz03B6TavJ3O8Mt1PC5pj/24mh4+IAQNsS8DxRdn93XrgNevcvTfNhQEl99Q
ZPfbh1WTQ5lb1oPmMXXYY2MpfF/4r3lUHpTRrp4Wy5d0ZUNfX3GuA2YamKrGcy97BbkKBuo7epoi
xhxYG+3BgzJtJd7NoEZEODcoyzFPvWw7Laaoz+QgCaMY5QVlHXeDfX5ZsoZcBPIAi1oycFlyufUF
3Wd9UJl5Vf1XbB0727RkdIC6uVcRsF3N8HrPm4z72xAl7LablyZ5mX6xbkWMeI0/qW6NHACL2xXV
1UwXC58lmKgIZ6gF929e8qUaDAji6LXORxQ6pI1gYaaFcm66azWNsgXLPRRxPkyIV+zvnMVpuQbz
RvDpmzinQC4KJw6tB4xAQ1M8+RVQREHl7zntyKE2yAYyGqBbB/7zFLpTqVjUSUYRxhngdMP4Io32
eNWfo/syP2fctu8yGI+0IW8gsh/0pWLjOUE16xeMw1r+L3L4uVAGOsXB8RZUwP9PPyOx6QgTlDwI
4/p1NvpeC0TJBKfDaMryyPWyrV3FEI8NwNdP2V3Coc80W1M7xCwQt8xFZqhxMWcOMgjEqSIbhSXq
UvIXOTZMfstfkkCr5O5Hq2zqpWdV31z/opm3NuwJd08sRBmBJRYtP41ngvjy1NEaJtDB95Qca0oG
iOrYmV73fE9kqvC8xB1S23hbcpvPf8PHq+r2U20tDE6FBepDxD75jOXSm0PKq9D/2yq1qKBPpmUD
6bDFtmngvAkGdg9LjB/AtyyR/IenqnmAoglRzKP/dHYPxNl/uq6j/jLJA6Xf9Aifj/e39khVcNHw
cZAVoDrV6nvM78vzpQC+H217lpcqVeWe4ZbilK1XCYnI4kVhZ11JapaMwYDCYELj7GYpEUTczTqp
g3+6vzOdIaJ+NIETw5O7t4UBDPMdfP479x1J+WrG0Q5b3Bj70d9l/cW9ltLvyKekKLaiyEUlcMv9
HbY3/7x351GwLxdJEpFukn4ZZ+P64Sjs1rPh7Ps+GxzuGXKfpX8tMfwMdjstKBlGCwLv9DPFktOB
yLmj6GXscyVw5hqzZ9YsUsJUS4aLEPQxcHvaieZ3WJqCx4mjdUYg9DnNMxElFdldq/Ew6npjaveJ
dANdJyFGhc1WNOdRZlasyE7gXMvM3ITXht8kQwT/mjVH73DqMh6iM1azutV4zDdYktrMbm1cYGLw
vFLpJitZlsUsccG2z68uscD48ZI4MvNQWu1xIIg3BJ5G2DdjyQTg1NamNOG/kxTQF4lRjsKD2Aea
jvxDY1LP7JolbLOpZSnyxUWFnFaMfhb+VFF4tmGXnEiEQITUbo+BrRHAcNsiy4Kr7Qwai7J8jqBH
/FgGZIeC6OM/Znz2l/c10CahXBoPzUk/kuyFhrhMtXqAXic+viA7+PgcMRqQmNqNk9ro8fgxGRze
KDp1myroTdKxV5czPrwN/PXs+cKVkq/RPW7t3H33WKjpNRUT4LP7yvxWiIoC+eiyLlD+aYuB1WBg
D+MkWNOVesYqJpBrT3qLfGxATsqgXB45PBmYMznb3ZGT5nwsF8aAT8AgoRanzxhjg1yJVq+DlJZR
8oS67RbbXRWN8HtELssysQ1OWdAfHCzzf1aTPEN/KfRJ/t4/tjgSxs6JudaZO/mkGKRTIYz8dQrh
TFjVNQmWlB2PUnxEDZCBOyMu2uX6PxzriV3dX/z1b4E+Etzgciviln8cW3pgUQV2tzAzkADuOpu4
RjbuAj0iz6hlPDFiCldk/1AeD7/aW/M6tcSGCASeEUDjxCrIluVA6PW2bwCmamImebrJj8jf61Vm
dRiTna30UU/r+Z2hppfic1j9li631b9j0IMLNV9diuOjxyjV1KpZHqqFIl/s7lz26rnt71Is509q
elvJ0m5zzCB0s7TS6d2VowHVh7BkLxqk9/VU+kva2wQa3alASL6psnI2s9R5Edv2jkRNBik8PDxp
XOhF2psaygozRMR0Z0KsHejvtOAYGUX+pVZcVh7JLrEhGNaG4HIXL0ZUXL568vazdSE3gPlUojDc
7CBHoBi4PjazRv8dFMCKJICIHorkuGSVdixvOt2a6/k8XtBuOfKRn7rYsgoibFhyEKo0/67Naejr
lS6VlQR/GnihV+EmOyebm3ZwxsypDZq4RMzXJt7Fj73Yx5BLiJpU/Cq2lt5vJcVNKokSeziylgXQ
HCxoLPRwPAzmVu0OscvBYDbCO3efG8+i7JoOmoaKI7b/NdLCkUuczmvxUY/hkoS8xT5dWpsQDb22
m6qsho+Lv8BdKHodj+a7OKNFuwPQRE2DROsla2ENGsQh9Pix7S/xASWrZBL9JPgfTEFts4qbpFdX
fjxR/4VJnhhXcF3VfqKspcUAMqF5Lbe4j//s/xcUuOGHeshHCemFLIE9NsbmSGk9EKvsYrRYpRIY
2D7eFWHFfjreN3eHnhHtYZhIUVGXYTfLQ4H8TEo/Pvxkjkmocs7GiZ4ZPBxcXt1prgCWoHe2ZQbX
oNGOHqaMxk2RK6P5lBkZpkRADgJwRzgdiQ+jb95jMKcyAvZzy4FusUtlwTGvu8qh4AoR95UNNnQc
EZO+WwDquSP7KLUx4po8o/0mzMjoMQtpOdkQaF6N6SApYPrukVSFbkItz0rS9Vrqr1bZIpK+SPIW
QIHcc75O1GJBYi5f3DUD0RTGWdJnt2MPg2UPJvgLs/qvNmWMsZdyj8fu7Gs4BLvYZR1RXiCS/Gdg
F2hZaZ3WA88AVXNEt2VO6460dm2raXo+xQ+BMckj8zLBisTsJuhzLux1nRkt4nRajUa3YrJcIPK5
PL4fTrVn4Sva3ZWZc4wiVuiy14CG90UbOFUGPDeAE78B6Imtn46qOMD/8R4Gm1jF/g2R+A0yG0ry
aanQscYIQfq18z3gM/eVC5FcntcT50shZHG2CPgSrJXMVQfM3Y9N0mshA0ykhGg5nhj/MgYSzZ1M
k01q7PBvQv7z+rIYcoyrgCp/yG5QM1v2VRwphFE83T4jS8hE6gPr5aUg/mjwyN7rVmXjXu22Npbu
rdE1k4dfYrRiJlhZlcHylXfUcchaP5aKb0Hx1XIz2kY35lJIaq2KzvR/kEDX8l8a/LJP1GYn37BO
O0iFIWGhP8OD5/ludi+VQKiUpK3Kld2ytvUTDHqbvYX5sHbl6KxCdKJd2hRIaP+lOR+e5SqrkpFV
j35D4SmTsmPhLqlt6qnm+6IT5sNH4PbKFq+72ytlNKphAfWAHB+7GsRU+LReIvaEByj63bdcyZxE
KcyLA+qKt9d9W7ko8GWjx57QaHxRr73x1m4C12/+8cWRwSR7GlacfwbPi82Rl5bqJpyEdp9RIxjl
7PzxKCBlqiLiYAHwYoD31fBLP8Gi+gO+QTQrzhQr7Qo9IyxCzMQ1m++Zn3vpB5qO4bC7J4RFG40O
AOO+tsJKOH778bbKDQGZbm5fA+u+VPD/yj7KpC3moyiubw340vLpz/YxnzZarTLb9IrCeAIri5T2
+RljTbEAYpCkpsWGQYAx8DT4DP3uSqHclPZ4pMjZWZV8AUl1E8TyGdgpVbF9qYPgrGPH7zaXtgCs
+cwUmMImSvjt6OXMIZkuhs02UgDm6AUBVtFSZw4UmA9EFxAyownaI6o9rZBIbZlIhwF2H7nL7Eay
AsBQtZvATglrD6Vxj5X/6skrFxUM4eOamWB2ih5Wu8kJ0DCvtLVd6ai5Yk4fyhspS8d3aFPFU14T
aUBO46sQvWb0tYA3qKcmn/4IVdmuYcVYWgqlOdY4rLmiLU+xCzRGxR5xuvFdi9aBCl3tCBTGjVWs
6FbCP3RsTPC37x7MH3Ru3WosMSYLZvX0KlE/9HQmBdIX7owtvXoTX6eGVCxTB2CWDI236ye3QBay
DCfI5wf1sop7WQD6ZbGbEJFT9O7GX/9/4SZaFZtoCCDDCYq7bhKQvoskeoEcI6wln6ynyGseYXHC
Xedkx9cPS/4Fd/neDCxDniz3svOsXWeoHUOdk8U2aQ8HjEwWQzwfd58u3J0/uNKIsqwZokm4LxBV
MAyqCusyg2xvfAJ+11hqKINqt2ILUw3drP9kYtBbogMm2LPsiW5U+9leGvBFtqO2uZqIyKwvi0Ns
Uq7lX/5cVysNzpN0dvL+a+30eF9TOR6wIXdURJP81bL022x9MyO2FekUdFfF5DtzF4viKmnKICDb
HnYK6W79NdKQ3AGytCs9QYVUNX1kyrzNIjvFXN5+RArghl2uBeGkb20ERlP43NatgdIuuY2saRTd
3rzWqZ6dHYZBGFxiQMijxfqcLLWo0yhqdsjyXkSU9ATRxqF8LQsrSo9K8FiEEgGvuqHqsK43HQrK
Ald6i4DW7D7i41B452Uvt0eA2MM34WC0WlrvW0ryYI72hYjtrNa/exnCAYk8h832bQgZZ33aZYvL
qRAoN/476tgmBtcgvwxvat77oSKNifztzOuipytOfRsJMYfiEvwKC2eJ3+ym3zJlBBhaSwWMeNe8
A/1R+EJPQ55PKS51izSn1QSVLDRtD1mghzLZulelCU0ecYCe0IkD/tCojOhdWzTWVfvPXUBDFpdr
nJnyi2KofDDKvojbDXwC+jfG/UmfI7zyxvMCBR93Ucy5l4lh3UBv6ssraxDF6FLYM8PuVF2BClEG
ZSKZ7pKBvC/IoHza1U+ZpkSt5/eWGiEgtl8q4sG8c5FnfzSqiYadJ4rNJ8g4ZRCLhEyq1pLZxJGm
ujvx6W2HNrec1lrhcCaw0jBjfm/DiZZUSm1s+7rpnTg49Ch3rwozjSGCQcaG+nFZFJY0E+0OKTl5
ST7cTwOuNO3E278K/VTLwq595XGR66ABurDCGg/2R2aPgg1LZwiRhzVUbQ6+Gqu2kxZ+iWSHHkrW
q3l+m1lIHxbgPjOX7ioyixln33jc7MB4ArU=
`protect end_protected
