-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qIgi+zFQoRsFSt99tjou7Ktz9TmLPVR7aXrXaFoDLVdAy0JZ2uAi+hjeVRJQOoHvRu+rwFDEVYDi
RtzhBJkt8SnZGzoZdgIR0Og9aQmEHIr6FDif0h+QJTkZkzq8vTLa0j/NKhM9tWZw++RW63y5YSLQ
q2zTL/fLN7ZjQDlSeGa9+ZQwjmCoSjU5yzC8Og5+F5DTF/XTCsRsWOJJGw6jouvTn0oM2xmm8UWW
+cwALm1Q4wzvQNhR4q8pL94Hcl4P1pNgDdv6vSxkXB8btAnc8wJrLw/irS978/mM+tt3Iu0bRwHC
gnUHK1W4BRfE/7RknOt41FBDowOOcG1c9YSt1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
7n3HuybZpH3tpizcNtjFyJtBsOUXTQU4wlWkJpSsmrTk1OMsBKwEu6cm1WPJ2ci+vT4p8yUdW576
q0I55RoC0E0WVwEvQ3Fc08wJk1Py7qhlQWmBA0nL4mmJa6SLbvx4+Us+/nuUY9brk4ZiashL1o8I
685h6y8wHIOsYUjehQuS5xhd3ZFQ0QhOYQU+CcQBIKZ7cnLLkBZRqJcfkqKLq24TaM/N6RvN/0r3
Jg6hnqtdX42HvaGJRZR4UgGWWkWPaIFlUx+QosB/GO/numyh0KdYsSuVDXDfvm6oeAso3PM1ZED6
PgomnHQ8+XU6P3ElFVTHMw1ydBeFIGGpRWEaw1Alat5iuxgzG4Dn0BU8tPatGOWSB68ICYw6WvCb
eIOxxu7y1qZ8KOUOXsAt5tyh90mci2/qxyiDV+gpEpwLTDFI7gGsCsKYalWrQn2KrXdcCZG8L7sV
bUHeSbE32aCTOkL4QalBbai/kil6zDftkqhTW/m9hK5QrRSp+Y1S3AaG2RzuoNditbQxRIJkIjmq
evWyHi1m5QQa0qeBa1PkEc+mZSJekPEsCcTgoHQK1hLIZRd4KEwmWCFAVMvvLz4JdEPFxxN9Semn
aDpgufFnD+WJ5miTPb2VB2hhFsfJ8u6n4McWRD/SCknwSdgjqpnFooWgZy5hPHJXPkXnX+fu+RmK
bW3NPDSrPTe2UKBiLIQvBBeItuCuAiXNHKJmhcDlS7cHXRG+KrK2kvm8WI3BIQ2Jr3T2i3ztPS7R
NuLy4NGt5n/tr7iaZeFa96aekmFc8SU5rsUNMQliUNvyAgHyzTR+vEZuMPd3nUv7psE74QptUCSb
gQBy5ifrbrsPRtxCpP0co5IkKhEstTLbk7HkBvq8YM8zisOHG2QgNjyc5wVSmWALT2juDSuJ/yOc
itlAYG8YEzKIiS+9jIJCRjIctiqqI9TuEP99BSyTiC6lUB167zyTMGGRXDSeThbOPtzb+EWHNdiK
sBLEmkXhDaMIm+A3uDAW62iyiIu+fWebzYujkhQEHlE5TBa7q1JrslWqeax1+dr0wn0yD/MlZI25
p0M7CZq9EkbzBHWWaKWDC7xbBo2xqih5cYqlCNcqe2Gmg1QZaisxBUk/ABxwuxdgG/1nUGfZ3BbD
Y+koz4SYMmXfosdZSFjMBYQeXCsD6tEIsIWA3TpuLhK7o/bDZUpYSm8+/MIWQj+ewyeCF1OXCYCS
lsupY7WAlC7nwgTLYCF7Y4K1eZl5h3NX5I+tUg4N24UKyPaMzB74QNzsT3Wm3cdYJVDZOte8RcCI
PZexeNxTOude71b5p2M96ybVkiY7uPm07m7RYryv626sGz8v6NTNju6DExH4ohtT5K21zKur/MEU
m+tWpFsAJl4p4Lri1Zw1rgwllex2fNjQXQwq/SNvX4hIGFZ+JddvBSRVjN0oMML0pLIbn+5mr39S
Gu/+f/hAL4HzN5kIir3RtT1dUfJ2sHs7an8P83dS1jTYFjT6xFokgkC2XyRLCLLR3jU44iRvzFo8
AmPRlzDgJqbCZ7Gku8blWwSPASRvZUYFpLRn0ESd+2+CIyWUUJWvORdG877TIEIa410TiTRa+Pj0
OgF0ZUcc8cormkLUrnwEGsn+ow+qlZbQV2NS45FEkMkz704IgQ3YtsTwqI5xQKSEyy2wlhnIyQN6
9uzMAGtTC43LtEu+XtAMQuiCvOBpvCaXleBL7GgAyAUOPPCqOxSjLbjIeAPBbgUk96kuI/ecVZ++
cpuVz/r6dpkuW2cwUKighlfKSjjcvEs+uV8nkRGDEjzNkncKeFaFNq+LsQFt2Vp16bQnmAHmnmn1
PUQroqHF9DjDAC14EvUCpIgb8KXPbNwT37roMBmw3yiq2Xsz4T1MqaRXVk7G2+o5uGqjjtIdFzfY
NA3G8ygzREb2l0PvXnPTKh6raOMnUVwAfCawBS0mTSPVlPx8Ygj7ND13iQo0FIfAu9fBG4XH17Dc
mDxFClmk2BTq7FLbhCjSpULmv8NDFTFjV05MWXBuFucfM+6DxwjNJ+IjD6b0/flyl6p0b5JZ+sMp
zroNsD5ZcjiWVqPCd2T5V3/YVUYylmVyuxTowit1m1tVuj18GR9cbDuNjErfpr7SU/oGeQ+f/zfY
DjeOQfuZmeDDOQVnkRHET6SxXtVc2ngGKFkCDoH6jXxkEdIx8Z8Wo773BeviPqTsGNZxpt0Tglb6
FDN07ME0y1giDQ7ygu/SRmZrO0a7OmQvqj1aqZqL2HsQQqGPjmfa5etfXzlOQJ1avI6kXFHZSdhK
sZZel+tdoVhvLlBpLuBg6iDu7fs6gcLVoL5iAh1E2x7ZMuo8Sa0cr1NtDrffEV1qom2vff7Tm1cm
J8oKKkWKO3t9Ycuz1ARC+Xj0kSD6IF6JOoESTm1U+C/O2pd/keZGve5toGhfHznER4z9aBSBicsj
7S9yhg8MfUWIscWwIop6bFAfONZGcZ6MZBRABCd6NNuYii/trcCVZIJNo8yZJLMbtwnusX2L5UWc
iIJCh35GUa+KaESvRQOJUVsNE59pBxOPBIkrqH8kNUXPitsBVr3ez0FuqwfugLVcfp+YHWxFMAi4
PL/8uI9eIO2v47nH543szTgo/ei6Ns2O3DVF27ye6lxPnq41FjV80P1CSWxmwHKSTgmtvW0L60Go
WlwCOVQBY9bHOyrFiLOKZy645iWYkJE+p45Cb24GvUCS/Avx9Pyph+rHVxJFbkba/mqstEaNPqEe
TmtWBCXAl5XHlC/qEp2X6jbzpMl3pFW1BcTfx1UrUs4rQ5bT3g9uc2ZiUc2/7XmY0bVsZ5J86FxT
PRRIqIyzjn4IOanTmA2qn6BUVwEIndDmye4sp1njZD8PCR5/VMcJbtBDtI4xkGjpVlCj0pKJFwup
htk57f+npM3zzLJBhPNCsLm+XZePczCo8NH3oLFK0tIerUtMbLXO6so6BBwQmJ7fcCLbm6oN6kTo
Y0HpCZyNUMotpq/g+5wRgWGiOD9nRXGiGvqE9vhF92lYn6uzbeS4vQioRs+5QqTWyetxvzW4qSpL
A/KTb+eFVHQWRfW23vFeL7dhQhXkXMHsx10szBatMPTuRXoEHTK9UWKjpyyPJHO5m9bgArM/kZUr
gh90KwvcpYKeilMyYCXYkYR2gSS4jKycYn04NAadnSvDzAFF0VotMakBIOx37StM/3huwjyhEI1C
bd9BYcnwpL0Ip/dmDr+aJFHrqr2SLlQqWECbSYUiZKlknPtctawtGnctxen8vhWZZjGvHTNiGvqh
mtGbKcGF7inIDBU4syhPJbUUVORLVTnPwvKJqU01uszTlQUNGbk5M3DwpHzFEzkolELesNBZe5Wl
TlHuU+xZkjogPZHkOlWVE9qvyeEWIlcum8QCx05/KeL7pOjbOpQecTOQiyJPGEycGpm8Cu7rDGfW
NCLsIQcxXQl4oDexJPka7u+WHsLu5wm5b9pXDlMjlpF8vkECxjjTjPpTnZ41n2SyK7CjRO9mKRiZ
tLsMuaSB21Pv8QIzIFoZV6BuSgZUNUiHXBR6Yuoq8rDMCuldjtj0+OL9if0MX3or9L1eGvMFkdsV
JkMi69b9RUbRhEYCI2UkA8y+CTzN/xqJTcGx6FAEoD2xCJsEs8xy0OqmbOLUlkAKbjsbnKDnXrG7
AjtMs9ooVGnwVbgwg57ZfuZIfKabi52ZVwOkN1Vwz/hnKw3JHK6oSXsLn26AwbKICKpbwUrj2Rbj
Cx/u/BhY7URKlV0PHGkT3vKuGQsQcTgH2oXMm8vr8H5bc+M/SRmbNJA2+LV9cQG/mzc8XnbVPncw
wB+0cIzjKyz1pxh08XpQ2aatUb0VYC4Dy4cLVa59zS+apZbre7YmTAIqwe3yrQ2/Qni9st4Jfi5k
Ymyxjlv+u4R4I35UvNpZxoYdOCchGPF1NxIr8WLSiLKqoOu+LK+iP87xU3b2H8nFegdR9EbdfapC
i+olL8zSgARZKXI23YSHcaRMy5pro5VajCkihV6azPkj9tSq4RZLaD73vr9/G+KpT3RfzzeMaElW
UU0WE2+iUPsyRey1P5fhKUgQFCXp373xojZk1cAaKjjjARpQIS4U/UIdbXRNSqh1lVebU887ew00
SI6TUeN8ZKiydeJMBLEte4z6kmA8PRh8Hyx7vUZ1vELTt+YIFTGxYw/lEsuXKSAiu5O1ijp5I34E
hSy/qpUuco9SBpwW98mzGPQU3P+AJPwoWV2YIYUK2W8Xc1ZxL78yYGTWv/XXgwcMtmnGm/CBQuE6
lLsvhe9ruAVkeLayalPL9wfSQFzd28GnFMOK1pS29CslygS5mNcAc2Tsx6G49yM7Vuo404wVf20d
pIoYxQn6rUk89SBYNAsbx81krmFMnTvtz0OsPYVzYUyQx6xQPD4jG6ERv4TNnQG2p6SZqGEqoxAr
+NbP36u7txthNKSr7U1RvznjTgZNyg4PC7y5d3Yi8ufUajzFZk+4hIgQKLt+QrlGkF9gk/RQOlqK
p9DzsMRf/Y9t1ispHCR15m2oIfoOfrJEC6QdEKxy5AM9V6CTgI/pCwPBx18YZNumNLrk1s92aq2A
Bcd26anNx653Qy9WIEDzYTf73cVURcGw6/G7l7GvzUXNiQVML24dGQ3c50NQNbeuSK5tPXmZipXh
0ylk7cwwnvai1DpAYkbphtdO8xKw4BUyap9es+B77xWZzM+AWpSWGqZTep6pWVX+YC9SxHiiQcyx
ZTvRUnNKLIHwNR4DCrEeavm26RMUsJTsDmL2BDHeqWZjlz+uKOukwmRBLK1mFGlqJk893G2KxrmP
J3K/mf+mRJNU8fVquzZhvtmkTCd6BjaHIYzAPZKoBTsFGNHfe8rEpxqHak4PNfGBhbkr62EfkiRV
E/2FOIMUlkTB90LDoV97eg5jhOGWIj6XyIyfyD7wgOhxdYLhIaslG7OeJQ2jC4spZYBGfUPjCVC5
atZl8qehVpzHvZR+1td/AGMLLiQAgbbr3RBnyt263HIv+XYoluwvQ6oycLNnrRJLWXphr9OBZIPP
4KJZPhWcD/PYn4c0B9xemdWVOM3SuWZqeuMrp8B1kp3stH82GErmx1lFjlicsAatdKzpN0vgci+3
6Mz7tmLC6hM98MDq/PAzkaPsPBBJn479R/ObZX8DCWwSmLg4v0PvDbA/xxb1Umg2Px3ab/SuXxLb
EoaHAtW+QpW+zKXFznJzSaqkN9FwQe4XcsbKhgNYFrDxpJLpsqdUyX1j3kE/5ZIOIPnpcaQIdMXO
omO8R4Z3jfMKtQEvkrFeHpCjPFD04vr6gZ5TpFzjgVyy5LYst8wI66YdGJbSNoWGfCoN58Yg2YO4
pREkCs5r09PpVmBQe3PzI7Ly+WIe/b/G64gCN0NSKs7fAuqcyfFK+wMEGXo633saGOaWp89YxAzM
KU8stIGF6AraTv90W1cI1CY3NJPA+V+HsRHuaxdC7cAEO747sK1Pvdsbnd4vohIi5CbjcatmTuec
AJJk4NWTFGkHQHLokLvZ/3bEsyxz7FHLyz6a+1nCUveAqys5NiKdhc5dZCmSegpSLDxUTC2IUxe/
YWbsXxBxiw55km+ygLXODNlmJHdBgVWd4Ej8nEQQb2QtriWVZm8gHhAhncKLaGbXacMPdpJLjhkG
z9PYz1pieEjT5eptryqnChZ4zK0sGZA2axWyMTCw8A1jEprEYoj8D5t0KUeratYks64AgUqDiRDP
ZbgbZ4ZuTc8T4Mt6IcESfxJzVL+bTqgQ9NVwqENFK/Pw5Gc4wlkNXbTAB/tFBN29+g3NXJN+Tne9
tGjt4iE+O5FmgbMslIHtzlWYqMPAJ73BAR6aofFJx0txJmXjqnGUwHj/UeWVg7J50yYneGM0CmCl
nGO2IT9KrdOtMmRMkvrA++EyBHXgKhG6ttILkMgc20RSZaXcd15YgvoCqWNfkEkpOM3UGiM06tM2
bOJufbMk3ne8SKCqS7jViyvcnJi1H0ovWG616QBHCx9hyW0aQSo3mNqpMZsZ7WEtuWn45Ob7wpN6
/MAtI2DiColiU1R6JC5ggr2r7k+ODpIR3lFjxtBq4ikM+EiXB0U3el8BN6mG7mfAHiy4xddhO9NF
g/I1uh0nXW0DSrAW8IckQApL37YYWlZhEKWv5XjhTqmbKrk3byIJBQ54auQ0+cG4R/WNp5Y1Dkv7
qqVqN4ncHFIhMxyKnAPM0mY0rC58kUrEflnMi/V052gIiQ8rUeuLv2J/FctoJexBbSallYZRymGh
fCk8j1Q5T1OLhhAkY4pKarOS/sQ5ShLvM4eYIQbmv4agPk9cJtIsOdn3wvfpnosmmgMuPIyvFq/p
7WsQIecfQq9BV+ne4sRe7VF7pZ3nCc2h60nwPhNYYZcDiFbFlcRtcMWX7OhFSypFwMqQDdW5PjCW
/wnq5NjIN/ACFK9+Bl8rwLRR5omYprt1j5jIyT4gGdgU0az4S0J8Gm97T867SYPBZtOIdB55QSlO
WxEleBzsXTysFiF7rgGosH+syyKJr2x+MIYuRUFpoyKOKQri+w8t7qhSQNuqrSZUO6UbUD/8ZQR1
yPOFp0p7RXxBxOP9ulhPUk9xgEX0wO2Luq6PmkvyuVgtGUyOR3opCp/EdkWBr5dSco5fZ1aCdtcb
5HWr+M29pXoq7PbadBo1YVlxDtJeetY53HurDEnlY0xeFrAeOnP1B0iI5pOGJrIp8v0dqCNh1r1s
2E+VyNbpUEBzpZeDPNMjVlJYL9IjGTOIGu/vvTqJ/RRuIUDfD6XY6je17hzBde91mOCOqEI4GVYw
+FNQlOv1zwuHAJ8uzUyB0xwz93inGbMbGAlpUIj5vkqcG8szKIHQSqFF4Oc6HhC9+4fF9W2nMKup
Azdk13ylJotemRw1wudUJ8lCozMHeshYMiD1tmmhS99hAUrkqb+ipCyksu5/tcL7KB8TvVK0XiAY
d1RqCB2W6rJb/bDYxf4F+i4PZhA5C2TvGwsWUj4lcglJ6sZ5ur8bVHu6wVVv7WAr/bvw40rd3gs0
zOFLMT5Xi8Tj0bCJJhkgtThlFd298aJ6O9hWL/4r3Qxa9o8rnqXsZO0rVVz1I6er3WQittFuwHV7
2SL8LWtTJ8sAumYzVt7mq2lM0+qa87YOrCGgjbZtYW6w9r5faXP2Q/kndUWk4eHqK34GRaNN6HtU
x+3KnHD1oKQJN4aWziZE3DkUXxMRbCIjU3u4ay9JuCFWUGQ74sSshupQJeZcL68pVeCBu2heGLdV
BJ2vVFmD13MbeRvkqXrSNvR+9FtKfiFT1yldI2DfWBNNDe6PLg8E8buXaZLpthIiY4gDYqMrH1NP
8EnXNPHpFzrNfJiLC1Vjiy1Hzuln4N8DynGD0DzfRNOke/gp3zSKf3n/1yUybmXd3ALkchIdjtB5
cG5CdpZGP/w9NHME8Pj55A3BXakDPCyxVPGVRcEg5ZM/ItJ6sl+zUEFH+EsC1qvPFGKGZ03noFum
oSJRn+VWkgY9ytjzVtk+hBmPfsLdwLzzRAl2Td/ntdtnHsnpu/0dTi8Y7RxNjYAvf3qCWwx/3XBw
YY+TOgF+747prTn9iaEHfIoBPxSd08iqJSrniOoxSW5LkgOCjK7Zsmovokg9sL0JiwoBRuQp4/T3
D59anrc2G/rq/G+p5n0p3P6iNIF142ODX+JSxoPvj5cRg8IK1YEVodBEHiPWYyc97ZEtS5qkbfpm
of3Tgvzn6WBcpWs1hLdqZP/2/h4muVn8GlbqyumWis3c4Cvdb1jkLvs0AyHr+5Z4zzQKQbWJcH6t
JXT860qcGGziZXEB9M2C6BUxQdjsRWcl+hqeEiothuP+vg67tUevUCKCPqiesB/W487oXErrNdqK
UPKBS9a3nMX65VeH7avFGTtjV95Apzy6Aqwg5XVQSLk9vMnUTbjNQ9ScyBTka9aZE5Q30rxSOHfA
mAsJ2+t280LST2jo+MK+WK5I2BjLnXzGJorMrkZdrD4sUX0SeOAjdNdO+epkpwN5Q+tIeakYhRW/
GhDYOk4p2m0rj32QOrlarkXA2Nx+TxMpAuzNH7zzEfZ1s+TzIZ5VHnYf4IriH1E7hEYbsqaVgmXu
0VFrUzFi/F2Stm48K0IcBrMHMQx/u92JykdT1qTKo4wkXN3kEsEV8PKaaxXR2CZJHz7wOFEHIu2y
KkbFyTV10hQgAfnDKmPVB6DQobB9SqeAuRknG4FDDg3UqRJlqWvvwGxvTTqRuO1OuDeguYum/bY9
8B66MxOe9LjAZml5V1fK0LRqfdGKeQKxwxYS8HcBthC4DILypiN0u5D2X/D9LEvuhufqwZ+qYEsZ
U7rLA6yMKVAkHLgEGyk27WI+gQzq5wtZxCqX7QdR7DoLB2xpqNSUqM/h4agAc75peVY3tJ+Pwx/3
PFZbB8pxZhKnUm6Q+vyzFBoyGAggNEoqZzGQylsi18Q8DDBySr8HdtMDbS3gZeinhWQN2hMqcTPT
MNPpQ9W1ZfWTvZbSl7uFNdjebu4rDeUcHG9KBxJEk/tQtVoFR/sFg0k834IePA+y2FhhWTnyYNPI
YBQD/4VXAIDj25UTohHyHBJcSogwU1/rIgBmHeoiYGM4KkpcMAoc6YrCghU9SfrXr6e6hktNci5Z
DIJYYPoA/qmDDyTORCFjCDtZ7EmWs+nuLuYjWKRZlQJ1w/epMuqzYIsVsa3jtwCCE548jJGtgFTM
gjZZora6U5mtZ8y0OQrDQBQYMfyVP9ELv7wTFSMr+F+GA+C/5xXe5ze1AW8JlfY+FSih3AH4lewt
5poUh51UsWHk1XA13SDBjANrORaq+bd/l5RDVaQEcDj3KLNlV+Ybm1iI0Z7JxX+dy1wGaUa91QaO
dxHqzx9yCOLeAOsTcdMN+ecl0Q7kMMqy/nr9+IHTKmJPWCsXhr15QIPN2OTT8WoHcIv2v7/hNCnp
0OwbOZEpqzjGOnrO6ZAZp4lnDoLB+pvO8KD43lnZ3Y178lmREPS7U1RlbwrldYoRVw+a4chGcPfj
MgZ5kLJ/hbj0avnj4rxM89GF306T32PPBveurTU5YUYOSjEha9DJr9wqLUFAwaMRokLRGgLVpwfF
47A5BB75gSFN3snYNa8Vd9igGuHK/QoX6b9/99EywXhnQkI7Bn+M9vGJ6+hPIr9+1Rcv69h+n7hA
zbmXbaMg3un2aHVUJuA3mp5u4UjV6/trChy4kMJM5DVMDAE8Z0es4bhKu46TBp1Y/OMsAG7hHRu8
49rodH2Ir5PrbPTePZ2Gk00s8ISZaQ+5owfif5LuZPesG2yXXUi9+sMHrIz1JPzNyApJ195UPWIU
ReFmOl0fyMNtOQ9KKspxBG8O/HZ3DvxLs1pLZyoaybvqCrjph0/6p8vFHRN6uufUCyH8ANU2epm1
G8AdHG0jy50btUrDVLrXLf04A97uo8/29Py4SuD+XHX/Dp9JCgz09awTXs48vKHpgoAWVmq+Pjcd
7tUvn1sWuwWJ+uQdZnYnR0PDsggyGav1im5mygitnS9IIgR5VpLBxw6uJMlWo5SOIatyC0ZBPnnL
JeQd85zjyp0hfuxlT9uikZHv7oVItb5WZB1yYwHZiZ7jrsgJ0J/cRBbx65KcS28zij0BdupLls+T
FLkkjRPDqEO5ixfbr+bFisdhBH7kGNn8gs0z9GWw3MgWJmylRiPGwY+OfFzj9KP2lZgKiqqK/ZcL
7cEPY/J9vGNWP13uXQcs3WUA4L59ZVbfs+4ZYaWvx2yp9FdBcK/8xXnwK0e0j6qL7v3trFRHcjTn
faL1Vn03kNKKPbGGd/7nMQE0+Z7kJoiO5FtZqHKJLxoOeDoM3AuDUZKL4rKToRnMpa/OUzzMnpdw
JocCkRaPiWO0/DNcSpjcPGaS9KU25WkysRdIuRC7bLokr7SFM6Mk/tMfx4YgJNe9fTqOISybBn9z
oK6Zy4n+WYnYiLziHjF4lymNK62KWS8seMoUHmIrpVL5NhxRcwqsv/TbWCFWh8y2O8RVXcs/Clt/
xLJ7xBAB8Y9sSFtRCrUVRCyJp+bQnxT7I/XcnkBfUpsg2A4eHT3kCFNedJRvpBhEDVQE/RKMDn3p
vJ45ncC/Re8WaMwVzKqH3LL3L9HhE0z8H93GGAAmjo1alJCkhLpyKbw22SVlb2/K7v7CP/6fv6TP
l69n0KFp2pmFDl2cBEHRgIwMdBdkuJX5pI+26z/KuNXSn//kRIwTwXcj0pwIWNK6V7Q8YNyRzOpm
XoYaDFZZqhm139iNs/66fgQPhchvV3+U8b/lgaX9CYBGreIQzC6muw1nGtYW20qe+FK+Towk8rVZ
6iQHKks9ttOrGpt0SE0Rn1UXooig4D4uY6MYDJSVf67ieq82inikycFR2cYNQq2j4cfE3GiPGolv
++zYJd5mGxboUzuYtBGX87zvQu/qaIQnGIpHFxYCSwNeWGIuSpb7H7fbkOTLWKi0+LRAxwaa0Nm/
Y0eQgEQMHMMktCxiuNGZJxvdUKKWboBriv+siAoKED7sQMfRoHI1wHCRAHXa9OOOuViS59w15WCX
p/2MR24dKCnrLWE28pHA6Jw5uFuoSGLTLXcUZFIbSJz1t9TNHCV+2Od4yrX0YauZetZOOe10KhDv
Wo5+XKc/ABAWXFApkpDFVfOI8Az779gMODq/5ax6jcNtEtLNvhcbsJfm1gHFUamKaAaBQHR2W0Mg
AWn2APBSKJ5I4iuuNe6qQ3opj8LJQtNoQm81mvbScxReIpsZhtSBKEkCVrfdQpp5HgC0nsJIjrBA
nnELV3Mj2y7tBj9N2TT5pKhwzPyeGxUDtI9cy52AXYngkInwz3q81b07BWHSoH4LyfMo51jWctTK
aydljvJgY/5gu9KK1fTd9ibkEJuDCIyvPv0w3NFwjZd7wFb+cJzVo4UMGOyf/du9f5Pe5lVCmNPI
8VG88RaQ6c7jRIEhRAK13vDSGx3/+P92o31tl7RWqvtiky5NfJ0OJYNjcFQzDYinAKXaaZAecsA0
jf6MvV5BIjCBEP4W38A9X7foy/CZNMtgs2C7DlT9qI0Pe62zZER6JyAV9eurws1seD5vGnRdqPRx
V/VCfLBdfKB9usKOuttCtV2pSAX/toH2zbaARspY7ZDcBhd1aXUkjbK4PTv1UlyfFrHdsUn8R1cs
6lms/CiYXUFvJ3ekk/MfiX2JidB7GTQUhk19Y9guaiidIXy8ppalhCGF3QYxzr+zwEMTuIm3sz70
wrr2N2w468lw/YqymKSLVFLUtIf2y5zSI+Ctepz216YfjqxzAo5yqcjNPiToJZ2va38GnZIcn6+f
+tVqYsv3jP//md62td+0hMQ6+kIhzcd94iJXAk0WGVbRUhLWbjDZaS+LLTubwNniDtq68MuBedfW
dBKlSHT6fEmGhprJDxp4gp6JdrE0eGbkbUvv+bEsWiUsohe8vM4R7Fz9jP6AGZjmqIY02ZHMtjAa
LEqQlfzSVtIhqAUWOuSsTbV55ElH1zvVMpFNIgUMxO7pmtcmOKTsHTbzMotp4YxRcOX69tNjhJrI
wxmP4g1M2L5uZYxH+brnxQamo//uNS5WyVps7FBcOEYsurEfUXeerA5g0oNEX34I5tUo6pa7CG9E
L4ESwsKJFhLz9FtCFQ4j6sgnrmdE0hn/9LulNO/98fPQxoiir5JJqxuNOMrGD5uMAvdwZBkvAElP
CD8WiZlYeBPUsxQoYcxwM/9q3+WarhzaDpoAjq90C4gXwgmIJwJ580fhr8PRaJvhgC4ZyYdXFoew
r5FSffQG1Wawdn0IT3GNMdFk6WE4GucsUqEvqPPqV3SKcRdgYkaSlKW10+umtfFfX5fmQUfNCmnB
OoS+1ssaYQHtrLG9be1bnrG3R+/f/pG0wH+aYfiDyU27i9KDI/ouygKFxXakWDfn9rdu3V4Cmlcf
WWF3HMsluwdP8Z04XV1WiCILkSGrQBv0U35mx3y6fINd8EWByFQyZdl2qZl+R79ye4de9oAi2QEv
zFYdnGyogfuemmcscRDBNSUTDyinw41icpiJSttvBKT7vrDfEHcSmyLHH8o5UcIxFutll4eMmap3
959PpAwHZKxSF8QFJv6D5MAUpVACy2JJDwyRwkAfuarNxAo97LWCUTPuxaGHbQAB82pbnqKEKCBI
0QtRQdm/dJLgDoYgjit1Kv51PZJoHM6HavqPIzxk8eyFx47c7ak0H+9ksz2OWE+0PsXa9Uwlo7Xo
dMe8rPZ05Cw4aYuHnKk5DIVpMRh+K31xEQcOIhtsufdQkLAFEbCVbWsq8/SoOLOnDGh0XIwJjeQ0
Xn5z7qa26xOQ8PHgpPcVVH2f9mORcXdUrqCCSfZSd2uBV5TUHJjNf3B9QFNCHmXFg8tXMyj5H622
HIPeFc2uzVg48Yqb/9ocf2DGs25edXDWZcSNCqNQE9PRZwzJLF8gJgO4/qSd+wFCRvuHqSnrU+v4
ptdPCWiz3eXwkpwfeNaRSSy+x2gOAr8KvhShoaa3QscJuss1LPpqYcuNDSI1TkIJVO6uGaLbYxM0
+ikhjb0J11Frj8xFep8z2kugMR/molv52c6o2oVpwfUhTlreDsjrcoguqUHJKIPiTSIH/jxI/jZ2
XpQLM7WWiViIJWh+OYGKrAA9rUqUl1w5p//7pYf4W3ErkRqkYTcX8jluzsV8P9sjS/9azyoiQJI1
k80XbwQSAg73eOMkaIbM8yE/LpYdAkK7j47xPGVIiULtQe3iFdtWle8BiYOa1OguuBfgdbO+Oe8U
059NVxkXNC72L/p5RmmbUbs2nLN40Km7krSIuE446Uq72s06pA5TrLh/zy7O/TwwD31qh1Gg268q
DhzeWZVHFGbh1K43eQOyC4+m/+wi4N30aQJO1ATYjWg0T42LyeDUtFNPEEM8auV4OLVy2Y1Xcimi
1zruLpusL8156lzDlL0YLS4t3EFxR9bizjouE77wRze4DfANW6Fd3yeyeS1uChwEaW8TdQpNj03E
k+KGVN5VIqNkzFF7K8M/7PvFfK3MpHkqqlFWOxllDgIjapZJsfbb4fPaGGQizS1kw6W5azqXCw9Y
mG9dV3SEkdcVCp6ftQ8pAKJMNHQTXk1vjHNFptq6eqn2Y0CS6FVH4VTCLnS57XjpHml4/ep1o/OT
QxmcZJ9kd3d0zuaqOCiiYLIa3oShNC2XWMPgUk6kbf9Czff0dX+qKids4QWpTnRsfGFA3zn6i7gv
i6ACS2xHwUSXX8Aatfc9lRoPYal5jxEA7qfFjiDKz9Mf/8MKzpi9x8gwkwp1bQ/ZaP4GJdBLsw4B
Zw/O2t72RiLV2vli6QqFOvmWZr5B89LAeBjWwX9D5xkzUDlb53ZpL3ZDngxE3w9M0bBTKHZrEgf8
a/MWTcXqgF8PwO/4nP8ZKmULrDLpqlkfzqialBCpH0ZxBORM5tog+bwgbLYGxp8JLxGp/syBFDpp
Lfn2IEp6dcgGxkPsoCe2IUcQQzfE4DSHc8QSAP0nO3qImj3uhisFg7QoI4fI80uc0Jqt1i0WfklU
fW47iOo/a9TllJCdeQTWZH8bY/yNDCiE+vvSyAZheGEGsQlkcgA6aqabvj9zZum0cLgRAll8wHSA
6aG47Huos+4EDpXUnTu+itTBd9ehqNiFRgR5hQf97UjnlS2jE2DAjBNqj+zoZhSScI5LLc4/lVMz
tpS1xePTLAwZAhZfN296A0KKG5duej9pSFZRsRbAfs2Oo7r4jMPY52O68zj7NoR3RkkmEUWPmXIq
yEAHXgwv/zKti/1fRrkWjvKKW59GpLgbVzgJsp2QEc3lR5cVjlGIAO3p6HlxlSy3hE0WD2JvHtgm
JFHJ0UWfyJLNFLWfM5ZZXDprQnLY4yFNG6Q8lC9Ub0N2y6XJkB8MtyLwxUH5oO8sNUEYPtF3oz1Z
gn3UJuByXaXTzdNQ+3zDfn7sRdQu13BSBvCWxf6h49UyWO1qqBWmxKIbA6r0O0xKvaEjrTgOK3vt
AK5p6cQzLKeMiiZTuKmkEcMJXCDjLkiQLPKk3oizNQK9Cd1xtts6P8CrHcFTXmaDK1qShUPhlYpx
L0sq2XdNT+2EyHvNErbhnnIWWZGSy9OxJZ5Cj/CkDAC5npacaRXZob4sAzVN6glkQJ1GdkL4PBAH
EMSE5+XflniYvI620zm2IMVjB4PA5I2KuGkKy8gl4H4hKHTzs8wl8waq1s3JrAZLNcbROfCMBvja
yvcFm+Z4icVCuw1iBDl8jzBLBh1BqAVnQVfQBe8qQD9T5i/FZvm5bUYox1bBSUg1mQld81Zx0onF
q46RUVcY+o3mngd3Kq5kC4vKKx8kqZqXdVLfJDtgEiWXoOUaGhY52iXOsDtac0TZ53czm0AAh3eE
y9MYzhD/IhZV0h25eqa/dYNj1iLJtwgxKbXrPwYWcI//yKZObsQlIKTudXOEvA29qeRL/91qz2ET
yaL+A997bSFuMudLrUzIbgXTAarE8rOXkmv4B0+p+lUy4NxkVnMmcmVl7GrQaIFiO4QZL6jx+UkW
eqyik6q0ZvALsArDpsjPyI+MAcjptXhgfOyOvRIx4JOd7HbYuRK6eizXKKgefsSijs/1cOZ4Lxkw
JGn4uIFI1wNSMupTCBVzOkM8eKNq7BLL9VugzPc1QkEyndjVkzpNomOKetsvML8OuAqOGkr2sJHc
M4TVDTK5/zBDe/ev4Q+R9YlBGn1hsuzRh+dXj49AzvJbHiHDJ+lOXrMc2PPuwbKbw2l67iZ5gG9h
FzLQJwMs9bfabi8hIciFI5QHJXjC+GlaDTbEhfQeb/yyEtmXujRpvp4uf4+Wbg5SE4BZs0jMQGdj
d/oqSKFTu6Hn47ri3sm5JQn1NJf753CQSId07tezpS2hdwtbKCo270tzw5XDa6ghYhJJpIMMVujU
1HlMOM57ZyNoH3jClgesGX+x/ia6CNagXtyRZVwLuRdV5bpxv2rToQuKgFl8j8xOY8J50ZgDuziT
TkxExE+JoKqQz5mIEzNJRE2ZHJ33pdMNrJ16DRfzJErcseUpLqIhWYMBGwtPZ5sVaOvlH1cNW2Eu
rV0bYZwPhX+kWe1ATzOrm4x78IVc5YfopMIFslPQvJwtcaCXKwpBbb/IWXE1QRavnUkeP9hGjUmb
hWAlPXxWnTsEMqdilBIYsebJY0jpSsqCnSl3jsvn0En6o1UPHK3LvExyM8BAWkkjc5kp0a9mZppR
iUI6dAkNSyrt0L4ods8jwe+l5nRcyaHP57czJ1s0qPKiedLPSvLHzRVUvgLI2xNvmj6yCCbV3f0T
m1Izw+b6MJw2YgIvROt/wwwSFheIZj1FP3FiLmbqQrvkxconUrK0N29uprQA/QxZVTlwb1yW0B69
pJOeeVfp2O7kFP41sU1x6EjhIDkQVSktpETL1iUHLQFzVlmAsp+PFT/LZRm+PQ+VYtykKQBcMaJU
F9wVBFhQ3FhYMlIU9ZmZPHhFRh0gB5rXfkop6pFDZS8KWIDxifkpkXkzUc14qH/QcV7d4N7ftPgl
uLi53lp1Jr1ldBGW776wKe84umkUZ60WxMA52EHrzjP3tCtHalZ4JzCxUZWLZdRl0T2VBfbe4Bcc
fRIPYLC0KyOkjN0GDA0CR543Z2nlTTAmjZ0u1EgLlZcealJO9NrwRdxJ68KZ+1PKuig/s6CVpLze
BQHpPa8PZOPNRNNnRoyvjERKyuBm9db/rzaAQVsYViA449DKgv0TeNybOSehvXfcjDvAJUhOspHC
wPogMUAk+BMQqaEHMyg0pO+3NPfg7ZoMw/6Yh0mh8TkXY7NSB0GjUbXYPjC3kPULOfgpfe55Jui7
11BCWUhfu5V4rrj8JJopkEZOXSE9qV/aK8J1nMG5vSMXuzEgZcmOCdVzuOCFYu02E2mc9b2KBck8
MxJCTdWgbbKz1W7zsJpuHy7ayea7O5wPhdbe9On8dzsIE/l+RAooUbbExjb+rpx6Jlx+iVg8N4d4
2nL3YADDV8etJGrtmyCTgvy89oY+evb+caXkknNjgf+RggSsnheh00dXhs5SngYNfZTkxPHmtE5m
mFKjh6fyGXIq8+mm33N/io8QXvdtm1PAoP4+qQgujBNXIde8BJNbsI5l7a3ZkV0KNn+uvJ6cDED9
LW3B9fkZkuawJ6naB/UbgCYUWKynftkMX0I4pcteY98d17tqeqkx0KSujkoPqq/tuJ7jKv1MrDbM
gMMeO4NF/v2uELJ+FFTMYggztAQ5MxYlgcczb9qXQsmjp8UiXnrYnNIxmK8ur9gE30YJyg14LW/L
glu0uPQyDE+OV+/2kUxtrIJ31C8a0bG0jA9vftFN86rnNfx/x+Nk3WIwhHchanEBqSnW2pRPgZnr
Ita/wA73nW1ZwuI/2B/eps+o9HRt+ljhkn3j4BGH5Sdopy3OZvo6sUo8vCiYmmn/FzHxLo0RHqNP
aO0TEcsl9Ji0cTMipudSH4jAHEJ3cCogvbnHa7XyItwXwbE2yjhanZyqomWkaKLecOyzFaS9TmdM
cJysicOB+AbNBBQFBDuQSXLhwkMfcBpvJyVCyzeGAUybqXjyXcydRmpMqD1VNsTNb9XNienGrg2q
ALYjwk5aKPynM3HM2v5264fNCx8xwWEK+7EOGMhMErPzLilL2Is/kBl6tmQvYp+wcd7uK03PUrGb
verYt7PAxOVTHUB29L/w/x2lX3rnvQKL3uEDbNG8Y9TDTV5QTbbP8tdioLptDTCBrTVMd5Xf0II8
CeccUAFoU+k7VfbQbIa9svCiWJUHDBiLoiN4tbHAuRww1dG34cYhL/z7ezTkC3u37/4EHbIY46Hb
ZUMFaOR+bGF4yZaRiTmiIwhiadUytj1INLlANaBCo0IWzEEU+EVd+HiNopePi5YqcCldGRb/MXJA
J10mrilW5IW/ojWln71NoYEBHku9jc1RUPEVFYBDOygS+tF0aVafGNDCn9ARbPAw9wz3hH0rFwmd
j/vlDPGY0Xd1UOCROMAOVbmomQxVNlBAx3gNCvbDoChsR4P9eo+pPpFAFVXktaOQH4RBqNzAFimE
uobTUM7rG+IaNaNAEYwpGXkUR7V8Uow+7NiJ1kdbY9t0DXMcFoReOhR1wOKlxBqtpCFr3uPVgVt1
rE6Xu2OnXV9PZsC107ZjbjInPEOZ9rjpayhacMTGPH/JFfyjQCBL55WWDVnggER6TRI8fxySXyrc
YTcWpRMAQr0PbIXyNyiDWWYOwf/58TVTqQ1ocOIKDpUAfpZM+1CyXg8St1QgPETIUu4N6YuWLSy3
dxxbzZK+96WNt6CDtIxX35gYKknAlfb/NETUv4MF/sZ5plA8n8eovxwx6o1ue243t7bnLn6EiWKj
D0Emvt2U8zZVNteSAmZoodQvJzyrk0xdifQB9Isah4qECBwuzdccX3uhQQ0LbRSKxM8tw+SxpO30
bXk6O0t3EkuAQvXrlTDO6JfTlR3mCjvxTm9TignbYccRmgUiSLAym0IG4udPhH3MDwSmRokT8qU7
d8bcz8eMo8S6eRke0Ol1GqOqjb3MFeDvm11sj9emrUZxwbgPNscFqgu+a61wcHsy5vX3R0L6tyqz
OZev3wek0xzjGOJNHvzahQIdkRB8E50i2OkM/rxbU0TexbSK3B/vLGcBrLsLp8d5C43YNmPgtqVq
mXF3PNBnV3IlpWRtkoZQwClEZ8bD4Wje+rU2c7VxLXJWdxMx/E5Pnrg2QWlnUYjC7Umlw51DAEBy
8ZRNydsncJGbRfj1HSbNl3casvrCtO6o1nx10Vs9pEBNrdsFLpkC7RvDx6yeWlCTOY2D74K0dZYA
jVBZQgQ4drjPk1cXqiFpKm0UvKKbjbyz9nQ2PM1zoz7p5ExGDXf+0Y6chzVDWs/dudRdolvjCu/D
iBnm7FsNhnPPCBRPg0o0jIkzHovstD9gCdze/YX580l9E39xrXp+hqxFKLDDx1xKInSsmjcPn6MO
Bhq/tjrqv8T4FHi8kcFTx0936mdV4U4hmnkzuyIFlaLrpNirhIggXNcqOn7dEXLdVnCGtsrtcgZH
BT0Vpf+BQ/lekO5WYRHoR6QtS46s2AvqG6/pb9yb/9XfPnrztHodVu/uVkFLNalRotI5mlPikZ0q
78ZA1I4I742+rmbzamBm80zIe/FBaopMeY3fZXVEkG61GVmI7NVWEf0pEAKynlt2lhZPLWlTDK5f
syz5mAyFS1WfPpG4b6ADjzymqwM4iADWMskTmyEOEkFD2bX6vKe2LcyvU5LfuUm/sLO3YGBWzvQj
NYfTCcOGKA7X9vcIb0myUSpB8K3Etvib4TR2DWNRAn2Fu825DeKrbXaVAYUN1a+c9toxR4KtwUql
gOQNgOK4NaFZQiTYcKUn7+FkxfmjKlE+nOWgWs+zacA1ZJp6fmFjLtXBiImjx9IbOT4pKWP0QN3B
Nrjf8O95m/5kbnIepte+h8XNW1doRL0/y4GSsqnd2mYGAcZkYKI++mM3oyGoD6XnIIn5j0sTWMnq
VKjNOc6cjmG6HlxUmf3eb8nzolKMRCZ2j5jQgq+3M14PBDRRr8igmmEY3qwKWnfewA/2oXYC2rdj
p66uablyw59IJ1NAaLDsuOmaUX4fbyLNksryveGeV3Zwnu03O5fxg8IDAC5Ht0teXULYl5ytOsFR
3DwaYRLskm24ue9cxnNaheJ0A7JTNHZoXHXlssluOW8vRHQFXoYjw7x2YtVuu6Z9NPEaBMYfRWlF
AJN6tXAbnoxXr5ABsVinao10JWUs46haVdjEXKw2Xjw73M4f121d1lelezXkCYSj+TiEjH2tK7AU
gnXOxt8+/94xq+spkcflh/Ajmlt1kiZMcUZnw6DVc+xt5uiP9U7p9GSCofiTguDIkB946mRUfqCt
hEyokMrp2XSJJsGRFjNef7v9vyxvFYgKDOm9AkjSm/zkM+T76lEbq66d4rixoxWKPrslDJpKkS17
bhzeKhC2erVeSazQZj5P320Q0dalY0+zivAn8L1XDuhavunsVHPNC024bJdokeBTKsiEze6JPP+U
mZOGOSyCE6iJluOqJjae889a7WxHyE8cNIQvqnsB7BofD8bdPT2c2nBm6J+X0hx7g0C2CvNhZR35
ob+5DVDtqhmyEZcks9jJA7RF1N8KkQh5/yvr3SDVdSR0E/O7jiIePklxxVGriPTemHC4B4zm+Her
MR8Jbdh1CEZtkb5iUStZ9os6kNrZIvJdzlaqN6q8P9Lv0I07wj83RjgEMGRNySSF5vRe8pTyCyYQ
WthovceUi5LRE9ZiwqQgvnTG/a6oxFGAZ6fqif1kea6zdf+l9SNB8xdXQalVw2oW4NltcrCnRxPz
7wRa8jXf4njG+ozW8CZp2nUFdh1h8EndPEMjN0aIBqVmGZWK0xLyLQDB3Ms8w9qKvrAKgEqsPcH8
Gpq3UfN8YbhyVC2Ekq3rmvnwQJWuDni4yqX8TqUdJXeiGuZyHy9ZDRonbGD0bbQFO6oX+HY42vHm
qbVEGObimSQp4QCtLT62wMue3/3uF3TB2PRQfCDo4wta8wspb4GI86CWbBdlbE2q7vl/iGLa77+P
L0K5AxAsdLYZw+B4LJ5z9b04TnltUKzTwNnX0px2EAknfCSDqskdhfHxc2kZq6nXqSM8bysyv2Wi
sjGX62i1uk8wcfvJbDDZD9alvEUB72kG4nh73joaY1IOVirhuz7ay51vkzRYUdvNBEjWONwTWVqa
8MYcmzTQcBHvukLVKmkOHeo1aADUqfeLCB3vEOOaAYIkC55ICCGgyr6ldS7/UellwRCsCPzPzqmF
12CGbtzdBlfdVnvLoCK/398TiIGMr0p2OAvS+JKSZTTAnwfqDRWxhDMllzigYfveImH1n1Ig27iK
nD9aHvJoQYy0RazCeMk8bCa9l1AOwhhMHo1+ITk/CRkzwtLGU+ItJf5KoEcEOenoglIqNXifbvkj
4uDJc2Rl6S/uar+92S1sPA8q/17saUiglseLsjwGImPDMdP7RBMvJDkrAQefsJiCeOO0zroQVWY1
OoBEznRDTxE2JQHa/2kmDqUcKUgiwNVVBV2W1kaAgjfIYc28sZc4AyyngcuWS4M9rcKfXSwTtdAs
VnNuaexc5JbnbFkQ73VHCG33VS0DlHNV/0IY6JNGIKiuXsa/i9VHNiOnFJs5CQ5e8FgJqrRwC55E
+ZZAEKcC2GxpKJEhlAbtukrUh5FlUpjXd9UEHczudVwoiY3LJovAmO5Fsax1ye9h3bc8lR3DVHpR
SPpuipiM7Nq4iTIKtFG+pKbcEPUOYY/16VAeKj0//Nfby8viH7FMOHAUWMZgaU3OtKAXOQ7KRD0I
PKwXOq9p4UPPakI4C8iCoRej9UFWkNEOn5fAXp2xVXywYO67x57M47PrvtnWPxVgpInzO2YqKnM6
fd5vFwsxNK+A583s5VJdDXUaOP81km5Wp2hoyPFaYdxnmo7k99wRPcY3G2DzFrVkrrXLYHhYeKsa
cH2jSzwIrKQR1mMEHXSHWHG00DBFQJXEzql2ypmxTEyr0Scj6xK54F+10AIkTq3J1gdWk1QPwJ/I
VfrxGY3IZvulQUsjQzkrLaYLKCn2+q48xWELLsiM3h9IY9K5RivBPwmXI1u78VxoYUOGc+SY4GS3
7JYP029jP+SGOE2nS4Q7NJhmj4YigUB5jBiftY3Y8JL4vYRLSyj4ch90MKFsqx6zSP0lbGAqxpgm
Nqqmar/Ln01xk/aKuShsftJZ2KwYey6cOtFGkYX1t7ZtWefsWfKdmGhh+/3hWcdrwxQriV45xsL0
ukZIKO2n6e2X2ReiaJS+G8ejXnxzAcl6vkzy8KLQoxvRKqJmDx27JTGgAN2VW1piZSPZ/U5Vb+/C
Kll5/Kb0wlxI5OWD8LzOemlnSbNn2PZ7MU8igk6RJc4QnRaokb4RCSN6JrsQiSXrkZ9P88GjLt42
/mM/M7/6oqI2WHTVbbK+PNMlnBCyabnf07sfvwIS9FKyoUpsYvfgzFzOJN/KcIDqrmgNrEMtsBgU
AnQe0QUotsExBPs0/XCMwJsO6+iDLYgL5XvSh+hMziBTgJPxQ26m3rph+43pIgceSSxCAs1hSFsu
W9yYjJU4iRzNg/Q/jOuk8C/6hCwS46U/fCsMS1VxsMRusScGDeD9mpZxV/a4MPNbVD6Ac4m0RIVU
6GhaB9BLNDOdtmhqCorntRskUIZvgA/eGwxxYTZVV1n8ffT1t/+SBWP0BhrIUzNA/X/GWVcP69Fd
4ntXUoOAfb7or5/il4Q5ruqO4aoyVWYcfbElB4wBbtXkJzejeFH9jjFI77mF6DGru3dg5eKssn7t
bVTKArIT2LpZn9y5VBI9fOjuHWzxm/+FluV9P/one5peD3pNhac212JvZaUu5KfG5vWCkMm+wVcN
eT+OxYKOcMeLNyFqc1aBQQv9wzgRseApve65b6k5jTzmLZx4PFeflfgbhmX/gqvaaQdr5foSAEi6
u6HtS+OL2HCxJrYfv4TOxRwFbXCe8kCXR4xu2UDfXlxgmtMCRLGqQ42E5aNBSi5IughOagTAIS5r
XHRvrqbvzww4vYlnTlIQcSMeMkEdSZs93gKfN2JTSDzG+EdSqI4e1di3WHI+fWEUMZv3aYuj0c10
irj+cyC3plLDm38vkJa8Yvq8bMvbCFGHrdz2JrxWinmpp1zNy5OQFjM6g5LmhWe6HzJLYr3YIEK5
JS3b6ScGgZeN7Gm1k/ammNCSOae/us1YtgyveQvYVF1BFdd+0hUfLAH/V0OoPL0i+NTPgHTkP1iL
JP5bxq3oXPSHZVBLtiX8dFOpXDHTtZuuRRZakaBnrcB/+BBijxexsUEoSt9wTuaz9pp3SVl28dZn
rYN68KVtRuo8rrCOD0/K6Ji62CTnwXN8ut5FLWqcnB4xN9zIgKeuNVmP/kHPey2ec/BlQ6EUUwyq
f80pqk2fX3gT3EnwNwobN4LDAriOCJIpLaF9WYXXkIxLB3rZdTYMSp57YCa6sSfxc/61SRf/YhqK
5SRKo+i3+HfTiXzCF7rzN+ZSaPCKeKTUdftiKLU59r+uPsGusNhpSzCypAZBsJ0LVLRFxsur5t5S
z41+zydFI8xyDj3hBHutEoZfihbJahPVgyO0AJRg7E1WBa3RE7bXwsfRvK66Ci7u4AMg44Ujli+b
VMjXcWPbo0NaQ7L2SrK72D1ox66mdLDsB4NGtvUlTt+0iItM0W3wzLGJwQHoM7U5rbmv7Q/SRKOg
vKK9aE3QfGDJJljkGK7D/dh2qm/W8rUkQc6kI0BY6i0nZdCzyJHZz+heH8Yo2OFlt3J3yHAIyPa7
/wMSl2AhtYHxPON9tUeCpZ6irkQea2t0R/oa3gZmvnidfZuWiNhKA8TpOt9UxiclDnKIdEYB7Dl2
RyqwRRn7p9o7yNFkCia+4f4bp5s1y4zam137OksHe0aTHqES2jkcjwRNtwjw18enNYzLR8mr6WEb
K4GEDB9ZZrP3plw3fI+MZMhnAcKB2Ct0gW+9tZHBZYiwuLG6OoDT49PLpB8OxeGlA3M1lzmhokH8
VPAwW6jy6Zm/bMc9rH1xludiVqawOuCsHurozc3jsbAPuIPraRHMmK//9U4cn+/64JFXo0wbPoS2
5DYzMYpd0JLXUUhyiITcVpJWIWHkFkDIcfMf3JQprXR1ScFfz31CByCYCWyat/D9Y24ZX3bic+cl
QXnw11oIVkVwGnxzy6GTEXzqJp604nA1WIWh00Fn4itrKUMRJHYFX+CdLqqw7BYeH0KDdoto9CtW
fUA6heYCnQ0/kiS78EoT6uTYAvUKk5F9h0p9wyagTQqFrGKUwYNH4OtXyJqsJJ6DcdBiLwG1zN3x
MELWZeaWpUtnZ+2EghY/ix0kvpSOuZiXDqKMDkQLZq0opOYutQ4+VmxAriIiRuPhSE153vWC1BB9
UzxZWIhYN9vWZVUeerjnRFS/9V3TiFhrvyLeJ9OvoCo0glDzt157osmHhig8zEM8PoTAI6sYnBPP
lv0nxn/8O7KjYL5bB8gCN5fSg8qk68XXUKkOOplv8gJJo1uwLdpCpUgxUEVCwMN+q6bJbkTUcIMX
iz9Wsxlkfg/yz27Ts+Wgq7WWPGE6GBNXFm+mTEjI/5xir/GJsN81jOZQw2wmol5wiggXvKNUXkMn
0yVvunvG92T4ntUCbEz/lfyQ3XstH6yrrnnv382O+OU50LyzZvpTn3xrifdP+JN1P9b1/1pRjJao
eG2qgv199JJxyQ1vWqtiGID/ZKveagB5n8C2bMul3i2NXjK+NJTCCSOl/yL+IfJTTc9nOVH8fctp
T1+srQAj52xzM8SyW9u12buixxh7H1tkcrOg2gextK2AqLQAyw5yv8SDIbXxwqsD3Bg8/rCTHRqK
vsb6ySemqPMOQqV04nUUpoiyq9gnYOjYzzN55CIXH+cSvxxVoo8RhcY4D+GYRLQ1V6kdy0K755LD
DXvP9KL922O0H7FEJKzYC9WrACpKLBPLqjqIJBMQ3/zkVTkGGVaP7y48MsNVeiveLxsJPulod9Hw
3RCUe2vUgHSD3FGpQEcyn3WrjUKOaLP0f1Qm1l414OiVAlgUM2gsn032+3xndT/ehIv/XE5rgu/0
b9smSB4FGcd9QIaaT3NuewDzXjVS+MOuJBOBYSvBbg3yCyFn+FI91CQvU+TU5budrjjLJ4Y7J8kV
kSFkaPnBb6N72QbZd/8lPU0hgwmUs5y3CScHBm0TyILOe8sn/g7Bw9B7pDNInNrnLB7YjVl2GXva
ZT2lsMq1BXmAiEpAklZfXtmZ2KEqt2qkTQ5aJMaUQc7zEzzPJIthU7YN/JL8ndH8fGVuFGvIIO50
9p58rC+GWuZbHU+NkJHRGzdljFvik5jz2EbBQZ/TJBm9co/pW5PKt55P4X1o0HLxPwXUBmNg2xma
3BywLy1qB2o7USdb8KqHxZFFCReBmNs7v+8yq7Jx6W+Hfw5AY9jB/Wd3w7KGpKYLcvPAAFuZa/da
mJ1jgW9mrZW6fLRXLqKwMG7f5Ymvk6jN76PfMb93r251lY/e8PW2DAUrYy8sht373o363ifilKIU
yXhM8lb/3gGap6+j8mdxoXE3qKDt64KYElrPkbdEXwGdeEKREQOVKwZoN9iVt5HldLs5tXjH3kvC
Px5KSBiwQ+tNOYK/LNx9SVVxY0RpOKzwbAVWxnIrQ1iSD4PuhI+zuS3mIHltiXP1AJyhw7Wv9Hke
JHb2b6bbE4Qgb+Zu4JCcMr4FrjHry2YtPmqgtEZRrP/vmORl/F7nvAaFb3bjmddujLk2+ALQikO6
7QEprC66/XUZ84GRQtmdywb/a444okpO09841nnGHURBupnWnb+3Z420PrWPX8D1ixW5L0ql3Uma
OOAVP/WH88Z0fcGqUiFnTMDInDSZl2kLHXSVF53jQB94fsvyvs7veAUCZyYbED/HPISmMIzO74/W
eF2BX2lr2uWRRnAqwUrdF/yzphoXEDoh3abeQ6JISDupul4qOozXhKaA7RLE39FyEovznDSdPx4T
dlb9yAZ4X3en5EwWoYxYMgGlZv/EwD1gOjswq6jKFUP32gT990nwM6sm2QNwdZsDgP8vADMwXeo2
a29k2cdfRIyRN/jgvX56Db5uwrniaIv5opmXRnAk/V0QarVEQ1gC5gfg4jnKlWzKAcHhpbnKKfkb
jGoY9abb6lOlqZsSCfYceSHtHLk6lkQzeD3hljMNrPrAreXPURENIw71+1wNufrNZkGWclash6Jk
jr01HfuIUU6nRY868vCX9XtsCIU4E6bcVo5ESMVZFUBult/iHdBr/9xqdlkfvTAv5u2AFsxcbkjX
fXSelXJC6uLzkFaCpFAvgy5yMTY2vudx90f6IhfCrduxepKbGvHvr+jHzrFwDnSD9V4KK6Jz+kF1
obcinD6AuZTRILI+6Uf7TO1nYoHvYwo25zeyi329J9M43BqPJvITUcPXMIBIv20hQL5LY5OY+G6T
VUaseNCCbfU5YgUkzQSfwTuR+89lWyqDq8LaRTHXwAtT/jMAA95D2tn7Og2hcGyFutj8l4P9CyAx
z8PAzRQCJCqJzqdDhachFat6DGTA8G5qA341nv3OFIjh5iGsrJf5sUOpHSqdAvfajNkMX92cUBA6
AU7w/g/xOaLs3MGMkTPgN1NRDK53vr1nkcpTG5qS5zYbGWMDjhzMQRVYCFujofMgAa+/PHeyZCTq
Sc6LlNZgzLVBwSn6z1Qc9QdDNiymQbUVsvFlQ3B4F0n2fYAbX68rPi4g1nAuq0JUMNKGv4Fc3qaQ
Y9ngZb4ydT9WV2hAtPClSpJJc1RdeAVNTFun+70dGdOnwcpfx49UFItMcRlcxzkwgU4lc7kG6i0z
QK2rREcAGgKh4ofAmqXAfq3Rh3UHTUzTIZlRzz4UiGfuUNw3OR9hw0Qtasc++9lPYgA6tU9e/7SO
NKHubslYmXBvlhDKH4DhQxW6Y8kNZgmZfbX55YQTDJL2u73iu1mXKigOPhtQ4S23fb9tgBfFHbpK
afnfzsMz6QGM+7UiNmBS6IO4u2oylxdhQ9vEX+KHDon135TBWM5jNBhWYM24o1O/jcPnMN9HPpZD
bWn+beZdqQV0eEKjz34ZACVFWMjdN9Z//tbUAUTeyHQ9O8c0aNbTildXvKZdMyLTz281exVAO6Xb
lLiujsOUBBrcnjG+3RmVpqxk7YxBkWwO5p1SoQXBPIjYVA3YQckm7sTimvagcTGIcZaNGXt9jp6o
MuoKBAmlkwqTIKqVgbXn5YvtlcGPXx4WcwRIwLJGQzq6FUn+KJoLpGibBWbAc7l/1MXXtRijbPuk
ZgqiJhRK/F06chI7TSEICicNuXHX0DHKt4FXr7mhpgzHx/Bvg8T+lQXvTHDoybPlfslRvoiuKwEC
QnOM6r2qVWUuxZ09NoZgs2RS64KwHIynDpJ3u+f7x5t7OTTJKSG5MVD9m0/MmuGBTsFapL7sDgQ0
aDQ23er/NcaHH4+EARP7LCyFgz4ppLal2LMFwl+ISqFAQz4e+CM6ibHvbOOhtDRF1/emNnVrUfwg
vdCRYxKJHQQKV+AReIZhHpgt6ZaPLwz9MdZ0URMNe8GeFwVQR8JuPUggrBbSBk5ZepJXyzQzoEf6
DykediFAXs6EQn+TP1ahQJFgoLC9XfFBOsj1hl+6pSyUym/t5JdLXDXywzJ9CWVOQCWtQjnUQ22c
a5Zahd2gRGNZ5xC8cts2ULPqo0e1Z0VJ36FdOMe7yWmQBizbsC+a5beMfDh+LliiWCTaunbwr7H9
2dlt5mjnnjDVWIanergGUdpJu32wzwEE3OIna68BbVTKpPkBfrnPp4TE+RJ9WyPlIcAmThZZvfQj
JztopQljIBXIDN+uJs7tcsHhQzVinZgS3j/UeSaxHO+czXwF+mwKXK4w7lspqfmun0leL/M4F7lN
kOlIEYfcnyf4qCyhwgw+OS/UQNCtXtwK7EyUDMsOdNyImgowf+XFgSdDbA0rylCH/5fwyjW7RTYq
n+JfYJKhF80QANOsZyTe0DIUq4meaIyOmTfi0EgVlr59H3bAwlXGkhR/u9kuDJIPI0dfM1uMn2YU
u6PLnRedB9VBcWyZU+SaaG9mRI9WF2GzDpKcg+ZB65J6mEZTKneyU/J1VRFRWd1HC0oI8C19LTzm
fRcbuboVN+P+sREpMl5bywa6y7+0rmw8RS6tx8piXTs5TTDq9PNmGuojdWtoIjxePxGtJR1sqWiP
B6ojI1UuISHWxmlCXjAfMksmjfvYtv7rSTJfn0Bq9nDXaqrPnxlwVSa4VrFNNEbirknE44LWpQ20
Wt6vgKoDDQYtDW/I3Hj/9vde9ghtY3qBaZ1NtTYWQHR51Iq3CK6iLtM/NQoomLA9oDjgQUHVgtvt
YEa4ZSDdoPeEUetk4Jw5+Lew4kOpK6FlZ6fijaXqFQgoOLVP0UhsG/7EMTkk7X/oCaSaeLAZmcpX
vuulgoGwwMX/JUWd5DFpN94S1C+kkWoEvlOuWQFJzzDx84quhEe6cVttfBEPPo6mGzglSLinKceD
jN8u56H32amrwfxQxHR5XX70LXmfxj72a++9RBdqgd1ycdkJJL3JDx+yGyj28zXHc6zxz59Jj26O
VaGsB444tP7DHuxh1vPAIMRZ/Vh4Y+xFWdxnnITwRqSjxd7lhHlCwJ3n5qhzaiQjGV3mzemvWnKO
xl4Z4JxIYymz7Hdb5eE2M48RPNABYEa6DOsqAtZ8HERDM/Nt7oNdsroB23AlIBSp9bE/sLkNrOxb
89edVdAb2/hxv1/NtfsBSrFUbUEkjNTgP981kmOxW0sUPw3hnf4x+bMHdCJMaPtKYbZJzslHeq61
WvYThXvaDeRbzJyNnQwWqx4/1LF4aK1H8H9/W1cyhAEkzKIoaNGzKXYA07AIDaopHcKUdTuAEwkj
DApJLUlC8tgQlkyqkpB6zWfc29B1ByYZRAO1QI9VA2CPrpR3zaXC1TqeJZC4IL35T5ZiWDAM+ZzX
KL+rN0wPWXQSVPiyxkh719mEYdNmxe6bfRtj0WE1DKSQg/kzRZPq9pMURNJvJRy8Y4bfAc9JE895
o1ix66uN74o0oPlBvAj9TEW1Hr7KzvMp+JyNreZXynsRKrafDsBn8cLi7WZiPaSO6jWL5FuulseA
WciPshIezYBF8Pe6zN6n7P/PC6qXUjqse94w++HGNRPnrpGXlb2gx0k+NStRgkrTgn12ytm11F/K
T/xHSOqHJDgD8I/ajvp7SeySExAfD9Id3rAVGrxeJu7Vq1ZUDz10ueup7Jxx6mBBNv2ZA5bBYXIb
DQdLbdmlPv8JFJHuKUdG5V9CIaR5726lzwas4J3YtK/IxqpWl25DPWp25EemTFTgSa5rNxJXk2Ms
HfWKF3THKniJSVGNBRrLkxbgrdlwY7wm05Eiddw1I1DMhoA2uvtwyLkC6nHiDqJHHGM0yUBP5R3N
XXcRCcec4ZFa2G3D3Qcm8lQrKwnRPArmYzRBOg6bugvwwoyT0A2PqBZXMNil/Hk5QawPM2CipPas
1RTuMHeTcS1FjFQBKYLMJBrLwuioSVUwZZBxjwmssRoWmCmqHfyY2B6npmcVyHrKgU6i4I9I74Rb
SzZPm94HVXwORdvgkI/dyeaaxFo8RYgWj1E/nmcrHhLrwH83eLm+198dfPdEdP333/dEqI1AYIk4
oGV2t9OCHaz3xElQDoI/5Es+vqg7jy8/ps8KqjjrgP3D1zOLbAJDnCe7O0AzKhx695a74SnL7JKd
JPZrHG2mxSxta5jBTDtDPOeyekq0JMVFxx1D6zQPzQ3zxVj4G66687ABpB5lrJifATuiOGsCa2zq
K9fQcrwdA9gVM14a2rApaSK3EU3Q
`protect end_protected
