-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ILz1Z+kk2OPyQev8mgHkKNZOYvCkY6msTrP7bFvh6y5LX2DbvHlFPG82lXJs9NSOlZDvJXpbNA4d
SC9ERqztZMkRN+WNC93nXU6kcHMxmvZoTnrOzKCXy/DoYgq5hcFbJfK/tld/oJsJhQwmaPnS6pt6
kk3yzwFrnQ4Sc6E5O0A91Xqf+M5U8qS0rewSwrlxNFoIVf8Z+oVGncosMQkv8ie9B7vTlB3WyZLe
W1E7r5PluAIn57WJ4lyiYiZ4xv6Eano2B8fOCuhjCUZR1Yj8sHkHujFvGw00RPtAsmRUpXmK7atP
8ric3fN+XBqe7f+11xVib8YUYii86+n5TbteuQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
J33t2OYioh4nMHSRuWT1zu62Nv3uFquFyL9TkHePCTYEJU22S6WZ7b6DAa0M0vEglyUmTCCp7K8p
74lkaaBWqeYtFblylDmy21qsnvFpx0dPTCWtQgxIJFkRR/TM3o3Uee/8nLyzX0lS926G7brpLMvN
6/lmJIgXGFtW0DktEa5k7aAIzir70shWlN1jF3XeEAfuE2bJ4ez7puMzZ/p+w4fID/qEg0ILXBUb
j20z47Gabc8ZuJNmUClIxeO6Pk03v4zo3z9W3Mj0lT+Hz+XslVMYPm2PsaZVFyItIkjruwMO3yxx
xr1qIALPu/PFpISKQq2u5D1cKU0HhvFsb3ysjEylDclopMJt0B/r/9wBZ/nyoJx+tfVLJeKhfxMM
FXtZTM+YWqJjJcLHxGW1HobINHMdjz/hRGPTHp5fzEOxHzYPle4xubkGZrsE9fThnbJ6OVrjG3+H
VVhszRzqlqj6T1Da/+nOfxaKl6bXVzJaoVm1pdLNbRfMJT3qgeSMOt1O2ipI88X3PWv2nXU2qDUY
uE67Ks+XTYemPRdl20ZvD8oxkv68uKNcg4xBNg7rZ2iHl8Nf4zL7UGOaAlpsYzDDXLBbVoglXpow
9mN4GF7SZD1158dsTVfA41VAMgUqymfcbWDi90LbeLl2UwkIhvxiHDfkEcIe41BSMKXgzX3heGC+
bOMXGN1W4bknv06DQ8MQdXWnWby2OaESxIiRaJpZBQ5JnzYbHH6hQIU9ty8HTqocKFi7Po0CtT+I
h90z9CrTGxUkd+BpG52GPlP/8wsiwVW+uS21NrpQQqka8gH5FqdVtO+wS3oyo561BoJJBs63/yD0
prExvXOfLW1oAL9FdilRpyI85XimuiodWbUT48noJt3LnFCQp2bBSl8nF9mVwCBGcKf422Z5HsG9
/fJABSgF6DEUzYVTLKaIyayrm4gP/0Ga4MQV8W6POqPPDuuu4RQEL+S1qwavFyGOKZbHxe0T5LfG
PrqH4NnrdUoF695hViEaeG6xQiNqJjU7JoAgb1/sDPzjSN2wUmS+k8SPJA/c1XWMZq+XeW38LzDV
1qN2FJCJMJZSqVfmJK3P5djJ/xXr+o1q9gd5dPdwnf8o9TxArM+XTv+F49KJEUfwzErm0bIGdS/l
dxzhtNX5n8a5DvKXJv0n3bCkvarvYcxFc9/oxN79D7W1Uw7yDWMv2JAA3NsoGEImUqsthLwh+7Jt
+L4/UW19QlKEQKzVZhmeB0Ss4XIAMFOYXQ3WKu2bCy51VdmzjLNo33E+fMgu7+9f5R9KnCSN+Apw
/LyOtpYz8mFZyCU3saOk8iQO96lN/OsH93Tp8GEGQj3LzS70xKaQ/H2dnpd3uslpfk7CzGVJxeXw
GT/npekEAa+1M7YYTG4Nwg7dpUJ/m6YhJJN+oG6KYHQPQtRcaFY5cAqWDlmKa0VTh9afKCQpyXyB
bqoi6wU47QEODq7rMmBE/WdenDHntMCOW59U8qWBbPAlfIuI82LHNkT5gOkUuoHEbQpPfbt4ClON
lTQ8OoMKvF1CvJ3HuBSxi/xKzw4wfo8EwD/f5W2eprCG40QM350mUpPi8OM5mKIQUy9/ToE+l9D+
wXCsqxvGQYCad2csQnEFkzEmge/AHH9qDbC/x/4GgdA5zy8muLunnHDQnvnLyRLVbaMJb8P049og
f9DVS5i2WZhk9cnvk59sTK7+HW0/rtiZqTVE1tKdBwfjoVBD51D0APQH6lBYXwon2IAra3vVbOgv
Bw7HPTbH1w03KhSToHbQ7WOdfJWe9HpvwRY18JuFw6V9p0hKx47szWpdIxt4ldYg89JynPPN3q/s
cywyj8tNuyBIfj15IMfzrvWDcYH989hWk7gxqxSarbhvarGeIkPrLHtigqYGaMtgJGwcrsFMzoYK
lnn7V63ePW2UJNyIzDri6skidc867gJVCWY4NTDmLB28h51zpTfzfogXhWhNkAE73RKjHDYQgRKP
6Ku4YTntREooIu4FhNuhoVOZdxQ+/9W3r5k0YvUKSUHsrSSPkDjsxu+rFx/tkOH2r1k8wfVeMbcd
CkQOZLcmwNNzd8ug1XUyKEtbLcnL/WSQhQSJ9b+bWGISd05TwX9WxDgcLuyjFavL/QdHW3+c9Psg
q0Hte+ugm8az5AgQdEMK49xFpwTLVZZ6+OR8XIwy6Juv8ucFmizRj49kfzModYRWJCGW2d70m/GK
B7rzkM7fbxKkXH+X4C1MSXEQo7DRPwsu5/KkexmytONKhM9gq8bapK9febe2gvD3bSEVWsxugjS0
qNTv3n5XKSi/2ZUr8kz6P+BF5LKLcIBD5j9pTBHTpPYyFMXWUld9em1DxSfwBe/y/BeweGoYHPwV
J/HEQIjhUZDoyozWK8MWhTioT1tm+z+5WtaQc3bQhAC5G9dj/TOz9wU4+uDizQNFZfbKAS+gj5ZA
HxIfx579AQyCJfPb6h//wp9iRJW0LfOX/l5HwpkULG0ghB7ukOMk6iGKdVJN31njIt+ZOoPf5cxx
BNOeHEARUhR4vOhGPDjrhoOnLg65kR6T57VyNalZLRj8LZC1iq+xiWk1r3Fy8aNZjlLhK3ooYjqH
F78A748C3XwZPFRHkq8h72UeeUF3ain1Ndws93EST+fW6FiM2KSO92BbjT5b3B/Xqd67/wJbAF9M
6CG/383irtPSCiEE3DLE7tEbHlas/GiTkhXET+9L6mu/7BfIXik3KOV60Qjm6c4o9iXHUMr72hub
Xz9SJzhzUQbCnY+3wnP3FTu6Ndl8iKIJXJtIgbwjp1T+J4Aw8Fr+XHqs9t9xHOjPsXAb8Yu27QQz
/zSNYmUYyoY+WM+2FSMKR6SDnqXZrtXH8I0J2RaFljBScwfkZBTcWMpiKQQbtpBogeS/UIqk1JeK
5HVvauPXo0MZPofIHgj6bqnWdk0Z1fyDkmNJAqRTiJ1OzcU62lcAO8lYBXLEFIVQMM3Xcu/l7eUT
M8kwUt95Lyv7nHwOYqDUTwhj6dLRyZfvwI9idlCO8PD+Xs+vq41VRqAmi+N5U1eNyvSEj3IPkEFx
Xe5w+z0vmNbryPmD4hlbDls7zVCVc/rTEnC9nm68kONSYpvNaXkZl2a6e231o/ZvfTgsEGminai2
2Owtsp4nnoFm0OEi1HV1qQ/mRVhYIV0l6IlrjA9G5ha5rOMuP7hMi95sG2GukXAHF/8RQwMkpn5W
gvIg8Z2so0OR+3bWTzQrIyou2sPVRWnH1I9gbHxTVHYGorteNKrB0647WF9jZG6AA+8rJRBbNQHC
KV4dR3oW3R/lTg+BHH1eZZNOyTq/QqE/ZK4BUVTazAiadkkzultL4ZtYlFqKdH3B6F0T2TN21v6u
NOOxwn953qe6w5UdOG91RHGyfErg0ylaWBGLHFUyFZJrxJU4RJ406tVlgfMJWHBiuwrjtgNO2JVx
Jmq5vxCTAIJKXThcipEwgV3Uw9/SsS4acjz1a7e8T0ftdlzeYSHsHvZzMlhh41RAuEfOH9wRLmF0
CYOHZG4CJy3QS6s95tU43wPJQSlNhea/V4GKeziS42KMAeksDKqVslMRmPsbG01BPSCKd1/0S05q
immKrpdeakILS6BccuB4ItKqDcJ7YysULpRkqA/I7jgghK915gaoQU1tmXSqhht2jD7OYvG2RxFS
z0DbHl1H7L0sGQDK5S9QwCdBDZF/vl2lwStMlKMNZVKCU2YNVfN4lYz3fTXTAdR8/mxi+hMWCBxc
HzRpysGtggNCI0kHxa66TUKKaRv/eaBEGcvHaW/dItjku/lhHRNys8ZEAEDeZNjMtaXtu8S5fjea
MvD8z+Db/1sUVfcDlSFbruCnAVpBR6QRlncGIx99mPDatoXcWzFdXh3/67B9Z4Oe/9Lls5jJDWc3
paDuLjkvyhjFcUTQLIpegtLBwut9tWYfj5RoX20ZaQYbanxgEgCxYj/+iQzF/k81mVHW6XyOK6dM
Ndu+488teYG6I/Dyh3SUzsIYfPHjWq7Z50ZGVDMCQNAX35LcGWQN540vJPlltzzuh0zjNhsBZFZg
Y881F0/3xnWV+6LuLMRD0HdPOoXI4saz8D3uyxxvvKKS1Ct1oelV3FAC2RXqGU6ePdU9nAWzJvMP
RIiPWmgEYbQ4W1UG5+Rkh0TgiImt9SfBOVF/vRuVDSF2Qox0KUNLA6ZL5FrS3gNRcANWkXrncGNG
Ocx2zxuLRMDFQgxzvjLJFGDvET/ClyyuWC8fbzXSp12IzqOp7XDtayfZugZGR/Gc752+oodJS+M/
5EQ9ySlklivpzySpsxvzzt5EeiqOyOvDQ4Hvr51XQIZvgaoWMBOBA4MYSzvxTOl4YC9/XDyk2yP0
rH94U8bYUhdKvMvvV6Yk89219tyl9ejPtasgSWJyR/CKTl+5eHXZqv/wY3M7ruFYR1w8HjWNgD24
fhO6ZaD/Yr83ssuhMO2OoRh3u/uAktyH0NZ3SOWYSohkt4o1+g5kY/Gn07j1AiqUT6qyMZvV1gQn
20vfSlkhRStruj++p4M/Ldwky21nXhfZOTPvexzfFBo5vjfV5bMRNR4iWRD/aJ5PFbdc97OVExs1
9kPN5L9nAXOHtXIGPgIFjycafc50uXFWi7EtGNmOaE5/EEPdvHk/IE0hBWD/9Y+1IUtKtY7C3B/r
bJg+apQL4chiQGcumTUIoBmHjeVuj9G+SY0VQQMe4nUSd+pYRgVi6LEC/qNZJlBh7q3nIO5+Mvhe
rXgPgdP9YcNW53z+Nl4M/BXABHYyD29+eYJM2kbd2gCCT40t+fEDpzpEVmEup5duBEWx8xqgCr7a
Y4JIP0Aoq6QaC9KvSbLnsNyTvIhfp/vuyIJ7uHjvnokGz9viaTixO85+4qVoG3UGLJWmpAH1uXFk
CKYq1sHWjhZ4l8jMWgVP/sVXfgs5yT0rtf/6I0P2a9bQlOUc6cfw1rYqfDrwwh/2FiQwb08ubyDC
BLHy1evvZXFN5oGGcKwxH0yENv1XVRh8kYoLx2WOexKlPn4LgLMgmQ4v8A0YmkFhHwFisu5q+rpk
v8fzX6O28df/FmTBLIJ2vBetkHVdDgBfr97/uVaZuz6/E5BXp1o225dPkwrzq8zM8w7f1BdHIsU+
b++RtdGg04+Ia6fGTAQQrc5WdyIIbq+q40WVmnl2+BciflxqB8lSe+mDKV8rJ8oVAVnXLaR2ZhTI
75RNB1CKQPmeByhTkxa8sxZMbWQKrB5dlaHvMChNHZKuDTYLLgBlOdYVOWa+Z4uI8ct3lEeVLAV3
DKUrFuJRC/fPZ8L6wfjemZyB7GwsXzLI++IzSjB5TfZYowDduLrlOt8Rklc6Q7tR7Zyg09Ib5Wic
WCMRbH3QkJG4DqIX/p0SaKSbHuqvgG45MZPAG/ZgL7SL4v+44Wh/0HfXN7rwznXW8ANchf6OomWD
vf5NKq6gIGgQPMrV5qYUw0jDTiBQZIC6peDDkCC7s02vRPWcFiKIAxX5r49zTmoMPISoQg6uc5FZ
kNfXr0v44Z0p1qpBgX3ujj2v0nSviIFOomth2mbYvAsA1baeP8z4swmkPvbmFLf3DLNTeZC209xw
7eGpCzLmw34Fb5Kh/pjVs722ZAXRumPyI2sSaiqce0LCrSQ3em6TR9jeH3fWPvLk9DKAo2YIHibd
LmOcBSZJJTwI9ZwjoBj3DMwmtNvEBSC4uvUbAJnN6BMBX/JcouN8fHstqDj+VVFp3EL/+ZBZ3a38
NnRZeTgKiF7Br33ROE3NffXHELbwHQ4MiGMtnt3S1jLh1HT605G94xBhE/jx1UtfRUlGISjkjKvZ
LLtoeYJypCNsDeQxMPfanMBs3EnD7BUh3y62rpvbyNNJiz86tlHYGySM3Bw1Lrk3GgoW3AAiYqU+
YG6T1JQQHbx7WS2dxSIqenNh50f19uSMKPW1aVXer9oyrUsq++IZN8ncB9RCMeSu5qA9b7Ze2mUP
p+eCQPIOssmx05yiF/L6qdWOVwf6wrCkG8hli2XW0jnODBw3oVCxyt9g2oP3o8dZqnoEo7gB4sAp
uHsy5OfDEa01tvdbz2ny/ls/bO/d5ue9+hDl8nJj9Gf1m4XZbLKvSyRFKIWenuWJvUoQ1Vts5+jF
cRm3q6WlpDNF9jvUuwnVTZ1rr9zvuHCsiln2GOUWxjcnnW3dTBJmJQvJe8JvLN4UuPrD+alL+gvE
uzx+woQlceUFU9tm5KhPE0qbRsg66/G5DLbPXXvVpraXA2fyUYG6o0rowdCodq9T09tP+RvWIcpw
SR9TtaBGX7yg5Si68TAWtY98TqGcIhfuucYw6cMxCNeWgKQ8koA3im6HZRPtO04RTEFyla9oDNFV
lkWNHfi2HVHRiGjdwvkUjoE5uASa6WOs41lnZN4lKTayU3Syi8D/0SXWJFN48LGQdnLx9/Xr7I6I
uRnRQOU34ohuh3ykObxZGtNatyRsgVsvXNtWrkU9jpkUqgzZ6JSpjZ5Q4EpxksjMbBxm+7qOJ7xo
2nmuCe5K7kiB4QEtM/p4jcNstyErE2Uiq70kb40ujZfwjqLItTLVlwMvx2usX3eSSCtMjYCU/rm1
mebsch7C1v+apB81EE07uDljlm4CJ6Z0iZcXR+sy1K0i/xfu3daOriT905WFORy/xmhSxS0ILhpJ
4ip7XbFShdw8s70yzSf81ncPysoZoHiAuz1LZn7QeS4fYtFVJz3gHQdrtAaPjsXY4bP4IJ8O2Lb+
+DltBjXw4iWVy/T9emTvF8x0vCBzsQsoG5icZnyRD1bNy9XIhxpQOMP4ztuY/9bxIZX7zJWTySZR
3a2XReyEw/WG+rSPNcf+ilU9t79dHz6e/2qCoIXy9MxO3vStaomdmIvTUdydzPn1aJdMeQnVB+mX
Xf1akoTorXFN9FhnpqXQOoUYnP8lT3UdAwQ+DIc9dZvxGMrRPChyxKh4EixfmAn5K2iGdo9e5suC
zkB4Ye9PrqKeYa6YK0jcaf5vHzzHcLgsSMDnIP+i0r3qELwmm5pAM46uo69vRwDVJ5q62THT7r4/
KEDUyp7LQgDDfLsa1fUSm92nqctobJM7URnmuOtD7CMnENK4AwfXtHtFSz85of8OdIIFDcMoLJ4d
cjx6LquN68kkmXXxE8Jfw5AFzmYXl63HDabSlJ4h1toC5iOB6yjabwigKNKF7WYeAgHft4TRu3oE
Q94b1dz/watT0qDYTzVw+tKHK/MQoUJjNUl12V43d8qIPnZjl7mXwcGzmckT7RCqzjg05Z3n08er
s40pcV9EtQ/9MxRxYZBzuUhSUOF2xb+cBb4qO+TDXSb1n0me8S7joX4Qin0CCcE6dbK6Dfop2J5N
7HQW1iRrvyA/gzIdZcZU/F5ykyVv+gEVt6kkRoBBR0cTVgfJf92H9/8EBwT/xx+j7ir6P/QiOfUG
MLfFNVAmsvkPi8SFexm5OhHq3fUbhG+SysKGIigOgqGrw82Yf/2fmbCNPXiaGg0GhywJ4x8xSQt2
w6ZaaLe7sGvbVExzrZd+zYc5my6Ljq4LNWAX1vZDuS+WnKjLv0oAppL+8il8yYrGhkB5dDfG+qxB
WZtVYdmeW8/rgcr3qO6J4vyDnasoJabJ8saevmRi1AEXleV+huubA6wbP9jWBCFUGMt/Yr12ISq6
itAb7fKQDKklZwWQTVZvmwJZdlHv4Lp6i8LxWQwW9lNTg1uWwzuOetFBK8p46zC29aJyqs3NB2Wb
0pOpUJGCz9X8KDNSjSufWYU5oIrXtwbpm+Q8bcoK1PxigG2tPRYEKIARJjWccNAHIZnRGgdVkCyM
8yWIMDfV3vAG3A+81OM2po0XfHpPpqdidgweQQ5Htz+c6aR1fYabaxOaEjo+gsiqv0VeaDvKrJg0
pNoe3ZjtwqQIf8rpyNJfmll4L2WjLv43v1Nhqyj6FHdSz4mkiyNaeBaHEXw0fkDwjOa/flsVMmMl
C0dXD/+Qkg+NapPZElAwmg2MODX90dtQvMaDAAeQeTuGEq6O8F4vkaxhs0gPzxXU5ZtaC6YMaW++
b7j9i9Hdf9KX6XBK1NjyDAyeP13GTHQ58w0XXBdtOnSU7BgOK2OgEjLmglJA/+tKEddme3YfI1MQ
gUSHu4nU84VSlK1VsFZs5MWu9DOn5WFnHW86646fJ0gvWIGP1Y7ZaEz3BDp8eSA0jusdYA5WOBn9
7Qt0pYjxGu+ZJfOuyPavbTwxcwX/5U3Gfzm2cHftpwmJPHf2v0It1dkGugQ6Us4M0vwLCbGeJRXe
1aU1FORwBvI5iD/PS4gvXXu2ZmWiNITVr6MMhmmUIMRgtyUHrTe4QZvBtyhQjVyd9UqTSmG9hFYV
Nslb6SWXPKUJktS6eHYMN2ZevI6loJoTvxqcJ6CF/yxxlapVKrdEJaScPkSN485XX5PVJGomCOww
pzTrSm9Gd6xz6iJVvyPt//xlE54YEOUmYBdn4HTWpvHPE0yoMwubC1Hy4zjGqeK/0iljl+Hq4cyL
0MmaVDypB8MkdFHGR/Onb8cRJ+bdawrm3cGFG+Ev1oIgKkyDMyUK76FiBo7TMPYifNpmZ+a4vuBz
I9nX44GMY077LtW8gbVQcnyLY6pZO7G7nKIXrA1YV67Wtkz0k1kbNhUSJtCcDNcWraXvOqI7TMNU
/CbIPIlVnXz0qx7wmLCRqIOx4n/S+SMMCRnOyquZW4YgOdDGZtnMFS3/wUZsSPnvEJwLUhmE37dQ
Kl/nKOMhVRMv43Y8ZM/hIK6nWCfaZ2Rq9zRKGm1icH6fuzPD9998cjrqDgX9hd3Hgk+ySOqeTiqj
gZ317ZXYS6DTq1a8W13Hwh9gQD0FRljHo4y/+2CYZvUsMrHLnUmlkLXYYtDXu/U926uglqUa6X0D
CD7LLPnKEqO5h4fMMoV0wxyohng2cwvyAcDWg69NmwoHVt/s4aOYeJx3XXT2u4ram0uLcgfAkrIP
dAB/cVjtE852TziIwW5FOYbAtaZbIlpRNAi7NEMx8BXnka30z603/3cjc8GcmjjShRJ0SVVTEiio
NU84JUTv9jKAytiSCQKiE6ARlrHXpUmjPLWb0vzX5MKsO/xR7pxDuLVzqWvBlk+aJYkzSM1c6VYV
X72A0yJxYI7WABTnG0+olgn/KZsyw4cI0u1cd6vzGeHct2m2XyVHCMG+WVoLs96ghS1OYp9Zk936
epnAFa9cZDvnM8BDuFbMppvgvW/prtvwzuSOUHpz1yfQ/MjcUrswhoqPf6tx09Ug+lhN57On0g8R
en5NrlNd16w2JsI7r6pvzDOR3e0eQyIJvoCx0fWYGfK1cjw3cyOWWBRl07GC4sWBYkiTk+z8a1vB
cHktjWU+scHr/+u4Oa+oueGaWQ+GvzU8cI1HJo90KgfGn1YPgvZNIUkz5wt3BizzezffPaRi+Yv2
DOGXV5AUWREmGYMYlnvt0YCQxE3DPl/9zGj9Do9NzGHSoS4V/e2lHJLmAoWmczoMVjRDs7CkPsjm
sw7cnxh7ICn5P/xRxCukdOsxgxEAwL6jqcCEv0brCFPPNF5It4DRePswBwYm2TZSDrpKK24+YTKy
YoHUSe9hE7XU86mDV2ieC3PHwLmGSTpw6zyZnNfE+Nq/LQRkFKMkhly7S/qQH96YBWuOq8SX4Awx
ylkR43fp9HC5d0BC8F4dacSbzufRzFVQDimxxz115aZz/emuehuAsPvNEvSitI8ZYzMDtX++NdAP
o3VyDlXwq/YcdsPY6W5EIHO1dVPc3jziGg72nAez6H0DHoWbM9DjcwGPhZPLejTpqikgoGzwVBhC
WqFrv7gvjo3O9c8jFSJSagz0PcU/i/6myw4bpM6Alxm9h1/6PJKHXgpS/bXyZZbRUJyOnyXLHK98
4n34pQFtCQNucdViD5pgRxAf31V/12aL12OHycJEck0/sTo8CCc0jxjP45lxc9xkpvT2YZt+OppK
VRodS5L+FAa7M4mnBWblDnoplUf6g85xUVywBu+hmEWBmqCQPEAQHXH4SjnP1QttkSIAxyExlSUx
4I2EO+XUTsXAw7AnB/xAaj1/hRFltXuHWCpWd+7yXz21G7thVPOXry2RlUiNmaDtIsBNEpA0/QLB
02Xa2MBdu8q4R8ZSjC7H78FWUhUsZ/filLzqb+WDx98eI1yod2inmUwK6jUnr5lQQBApXIS3Wcz0
3hGrVBiF6i3w5db91Jk4nAl/0LMFrQ5G6jRif7m99a0QH0tZLzTcVF3HdofSq35WiV6ixix0vrgl
Nebu0w/HwBXy8p9PW4lDgR1Fevp3YhH8E16BoQ/zf6aVKRFvSFh/040QX8VXdyeGtVGd5iLQVXok
jZhU91uuWwfk3fcdxqHYrlw2vvRaYW3behIrsiOJ9hk8DFLVq6MpOCRcH+Z2c5pESldOoChsoYeH
ofMkiEHnEK8KhxCP9J4EcZnMiYeO3Ba+sK4my4We68bnFLGKWDe1MlUgpAmIrwrdZ5qsqenczR3+
iGYoAY67HtTR33iSlbOi6Bkf1wePCDSsiHkym7ukH7Hwc9Py3GXUUc0ya+P91u4Y1Oa7NZzlLZd+
yXA/WCpWNkMXxZQJM2z0LD3YyU/7sw6BAEt2e6UyEcgkT6FAs7cbBocjJtAxWihEc/FIpgC4R0EH
iPiwPdx9Tl/zrDfS0LAkp+lkxto9iQcwqHh2QeEKiFAoUdgW3UeHTRX9RcH5+UrUV0DSLEkdgC4s
ju/EO3MJmhCe9b8dy1s5/h9bbeQv2bIFuQcUH20M3bqqDzFKTKnnHWoRYZxCoN16AtTZuNpXTjAy
1tgsiTpoOe+XdaR5bLLTQDJ2xgs6TRGXg8tAU+FufRuBszW4WPoHsNZ3rAiJ2x7nBtUQDyKNQv7b
oaHBPZuNjvxXGYOKQDhEn6q16ms77f5JdbUQJNdzwro95KXXlllzdmzgIhRo1vNxEo83yM7eSMa7
Gm8f8tFUAczNo3uKSxbwDIxSqvtSfdXNyE8R+9gDWPH3Jcn1/Lo23wVnhStsH0DEtt8UO4TQdlIX
NLqY8FYYz4rep+lMn53fj3XBm2u6D7Y7R5oVHC25tOpRCZ3Nbq5FniNEY6Wtzv+OtePItXSX73O8
MlihNY+J3u7K+byy+gETwzDv6874OiNj2mJIQFF7+hyBzmiPYcHHVr5MRmSxqFgm4y/rBc0cqSW6
tSp6jnbrMnKfJqT7O0vcpc0VCnQMNs/GtCf2uvIsgGBKNMfCidXhbrO7D+26nT8D6x1YeQsMVM5g
8/Cazu/+BZAxRmGFTTfG1BQ1BdHkwcgSLXIABVyJsqJM+AlQwqETGXue3pHl2vxB6LW+X3zNE3cH
eAFDfgonM3ROa1ZH8sQO4CiaSv+Fww1i+61Ratg+4ZSxLHWZVYgjD6VlmJqp31Wl9jkfdQ0EBeR0
TndUvPe7NE0Xu73myAb535nTYb3TBbNs4r21yjSGARCisWJlGa079i5CfxHHcTjKRqfKEaURDK22
K9rn0lt/ayIrBnJulr0R+XGNJ/hga4DkECXH39fI2jWgkmYMtFIMw7Cbx/s/exfM03t4ySEYIwQT
M+6xpP6JoMTbiRc2oPUJkAGXZcF+euxsozsjxS6FVb7A0yeu0a+ALQ/24jXRTIdVnuoqrtmHOFUi
osZ0HX4tmnGwBCrCqbJrclocROGo0hyiMRbKbNOrca3ha0OmihCQq32M2+SNYKsvQppsVihbw8Z1
gXhZz+W2uzGZDCesoBhSlrm9aW4LKB40fYCyGoXgwKayepJlLLhRlWAD/bxZpiBBB+qckgMdyXFi
YgbGYUYEx9W3kJ6n9hRvGJiu8DAWDdwYRp1jtO+jpAKYRTkg735/1FwGXzbwM2ezW9h2DuVOJYFW
dx6G1gdQNdgnzpxQDy3/DIpizKuHHlJWFpioIuOToSpRK79u2HxEubLXGhBjE0Eum79fyiKs6iOY
ibqSerLnli4joHOB7NkYJt9jvrctPyOmkhEfFUX6yNjTz2rZJ985Nus4sRg8zfs/ywHZZobMvqCS
34DjSavCQAG+PN6S6Be28oO3s+tiwzHoCY6PdcTwMrcNBpdZNY/ZEGJhAwqTb799HuOwpKbKZzS6
BBvRpPzkre7/A/aTANw6hOE9rdhdV6lYYmURKDzWjqEP3L9mIEFzj0qbi0pk1Z6+ezvh5Zs5ikUL
ZA/yvTLr3FIIQpOMYQRW6qsiXtQDw8WTl6i24HzuYJCGjtJvUaGu3SQTRV5fQOA+bS9XUqRVIP8e
GK2i9KcIlUKHmxlm2fiRmuDdptrDFZ38qBCjiaL3lTzva//dEcwFFXzNALFMSyN6CN1GIzKsbhvJ
Eod+FaZj7neF2qC2bPhrgr4E6gqxKlvBQ6763y8WDQhNtlm198IuGfd7EfyTUC+QWw+hlsXkhk+g
bWZ+rlL8uKhsAtLv31/hwPkXXzQJgPfKFdK7gvyIW8NtXUEcMuKwBEeIwpmMRLV3cpyJRjXX+KM6
lz+aQYWylcnchwFJnn/RShluJuJTtToQLAyOAy9Sv6Hf4lWl6SX+i4fQ5dnMzxKOY4X2LVAjbJTA
R1GyqmJNsRP2IsgyZ3nq1se+0nEAOM5TXK/Btg/AClQ3xRqqT37WRiG+rgYOa1r/WbK7XtuKeuvy
9hEGSIuCURHS0Hn8ohfPTlOGAeoz2pIcxv4VRp8EKrmM9ye5KZ9eB1/szvpgSx6gZOnXqlaakzGj
HqHepRovlhckIKKJ85vi+W0SH9RajSFuhJfUQS7j9Mxbgf3rNXwhDIsSmfkfZ/9+X52iwSyCUTiv
s6jz91G4cNrWbGNagv7fWNTKXQU1mNb4ogMaFWEh8tslJUYDrDnUIqGJB4FS9gQJIN+jcfHaQurg
LW6PpV/eEyM5mdQqF5RN7IqtgvtyfwucgteAQWPGRE0ZUUr/Q6uwEQ8uWdSjqCJbYhoZvx6se2LH
Y2QSLQ51IiXBMNdUqtJ5Ix88SlDVHF+wgFS3EJXk1IpD8uRz6yaiQBDIyA827NUXab3mX3kwNu8o
8UdboPNz3DAXNBd3eBZa2xNcIxp6Qv4i7LExEaqPHDRXyj2aDdMdnCNAdsHVQlO1ZmnaaCGZ9yuE
NIZ8lh8ck9ySIChT063X7zx9dwLEGB/4FTRWWlVdn0V9BhiHWl3m6WcV/9kL2AmIIjWhFAY2AUt6
lDANcnZbzI4ojqGdgu8GKaM4A5feISF3syKqUxadveFbex5TyWh0ZwqfV4kknW9y6S9IgVONOHbs
Kl9k2PAuS0AGfHhLGhUpTKDfrFKLEYUGvo34rPos6MmOKppyWlu79hcLti6+6BN+ROj1Sb/8zbe4
A6DFqMExlowy/FS6vNlYt5o9uaUVE/ENeof8wH/SCa5OKfCNZTQvAr4r4XheN7++lLrJzeloSfCy
bmpHLdppAaxShPIUmw5yZKuKneTkuV3prRXD4bp5zQ6DRdHno49ALH98vNkHCU5fnEXCEqvk1XEq
PgUO2/Oxv3hBG/lCt8fPFbw4xmygt1TsbWpsfhHOTKAnqGVQAptkJE8lSp3lrQUmG8clWK50mdoa
Li53xDqvY7ohIjCy9ed8lqpNoELhaNLdYEgxjbTt5lEKLr8x4nnPMrKcW2i4IQEduVYFt4gntN07
UOJuf7aN2XDHHXlOVIYJ0vt8e1xGsrO26g4F8GhqN88UNUplr+mNiAOsuhJ7gF7c0HxPZOomHNEX
7RanEeoDYs6PuxcHqK/T1g1k/x2CvnnlGMGG2h+UmEOZwgO6hsEsWmBWtYkgAFLXpFrheMtqeg6g
EahVCC+f+NpiKyAw3fpt/O5NVnyz/+FzgshA+F6eZKALskzWIfuUvf5TqZbW4eCZdBu8uesHgv0w
d5oAM1Xr83Bl+ivhQEda1/BxU5U+YAy1dKi8+gY/wOctafzhfUpSePW1uCGMEdyrYdQy03sejYOG
oCSWMd5LgUgR0JMUWqEYSsiFsl8mO55Ar12LzwFMvas4DT5T7EZWc2D09Km0XdH7xx/hoqO49ui5
KvUuScWVLSSyYxFVEFefPqHL3nctbHhJcvuOJseqMdaGxwvTWy34eeILPsOaJ0yo4cs4YWz/RxWa
ZXu6SFXZYH68ldrSncR078fL+Wqln6ZL6n68fpuO/iZi4b60PvcQv4hnFgIP5fAbwhR9gPuTqO97
BiiT1AB/TzW9Jl3fjbxYayjcIGGZRpC2ElOEwCrlQEVMs3RsyzzAvezT3XWpeafS4oDkn1YCUXu/
JKZkfjTiC2jO44Dz8bx9DbFsB9H+QpWgzzDE6wRA3XA3O8+JO/0KpouMGbsDLyvvQ5rg6xjUidU1
a8Iz0j337aj9BL+i0dmtGlENyemiFWd8AbmyGuzla17DR2ScQUIfKXnZkJi2b/obMaNJpm7BfNph
a4LfB7GCLYy1TTuJZILoU9Ib1jy5upMP5clu7o9cSXBzoOTqf4UlZIQMHzgwpAi6HF39I7GQE6ZB
nP0B0Du0ubaosQXjD/OIH2YvXExupHcC34Iwk6svTTWvKUtLbbyM14nUFOzN5Wox/EGtM/rVindO
bufDOZioS+RGDpebfipQ/CRT25vfA3u30uI5xV73yLbcXFfqEMf06e9OYOVXVnDls6u9haMFTIqa
9ICv2MGHCdWkI4Osu4ObLL+/THGTzQYi8X7Yaxd7cNvWXwHw/tV7InLuDqRRG4+9H/tIcr7DPwt7
lmzpCGvLWysyVpnz5oyGryLQcZJrobauMAaRSnK+O8n0shSBid4zcctO4LYVw6ZPNPXJE+J9fVs2
auVIlvozjQ2/TZ5mm3C/Alxfray889LK3SXW3TVN3rsDJ1dJIofeajm6kWObOMc7HaoU28wi0nzX
76v6MOM78rIZRnIDaKocpQGOiMKb7GZxp0vALfPndB83ZZ04iZI5jJIm2nEm0yfivdT7HFC8yVRp
5ojIP2xEJ6/GG0ETkq9gBU0TEZHwZQA87Tl+47SsiAbxNvPa8oNQQbAlECn32mXENTaXFIrrdh0n
RBqfLZ2wCbBsTGZViP/8iDqWTNZ5zoO8X5hKHUUgJPGHprQj7wvCaJSoXc7P3KZuCuIQ9bYkwROp
3Ucw9m1u9Xb3VkfkJKB/t56MR2m2D+01fz36oCag0kjk+wWmMiRAt4C8lqkH1cRpMY4E/ISypUJT
NXyeVYHUi7i7vytmxOEDC14n/NdIiJvOKiyFnde8xZczlp1z2z5wEVM5dIOjOBbgNZT5frtNZta3
2exHc40lXpwLBjlPrxdTzo7l5OwOmAqMx0ZaV6/eozDed/oiO38yO/Mzy4a129fxOBJsgPzcq0q2
4JSAwJFcCLvgNZZcF34Ioytw5qNEeSz3IxeklIadc0kyEG+gUmKlF0CfFSxjjeFrJXxM+mIYXZfI
FiM/5kTP2uyq0d9bA95yYmHySPeBiyj7lGrs23oDeow13zTbpXFZt1P2AAnf2eglbl2qfudxqXId
Jd4HSpUkCuFFQtTrD0QAv6q6SCzn851WKf/j3M3hkl3Dpiiud3d2Qy5lGURgnrc+YD9+vYSTUJ0v
G6ZCQCntQi7fws55HGPbPazCAeNa1FSUtAhAnGfcwEMjqsjuJ4+DKe2Y6S6ySo9QfjSlMx1Fp9/5
K88EEUG+fUa9sxJC01C5SwviTru4iAMLRT159VcwLMGf5OeVj7JplTD9vOuoOMpWzjAEmH/c8ux5
WxYFxMY97sno0LS9hPQ6ykkMXqNKPsl+fiuqXhmjlOfpGsqpVk+p2+//P7dd7O9yldqMDg46ToR+
eqNulxBgmLH1QAR05GaWdiKQS5qQktabs88OW5mY7JS+12tGgV/RSMLAhbtID2SluWEY2CWVDpER
6mJZn8HSmkeHDLKJQwKjZUL84aPsbTnwfDTLtbEFR4mEAdUoh5mcFiiGviF3738AHQlk3hFd41fo
r6KgUje54i64kBU4z2qgpTBseXB4rW6NYrTnZ0zsKALvY9oTZJwrhVpIw7xyFgQOfVhEm1rByUtx
1NR9F78DKKH1++nlhHSf96wRBkRf6EypWAsNY7UDBNEZdA+qLQ3NR6DoN43jJRzCrH9c4GhIPTlX
UUML+ShUixiQrA6DRObbxeDSOzFOoew8UlMTMyOoVEysSfMMFst4AxDg1unsujBdkUdWKPqzjrig
NcStTRTmULvrISmt9IBDXc1eaucNZ+h4c+r8d3Br0tXNFicP9yKlQ9j1tyXegZSLPClE3FdsYAVJ
FPw7OdABFgUw4GSUO0IdsTFQiufhNjlc8wt84Xx+LezACIsHfSDjjGtPVyDpb2+zl0mUfsp+deNk
NRk12Bg83OVzrTzPXWyGPoGKGaOJpYWYNcgTttcj1Bk7a9ytvGsqNQgq7mIOlPiB1SVi2FPTlOPt
yCoWXJKmBY2RgiqsBk7UMCt8uy3yLnWUcaN3hbLtEqD7Ej2t6i17pCF6PS1jRlT4ZyColZ8uHk9c
MVvhIbmSRYeniZxSBDkc57+gY3HEs0Twx/Xlq1jJT744Oj8zrJ3g4FpuvcbiWicFFl16UdsZ0Yny
+eYOIIO9ZQfqEEfyzCNb3wL9yi/muYTfNU7sobH7Hb9SgO4LUKmH8ZELjN5oGWGkZZkA9MWdCW4K
VmTIOat6uOqQpEDHTRDY0vLSHBL3OaFXKKJrxvVEcripl/3/J1QJY0a6i/g0zvKrV47lJTlIu/c6
lAPAOGvpweTDetXp9Yn7uEUWclspulXr1ycg0pBuVJsQnZIBr5neH8xvNnK3NKZ5fk8mpznB2wND
HcqYoBxo7VXSr/3A5m4iZzof1MZxxCxXpoLVcbIzfhT8BL5ZwodGCPnGsOl2UWmKgwolHi2gO19d
JPv/4t/l2vrJGvrCOwZ+84Fl8O0OLWtlsAgj4cXYM3aULC3ZWg5Ar/6sBpG0xxZ3gv3F7JZ7pkf4
x/I+QGmjopDaERnHXpZ83h30D5GHpaQXXX8XQ/YkNxCkt/fumNu/aRksFW4EKEB0dgteGl4ww8EL
n6kPloEXkRrtoV1H8MfrgqWdTRe6M9XzbcdvuNMwZA8HxR7baDRDfrCB5dy6xq3EuqQxqAcvWPOO
NfveqAVTLkMwRH3wDeaHg3rWuMXhaOh7zxCNmlrICrMXQeLTraEuKq8OlOKwzUeuiqIjNP218rmF
1LQrMDp+pgckeHpA43M5Vefg5FgxVcyHxDMSMnj2Ea4PD0BT3sseuJEHM01T5WecZXfzKfiviofR
coWNvzBlRk6jpGCD7NztBP7M5A9DQqP9OKQsu+3z6bhL0mJK2X9T4EgbvCjnpgkEBLeCxJvOA/K4
chwu8nB7hdMSCjwcIzgJoWg+2p7qn0AYuYk+MxRj9phkTuTIFAyOU2F0ovAXk5SEqITVUuy3Wil9
8WOOjY+xiFwQHgmeGQzR/uAnk7rE/bdQvCbCxUMPbLU7h8gGjG1+B7CzxcaBTQc4NmpyEamVvJWQ
455CR0BH+VOfpl1gJHtGG3i0+zvrsnsZhicMxrSXF8SOYdHYkOanCtxDJ7aXRdiq1PPO8n6fjphw
E1VPAeYrTziNx9OrE8C/PksnuVxomEMLpN0peChod14p8JO2L0PaQrR8hzkA2HxGApcdvJOxAnXF
yXgHv5cpz7x0FH+v+jgEOinACR0gGdMbA258t3PY2heMCG+RSvjQ64Gq0Tkni0zLRajtzkujw01g
IGRHjMjq+buCRHJSOuo8PkNX36GpkO2qFRfx4togH9ewpajgRb5YLSWgkMLLsPrgfuSFbEh8aumi
r6wuhfW9YvW+Zz/GbeclOMjmXJipRd2u9UwR2jhFzmdZS4jTsYK1kdT1yjRMFusCY9+Ff82iuKlC
51MPfegoXW4tSAmqDgQ2Qcz0aEcDn7AxXlA/Ekf7wP1MWAJSjBzFjALol2FCuMsJN/Et+CSfAtr9
1z4yU3anUl1ioTu6ALm6V22G+O5NJFkVoCvmW9Eur0Civ7iFwYb+be7enMt8Lh/g9oi14huscMMT
4GgcPwG9osDHF5z9xBbffsYADB2Fa4pIp4759ixfwohpdoJklx1qRFQ/wqikzqJnNvf77R64fYdg
g6cfi9w4OQCEx1i8HiGDyGazHgr/AwiydRt8UkaM/cxvLmNKLlVPoGyH/UmYyowIvFcjb6329clD
a/lQY1CqerrCPa25TwGdWumPAwPWVu4IeFynzC/wRBUL0MtZpUOuAu4uDlzuzvQ8EfV9Epx/u/uM
WUevFoZbVK25LK4FUbwaiHAV3EZjaRpPkGdDLZVuGcpx+1YvHaidWoey1zlPkxJabhutJIqURCxT
mmvZTUFxzGdw9HdD1ku+mSLat0kUveQ1HWNr6BcgciPVqbRbL0rpeNbj7RC6dbPZ9aXIdDNUPo3N
OeJU5ASKgkBUsFsk3ecuZceB4AE+tWVryYmRpLJRoZf4rwYRKWkmx0DDnq8+nSjRcx3+TSRm2So4
To4QeweYOGRK/eBAZ9WiC/818l4V15lIRU3jpab/AbVc1g0OAZBntQB1FfGC9nzXTNGufwzQ5kMz
Pmg5yEiR9+N741pHU0KFoldHdpivkSuxShoaB7BZds1GzFqqtXXCAfgLBp22vsgCiW9YcyP5lTJN
W+ZKf7WDXD3Lku2/QU3699R5Mu5JVUty+dzh+TH77ajYvV1eqKxS6wpZVz+hz/JpSakcKr1Wdh72
0tjD3nFBjreUK3ITfCkdp9Gwuv24WkwsVOdgP8FlkuLkLvKMF9UgCvNYDLTXNrbwAX//KysUJw4f
4lhVQEkhcyesnbdwMtel4wE3XVk38jX6il2iBMoZnYhsIlajNIQmFCYGoEEVdeJXNBMgct0d2cAe
47VfN5544TEzXVUH8h2J9WSl0EHoUDNcGTz+Fi/CqOkN70ug6CRnzmMPC2k6rk//YAZGx4WuK++H
maLunxa8uTScAvEGymga4yNKDvBHHscZKMrGWZVvAdP3WSP6LU/BFDD2cbynZlLI4sA/37VoFsdK
t0MRjoHLzFypTBe4NWhorJqgk5Bmm75Acj+YprjKMs59hBL9qB5uLLH2onCYndWcTGClBYiXx8tC
qODP/yGXjY7mcIYtSBdwkZ6AQTn+M0WmOhBuv8cLRmfI/jzLAX21sKvQ7eASav4kSco5IKkLAoHf
FP+NEEUQbFOK2YmmCVTgVF0Hrxv2n7eT/2W+pcDC85RlW+e+HxdQC2PhSjdNJJJsm2lu7cR9sW9+
frQLh18cCBiUAI+tAC8YVx6yhiPb9n7/yN/pnKE3/u5SvTszVL1Vjpa/Pezpz+7bYHuYOmlPH1IC
TtgFnnTptJgvI1z3avHEqfMFi3UGgQVO/kXOXCMBZPNnHAG5ArbkZM2cOnIYUOrgNmaGoREDF5UJ
Dwnt1umOlvzmDcLONit2K2w9Nz+ZbUuqxlAj87XHgs4NvaWlkQKeoqSUJkH+fUG1/iUeSbQc3jIr
FAbBYVE3Ssd12Dk6PO6QPs60o7+VBx3xwaMXSt+u0+4LXfigxGYwYfqURPpQmICxoGJtBZtP2iGX
nXgCcUFgTUU/kWDhoKTAHWKSiQGoiR2+Js7gTd1uJI2/ba/+frgHwu8FWP5sX3VkxDbRDyfobYr8
gOcRJaGoSODn5gIPpdhTHJyfkxWxwyyQIzB2LvqeZSk0IfYjU9rP0m3kII/PNOCgLB7okar9v7Kx
uoimvmYwmWnzsj3TbFkEbShGBt4Z75PrnF0T3hQVRiYANDdP5xpWiVwKmi6rW2QyXePUI08Q6+WU
VH3Fx2ZELM7RN2g5FDHc2s72zH8c1nfBZKw6GXcRUcL3uSJcW9c6xvExvo/tfAY1bkXHC0pmEBf+
jBywCICU2Cl5y7YDUbrg0FScNNoL1yeEImYBhozY8liTkx3uTLQ/bTQf0HQwKWkAcpFDQTdkdIrg
i1mv2MauDCRMZ7sdpfdD+x6HCufvRu+f1jYhbuuYAF2I4RY4emF6C63uGcV/pEtPrCYRZg7E7NiD
XleqLL/JIO5w8RCbWZbPZyMwUM/fRZBXPz/n8um0M3LpKmOn9qJrmOXA+ZLgaejxUV/r6TfPlrEO
MjD5dMHedsUuKSjwz/hmEEEjQ2P1Us7I+bOHCrQyN6eBNNq5lYqOnrgr56NZnFoGoCauy3ov2IYm
aBCdfkyuj8GRMBewlw5B9fVkWh8MeeWK8fwbZ9fMTiImrTRluJehAct34rlEnjqkitl0T65mLioE
Y07yindM+aBPbQqWVXA5dygUV9fTHVySLAXqensyCnUzkagUt7mlHDrQfkwDzXxjXCOM4GLo8i9t
aVTpUZJEFIMhvhMrp5uHsPEl5SOsCa3Fxy9hBSv1fYVSdxGltN1m9e3RlaKkj2fpFqeR4XxHq1Rb
0ZF+l1Otz4FAs++En3Kk/at8qoGpwolVJqUkYbjuQaaD1gSFsMR98189AFAnhKOM8kijN5e7D5+j
66lo22ITNEPOQiZl4K1pXnWNBbY/8U29tMLKHHuNRBOzZ5tv2oi6v8kIdhaBe4wt3A2tS0FRT8RF
URmbFeYhkI3eyxQosxCwX5raLzzMH6XziVadSZkN5N0QtWHK52ASVq61q7+jHk1F9p4GREuCt9y2
7WRg6M1hRc7HK/7JVP/j/NfEMcWVBm2E+877PlGslaklrBjAehNPacD/eB6Wx70M61ZdofYpywpy
IIE7MHd4h1DlpLtWngEXLhsZ2bzjiPGl9LbvuT8HdzP/Z/9mm8cygnP1uDpCuUtaLNw72h35kYrN
S4/rZ96vKrCZt5ih6uAyHecnV7Peyr8MU1nm1K/z9NHkFhyKjSZ8rkZRY6xclr3eklaag09j1ujC
SNgBLtYx97/A1o0j4RQv/Y/xUlXUZSqyxlKHk7PYPuU3najVPLFD4djSev7tECGZ/qDQu9YZr0jk
lP62gsz+oFJhcxDw9HI1zeZYRRecXOZRHt7cwjGs8Et7SGVjm3kiTVgrWsVIfqgSCsxvMBxM7d6+
tIOpu6C+aQEsiWUxjp01J4PBZtBLTDwFBSUaL5tD7HxjkjY7lkNSVAcz1svuVyVGK7Moc90+FDlQ
8vJXcRnMACn80I9d/hgsJIMU8/yfEs2YP89W+PW7LYepvnfzjPfG8Duw2zLwWCVcp+8gM5Gslc/n
SXqwHwqQBsxGGYzYg3ZQbor+dLnvxZyhY1feEpURXUZCJp6/kgu1Rve/dB+qL23AKLRQ0bDPZ1Vu
6sVmKc5XGaBpG0qHAr+EcNh37Ou2F1FS9m7f0MAsPkjoM0/ETzCjPWqMiU6YWvJaW7SfRKCNHSG7
2J8KutNlSS5V09N0PV0Qm3UhTLN+wwuuNSzKxKZwozirONXgoy/7OZXKNE09t1cDUmVFXaAw7etu
fJX5LrqAwVBUTrx5nsbHP6H5h0Cs4/QT17RIDS2rxAYyCCGrL+Vy8R7o6bPNIfCkmspcxF79lPce
sHe+dsbvgzC0yDVWMDzz1tj7fG4ic2DpzsTQasrBmyziwwyQbMvOWhsLe2K5vbZH/WNOseTg4JgA
QAb4/x6Ai3Ak2i0BQVhbeZR0iPEjV/fs/QAhkKEnKSa9EYRdaP7/GMu6wHcH7F0alEvSN6hiwDyD
Ve/fhWLRALrf9DHXtqpfOISc5VevEVoqKOh6xQ/xpY519PUj+SYTmrQyu5AD75L/SK1pyM7zIZKs
9N/6hkKo2RbnxfQ2LIyvvC3mqUzHyAXEgA2Si2O7VPWQlRXnpJVIUUD4pF0JcDR4NeRqPRTJgqra
rZ/Qq4Ly/Vq2Gd1ttMGzKJ3hpRKsfCHC9uiUfQ6WcEXGwbJSE1dFzSXTe9PDBcWS9/VtF0YkVN2i
qJybwfKvmKWOHbxH4RSeI551F/ufYcLv3NwcVeAaccMTJlKGm/5yEtXpcqOeCYIER0ijUgS81/Kr
y7LedGyaEco9iOULLXhvaFnedTJ5eUpulhp+1A8XbNGIBLL2142R2Tetq21dz63aZRarb3f98jU1
2P6laPMPvtua/sMcokbGiQFkONlFWIg2l4kxGCmH4zP0lIoRE3reZ0N2NSuGW+nxZEPPUGzuksCM
DAj+ESNJkK6UcAF2ISm8je7ne4nd2L6ALrZ8WSpAFiDr4BMJ1e6ZJBSubzEPYSsjAUWxMAvbYzRC
bcyVnaVwMtzlFd7lfldKEHhLDmlNaINwqw/PkLlmVxpG9nS/xJe/MrE/CeQ8L6vTlSlW1ixHy2+X
otTzpcWp+H0ssvC86ted5Ykgs+IiyphcfbqvKMzupy2pCB66bUB1R0IXosB023M+yKUw4yJrqDUV
9EjalL9FNUg3E/dFR++EkAMViK/Z2o4dN8j5sUWdGuSmCPi40alNnr9VM3OmKysoQmQTXlSrM0WD
4j2x9NrX9Aakl19cyfEwUMHS5uUezQfJDdCIY5QUZG2JdNCH4VmgRfjHM3ph+zay9gNRkNQS0kp7
VfA/iKjdmViB2xCZlKZjFPS7nyEegZF4Qn5VGY2/4uqLFWJsyPajmcJ9uOpZGyVKnqikTCly+bF6
3Y8Xkjj968xo+1eI3AVKzh8fpqSwZ/QZazjRXmhbbAeR5ltm6qSmylYq1XUDFYdZrW+737dt3hDR
QLD6814WdmmcUqydYvjVhYfK0vwQlx06vbPrDt76/fyq/GrWnwIl3DrvZP3sy0rxxwr1jXLHwhTB
YX6RfXqQ3C356ti0Z5unlqwmoNPI0g+oojkIll5LypHD3hXv53186Ai8aW7NDL/MmkbjQOe0yKOT
rAhEMNDVexiRiRpy6lJYp4ykS6CmVLG9C6KdTw7ZqtA1K0ZYH1rerOC1fzz24jgJOidHlRGbU0yp
MkVYOV0h1b7htK5LTLTicQ5o+rfRDIDK19W6qcwuVOcIz1PssstpOsWZMUPrM5pW5V7co4pU/eDw
xYWwt4S7VvAr5jj8dfeGtd7sjF07J47YqvEax8Xzh47qmIMXMAxKkZs8uTpeu04onC4n9xkhjc6l
Ynng6Qia/NRmHv404XbGyGdWEy1wLsVt2x4JHi6ZgfUgkdOOQjh76lhyo3eXqbHrnTlttP5/s66Q
zO7DD+mqnxEmkejLIcTf3NdyIHPuDVthHkTP5VDdYXwEY/+vyg7YKM9keM3nf8d8wSPKW2q5x9J3
drb6PnI3fhtGbcik2zL6NUX1NMZf9mmQ8FIH+08SKkpkW/25h9J7AFhiVwGBnA6Azxc0Shby2YXN
1sAl6wAzsqwfqtxV989qQi3aD4z6pCKCTbnJgZxEaZ8vYsMHRoSDts7XjQlPt10cxIR0H2eJUWp3
IKq0cG1DdSMnFCmNxiRSL5gzZNpaByBY6CWkyRaWMaIoFuh4/RppmKjULlSLgG96Lwst6SrapFbO
m1VNQD77z3+vH7mlgeC6KAoHq5KYHEctDYHod6T6/ttVc1nVJ8E6uBcRx4bfS5KkHW+2h+o/hwgs
G8y276iRCeKUv1paCV4kPfB9quZ3EuL4x4od74OZoO9UzSd+rj9vME+n+CwupjQWFsgpEv9aXa70
MX3Y0tHqn8e0iazrWMQOeWmALYTvv0gHhz19KBSLc+spaEmUqdHnh8mhyIX0M4wjK//of4BzHQjE
OuLxBJZnj2ZyYyIeS4GhoWGJ0WH6N4HirLvdo+VRWuIyzMFHdcEhz8gVbpGKBRCKjRoSkuRtuf2x
YUHC+GE9CaDI5GGDUleBpgRxR2AGe1ZFz4xbKhCtvrQTHCG9469H8GwtlRMOm4e161Qoj/UlgJx2
f4NcpR8h9ZqnNcjKC5iy0/JtUuZz1rU4mT4zS9EiXl/mZEDUHk+ZLWO3z/nq3fQ8HaPYIec9o33g
n8jPk6iSc0BvBHdwpYfF2Qob6jC7KCGK/eKBtyK2qhqbKJT1clAMeUgEkdRyJI5BI1QHehU/MRX2
neYkEJN4ET7Nzq0+rEjkouImBtZ3NtbynDr3G4xZ2HBGaDcJg6iebs5SOiV/CBZ9T48a3ZQjIZMv
c/WWQVGmoHKGkOwVutcJS0HlL/glWjetuPHWFXHZlPdk2xZ3+UlIpEmU5f+0BkUZo3H3blXpr//G
SV58eHgEGFNy8l9KDYbLWdgf0/r9B9OodIvsTgwRKKEOmcBO2kSw46xFAn5FymJZqFxV8yaqip+3
9luPtzikhPkcrf1RJBbCDE28sQLrSkYcTWGV7qaYetkYvYQNGnj8D+KMm7+WY/D4d+0xNA2RySrY
iX3Y6m/6EboKiGg10XpzVmg2zxhwvGSYaUguUD8fJfEsYeqJ9fyOBeWkaS6wKXdUAB83hxErbULW
3jmbRbbl7ZJduvXuVOGsaOPiy5uOsj3R+2zJdDmgzWHtcrLeG0xNKys5qqrNWk3tPMD+3LgJeLzR
Xb7N9nOZvHmjp/etEGU9aWchQlohmeG/C4qFfHWJIVbBcXVya6Ni31maG6wpAQupD9qKv1PINoWI
1weuScM4LwzfsmDj9BfjHH6PbWRuZyfC0Yj13qoSU+oJ1gB6x97meIk0hYqYqu+LIst6z7bgtk8p
LS+k3M2S+gB0QEr3o0E5AfJPQcpRooEWr/H4f31O6v1ew/DZ6hrNO+I9h4tFRwTjR0j590TAJrf6
f4L1YTvoD14qDunjYxTN2LZYdj+XnLU6NZd7slrMzTArc/l3frDB3GWBkfJAY64DQaAvS2MVpbsN
xaEcod8przIGizaLJez4r1Ch2piGxvncdVINj8x7v7v4i5OMJj6Buws1i39sZEHw5SX6v2c9CbnO
B4xL0M+5AsYKb702Y715OGfJdrcG+GgCc0sY7i9EJsj7Tm2NDeKGl8rMO4/khW6/4v7OooIH1afk
C1DBx492CP2XTw+8ns+F33DlXSnvHqVkZ16Ow/3c1gHerEgeFk49bd+4k4nITcw/Bfk8QEjAKPPT
nkSZIu/ArTBHlVABgdcpU1Ez9vOsfbriAafAAyrYEp1PbpQaB4ILTGbI79G1iX/z6Vi+UdmDL5Ce
lKB8PJyBdPCc2k1H/IotJ3D7telyDNceUoTm/jqH5kOwpAUWE3E255DgCPe/JfI71psfmA/nX1mJ
OQ2SEdPZjrKyASTDAzJl3cxBjNOS1U4PF2JlcqJXDbVTC+B9UpuPXr8Mo78RaJU4Z28F7wC15cmi
qoatjmiYyFVB4DeyTg2dlfo//OvHRW3oH5GIcH22RfWsVv+OV7Z4rh7Y+ysBn5KAOi6Zre4nMPig
CkuZpkD4LoYWfIZU89LLIAVMu73MsjDO2auPB+HPbgB2Eqou1qG0iHe487P+/d/blyoL0FTFiigG
GtHt2NipW1NIXTQxCiEHq3C2lidyInMALyM4pUb+tRB9YqVMEK0vyiIMsWy2P4GHPPOe3Q942rpQ
irEP1kVTHDqfgeXlRUnlxZIsTbxONtXTRePBoxcZnrbnqNCu0fp1CwAgJVyph2lbDR3KRvdrZviy
3YUFbP89NrEaQ/U1OdE7URK9E9tXl6mDwVR7gCDKiTgJgC1oNOEJK7zrARLqnbNGy3rrUERKrL04
jbUBLS/uUI73bMM80G+l837hI0XXlOQDC7yi2SZ6wHuQxoTKuLQQIENSjIOoBgSHMC8t+1mqA9P2
HvEyxop6MDcv4DnkWfLyFCGendwKxXt8IDL3w18Stcx3ZQYXCD3PMRnuo5e+XN18RHfZiLNENcqc
DTyGQ2XIHGsbW/oaRkaS5U03BC86NlSK2D69l4009zwXbTYLnT/Ovj7tIfAXWcGDDsT5JDx2sh7z
dFN4hZBxl73uYsMTnZv0dAkej/cEIucHrU1204Q0ur5vDf76uxp8Y9r32OFWGAQEyA4Ir9RW2bvw
DxE1p16Xx8nHCdUcw1Twhx21VejAVsTSJfP++z7vMUre7wx9TV2CLrCXWvaTJKv5H+w6fFesyphF
c5p0CbeQ+xIi95lZdaCzSmzbyi9/WsEC/9y8zsZRBngtc4i35QvdZJ0dvKuJ/fuvex8/X24fXp9c
xdmSBaoLiEPYTexeKclEEhuFNEuUUJwokQFPXVfVHO1lIYrhme+JuWD6enXiMosgGcVokJQZ3kmJ
9ismzvR14QugnDykCmw7q97tTG7IyeTR4Qqw9RV5gZNj/s/EIdrLlCljFfuO52CH31f5pV1zL+pT
dGO+pDO15a+zSouEEFR8oZ1QDo7ms7azQG/e8JTyK6kIrt07A8HYByTC5U9+WnbphgCE+BFAoDSd
Y0ttOFiC4pIsZCZz+y8FtEKOmszSsuv2MM5VVm55mOh+cKhn3yjXj/I0teNjx8CNiULEKnG2yHYW
tcXo1gsP2VdiDGF9pGnSSGb9JW+jOH66jivOY3LmpKjDGlEoDAp2gebsmgmwF5hIt6jiDWqpcPhf
MJQlgYJnP8tGsow9vvSyoC73sqcIWJRlmQ6Y/ZMTsReLhF8akF9wYeYS+RdHg947WIwhg/1+H3WN
/ULmgPprZD9BP1UNCN6mfU80Bix6Oi2LKfqN5z52LW2Y+tMRXDgY357TjIoMzw+m1ej30+bP8HXN
po9d0/lfVXwNoTuvF6dVtbgs6Aavm9AqYby/xd44qadMYfSFOUItDwN+2AfcY+1sJ7Xm40VwLqwt
lq2TrhbulaJaVGtHOJ1cONj1ImUWsopHfoUwfRobPZh8ImpsDc2mHWQVFOuASYGvSNolAAE9RiYV
lfY7UxK+MNu60PwGej6KjPZyIPU57L3FYr3QGp5PE4gX+9wvY+BtpSyUwA2ErhLD2HtWER3656je
24O5SIYrhfmCY4MIGhDdBEHB8OYZ6BRGZIJn2y3ik/3aKMexzxHQS12epq5ixPUcHW9PVzL8JPkG
HI1krYrvWqW8NqGLqQM81guk06X6WWO8Uq6Boza0kS7A/iM7qJAZK56STl64q1QLTwIXuC/c222P
6bRaL/o2bB5YFZlwmZuSA0BRu1QyvCLgQfaWxnBF/TfiEsSobs6+GZe5JsTSysEdcR/KyrEGURsC
OJjFd2z8KFaZLnEN1c+AgzFM/jlNmumb/yDNgwAdp4ZciHRupxsSZ8dFt6AqA5P7pDuoINGynCEZ
BfFbnSxXN9fJDdnfR2wyOhNCv78PEZLDjPrxymc1zrZwnlPwh/8gS/7UTwQ0/16eJUbCadCIPpin
A3JpTmSaO0BwVoWNnHcF5WoM2Un7942s9gQIEAdeiSec5o78rBqfvOByzv1/jwT8KWvfTj81zX5S
ZYqcHZeCFUs+6PUvFDCd+Y50ZlCzkhEaWUQHgoV7FzXpglIl0maqojLbejdcc6GNn0xq9zRbkDlX
uYo5jfL+pvHufrtPEvYSx/0Qb5kNYRBxYy2wIk9QPRl1OExzKyGi/bKAVStNMpPXj+tiIeN+TqVG
vL+Bylc9qlbKuKN/S/J4h72QaeZ3FJMQKxuTSR7xXZNkHncbWnNR02Jt7kwqCNH2k9gH+p1xqWLQ
omuzNvtRXpIlOSFKL/r/wdLfiTyk0scsICUtLzVu+rg63V0o0cxwqIAylBwlpzINVYpBXloxFT2p
qKc42KA+29bTCrVfEQYHwntV1H6FPx+ybtU8bFWEdbhNhnsoxqfQTlwDrLpBFpA/LaaqE2GlFvBL
OK2HWwS7DYgZNqLJlXRGocGrP60mep7DZoyD1JwtcrILOzt13oc3AyrGJ06gQHqPRW+WkXnPtP2Y
QozFLzSKaYdqDpMBeyjlu3EogaL5guX64rYSaRPDBymbIXlhNrXDDwWyz8pWvxx8iTB31Kh3JkKM
33Lfq4RAAuttdEr4wqlPDe+d8rrpFmpMsoT5jVDn9kyY6fnzmZjPH5vi3T6294PxllwOhxaxJIrs
7mDBaCBtmGaHzw6U3/8NplaNz16u1yrPP9iwWqp1N/FmM2d65HnRkOCu2ZL/jJG4/43LWXsBObMe
7lk45caK92pQPzUB9ztcVe4zwHrZ775jp1AS7wdHQiTHYqwqNlF61mlT4eV84UkhxlEt5iWi2qVl
dP4My+6+O4od64INFMQCo2BnvDzzX/6mruhqtn3dpWghZZPvN+oFMAZ/lI0+TH7m8A/De6ORVMLJ
Vc7EkrW/k68oxkPcr9eapX8JgYnMii+z/xQkcCqPfhSg5ZJYDlX81mvq3V1x9QXSOvlszkFsXHWB
b9Rk/oDFNJ0FWN8oHz5ZBDPNfHVH4fRLBHIkmrsf1NkYPFV20NJnVtvrqvQQPBh20FU7zE9J4L7C
Mj/P4phnjnXcbCrqpyVOwyXUuKABSmcT7iSStteVYmy6JCCyG+X0/LQAYdmNFLJd1P4ZtM6fvf1f
bW4gAQD+JuXevqzCqgL7FyDTFTbtExsi1PgaDdVymx72ei2I9lo7rbuGhusVu3mM7lDTo3BCTaps
KcZ/zlng2p87P7BAjC9GfPnCgccdpmdMdJ3vuvE6nB05oa8IzIBPml+xfO6SU12Fs3/bLn/qXog4
4/t0KS3wS8GO/lW4krVh6fHUiwQ+3oBW+/QF393Pc1NKOMG1TU6z3dqB2SLyb/ZEIi0fNKZSFcKh
DDpYpfOXhrZfr718cbRUlGk+GPMi3jx74Uj1Z7qsrr0YGXhqGrGPFkZWgPaBAvjnhGVVkrYplGpS
qGlcA9abAztJMzHgNyvFPqzzVmSf20mQKXro46owmVUEHIpcOrBffmGetEvdDm8T2HGSvdx8ihqM
vdx3qL3/8GyIhtsXGGCvpz2dCP1RV/gS/8dUmjiHH6CuLnQrVnaQawrkDiWKxDQn4KF5VbYd9avk
r4PtMLBYxVccNZlogfaZkG1531pAz2dHNC6w/05iLsxFil+fcmlkUsuOXieKmAPdasorzFdc3eRU
Ro0R+ssQLRlFEjjis+uxQk/A9RHze5RWP6wn5xHujELPPn2qFCUCBPiFEXzLmHd4ewuR8yiKkniG
wOVhNRHsZ2mlHGv39CykD0UoN9tXn5Seshjmc66jkc8H5FBW+WrStdcN8RVyZNE8hHZOGMHYqW7f
gsn4fueZ2sf3QrJThgxj3g90lNch4GfKvStqUD+170ryB1pvbu57uDMEF/IqGyVScof91vaGWiuw
bNsM9dnPaYodRLk7RLuJPUjE37FlQrbpqGWxDtO90+BcoUUHm4+BwmZpTQtwlC7MkJKoMjIFzexQ
PLoyGF7yXidZnKgRlR2YXbSoUyWHuAij81T7/mfF6lGbBTPZ7B2Wu410XUR8TSvfdPuyGvqW1NsS
GrqZQydaQhvMOREWMMCi6E812gdTcPw0YfAYEeN0jabBrhN08ym23MyLH0oT54o0xeu7WZjyLS64
voeHEWgTYP4r+Wwt3Nc8FY/6nyTPRd1cHzryLKMCze0WF284SA0tIQZ0zfUV5/OhCtLtZeVeXABJ
TVqX+U3MoECE0PArLEvLvWhMEX6YgYqAFkCaBKfzNHzCU4feEnGOgVt+LcEdgZ1B2UzSQYr1AG8c
1ro5prkCWwlWa1Jnf3VyosOmtcqhxPrE+TFv5kofeySUs54TCoRWQvoRjYfgVM4pVLkS2d2wwddJ
g0lUY7BNHcyt4HiUTxyrIF4F+g0pEM60yzFzzqqEnJzkSEWpZDRtpY4fypVPq0Lp+3bkzQUORLVB
r2vXFW5d0a0xd8PQMrP88RnuhN9LoLiIiwo0O2BwueyhCSBpTgfLipRAW+EvBHPnMplJaACZCCFG
o1wDKbowXvH6lXCA6vdRV9D0ABfurmls7L7FbbLrFXQA1weferSuMXAXHiFTse9uBy59i82SmIRF
/Nq58XjKBQKd357eAx2uIv2gvgq/N5OlrRiPj9YsgNhu7mdOqZEHXkjL9nBLkRDwS7Y5OUgh/1FV
oGhdxCOnjZlm1dzeyyCoUZitWEEW8Fn01rbSQKCoNnPjaZDja4XtMu60C0S6VQqWhhMI5xlGPH3E
+1BXa18123A7+raqJd5j6ovTAt1BRHAfKyBeB8ZYjBO8lMbUz3F1EOhY8zieBCGEe5I1P61zpTwA
OXeSmNhQ8j2ZsIvwHJQPlIKK1B+YmBQ8ULzKvAP7bQlxeV99Z7gllDN/wnakZ/7jsHnxPE86MYxg
J0ovFOAfOlC73geqte1QbSA2do1x8iwAT85t5IwGllfftJjgYSjEqnn7QsxQXJudjC1vCnA8PNTt
G7AwZst0ODKg61DV9PWCq655XCWVHYSNbZmtNwmy5mu22OPnZ65vh3TlxQv531joIAfrsvYALvR2
1AAOLR4FWgIsslIu6UVu+WBXiJNKqWmXm7g6ABi6g5Z9ECihvXrbFwECyjvJJZenNwheBHhTNf1E
wEvRCgo7fje4whGr5F31odL1vJ2jWqd+wKj8tvy4H9/zszzmb7k1y2/QHkfwYijXDriq8zWr66qY
x6Bf1wcPTzEMTrIqw4eNEBZQJgW25WQtx1zjXMSD82rCJfuxBlWiLR3avYYE2dKp2OQ+0f8sSNDn
jHsqA9r/rM/wDXJCR5eAd3fXgWu6G/L09r4SGVIQ9iZSLvTEGoYBSJiCKDdqxqqaPgOueeSzHeOI
lDD2hhxnf0+/YnJEEeU8jvF3dvL0nKHj+zAHcXWRdVFzWZEmo+p4oC2FKTNL9uCGMGdRWGMY7uBn
Eub3BXPwkHzatfTlR9xA4RGdk8+BPZTotq++GaC1vFfLVqf9ylE2ogPsnIRw4wsu5cvWzCBP5h9s
Gxqa4wl0cWmz4vWVegY0OOh2BQowtehg9ZBgYAADKJ6/+MkUpsToUvv1yvErEO9+G+x53YDHonHV
z+x4qP4GdnSO3TtDUksCR4/N86OAnVyoOA3Xaync4coZCdlgXXkQo4xsy25Yx0UUY/65bLWUBLB0
wdlEl0Mvo8RcvDeVOh+EF0BOgKPc0b+kaHVENfT2T7gZihDAl+VvPbLHdZrjfN8kDAWZOX4nUbOr
+dVzwq0jA1T2v6Igdof3x+sMQIA0X0Br4z8toR84wXSfZ+5fLj1zigP4F4FIoLGhATdPc8YuTCrX
tszbvJ6ipeebaaqL7v4SQGhSKEZDa7ZpEnHrqOk17E0E+HLBU5B7veu+o4GmNpVglpck0QxDjjgI
q2p+0U8ecoDhS0SakkWiMarMUCsACf3g0rW2BVzCM4TC8pFJbSaapHc1PxVwEyZvUl7afTDys9kr
Ntjw+Ok5OJuPp74/kGNodRBxx+ekt6/cL37rLXKLcR6ARB5XQ8PD8mzcDbJ090AKgmxJgixuRXnM
Qy8INAeuB/MT/836Ax3OIUgLvZaZdRSR+yTQ9ph6n2k58HLwi2TJldurQe35bNpibHw6fvPqPVGe
UbODtGtizAz5IMygUt2WCGS2OLlsMbf4MqY6agGgVMk/a+fJymwxUiDeuwVOsMokAAZBQezsQYX+
DcMyxaRi6ZnT2z/T3rcNABKr6XLguY8neG7ymeSRylDQkebOGokvWn5cgIEEIuv3DCcCiLv+NPIi
oVJcdhDlTLSptFfTalXYa7xXexrtihaWlIc/GQ6MgZcZC0Nfou4aKljxkdd58Q744XHQKX9Qp1ng
sOB/nN2lVxWNXnyy3/5NDzap0Iha/ZzUTeBqGqHxH+EGsn1UFZKDYj5VZf+ipHNXjdiqM/PVOahL
xAxU6Wu5FITQuiR6qBcGyG/Yx/ol3Rb1UiCgivGMml1jSRfz69q3W16udWF/C5dKB7VLiWi5IN9Q
zrbFr7+zxbwqLjlJA1GglJL+EX9hbgySTs2T5WTFKwGBgbeNt6qExuEQLN9KSNe4OUZs5dvFgsDE
MPX8RluwaLFz0LBsBGgYQSQpsgJwr+Ep1Yz8CxEYBjBmKXYUeeCa7lj3MPa6B+O4FFXhM3HGRONi
WRvZGKx3HYcGrybog5Z2C6LD2H0xQbuIxivkp3ot4jKsx8tWkwQwc+FjqMTA8Iwu88jK4YjD0ngD
Ds0bgXpypemr+HkcB8Kw8gPQzX7N5ZTBHTVFPiDZ6bi8lOTUT5hzu8hZjD5dAxIR8uB62uS5yBwb
7eCa7hUj3VLBTkZKE2t9QLP1AKtXkQi6DpF5YxhHv6Jm/Rbu4jCy2L1/uqRr9hvI7+XMhIfh3cVg
xdMnKmClZvpXDhZGeurZ7kL63xH/Iihwv0G0MvjjJR1CYqBV35j6h0VmiuoicYl2/p9uaVxJiszk
91mwY1opc1p65eN4Lg96Qrlv1MsIe42i/2mVXd2o4RB2/GIN9OjMRe+g7Vco0ywr0sfQ0S6hckf2
L7DZpy1hfTr7QJn+kB+bqlxuGt0VLuEBzMsvQubVICdlQJd4hjzn6x/ttXFkBfZFUCKnhy6EwGFb
1yqJI0RNqLjgaXXA5mbUsuNgWHu3zZG2HCCKo0t1M2LaaVRuPQ1ew9ZAAE80te/wsH3mN9YZspxC
CYqS1IrSs5vJbzSV9nZKb1+UCCLAFYIYIIWqD889I3c2j/HRFET0GrtjvAQi2b+7R5/Vyrm1mp4Y
E/pOq7/Qm2RXi5tHGc3u2moY62s6L8ullEpr5MkC4OSIBZPM0xu/9NnkKrB18y3pPJK0r+UcDtq0
t0+ByIijyov/IWsnFNtxY+T7wNJDG5YQ6jB2YImMTKr+tCEz8dafMqK+ry6sJ+kGWADf7/OPUr4y
UvwEVeKJdPtEA3nzNuVwJNS0QwjxvdxTHCpCECUGKtoVOiwIuGRbSRHk96I6htHAhdjzcLuA4hbq
Wj/zcksoFvbVP+7zuhPqPi3EVCv3gsxFVsuW1Q0OP9KklweiAhxZSehDLd3kFn57zzXRWV3r3rSa
8uktEwm7qOPuUilBrFZFoxIOz4z/dn6EhHeyM/jnZZKgyE9mSvaqu8Jy9Fmy98PhVvJ0HpwWy/Y/
YucSJGufUCLyFjTz7T4u/2Hn8EWy6LXfeL7UMg+cxgd58sdrHypljQHpl7E3bs2jV5pX6X7J0bhp
J9FObSGZbHEPesb6LTBPX3cFd/Wk4x45LW4Js4KEHrRqROO3PiKc4rlWm+f1FetLpTSJa21sPq32
rKMCYQa1127dJLdEz7VIGVKzuOHQVjE28BxW1y8suD18/62m0w5yxUG8Mt1TRs00MVK/VeIawPDp
f2v8G4B26Byzuvkuq/xBxozh/DSkly9/iQDL8t4k+msvZ8oowd+562FX+10jZ78w7Woc8CHarHOJ
UIRzru2LWLltZQPsMkwjiv+8aaBYg/izaw0q07kNH01c7Fmf/Xw3ZkjTPUKHUqbHrG8DU/b1ly/s
gjrn/g70YgF9NBwSv/PSc9RMpT+Mr7we/J7IjXX6ovJFI4OE/086ezf00oT8bvA3arap8oRGt8ry
NYUn+5lnmKwH5qrT2+/2pMkRCgyogMB/XLK/hDCd4QTUR+lw8zxId86wnjwKDouIPBCoOejECE4J
CNOq0dDLnZFH+znXzTIpJKKgfZcKCU+gKYSZqebx2FISYVqpyyqW5M1cRP719V+l+IZcR0PDDJ0F
RMhyDf25Vrla/LyQjmsPUS+rdIxArCaP4znuSgxpp8MWg2KLfaRvXi+HRvfOJr0UOTW8fzG0s6mO
kJ0VpkbZ6+kmtcyiB8VpaOoTO4705Q+7KtPxfB7XhBmszd1H6NuoAK8XV6IEqztkk73HvY+EUVNq
6x64HZsvbGgWDVHdmKTdvxEsKcmneF9Gkdwh3BqIaexxQ0kzflCJrZ9U5uW49HcSC2VfS+NrV5ky
EY/usL2kf3WjZplRgQwrgEkbXOWbGR5Fn9QPvUdYbTVcosx9Ic8caHiy22UgqwioJPHCAIS8JIbM
7UAaNWjIncnfcy3dAoUrSFC1PCiL8wTlcB4/qNkyxIblHDfT0oMU/yfLjTEZhcLoXOQFgMjIQn4=
`protect end_protected
