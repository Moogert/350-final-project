��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅRۥ����A��I��jٯ�S�s�,<BD�2oZ�)����Ȭ"����[�n2P3v8i؊bv�:�4���p��^p^W�Ga�8?OH;S�v���������Ǚ�5XE�$�'<�y��Epb��z�^���d*�`�6������r�D� |�.@��%]�9<�W��v5�yP<6ZHa�
��� ��e�K}��q��h9(J�G}6���O�<B�����W��F/��N`v<#wに�gNq5!"�SI�mF�75:�z��&�-�P��ͻOR�_�N�������:|�<��"���}��	��9Ra�;�Ԟᜠ�5JtO���K�T��,u}�:QR��?̸��{�ݯ&Ħ: ��أ���w��W�k�
��տ |����׿����Wi|R�drҎ��z��!��t���z�i�Owd�t&a�0D-�词��(��"��VH^mWR�	�AB�=�9k�]j�fv��^����BC �������ϯ�&8H�2�����P$������!v��.sf� ��A��|_H��P��As�n�P�s��9:�!yK㠆�Dv&$jF�pt�m��x�4w��6Y�Hod6��A�,J��;"P��m�Hl������ۚ=�|y]����KQ*p���Lgf�ӧ��!f!u�1�w��M��cdF��ܙ�FE��`ޗ�x_���{)����a-b����]��Qm����v-�e�;?�|�ҒJھ���q�_qp�A�j[i1�;��e�$(��S$�tt�S�;�ǅW�u��_�)��X�`�*�|���#�IQ��g����:��{��2��D���P��i;�P8y����ΐğ�?��"�>��Ld*z�j@��\]��'�R�q����4�!
�E�XY�`T���ߩ��PX&yN��!�%��`���,-0���M���81X�FF�w;n
0�a�dF/���I�=n�}
S�xs8��8eu`���>1-:;���7��R��mgjl�����U�ڜJ�����E%s�>�g"��B���'wKy�-����v��Ĳq:�!BN'��'�W*	�,�J���#�`<b�^��ph���S����uîg���ɵ;(��cE�ܼ��<���(ٷ�	mS����]����ǫ�Z��r'��(������*�U���/�`�r����7jMF��5FIC�Y*����g�-��m&4m~W(��f�0�O���!Hd'1ފ/���7,��:��~tn& �.֢�E�wP�p�����>��xZJ�F>!|���Cc��9����IZ/�����
�f�³�*��*��6��t��NM
/�a?��L�i?cɛ�s���g
�M��
1��'�����5��8�LH�>���[z(a,���%86��y�^��Kq�\��P@s�G2�pO큛35�n��B�XJI|�;UJ%��}!������6����s��� b��<R\R�WI0|�,8���y.��uZ�ق>\0灤����ʽ�k$��!�n�/��bFd��zܾ&|x����W�w���N��P��̯	�I�c����Ԃ����w�Ϻ\���{;$Dj���cMzI��h&~�#<��w<���	�.r�8^[ӕ�7<�z]��Rـ8��g�s��z3�m݃V���)��&��Ӌw�2�B�Q.S���,z˅K�����ˏ��-x��+:ş�ϻ�v���� ta��ɲ�#ZK���oQ<��$�]1����L����C�so��;E1�A��,��t��}	}9�\�Ǚ�b�g��f��X/�*z,��񢤿Q_M��7���G6���o�z(�bCпq�G�
*���0�_���27�Y+�\�����RaW��a1�|b*K���֣f�0l��s0��w���g}�@ɨ�Y���7A|)ߎFpl�%t�J�+j?y^��e�Q���v�����mB8*��d*M뚪�rT�,���(���(�.9�R�r�? o���*�͸Y��	�fO�񂎐j�S��/3�������G�F���"e*q����e�Fi����+���+	ʰ��0BAo+��<�Y%�UH��+���;��_�0�/��i%\HXǛ5�l�Y)??V̴f�ol�����ƞ��z�%���	)~�RͲx�P�����!R�1=?�\\��C�R��.S��7`G؏����K�n���7_�Z'���/��>�V⠔�
rc]���SQt
D�Ը����RG��o��@ѹ0�?�sMM�~�?2�A;ĕ�ȕ�oK2��
��y�B˸nF�����c�(�n��9X3�+MP!l�R��Y��J��?�L�����L�
Ems�"~�E4������,۠��y�:3��E���=߭n��3�ĸjz���<2�L�@vZ���B�)i�y8���v������g8�T�Ra�a0#&��ɀy�\�H�!�f�].ws*�~4��<�7�!�ɵ q������v����1� .˖F�q�a�{O�|�/9�Q\ai�!����M5.bW/+2<����Q�:,F-^g����Յ��%ѽ%�f"�G�#���#�y���x�Ot�'� ǯ�%5i��W
e��ޤH�F��7IHKF;4]b	��4�����(7B�y�����,6�'xl��+��O{�|�Ԉ��̨�L��ż�	�I�M�W��\�G�����{d�M�\�OHwNor���w+Q;@� �%���b3�G���f�����.�j(����\lZF�[�췋8���~��b�l�>U�ƍ{��ڸ�nL �b���VR|mS��."�6w����jZ�Pvl���ˁ�����D�!�%�9�Ipӯ��߈�������p�^B�OA����u�pxOH�כ��N��_Ɠ�YM$�F�i��m=�V��Dt�Ǧ�Mׁ�i�ʂ7�a���G6%	P�_�<�I�6�l͙ ��C"p��"��Wu�֟Ļ����0��an�i_�u��I'Zr,\�xN3�9���23�)�e��Ժ�[p+�m�[*Sb�1��?L�F-�^�S�I�3^lлw���N���\x�ח��o�f�u����~�����VE����Md�fc7Uq°��A�'@Ge�R\`нy�wJ��k��X�ګ�|3���'�_�=���<�jQ i'�(�`a2t���p�F�����o;�Nr!n� �x$��P�����yM���L����d�
��5nc��Y�2��ϩ��sh�I����WJg3�-�Y@�(���f:#A���+�S��jMu_��(2��~!�[�T��m��	�u��+����RP����1�a��B�ڠ��U.gP�Ĵ"�Vw��Oe!��A������߿�W����JڧQ��X2Sއ̮e������\�hy��d���r]�a�;F/��wT���䱾:'����+K2\⢉
�;�5�p�(0\�7s�{�ʹ ������.��!�����AW�]�o��htL��=Y���L�J�%)�u�Ǵ�) ��x��|�[�)P_���Uc�č(V� ������ͧ�<"�F`mz�7<�ʡ��vd)�F����CqtS�������_*3>8�vb'X SX7�ʁv�r��)$��^���Nb/u���_s����cj�N�=�d��Q׎q�QP/~���F	/D�Ӄs,��}��,}ns�\Q�g��r5�����?���t������L�O	}��lgv,-�K�.�4�<�M����y�c�9\�K))�������;�?��8�*�c�����z� �I����B��6���R+}�Q�j��%��p�CT}m��;��uj�$Q��q�DG�Җ�w���� ��T�v��L�x?��|��(x��`+^���|{�U�����P��o�	I�����p@+�4���a�ܸ#����_ܷ�j�:mG�*��2J�0n����sP��O��l� ��6 Mj"{<Iar�Dl�J��l1�7r� �P'��dS���Q	��ܥ�bE���E�5e��z�1)~�⇷Z�"�MD��ǵ.լڸ)!qdc��!�eD}mx�H���K�BB�M}yǐx�&��i	�$O�"���zC�0��X�܂�ƫk�g�E+B��)k7ÿ?����l��'��jS�9�%k