-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CLGdGqgROXwJsOtj/ZZwMTeZ2vi4w7uFO8Y0i+zIr/iq/+w/2ClTxVwz6ns6NqiAmEE3Q8fDGE6k
oCbHE4wf+3AfWfkWM1l9nCk0WtGrFkfZ3FcrUXBCJF11pg6zMT2Tjk+zdHPk818su9379O5mGZlH
EfzZXwN04zhd8KzxEGS/Sk4XtudRqA1e7iFqFZDTmgIghuFthvT9V4Py1mPvKytmI57qJfJNeNad
mcXM5/CzAF2UWGEHlaewHorJVT0qeC+FNL+ldwCqce8gZI/4cvlIHMmeV8dv8DM9TztHMGxsPQ9G
6nBi+NYofdIkLc07wUL6SjBl0gvIt1VeEMkN5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114416)
`protect data_block
ueGPFyAwnxZmPYhXFaveMRHxe3zIArquj+lJL++BeD0E0le0JY9HMsJrwBpCapHtyTG9wxixOKqM
x4JFJfMVYZjvwmybt8PRQJdzwx8pI1RTsLK9bm7TqVRaV7izqVbJ+oz08dwDLEEmOyjQCaI5LQ/n
zTbW1o5l7105GuX4ExvWzmuLd55MGCr20qFyfXQgeVNYYpqGoBszypOn7uOC0EHT83vidUjUoPGa
vyocJrADedejvdZfQncgtInLHHZdaKFgmEHmbZ0yIPSMcV5/dsS5WHlyCr1kDDXBFTmFfueg6Flu
q+GkBpe0p08hq+WYs7L/egL+dk8OqXN9TWeiIa59KkLLFSGs/vFMH6n7xBxkPzAu+vapDOB/McXE
49xPgD8DyVCSTIh2r3igetk7bU4DT5o92ItXSaSjy4qxa44FNmqWKzlPEmqrhT/oM5GPG9Omb1pR
y0RcEwaEHyfJ1LwDDOESo9k0rN3IN1eZHAuxKHJ6CqMZeleYGB9eruwKF7xepa8i0sHv3pg0WKtD
xhaBz3t4DPDgzqCTtMbylnMIkgxFrnjeLnK/ISDGbt+TR/eHT3/8HXHIzu5U+aMpVkMNySRft8Mx
wKZUbNRJ4l3j4yoHiOetnSDT8aKvbRKaxv3R7YC646vabn57mkrcAPFN4RKvvJ9Ajs77rSnDAaFA
bh7++/0Z7Gy7yPz1tOnICAt8mYrX8UwXqYQGtk9jDMFpFNQCIriFQYfvfmRV9kmzokHL+yO1dL5L
EoAk2JIC3Av/hXEQP+itU6NpK011bKoCZdSUMNFV+F69UtALAK4i45BeY5SAa6Vsb2jDTBbO01W1
7OulLeA33YIzn3YbxjVWrDNtqYHdnrQiVMQNBpXX3PmPWzU7xmnEWCRdiRIwO/HhcfoetCiXx00P
AP71yIqapt29vwJoDC9wru2vR20DNDxWDPV6Vv20uV5YsEjo4p914YZ5VdWvU6/AioDkwdTM3fvz
KHsyMAkuGGuf/Zn1dJjNIztKHn5Lx37u2NY4q0YsZFC+JkcLWTcWXnVW7x+6cu/zDUVje4Wxczcj
pmD7klchxEqvigjZL8da1ZGJhwYb1l6ef3vthCbyhD1f8E8AE/KmLJxIhJRjzVXzGzZa9wQD6svo
EAm0aMCJ9gzVXejg1uW/14pPPGdsM3+z+lPiTSDxQjnxl+yK0kV7/tNh0npHeRMRdy/fhCpaDmHO
bwpm2GKqLSahzQ7gCSKfzhhmC8U3stK78sLNxS3xpDyNMj9kB3jR7ee/EcHbB6HgaMVyHGUVg4rP
oGbER9jU0quvqBfI2Hm9kcFbmzGcIYzAQQxHmCUF5FHQ9bPCqDDieWf+wTdF69b0bJpgYVSuKQXi
qhZEvIZy6dmAgo9Wc8meJ3OO288WmEJC93/eiNLNj29k3xhXPHtV4HjCPjdeErDJyUN27zzGka/X
VdHE0A2U1Rk7WIMV3WrfKWSjfMy7yYC+WXeitkg7iBcdBY2qT72cZoZ9SW7w0zulVI8piPa8clfQ
r7oUr1en2chXRJpyCUTDl8mIWoL8n8pUWNziasNokuoY3GST8dtRvvJH9oqEDGTWpYeHQWXcr4fZ
QQ+pTQS0UBoHaXSL/b5s5K9NJR9+pPO0rEri6uoFI5BvyMCqMTb5OxT7Fkt5dnxDd8KZSNeVIVAQ
/2YAXy/O+1dnyL4lf7qQ5zD5twSfb3ziQLhxwGIRRP/9AO/DJumR4yPV978RTJTrQ9cbdItkI1fT
jiKwiw0h6otRoWZXSlbqiHexSfFj47gN766ADCrjPuRk8Z96Xgm4YvH/v4JpA8ysecVaCOYElPhG
U18GU2ukKl23JiCQ0pxmGMNFTSQ5V0QDasTPAT+6+nPEheQ8z3ZJybNmvatpTmGmvxPeFV7bbCVF
1aRfMV6gVd8Y5MbSwaZbGZNur5SyRswCoXTAa+g+6nkbxyWE3/FH/GpxldMxjXtuPw6IbXuDqymw
3BLwsA527xnczsERAObp9UPqYHw9SgXMuJBqPXZ223gKvtH7i3cSGxPPlsBGVhXVaPln4mNPI5/C
2LX5FLCxpxFz6o7tyvIG/osYfrevid6JacnCG9Qgk8Y1gMSmhCLJ2v0QClaCC18T1Yahc6Z22Xct
WaXNCWf2GZ35fwvyBzB0gyNRPYJuBDRXg5UDeidxsidoJahXfCugtY5ThXQfGCnGAgGJhjehl/Nw
pjCqwL9jTd5PAq9mxTuv+yhsMZ72kNuAvnxEsCl3X1FH2BIFj/F6b6Vk5zIvKwb4iibMBynRqdux
BgDO5yKgbhmCVjOuMnRHmL/ZPT5bUgaF295Dbwt4gwWLaGwlocghWsEQyRSvP/xlcjQmxVBE5G7L
4yu1WSLV87sqOMx9cOg8O3qzrkQigup7H0xwd5LZ8yAieH7tRJbdCo8+P95GF9YJRHGPDG1xTyUc
d5ToeE0baBYe5J1SfEfdaUEo2PxavrUANkUgsKjBbq2TMYpWbNEnMPvMMIjJX8QqHEnk9cxMkEnQ
GK3HKezkzRiIVD3sZqrQxTU/6+LspdL2X5lnyRURDa4K6oDDtmAa0dfA5M1ehotHkdrYIZK7lVUa
5ozUiwCi6RUrplW3hzPEekmzyYHU+arBDFIHN5G/ajnZ54bcIgOtywXP5YH2MDP3QCl/5UA/wORs
J1RUhqfPxu52HHuoWglFqpTRNvQ7//vx2bDL134Chj/nE5QCnTLdLDoEWlbJVjrJ2pCYzMgH2K1Y
sEwjK7RqGfOwtIpUrhg5YhR6AO8iQCWD6LwNiQAKRt6lL2z9+wEDkMd73C/hOslBMrOW6nHo1aW5
7sDUf0jCmgNUwGl9z3Tfe7kj0aMz1/eVGB0h/3ctGHSs7opaRnWN9OKFpZM9Nu7mACN/Qkz5MCgP
LDOLsrrVfPzqSbxWICRTWWq9sR86anHy3ppDJHQs/OsDjb6WeQZ0zGiyRWBU2fj4RKq+ayJVz7py
5W9Wj/nc5QuikFCc01hti3RvFUlLiuVHSvtFFS2BAvIYyk7Gq9kAe8vUwZbHq33Nef04sGFNPdH9
ZMG9lwXDoqHPLH3qRn4bj8+FV5fCy2IfiMxD3wfAunTBqOoZ5D5eUdgG3O/fJlwFgKKpUkJB54y6
8BNvcXRNVsGfzVIxa9wQrCnTYTx8NAFD+6Wht7sUC/EH52z+tZErMqBI7MGSC4/8lK+s7KJLKOhQ
ldtv1B1HwM4HoYWuXg4PYKyTh6yCaSjhG/HgaYzPvSg2+1mxA1GogIzXQJi0IMzmAsLBG3++wuiz
Zg2l3jHj7gqZE7or03YaB0F1zQNaVWcRBhMO342P4JEosW2YwJF1hXVlFALi4CtuOyXo/GurdtC1
GpXF9/KH+K82/WojJpajRis5K0PmHds689J7OaUdSyMOcueOejGNi2sNwMktWKQD6BH04jyM4try
3Ng4MjnZFAXFzKY0Q5PNtaVsK76qBQWk0nWNulU6n/yiikjGjMajvO1V0RmGCCDr8sd/34rfFeqo
DYCwadJbMWCNiKmdhc1S1/v6+yKp78tQwb/FKl7Js0loxyp5kF8nvqSyo94H37CkAjXLJWJDa/Ho
mgDLlM13Abrxo2ej80M9vaJbjZfE32lCriTVpM5PpVZf0NZQihykDV1krLbk8xb9FzVqnTTe1/Qb
cH/FtiGl2GxklWMfYdopqP6OvMbZrV/3Mkbpmxj3rn9EQ2MVjRdU6k5sykLJfix1FTBFK+v9gvWp
TpFpSYiVh+Ac8WxKZYx/pI0bkWNpajVWvhytlZpSb9avD+PG4bnWRmf5nHtsIkA3Hz1i84CF1AxX
LpoqazipFf0tH950ctUCLb95YVLNyLW+bgHh33EM86a6pYvUSPTU0+u4E3BaLvtKv2LnK9Xn/g2H
qBQwuFupi5vnDVvWosV1pLnkfdCfcgWSAdhrKGA3LkX1TnD2fA3RGTE5ZGGyA7DKtXt53jmpgEms
9CQ9neayJmrSaj20CwXUOTIOqjG/SVcWUTwUrvxOTJjESN1yyl8eTfkdiS6DGFWHGq2GwxQF+dfb
sGp0GsGi1PAOPRWTjwZQr9vQSJHRV91qGT0oaJrzfwCWJdNAb/u3F29hy6noBlG5L5tojeL9W6WB
u0Lhlk3296Y7zOCA2SkCYGOyZFEyDOP6DOBZDnw4Mqe13E11lwbWveABpmxsjd5QvLJ6Y2KT1lvQ
iMG4E/hmCVf4nuGnPKWWZ1br+2K3Vrx6jRH9uEeplJz8hMES3OE6NsMpQAIUSnkCLrwCW3oG2R9r
XgIbpoSh06pZv/ZWz3ZB6a01m1F89g810CZ82mklf/SiLjIfTX5QglveHlfDGo9JUJNuthXwZ8ko
YAtOkcA83o9BDfwxZwAHxFnwygLcBFkVoK9ddmPDejns/g+LbCrkEzag2xvUiCckF6w2XkDx3Z1c
0/VEpzisMk3z1vNQbaBlKQWu3lKhGkbjCvUm34+3HvgnySW0lzF02DDhzGTZRBu8B1TlHARlrnrU
+BVTiu7KKKwgVjk9o8znNAMLVhH8PVpQ6kPVbN9f7G5d14OX+ddBv1Zubf+bRE4AadZN6K8Q+xXB
Pu6JlUuWZrJznfkPwYfV5aqskGGWITowMMaebgClN542rYj6aJkMo+udMDyfg+DBMBpxC+VmjDcQ
akbgPH/utNYCSF2Tj32b/Rp7jFvhuiNc9PTPT6b2RA55ezKLqrTM/HaVIQvJU90bny1eN72Gcut4
m+aYgUaAwnGx/UHb/BFGmPi52qVXrlAvJNzpcNjMmZW7LVVF5RuaA/zzlAQXHaW6p1IF92savOM1
gkUnG5HsJ9qrIsDA1gUtlLOHixKC936w/zbkRmKiI1ehGlONLa7CPoQ3BijuADYumhXXuAnOrRJW
TLfXNZD+NTZx9qOe+ILRQNDnw3sL1i0aHQ15lUUouXsOs9121EbrVSTZRPjRNoPu89p/3cnz/9FR
J9X709hzfvGQIF3gA4ozE4f3eZJxIDh+S8u8hNsM7NDdMFr96LZhQLwwopCHUKL5c+AVcCxIYhN4
tEi3JAURsP8Y6Hsz10QjTRnF5A6c+brf+YLAHegs6MTXldIOY/tyJoiilW6V685O+6EFdoFzwcTK
l6UuD4oqO2Nxr3f9/sEeww43cN/R5L/lX6ecV31WuW8Qf+jOYcoVtSghkQUOxLZ+IlhMQvqOhMP2
bQsBUEnd5G0LY4ua41fhM8SU4+RkVW4N3Zpcs9rqNXvzonsin8ZWjvwfmszaqiYwMdxqgb9gam5U
41oWJzBuV3GcccuoxlyilfAaBl1oxIiH9oaqAE35BIYbTSvkNetOGlPeFHAQxJQmRRd8wAcnJwEu
vx6UY7AVpTRKhXjMmLUW1uw9ZHrk0i38Gh88A3t3SkF1D0mOIZkfWTWXvv0K+CN1NwQs74ciH5+s
lkujq0Fj0vFX5Y1A2Vrd4rR7T6HPnOzjknYkQVz0MF2iUADe0DadcAHFSSuvTMf35vSaWMp56cPG
X4r/tVtWH7SY7WT6tO6h5HSjv01WWVMpqFy4RslRnZ/UI6Q5kHu2S/dMFFNDNTdIESJMFhNPfUb9
/bhtUTZV5EDg6JTjviabyJ1UElKPSWRFL39KoMpXCEIeYlpi/Fdv4/Q0fm8KRcV8GDr4STT38XeQ
yUrZdkfEtebpGMUcJzNVQ8t0ZnyKw8ZS2iGGJLI0vVfXfrUQQu8qkz/3C8RQfrZYdRnL8/4ki038
nzoMo4mI0qrlaaNTVEEXMOOOj9Suh3H9NkcGq/BEinEX23iutJQS8PgKudDe57d3BBJJhtDs3DcH
W67Xr+9mhygpXDk+bURcYXRp5cEjCLNJLheEs7GnqZKsfyb1sPOFyRTtna6qSjO/i9SY87en1nzD
DIAXeGIyCZJZ6vqmgt6eVvR+2gaEVBTPowZsNqF0mPZcMqBlQTs+z1D6FuE+2o9x6QafWE9yPRm1
3OExJMOYdGD8GlYhd72lipP2nvERWmnN5LmFOjfTYsy9VPd7bfohxwYO0IC/uRRP/dujWqPk3Aaq
3dKEj7A8a/mv+qjdJy4IEneEhHZNILeRm5QVEavOwlohjt8w5sZkUX/nFos+SEsNSHt0fzm711dH
PPEgay9cOIlA1kl/lPd+b0HkIWvMGrlwNl0dQ/iUH0pNSgv8q8TVdc4q8puqfqxUXJNjhRv0gSPF
qeJjxIkhOIwaictdLCC5RqftBj3tuz80QMmWW5f4mo9m0k+kQieZN8+M5DsE06Yx4NBdwbrKoIJE
UTHLwxlA44uf69GFGPUwyLVRtKTzac2ltW/HITLgz8Ij6uDkkxElwnZ5/LMLe5KMLJCLy3FykXBX
bI1KCH11uBPrDOXxNfrZ4jcU9KvCYrtGr0dCi0J0XPwxkk4ofL+9meybqjlXPhDMwjXuyYrZ+5Kt
4MjSK4g72C2yk4xJnfRAMlI06LAh5E2m1wQtXQsc6ncv4PrhYCBRWiTV6+fIvPumFtdNnSN8wkIE
TyKFMWLEK1PYaJMAu4RlLN1WMayUFe/EhD/PV7LPFrignN6FPaatAve+nDrELayXXE7Syr2IGGPV
0zL0Z3A2hkTKmoA6O/sXHO3pXYzHGT7jX5cA05Hv2tymjE4i9i24p/BmVQrjQz/lrOKjJelpkNIg
4zjyYtX3yVec3pPrpKourRY2plCId8ftL9vTHqq5tTTIDyoQf3fxyzxCy41dPZkp6vVYAcDi2G5x
/bNg9BQlDhMRdpJGRNJQqBnxYG49IUEcaDqXgy/SbtGGst76gBHrJnRjeuX5D+ntomIIykDM3zJE
WWSU57FAl9qmeWGfd/GXf5yY2Lj7w4w1/sfdB3pQQjes7aL8flKKz5N6eJuIhCZXINOEBqHL+4vS
+syJ4vsET6PNtylearSWttKYNwaMGrVHcwbkCTQT4OjRQbn+8YVdvMPkzG8U72anOgFJHKGXezLd
j2msYia5RB8jc3qGz9Fy6YRYKPr3Aps6j6ih+Lx+5UEN6R4TGSKW17J0demIiIC94rKYLD7azo38
MS7lLUPY6ba/EOS2WF2jZm5bHZW0eL5w9a1KXe+XsuFVJfuXHg/+oYPkLVDHz2s4r7v5QxutGD5S
Wtjl+pXqS+HLeGcW1EbdJqP/mA1yMIJA3AZd8vmJ71uhZbd4aTvYzchlJR9LI++WStQLDhc9LEur
/UTEXqslPsMi+HbXVBe7eXqWe3x7JbtcOat52g4q043qTacUWBMfLr5TLj0A573D+m86tWm9tgbJ
1Vk+gyaOIXP164AQRKDh1yXbkeLWDiMYNyrJ4XCrBCi8uH6DJxKGgM7RKpQGSZdVGXvmFUb67Nyi
mQjZTYjl1IP35BPsq0X121VPqXoiqUlZhZdeZW6vGVBiJTjqFNUZMvnPTS6or/GHQ6ZKO6FLSBNV
HTKplaNfRr386VSerjCtb016Of5tQf3P40KYoKPc4J0P8ul81ykokiJcPWQbesb5koJNqm/K+jtT
gu6Abkt4uEjSEObGUo8GO4zg8y2VD5IMPGADaU22X5EUek2K6XW36VgqZ5/lMp5GXx8phL+01u2c
JYqaJC7DtO/5IoSDy4jW82/xuw8NfsKWw0yQLT/CxPMxQe1N5vDwGZ8XWVY2eagu3qvcLOLQpOwz
VE5LdyrE76q/1C+swCqEgRsJIsrfpnnwbBDVpnS/pYH2WE8PFGHQUTeaYANYChC6ICGKLKW++dSD
eXHOVZTFNLu6M+PQgMFqZjglpy29H32Ltus5o0AB+caD/6yD8vV3tcc9pCmfshMo74Wl0bzBK2Qk
rWUTikw/6b6A/sJD5TAmMGII/q+LnSWcZBT9D7oopcW1MiHH+D2aRhlkbnh1odb7GjwhJvPrxm7z
DM7a1YjH1cYGD2EYNHMP1G3+4hATP0rAYOuGS5U0T0z8GXFx7Y554+SpuHcu5gOp6GRG+APjXXp3
3J/Sfs2JUyIIJ18HpKZF4+RSs59LAGrtrCaQ20W+YCusOqswN2FKKag1vo4g08Uej2Q1+m6s0GTm
i3zHdmmg2d5v4UzOnVtDC4mrnFykcAlEmwHqNVe86FdSCmutSQ0NNHdt8casnr33Nim5H9geONjt
LgkH60sfzdiRhyjNCyQNnnjmruFEoDpWOG6fks7wUxAbtn9QqK0Qa0Eq6afat2YR2VXNmV1QsoW9
fzZol7ierTCNCyjdri4/whc2uQWXB0JT8UleS2wfVsVvJRi5NXpiNPgolikJyUVfVKvOEeh8CWG/
zgvRdcCVu+treUtnGXvQB+ZuCOTXHaWaLGDhTvWAqWjGky9Uv+ilXWu+BpygMGyqQCP2aWYrc4ui
z6Kvf3Yk5cf1W5t1uhsYbdl8/C0ScfkZCc8F3LnoznewDzQBO7OW2Rh7AlUvC7GHRxW4yl5jkkLw
sq0gSJ+taOdmdLOajl2zkumGCB94cDAhtRAIvznO89ptqL8bhqohGBccWuVqEJTykFBv7tGOnm7g
ef3ifoq0ayS6H4rYrmoLpdXD2TmERLQkHOs9EWo7SXT7GB4f4EJQrynMXCAWiiAVJelbI3YYn3e1
FXSazBuwRm8BP8f4npspWq2yIGZy7+j2bH9nFdiRM1Aj7HHYdxOPhE/2w1AOmX76LDJUNdlpftxR
PGqD2sSSNmhRf3m+HfEeAMeJNS5lS7ua8Vnh24f1/Qr6b8LbR4bxm2up6JsjBZNwgCasEaw0Dopf
nOAT5H0Dfyo1WorUh6F4qJ8TxpZzXSs7s77p31HlflHwOEt4S5cGifhh1ngfidcn97crGnvj9Y1K
57T07i3E7HbIUA+mMSm6OL7xlKZq+6zLYJT+p+hnLQoqpni8Fhj/t1cbCErg1XEtc8cJeZ3yNsxB
KMsfx8KxfJbPKWpTbRvVAIKrV+RiWuI2yReUZSFXbZetoCqYap4BjbyDD1GlrIw/vkQc3GfJ/nEl
nfpFNJoowgTqZsQYOpFUDkaXXA3RXnG3Lg6jO/9xYb+GrR4sADTIay+Ajrk01O1EMOevidZCuxnk
LtLXfsLAG4f/RW3BiHR8wQlZBLXyDsCtCmZkP+/wSScB0qVNx9ElLJxs+V3A7qZiFFckM+phN7Qk
VVQaRlvY8kzDXsnJ/1HsD9IqdhRCHTCHifJB3AJXJ/wwfNrXlOVIACOMp0zafzZYpbQQeLJyBLa6
t/J+Ardch3zG4vlVqqTG6zZQLNyjnFLIGiQ8so+Llp/z1LzppK2rwB3RVHXhiO4NiE8RoBAeykzk
S3qNNAb1k/y6f3MqCY+wsGTPGRwO//iWXGOUTawJ/HsLSy5M5YHFcRNnw0eIxBxY06FOd5aWgtay
DqVAIt448vL6NX3oUULj9W511/jfaJqDhO566SamW+SYsw/sRTEqJK0f9uSUZjHEqnEpem20R+AI
q1refm0jzMirt/Dau7lHkoaV2eYkFihzVzZJpL3S8XxDDY5Xay1awbSMpFm/zHfj13qYptYcq3HQ
15AXO38C0OPvK+oHfin/U3+YNswk+dzy6fsHTpymv2qxMSyw3Ngh1wELAKfQjTWJr1Vc48O1xGn+
oUk5uSe29YGBZCrU1yU25y2qLIcB62Qq+4TMNuhRoUwXXQXFzidGOXaUUnrX3Yd+7nKPLwWFcumC
7o0el5FE49OKrFC35bA2Z5K5/A9Fxi4EshOKqQ4eJWOq9nLVoe4R46vOVu/xrFI5wCMMQacWQRgI
lCopOp6lA09Yoa4D3ASYHZ1Ema3Dl8pJ9cH1QmElJWqKeYIEXeylUA65q36yx8gOLhwLZEaFzM+x
sYShOeF1ez30jsMSKi/v8zqgLXW9dMK6tIUhdh36gVnOYrSUUt8IGx3RsF2NNIXzYagJYscA/CeY
0v//nDKiGMchpFrhvMdnf3slri5qQVOud00GxU8tC9mbU9lSwAvn+IXg94VU8gy3rByVNSE9Yh9c
oDdm7se1/IXewhOfCY7DqMGAiOr4pDa0fL0xlvBGCl8QcA3EglYuGN0a883xMuRQesLzHV0PvmFk
OtlNCs08hi6ybdvUIaQUpW58OxGXmW8qj8q8RkwYC9w7UqiuvJdQXHlGx9VzWFnD9pFzO7XWhGHc
Ep4FxIjEoQbcMT68+sJxLaAzNK+x8q4HTnjJNvDvWSpAFRLSqL+gsn8+Y4bg9LKN8gkLWgVXWatA
udkVtGCjYrBPAZ18GLFlnDm5bwRxSeiIDcp+sdadva73HNuoz6nrYRzsnF/8aidK/hUzaBeHSmJb
5nYSbJdia/7x7460Kmbf08vSX7rDrDiak+R6ouct2dfvHjl+nq+cyQ4QnBlDxndaCFbsWdUgBjoK
EyWJ31L0x/EY/TZ19rfPxt3fUquKZei47PD3tSmWZ14t5fcFKukdVMZVBVy8sgXNSJrkVg4bhg9E
2ucTs9YR+qNOysPpObl7Rj6SCqQtFDuL6Eesz8qtwgqjY16WzJdeA09aU9hOQbJhPDQW4tND7E4t
5zyBqmeaky0kBzx3sNuGDprnVAAoZkbcC9XV8HmV0ogjkDjX8yWN0mM+H67WDG/sc58JREmxTO/J
S75ZGi+hkk6AoJgZWqK36aV24ScuDGBJ9MOqY94Win85qKuDRE3c58ijz8Ckq1l/nlV30XcI2hUP
VZB9Z4e8ogE+/PBY3svTvRZkUL3TLlJqORs50vE4A9NQ0oWCG6Tlb0BFEDGaVsmjRDUnhlmX6BQf
66G4jUsl0mZ18ipW92xeFF/N9s/EY3SQ2qibiAY0JIkdgwxp0EH3VMKEho42+JR0peNo7YSRTfrC
5Xg1zqBfqHt0xVXOtStFVIgrO4xgOlaRkh/059qQLm+lyMfAJrrcBf4QRg1kYLoA2sUb4/KdAW4L
uqiF2gv87hYNkLHOJEJV8QEfJ5qvzrCokI/9HPYtb6Cl0y7t97loBRxsOaXza3AfSkYCqiNJvAC+
IrjjxkknUYiyhs2rgSJ/jxgzSxmdJnSJS1Oc/J/y/Pn+4wwCM8sNEQqPJAPfmpwlX/RXR7VZnZqV
tQBsfeowgr/N9ciCnsxyOLICJg2BATBTcxHjezsbPSGv7IsCNKrGpQL7EDNjiuNq5r+r9JTPFHws
7TEjPrDrDWIz+IDp/lUTwaxb0Cww5HHyqEZsHwJo6TrSZKpwi5N8q4eerurLipBDr7SjmF0vRCjT
0FQeSQBv4Jm1gfn8+4scyFOMn0QSEtjdTHi/MkHaIF5kSkZ4fRnJ5mtbNytReYreiqTffiJ09C8z
wsuMeVuZbO+ko7ysIuqhJk2Uz5B8jeq/xFttMiO9uxVBvOqXZ8tJAZ/h016WbUs3s8vWHKR+TXHY
+Hn3+bo8k/6gxPyk+cHLf7b4HgoQA825BGr0WVV6h3oYpZLWq0aDgQMEByZXCCrL2ktGBI3jF3X8
ysvTySqUYsbWx/VKXGUONmEDpMa7XnlTHaLLWUHhpmsyEkzAqqG9IPv9X/WgoRIbTOVGs55bAqtI
xIZG6igprgoWylTT42Mo+MQfNIAKfbTfpCyQiA+GfSNQCxPFOMowrUPr2Qnhqdy83+EsUKpvNIUV
FqXnuGvNjxSEgGZrQ7jhmEl1Cfd6qZWOq79YkJXdG7hejfnbnrZ55wYve66WWjGWtbjfe8JGVLSP
3jIl3KxAYrUj0L/qL/M0MpC6fjegD6zduRH+IHojmPFRzml+yYwrEH4JwjvxH+AfRjTyELnWrV1+
olu0iwotplQm8LKwscalIMpnJCit++wA8/mMPgq+BjloInLSGMjOEtUirNyXXVjDFLoFYTo0w04v
qm24WcW/zSdcOyHrW2Mwa4CrUz/syIow36f4W9v/f1bfpRYOgeg3Z1ktE/C2kfaKpxQ8q0B7kOML
KTUqD8wOVCf1+xC6SuRSQPQuwlA0IY6vQ3j5vvQOoSYsolrhDGom/Df1pDU0nSCNkqtArruH2FxW
uB9L1D2NGFFaB2VjaRey5AL7wp6I9NBp2RXqvF+gu2gl3ezOkAVMYVudKE02CkPr0HQnGiOOFCMJ
hsAZVhpEsycpgybolPaj6zRTxajfxFgq3EgomILNANI3F3uPqrJ08XRU7q1N3BbDf+ITr88oMdLW
s71HIwDTD+L2tGpKCvDLLxOePAUyR2y0NhVDwVxfCDdRQXGYRczk5sT/pE0NMxCmLTZpmePHLApF
gpVDSjUmJIHQhudYQJIJ2BK0rs/rOVYMXdi0fEfSw+s6UK1vw+/9nUihJ/XxcPb8jUWc8C/2Qwxo
bjEQjGbCD/A3F9/7+DN9Wwcu0fGRkTEsz0LGRfg7qCzs4LLmeEmdI4SEGrMPAydId0D2YOPPz7QZ
89lN1t4W/IBunlwdVrTvBtWA/ZfBxy1axYGmksEe3kUY3ftfj5A4YfxUdKQjgTS8SSHNWatG7rly
u8SRn9sVGRKDbHyMQJgScwLwM9SGSKr03gCfbwGuNSwkxMLn5clwUKFkg+2ilGoHJnWcFejA3Fx8
OM3AZ/b0rWVNYVyQG/ktyZZqbJv+xBQth1b83lBXwKzUF63cyGlw6wNcNaBCPthIKjgyPIEEUBDE
6yB726G+o01qvRjoi9gf7T4qLMwcElauVNw6Mdh6gF5wVFhcup4pYYYa/1GJ94Dee7u3aKd8025p
+Hlot8uWC6zjHcevofjH19sgn+vHyvAMnRsKYnEpspWmQZjn7hZEKU8+YktH+di2vpdimVLBkvP9
Dty5WHgJ8s7BRtiXLE4slhmgITDgo48ZMoiiBL0/6EOeyOIyNUMajcpq87HHIAOWI8FKn9BICWye
u7wlv6m3omERKYsgS2e6Ra9pahwZ+cOG24bdSOxUomhLrx4YD0f4fnUFShGlr5DV7PDu/SGkryvG
griEpc/AD9iiikGP1LNLaSmDJw7xdEPWZp0+LR9oLn8f+YqJpqh+5CwJuvqpGRMwtPtHghv52EEf
4OoFdLZXbnfdkjSw5w2hUERPxoBHoAfbk1LPcIMvnYDcjCX+2xmu7fN7tJIq5tRT0nMXx7NJQgau
L2foiBYyvgSVACCZd2zo9PLd3Sjglxl+NmWoHoLuW0Lo4Mh7ffvz5Qhi08+cnInqJuJl/nZ3yeCi
dvUcjD7xIT6lXm8GsP3E4JzA/o6SLOKyYo4eg/hTnKx9Z37ibGx8kwKZh83Cp0SYBMDZFtKLPm3T
Djl9YDe3pOfaMsI+XevdkopPDotBm7YIn//snkf0dVnVTbBOWsM675T0fDaQ4t54iVIEbg8BW1s5
pZll09PAwRvLUWEBGiT4mQSOkhyFlG0Gg+StOD/z9sNkG5ntA/3YY7peoJUTFugIj/1PM05EMvUL
T+d4jXGE4tHX/sF69fuoC57UpyjqzULrAEYvAoVhODNqDFZSmggnmih0f2DDSY74Wfst+9uV2DaT
O/gD1hOerx62wHzUFe96Ul4+RxUGM/svoKqcwl1pX0wBau57vhUY//KX1qdpI3MxfsIiptujnCt1
nUXVzNYK9aR6iTuURk0lpe4edrq+wQx+eC0TIU0RBzX7LMcKNwwMWjT20K3zhezXs80TlgDuNsPU
MDhfTn4lLJHbe+YGZ1ELHGtbN5W+RRQmgLjvkpDlRWkhNaDTQJ/oQm5S+QpRFS5xUrt88Sql4Jtf
vQNaFg1VMk5oWPsxObEl3ylofRhvXXUIrjfX4XAnzvF0KzrEzNJb/eU7tmMoUKWW49yLqLWG9xjl
DZGZDb0AmdFpvy7xwXzJI7+76Fu8BhL+6jq4B4yyk+NwOEUu6Y8ITR+lPB9lE7qy/5gDAMQ8lWQs
Es3F+lb24UcVI4ce9mxbjT7Ns16JxHGFu8s/61UFNKzxOydQx3DQrOc9oBHD/6HfpTea/KGxb+BZ
wvkEwZm7iLJVEyU2cJm/ZeYE6XXQIAjb2lang6JYlFX/JoHKxUURz6zD95A4ENHzUym4Bm1bf4NC
5P+HWczsno2NA6gbaLcUBvPbpI1hC6dthOZyJGZDYNzdgIKOXCC++s4oNPwaAFJ+FN2bQt7fJzpS
SJxN8i6ylzMRohR7+TOjhL24gUlITmflAunGpMktk0lIQ82CjlgtXrUb5bv2OXZmydoOKJCmk4uj
HPK/xk+bhrZ+XO9QxI8KmO+N5wFJThP47q9K+YY/6s9DT4RCTsa2mapQROGAc+PBwwOLENSdpmLa
KcQqug7D6s7e4dhJ5v39c2Xibl6tpOOJuUMN25zbdZLNfV+xdan67GQOEEnZVSXKhevn5cYgVk3+
nDrlWOJEmigs+v4VmDuHypRBk1Bu2GLTAtWbNwi5vbSlhNZgrBoeNQ2UarZOSJIlxcuxVRpTLpA0
JCT/YbC6Ktr98r06JfbjLMbRmI5rANpAVOYWyZqppbFfv+SMluLIv5Ec1UGQT4Lq6MJWyuRJiSCx
ll+YrOESFZOJKeuicIrFLPX67YM2y6AYSY2hAmzk4TtNQmyu0ZSkDxQFS7oa6rRpyP89JObF0RxO
F5ZpHgka+rlS1/0vVHejPsq9sG+NN5fauxHFZEvYtqL0TScBKI2p2DWsUb63UxXzRqyZyTzlTzhJ
KIwAcZQxnJoBjuHzF4w8WZ/Vp57EiKo13iho5k/a7w6cQ/x5TNqL2Y6XIQldwxLCVUlI+id7GJui
B/2g8tJWjdbG+D1MzoF909GeFpjnDpIzWvaC+Tt5Hcch5YpAqbcoztzoPb2WyvA0Z2cGM46BCWD1
w1ljs1E0zEgiOMcgt7enQVic2iPFAKYb07nqQy8IpVQlrcLPmD0vWOKai9ghQHhCTbawwAAJb8Tf
OsmesiZdfWPVJlX/SJimDeJX0EK5NiqdZw4r1DTs6LnQlpIl1Ck7OMljCyBds5KsxWtdb+kDkbPr
RGnjmn4+8umpDU3JB0aXZlSDZePxv3LTIUSKQC57/DqcMTnUQSIiWiKcou7UqAdKZfEdL6mIWu8D
pABVexpXOQ2j1AILVbqySDkwT2f1R6w7d3eIYItN1FnrHvq50C8Koc71zcljPQZ9C8D0cWsrYH6h
xyYCkmjklKUtiLPRtTV61ua/22vRFE6ztnVcf1eiJL9knh+thxXejUXDdo5NEigeD12Hqx7FguIk
0Z05FpMzzycHpaPWNwvHJVOOJosDHKJENjkTNNSW2ap5p/VRhX4dYnWvEPm+n/FPHB6mbbGEkUbQ
MJhDLvJjljVa0YLiPyeL1V1seDzD3PaUJFcv2IQpi0DYXRQKjTj3EUNmS80WpP5d0X2MQjblqxBD
G3n45wBBEyqHTv2vYfptsoksrVLyioKlT9dy75gbWZIctg07vV8Jdkl49fWu0lfMYoTRmXpN842f
Qug7w/5gMgA73yghb/Qo3lbmXvVOdrKgOVn91c/cjh/vGRk1oWv3q/DxzAJtekZWN9M+vhGheRu+
G7SlRgGhueuhW1m/phLorzV8F8//+vp2m+J4K+M2zkXP2PEOXmJ3cV1fBDMg37M5k+ku2jxfw1I/
X0T9gJyyjN4ZGVEnvN9c7l9gXFp3k/3cJfaK+bE5COrZI/jHVjN7FDWjIrWbJm8aYk+H26UzELld
aheznyTfNXhFhPwvyPkekKKhAGzYdU6E2zWTuvkQK6Reiotgl91lWjNlVJU3Hmyp0ThcX7kCwrnL
QKnhWY4HN2GR5uw9zFzwQQVpKXvMnBFJxFRwDOGzthJ3RxD8xDoja1dDWjFl/19m0KOKIVorIeLF
EJNWLuVLgryNbZa/Z+j1V5a+XYuNG2Y2U5jmmZ+Lz/rjO9mZlZhgy65VvWxmZ1Uup2u9GUkotxNH
AFGZLZxFGDYg6XO4eHFZQZ7p44Dswn3ynsRuV8OXXEiY3e7AabavlLsH7/6K/oA++oIjrMLlSqml
NnS69KdFJk0rmEJ8hS/uLNsstCsJCVbh6PXkyXbnycQMOGHElg82FUdFxIso5xhMfjJe9ALk0elf
nmkJBrRKa8pgBPvvgmiomd7llC2XmYM6nno/i6gfrXfg6QRsIZV5ZGieZadOTti5Wfk06qP07pig
hdYegS+wxwrhcYg0AFmcmjLIT3L3l+5LYD6tnpZZ8xvql8yTJ/nzIm2c7lMUBQJIy1w746+hrjcc
HZfXqvxMZIQDu5roOq7e9xgOW1n8OtDulAZiElfvY6oNZWTcWvCh2B/619Ml+eSmG5YOyJzJnDSx
aWGN92IVaKAbXZPDnaeZ1sorPac750WsVg8e8O5XxKLVBPgCjUf1vANrVMPVZoX8YnGbjtlw3R1R
FnKHbNn3LTjqpmufBWhNSe1nSj86SctXNEGHj+74ZftHB8dHf2r3V+39eXbtgIlJGB/G48JGMGsl
1UzlUaaa1w6TqO9OoHYXtpINH0MkTcww1hcj0WrZUUH7dh2PF7esafQAUSocqBQQh8wxenVyvz/N
TJjtulHp32tHMmwxhVdJvRAOycWRd7RdwAjbtSNDotH8zRZGrRspPXBIyjxlLtubx1s/UhnYqXtx
rvtpB6bIIxZZirZUovQc3QTJd+4N/rhDx2hC6lmd4/7g1nnyP9RTBCCYGMmGV3liHVy3tTnAoc2h
Kz3jhJqXAYroju0FhHSxNuUjF06wQnmN2lc6wnlSvrSvtzW3tLvR18ZwrgXRVngRgpEAjCqk7/hp
JDjRdogxlzbWsdh+1icrBa2D1A0F5OjGt10cELtrg/7JyyE9ZWY4JWaeFiSr6hxlCd9O9a4+gb0V
2nfNbj0YUMXW8UdMbUJIbj1rI+hjq543t6oXiovE/9fitmHf1qdiCh+3mfxtcxBGiGJHaQc9toMq
RIhfg94S1Hg5pFgIiaMfvRafVno1RO10iTkFAikp8f52Xadwb/ZuH3lSv7tn+qmTvhDhXZJp2ZS7
yxyYvKMSE9PUcm6YtTtVvjD99or1YA8Y5MqxmWvlf81gW5Wrar0ruzgTGPA780sdKiwo4od5sw6C
PQG1VXq53dFUaafaRPcnKMq/pOQVsfUbKdkr7TK+nYjJ4gQ9Hoy+mIdqFZez51W1R7V3784oTbY+
/Nxzi01I4T1rp1WxVQb/+Jm53QhCTqXGKmsnL55uje6JhfAV8M5KHgI/7QFm1iT3aiUBCRqb4o/z
xm4VK1GFYQMFdl08N8t1+TcTEDBUZntOK0NaExkUCNICs/Ob6W6AHAnK8tgis6BV7kHgKPeH20Jb
C3PdKlAFcQaVdvPb30cYhuQJU8NomjXucUzEJXaEcA0H/AB1RhN56YCd7BWkBgkqcMGHTk5my0q0
Mbp8jsdbr0ao/FM+F8N0YoPa0/X5XUyF7egR+fR8EDkYkPoGV8mVE0VmHfcmWYKLgsJ8JoR2an54
nRXaJ1M1X/7mWKWJ3cH2oN32e3/ldEfRdHKdLt6Ga+hOWftvcnnU3Q84PAxEbSG3y1Y2Hn2iaTv0
abXiiTe2/GiGuSA4GSZpuVRddQIPG/vMERNZlkk5m48+Czv4oy7v6wbpvj8zn1kfW/lpVIxHrHnr
FNidLC88gGGR0lT70Y0NoSWpHHlT7YahFodchviIqXDCe8AJxJrfjWZDjmaxRuoKnBQAO/6UDW5v
OQzIMiTrmTG4fQZfbs1RJjiWGs7vk1Sc4NQb+ho3H6OxpNvF30B0uc+CwqBWACvvd7AeBa933chU
v7gbtwOqNQkDTlA7HVqGBX5gKlwvnQVjAuVYunM3u9fIPLvWSHrVzdv63acMOgPguXaZtrBVrkOk
EBD2RwIaiCrFzIJGocZQ7G5tWQF8tAXmo4ejnJEchkRzkZn9NA4AE2r8LPPdMCo+cOxeRTlEI0g4
h5umIG9fRoS99GU0P0aCIp0m5ChE1YCIQRxi56/GN1taxlwW9QZn9tIXGot6yd45nHh2yB1+fSY6
wauJkLAdsjzg5DkF2cLRu1lm/bvPt9hG7o982r/mUVMemvsolRMYdDTg25AdZKvNEfMH1gBAjH1F
ZGCoHnxP65Vp574VTzJh4IP1ysyzchKqriVHPxsPcdCjXIvK2Pw0kHYOp0tofcOvnXUh42qr9fQG
ZLZg0Wg2os8mpm7quKtszxDAvsdZOaYP9gQp2HON3F9ml4oE/84ODiwnv1wSDhupwYP2zO5vD9Zo
8IFjqJRmVqCiPzMqkttYZp1XugHTDrltVJ6DkSJivjGBnSWE1KdkO0wg510MNIcFVJykk6GKk6IH
i5o3JC/OnzOCZC3C9UbrnelvuvnKsW73ug9mxKyTQ/DvV7TjgZZyppbB8HZqTznde6YnEKmlSDFQ
66ckLAHdIFrhRdcDVE6RA8XYUTAzePoT+7AOBgy3byaXizoHnhXikc66yDIyrRA5vTTtX+XI/Okd
p7bLUskJWG2UTzCd6kK5+hrceu6RrnGsGQs1JMAoP/ZF4gVcLS3uZL1T8t2mEtN7BJpukvYpMDxN
XUouuKZDS9co0S5umLLmZvT75r0OVDjGMMtukzSvU3HpGzuwydKaLY9gW8BoioaiQX9S6lrlOJ9L
ktUbR9JPe1RG/0Eea6XTC2TMUOydoFRN7dbinTjLJprFp7Sns7OqSN39lR2cBAyLEUt/RnovTbk6
chzVn1lL8DyulWpEZgeLGKovPlvPZdb7Vk/uCVFmPslaVSWqNVqvniuunSWfVwaZmxULDh1zGAA5
Pq25r2/YIjUoV2pD9xza/s5yb1FWlinr29gYOM4d9SXeWRh83l4vNzMOUkf632z9kPY7Y5EZ971a
5dhHvUEO5IKDSOX7LM3Xsrni0087Q9vnJpKfpOayBPyLWT2s1UJpxSYgPFOBCDRdIz/Q6YAa0Sai
1LxI8RW6IslKzKYuV6VmzR5gjuR1y020hzTJdYWNPVIjieywg7rINlrd3jxLdrCXthpie/5r+FD+
2AdxUXK/RuR4fqO06bVErE12gFIIHexcCkHhJhXkYvKcQhFPO7f5+DgLx8fFHvRpbL4Mx0CgGQ8a
G7o5VNtgv0qiukejTuk7WD8KCLm6F16OQMOvacY6ditDptI2SZwcNaQa8aKPyuoqeIRcVOjJQLls
3krwnkfTskHurXqYachEti7Jn5hYUtlfzYuzSm8pSX8lbjYxBFbGV51UBb2Zc+az+l4fcypiucjf
TpKWw6APQbCvHM/AplMdK85aQnuhIZNcOremSQ2oLFnOav2CBHN3nOTTPCElkVjH6I8w1wQNXX/w
32hD/VENJFFpJ9maglkgH/xPSYcMsATmro+ahfVCz01OkN7TzLraDwFXE/EZpsQd596/eeRlZgPH
MRQfTWymsTmG4pQsLpPKHOeDth/WqD9EYq1R3QXf6kQmXrrbceUaQRlDO6BKWMyOrbZK0e/Z6eN7
FnJ4nmNGDLOCQVTwMRp9OzaYxg140rFwagMvsDtFV47eBb9g4iuWFLBEjrGIhwXJAUtuwHcT0Xi9
zCj4c7G24SzGbkDQpyig041EMLr0kHaUtsVBrptXeyrIiRYbz+KcGuNzPLOIqTNBalnZhwWybirz
X40oHw2Iw3b3yW9DDAzcBCHZv8ErbINBv8IKWQ4dULbqenLiKFqIBUVA6iNGpD9LUAyinsdY2mHb
JrP6Ip57MPQ91BF4CgLc3B3qmaRf5XXicsG3nyoNloB1lRLVG0cZ+jcxXlB202aAydVNld13GMVk
O095CKBXX7o2UHUpB30MEwi5fOooN3CorOP73Zun9rLhCw9ABlbFd7ezi2LJjt96Vut9AwVsjWWO
PjZncxKY8argOGXyfoVwLDMpQLvIP2e23t+OXBPV7STEoI0q9qjbUS49SuW9CBLpDJPoIZMwYSPK
IBjT5OkPxYJyR+ZEJn6oq91N+8ps68VIyv1NcpG+pLauwfm7NE9OFnifCUY12DKhXmd5HDzS72KM
nnoJ7seF5w4+rFovq3x87xYa85+EJqN75HfnRg9qkk/+FLA8FFhQZmdMLRTNKyPGa+Eg5/A/GY+F
KTHAmMj7bCX7YBfpzec9DO1SOGieSS4at1B8h6a8g/m+gt+niJt/j+A3HgMJX22OFBp6LvrlFaU0
Wbl06pc+WPOORrzu21L2IH1Fc0zgLZvbp3x0stWSQwIVvVWGvajNXsCwQX8my+tOkGGlzdHwBkr7
h+JsJtUzJMgHnS/0z9EI+HG2hFQrkvfG9+q55gh+KRaI5/vPpNCIcwlVkviCJoIJaYTIu4Fu9hiB
Y8TdQo6UkOUoT8dXvvp5VN8+J5iRnsWWIfFPONf0AYEHOde5ie5OsR2YBC63aYEoN/6fAztU1hCr
heSLev9KPudXVpWU/dzdmw4E7eemnkSLyUbfAqvDkG0Nl90lnlvlvRH7WVKMWv/rM1P6vALNkOB7
oMwlDvChhBDx4dYGctfym8yPX8FqLsdNiLCqJg8T4MbnwYMCk85yrgE4YIVnlP2bnNcn2DsVcZf/
G1LDe8Q1dXWqzaSPQrz35sNaHg8AhIpnHVUzvhkxfBHoxloG5mzbHxMICaGO71DRL21d+QINLPrq
cwi1JAXbr1mFXMogOyIPxqpmFb2YGD/gYzJXPiScxAS9In5ezIy4/MyxLMpYhFZ73SgJ2YTgFx+9
DcUCqZy2uQykFO7N6Spscq64D+mpF6q8EcNeyeIfEW48CJukMgbgQ9knEXtZVNXAWdmqZAxfbM2W
0faNzzmPCsW5wLLUstaNltqCl2XO30+S3K8yuDfqnCQYPmRVAhTGomp21rdpTgeDJe6TbznzmmIV
d/Eees8O/FoUFCiODtkGam87lQNC8irhz0P9rhbGm1BOpcKSCYv7EpVsQLpul5Nnxi3rfkAZZ/MO
E9ci83b9uorekg83wzb3d6US+s6ToMu12NsyvZl7J51QD0VNAK3Hklj0K48Rw2Cg0GN8ptEwDnuX
84jbA1Quz4+2jbIXgQseiyUz0scDxughKJ4inlCW+GUHCmoHYzz2CSgC4Ua2T2L9NQcfPMqUUGBV
b6loyLKkGRsd/oSwwiNW/CMqS0BpTuJRqEXFuFwv6Qtw5S+O1WOHIjlhZPS6JF2FG/AtL9HLgHvT
7XdCMaDTafBueOaodBUIpSAJETIO5K2udoD5vYQytQelnZNKkOVjLVKBY9tbNzNAiULgiyReFvMF
LIDFhkMqA3FrMtQ3chetmF/vedlRU3rzaU/Z0j8DC4OCePdWUbAE9siNjKULlUO/RMtnJaTA0lDt
NfD58iHd9JI2yCytllj6swD9f20JLw7MVcMFvwE0duI2IlarlEW+o+X1wJzpe+LoRBGx9hwLLMxT
7w5X9yYfOG9nWpjV/Q+Zfnq/do3am812WMGa3v61Ivmw/DMjc6oKp/Qsxvw559tzu+xBx8ybaud5
UbJRngats67NPfEg47Vb2XWb5cYLWNCIQ5ael8JoCHKFjp369+UL1kaFqFi4QgYFkSY6K4bmjHyG
V3dFAv2uuzAbKgNLc0aOkH7cyIrTJXB8L+MmCKqeD8SOpqnPoAsgnZ1cHrabWKrszeXxvsTNBvb0
6GrMGDXFaGUsSQuAViMCCiwrGfK6GmE1Z4jNkOWudBrZI93iKXIxseNEFMxRUmaiNA22pMSOqT85
RYy7dTL6FAM3rgk7wtb63WaLf1UTJ6WiQbkgcxJccKYZLRrF1QTESOXmAOHIMblSQlMadH+HkHjq
1+6xuC08L5AtROM483dkveV2FGwRRfEEiGteSRxCIzANA22/MJ1711p1pjVu/WyreTCHbHtj1UeE
xCg1+X4uZ5GJFc+9rfN2HIxoMiLdvHlYZVnvPJJIElV1JWi1zOsavNfx6LhSefFz75FMfO2HhfQf
6zuGBpb8+CVpAC5mFwfmPDedP1dgIq3jYr4LoWepx85YCwVrQo62p2Cuv4sbGzP2J+JX96z8h20t
ef++Y4BI8oukbXT/LfUQZ6iwFy/+fA4wF5JKvqtXrPRz4yslzOt1OlFwAPIoCKkLnfWXW6D6o5U6
YPgaNMWJeLiLuGvRrjupIE7vvqnF0dQhhjhpFAWn7kiw2owUUfWhkLgLltMoJAvrqollOcdULMXN
Puu/Vq/5dhbJ/UPnA5dxZg/DaYaFRkDLDq2elxZZ22Zw0reLgA00uUMkbOfHOiUBIc1bpH4S9BMB
2ECQY3YaZNGIt1KxtN91NfgCipJqZt5acMklACHi8YUGJL/wprgmlZ7cN8UnMkxDc9J9jyQgGjvO
E4mPowAW/dhBBfVIqcu7Zy2cJx+FIEBQV/PLEWjFq1abxLDeXTN15DVN8GJAMsP7T+MXwhx3w9uc
mDjq/rW5nHK3bP8fNF1rzaSpE7u3j6/aBhd5Vmz4XXVACKrv/+GRfOoTEYXXU/QZpsRYK+WuhFz9
tWYX4tK5z4a78496aSQHwChveCMlwl1n8CUQlfEd3Gsnuor3yurXcMUwjzQUKvye1cJY+6zinO5/
nN1IfW5sU+vUFrcZ8hu5MVIQ7z8YnswPRENtqOrkHkPW9q8WqItoSTyuSd/aOWaSJ3HLbfJvPZzB
n6Y5damJveVZrIGol2cHjV7OOoD03Wk2+BGdl9D8Gd7hf3IpxyFqrpcSYXBzN6aiqfcozB5JPLY8
zZONca1LsIu+FFxMKt0RcHdvHP5RThi4NYpgTV0IVeS1MZ7uaP+KHYxecU9RwSm/m00fAeUVewhN
TMgw/BRjtK+yW2BQRoYkKfA6LVJmeqJcwRy48zSxeAds8BMHwRB91neeNK6NvL6CELnfVsFlcjLu
2OpWzhoQIiGt/gFCIFHhG6tJC8s81v7JL6hqT4AsbECgDCuQwgWGnGydZhxMsbiBLqUgmeZrInvs
fKGeMzvmj4qB0gqOkKD/aaQXL+0IHrMjW5XHRiNtyMBlmxYqrHcDc/bgCMCUCk/H3a5UEA396J1E
1xZyZ522dNEONu3mfJfonqF821Tq9zfrFnvJYC/Ka+hLTMbb1/gM2TFv8rcwViBvcKs5Wk6/CX1F
Il6XO/vZKt2VmHRKaXRmXqrexcn7RsK/7y0n6OlHx5Oeg9xkCzDhuy1s7H8jQ096JBXKb/VqO9v2
Wa67cSGpsFmEDIea5I21AOyxh8DKT3VqRk05v4oJ+GGIWddbwrQLNWoohzZvXhelHziR7XXqfXqy
NUTO7mEHVMtqkNLDkhnVEYFXBDK5h5+DGqQ7vdfsWlRp2qtXBqiUe9f8Xt94zGrERRurlmhpPmDL
2pkQRuLnwWRrQO8LGE7jo87BuaqxpfqYR1T8K6BPWwnE+0CsbTVf8vBNOhtiXZTitq65XbuYuTMz
ba+8cr1bnbCh++HR7sPhsKTgju07kBNbV51uR0tqADoYSwINVmMqDrVB2tma1c+ZvzNKY6nTIgXe
/ZQnRjW0aOZuip3OXe2v+frrAM1zK0IIadqZz+ELfjRRCBmrivvcrlOYx/75oT/bykDKt+CaepR/
fXZForwMreijbIL19jNLutlGiOTTQYYOgUqK8tEVJsmfDiH8N1DlX5xE54imMAMAhs9upoX9ysZg
P0ob2i7f7cBhAx9c0kyvoJE1kxbDDUYgC74RjqW0e3Mr0uhlm6zpFcdUW9BYwhLnZx/xEfnADtd2
3uXxR+nSdV5hUe2yQ9dsmjK2ELbg0V+xthaG75CoQfV1rqHMeQKdDuMuPahVsxngtInDSta1tr++
QuVbN9gi8NeTZw9+2o/U3/wpW6Mcp+11gWAvwgygGv45C8uIFaACVk4pjvcApQW5wezxWvZr5mvY
PqOgUuZHfPPKI5TCxR/jiUugMqPMYvT7O1Hra4/ztSn8D4XxzGnrfM3sp3RfOPf455L0RL/AFk5H
LunjdavpKBhDzEUJOdhUIagZOoCHaKQdIeBxahanXXOFdqAd93v2UCrhoZr8Zg6KBM7gAL/+Ovu6
160+jIhxNrNqzal2Ub2OuKSW95dP8wl1QdRCHjxJO+U4IfPyty3ns4EsN1bQy25uU/Qkv3BwfOIc
EM1x8HPeRPb8eXhDXs4QByPVsvt7pJrlcwQ1c8lsyXSylBZDPY8L0yO7w2X5FgqKWPXVTk3jjtH1
tsNw86F6tYWB3bPl/YGko/YZYZKguO75FYYPd0RySE3TR3c/r0MXmDThhvXaQdPNuY7EBxaxBuqI
o5OibIoRdxXJLgccrYwyWD0GE50/yp/s+dNqk1a97dVRdTiu+SU5Eg0AbWKXUdSJ0ZcdatlRTor8
a30SV0nbBJVYUEvpsSQviqmhVg4f2wSp9Y6bDBoXaRuWMIxU0IPLXcahWYKV5c78SLX4PtmHcHgn
gqWoJ3AudmfAZc4KI8zl4n9LnqdPEKgW76dJeT1ZXIiDYjNfhRwzLjDcY0uME00KcvIGAy8+BZOl
fEJKKMHC1C3DmJxzc5opczz0IvgOvq/PAd14BTyJefilTvVDJsVwavyhnEUzN89S4WQ4qNvjAi49
xYyI47jDYonWnhwCqhMU3Pof4F8RYMGFjVzTIgkpL/VPKtdEl94qjUNKhZa4O3SCB963Ai/l+Q7+
5vsCjw/znoPfTTiyrAvPIEtcUEld098K9IIQ0D1en6j7zj1PNee3XG3Wr2n4WbLOa4804qBCa/qF
gHGut5AeCa4Ks3AjL2d72NFgRbJuViM+FxABTz+DL4O3NRC7mbUr/8F6dp6GpZT4w/r4KbuHY1pG
VGQkOkyBku1R/yaH0/HfFf9GlJpVmTYzENt+IeGz7fKCMDvdBuEWwNur5o1mghzKph+l/sYmrnlg
H9IbjYOwResXWEnbBKALfkntrVmRBf1VfFCIaw2Bx7byE8BrnPnESO6DytdnKl9MPw84PR4ShqOk
ozUhVXQ70ssDQNJawq5nhgXUp/wefXnLrHJSxSOwVQnGEXVqwQisYai9SjiTf5MipoRTFzRoCVUH
7PH059Q2ID+BFjr0riRxC154dBLJlUYlVQDhOFcdVTczC/181vNJ8RRfZa3lX8AlQzYfEk0Y8hP3
agAqgkFVEN2bhRdvOzn7xOVFqKVfKzXcPFKUXWXTMHu2jWqUpM2PO4OavA6Qua1QoGQraypeLynu
EXLz/9ZoggzplrddQR8gP9nMk0T1U0ckvLwH7WL0mYlOc+4d2CxNLhlJK4bzjrLmPl5c6cz8Acod
zRyfFV9/KTZtklHz9hw3GA5fMlv1KfxWi5hEnYXYXCbCfquIk/igeTx/CFzuVuXTgGfHcrMMMMSg
UaBLYf+/u95LbgV2cKNBXPeego0F/r0EkZq8QPxoOYBPUGXx34qSuUNHeJj8sgw4vkRt92KBLPWe
O/qKB4fOmW/QklOqHIBm9NmUKe3d8iSADvtNq+ycoahgXUKPvY0fTv4xq0SSRWvHkQgom84xth3Z
0ZQH3BSssT90StmVZ3Zg+sep6wrKUiQsRuMz7gp3nIuEgOLR6I/g84ncSr9KvCeGWTzo7iB3ZmQb
C4XbVJG+Kh87FpAmGiDhnZH6tRQ/YKLBxgUZAMes3TZsaCGEcICkuGs8JgRD7cdHxg6kRDO7Ckke
lJeS0bJeTHscw6E/1pg2o8eVvRJ2WDxIOx/KHa3DJqk2+rEMyhSpXx+rzD4iQNE9a4PNyUtB8oED
bx2mHXPDbm+3SE54+a9ROANufCFfzXw82WTHLPQIH07zHw55IhpaJDi8cHXrPhqghmXm1M6UPobh
cwiCe/KvCfZdio3eweymoDjt4gYHDPiFQ4sQKIy6HTCUIuVoEzLlXJ1MsQoAeNboT7kpPHLH1sj5
/8EY0XbS0L6Cug2PS7l2hHESTKMxakD/JG7EloelNYxLS948JDvLehIBnSCBeNusKaY770ksGJf8
OyLR73mvqgLMLPJfnRxbnMGJV0sZS+lTAr0k8frLXtYyP5H1cf7YLOxkNgj2jZxtpX7L2pXQs3+t
iQzukuy00NeK/20/AXepsxL+kyGgBsWfDGjsqcPyw65b750BMWVVyho1nuPvBU/l0svewfIYIRMT
FLmH/E8/K0AQwaglHFCfxy5OWDHaMxJgYrI9TSpzG+1CeW2j5jIj32/erKNWZMuWuTye/3O5ym4U
YH1YT1LwGj+8c9E9FnQbOG0F9YIdYIv5izYQYTdcGCJz1WH+7lHP6QhfPf+6T4o6N4/Md1an8kUH
QGQIku0V7V+WTYPw5zD3k/uwvKiFuItU6LZm8BQ2LB/ZW6qtCdVF9e8YL0vRtTpkzzqIO282pQ7/
wl04Zg5WsdFv2HFueSC/WqdO1Aj5m429vdkV4TTrwO6XdwhBzKoll3cNEQCafsnIhK7ozT4ici9S
nf+JuYJGHy0RsNTQtC32sz2Hd5dOcAEwVSBkClbHr/VIJtIhHy4l+V0Jr7/o/Xt+/iPhBvIcYCmc
0HeIRHmMvl7ZUpdLQGZoHftvG3FqRnZXpA6733mquw0oRS2Jp6ahreNM7Ax0Kkd88Lj9DMglhQ8M
6bEeWVfstLbBJQsdaL2SDJfxRrV+QJpxXx1hHI8/hZppfwj7ydWWGoDBqAJAaDgRxTuAw0BU4dmQ
xKMpxG1Hc6q1rUO5IHUE+eHNjT0tIyWkp/ZiZIdV/99kEIVhQr4YMDw1MJ9JpfgIU3yZzMxTnFnl
x/+/gIX0RLm1ieYg9kCh67iTTIbDhhQr0ScGGqKzhjwab5Qb16/qde/xWLAIeKgNWyV09vqQYbz3
GyYWm7jIR1+wWtYOMjsR3EYlrLN/gDt4hLhdA3x9L9glzrsG5hv9XeqyEhksMIa0Yq3F3yQQfRWQ
wMOnwfC6+DkvlZ1gK0mEJxxEEa6QwjLZ3EOj5iji+rzUtfp8EPM3vwzFb3q6aHicXU+l8DZyfleo
i27cSO1LMuyPpUP3BXNb5nrJ3W9sKsWqEgJh/xPSlWbJDCFkBgdZMBSMHksXZW6pjj+QD4Oji0PK
m4jgsaApvuv+aBrtFj3KTGmJUDajvg7f15j/jddosdp3yydHgQ50ZRBonC62fQmLW0+W9i0dACaQ
KIL1EadXi6V3rF5ooYhequN+geCu8Ka7PKHVVSUz1Dh+1f36XRAx4+7VnO8c1VjWGLEp38N6wdrd
kjuB8zmnOcmDsFSOxB6HfZoRAJTCE7YEJv8lVj7AQ8j05bQcnM6hvTR+RgKo+BfkZ1XU2KCxxFgU
aXXjzeIep8ysqH3uMm57mWldNKbW2gku8ouCkr1UJBeAB07ai8hMhc6ThNehUTYYmJlF/EDNdVZP
Ss29QhOcohde24hKQ4zVWjRMyYPf1aGbuuc4w8g0bDBLcWeB0H5IhpopQq4Z7uvTJRqjQQdsMElO
xdO7tYGI0VNIIkXRpR555MVlhZvWV6ZCsfTiStwdprJ+gxsasy3np4y7zgmw5PASaIpHQ7uJ85IB
1jVESHsNFpN9jg9QAJ++XYw8+oU5/RvkP7QJp1eZrLC33274xxn/0YMfM9zMZUer8eU3ZrxyH+Oc
c7tb1/dLmPERkF6xZV0bunsYS2XautNgvNF2f/83J2BVPOtQwkIxSPIvFj8lVoIQeeg1OSscdLmd
yA9/LxJmjsW6Dhtanu44hZh4bvQYxohcHi2RjTynRrc0tEBhwd3hCD7S59FD4Ikx2673YqHMuDtQ
hJWlbs3A1o7M7Tgwl7n/rgAZJGJhGlBsvJppx8YvksVYe2J6nqwJL5SHN/Bz3v2paVBxzu766mSB
z3rSgoDM7vswDOd1r9j85K+BqHdw0VhlC1AGq6WG/JQpkBokGFQuuvJaktzloEkShl6g8lyM3xZ+
Bp1l47nUAVd2Ulq7wGRGm+oQM+YBhI2zyolO++nlABIBPH37RbqEZv2vp3CAJYgBhbQQWCypGafb
F74Ze8r786jQQrzfQUCh8DDMBl82w7yIVLO4mAi3wG6nKuNFLAGPr7U56myd8IkNLK+5JqdQtC/Z
/7ttyC5KU73gYUzgx50r4WOc4uT2hX5NPVW4qk+1AYLeACUZCmmbhyFmzTewR0QzGCBY7Z55G+Bx
49MW6RTMAKGpW8IsrsK/0EM7OZAgLRX0CTuqM+Z1SGGeyFzv3Jxc3GKgLYMtM9gnQCUoilJsDFsU
Sr/Xda2VtINFT/6bKM2ECTUL37+QjrAzQbgff3NSN3TBMkAywMWwHxBsQeKW13iKmZCrZlaVJMb9
R453GLXnFlcECoQ89ApJ7DCA+30usX/KxABINWrHNlo2wqPUQ1I2GZeLOvaky1Fu2BdtoSZ8OVRQ
ucHBlCVxBW3gFvCOL8JMqK/+roYcRe2dLH06VHwbyDbItmHD34GH/XLmATU3kxMmaguz1XDesdoD
Qp9V/WBAEum26eOZVHf4M5XierFXClVw1Eidzo35Uh7Q0fAIS9YCuGGIt2xKZSVqHaAlbLv05tsj
Ujcs5X9kjkjOepKpdmpq1SRPh6nj0ShmgGjiYW858GUlXcX/YXxMD3aMuQonzZOuxf7Nd1tuAW/6
+c5lgQ0WuvIvVZQW6OxwYxiJ9OmMwq5//9LAXPk3/Nb2aP07bpou+np/r8SHCRbQtfU38cdKxPxT
Pn6TCv7xC3KNhgS0ImoQnllPMwFlwYXfxiwCWBfoFce0DDldzUnqWpO6KpSrt/9bPObKgWjDlDMB
9lxtuG5M3chYSv29o7cMFOyou6tDUAWvKWW9a3BIOjZshKVOaKviCXNsKdddViXhs/uQRZB6tnm0
Iq8mkfgpsF6x+D0xgCHY2uCX3fq2oJmxHbs2lmsx8WnZGhAeV3mywAk/qUf9PDZELNnoZj11nuyy
0Rh84xQcSiD0MoazkJJmU3camomnKJm5yWjWgJrdhnCpMtf4xR7Lemf9JLSV+VEdJJEMZbulcVR7
1O7pgAGryFZhS0y4V+EQSY8VA7COhcy87Xi6bYsn1Kd965kHXNu969dvElKpQPpYyYzXoH8KwWUi
L0XhDPB2BRhd2fSSgKLf9/k0Fuspt1TWB34F6JNdkpXKDpDqp9D76GGjz2sXcXyO6LS3OYkclGC+
I0St/WfNAnI6BM8qmbFrryguPZvDi72NIJ1dd2E/BkvzP0K/t+MdQDx+mCuEj+unGIy4rfPQYYt8
B3FbXO7SVLp17lmQkU6c5UVvo6k3/eYaaS8aOsOZMxUD8TLd/HvKpj+aXW2lHZN9tGOTYE3hGndD
4JpzUK/VRUB9gu+IrQQ5QbWIBDMWYiMqJdI6+rsIdInaAs/pxdQgvjJl0bi/8YXdu/2C0Qmp3BY4
BbERYl1aXYC66GwqwWVMARHPMaHsRFW7gE0Jm25QI4UyTU889egTRV1HEeSqaadkoiA/lq3St2np
JC2v5ip/+yt/IeJlGGZIVQ+mg2QIOyNu9o/kynXyxgH7j7klVCLcm1Ye+4gR6+EZDgP/0UFsX4Rn
166g1IU3EW7J6l9nQ30n4Rip+QCzfNsyq7TWThBZCYiO3MP++xGSD3NYGebotOEY9MHbM8QvCMWs
rWyF1YFJnRvN9sVhOKrDWJ1+UmHUsSd2GVqP1e4XDMpnamMid5fyRadlLZMkO/xs0VshTFj15IaR
0WzMNHVbsB+d0P2Yri2wTg17/CEYmA9ttxyuzcz5VZB7IxrE8fl0vorDecMY1g0qjiluE52DsCXu
6EkVvNB2WhEsTMcW8lS5Du1MyKYbQwZDkTuQ2hw+yM3InV40Ne3JuFzQyLQPUmfeUhYb43fgUbXj
qVHckDUGhdxyiM7uwz6yF6W54AL8pgcsbfQNbuGyb7Bpp1lFhSGuSI5CvNEUSvEWmA6/vwcCes7V
oaHbDjifH3TgQYLlTAei/wAFoBEDaKFMd4r7Q7usNij9UAxEtT+zePleQ740tbW1+VmXkFfp1Cdn
hWpVFP7btvoNBVQ8hB+9Mww37HAGCVds8GCpWsn+D67gZ8+a4q6AG6xupSa3qwmM0hjz56+t0pwP
c43KehTCxvl50u054WJt1PNbiKOYVeGdG90ABbQbIIfy65DMlqqedG/6Adi+Pedra4T+buTj++j1
DqkP0EiQ25EK+BZFsOl7yzR0CYXHtuS7U/2mW1Wn5b0zBbOoTAaYRCXyrHjbQxey9lbxeSe/l50v
B50xirC10e3hUwSgFRHD6KlH8Wpi4D4jCvNyG2LQYIXyPixpi93fHfGbLrp66DJS9mUgSKQpdIJI
gfaPF4CGAnLnjqkeKaWeUqmeyKFk1ebDhBh+F4xS+Ab7uegqRnVS1gxCq+bllKmB07m3f0EkZz9n
XqiMU5xoljrd9zk2YEm2J9ajZV0LenrFdSkst7CKet/6F+71Z64gidNYA/kaYCjnNRDPyN1uwfUO
Ef0GLPjR+Z7zpH2p5UCMFuwaRqPCPnBNI+6+PXfkZ+it2ppA2WPQAihaBqeKhkDiKpbyhe4mTMtv
vWmhVPjbZzEF2mIhWfZ98UraCpeAjQe3zCn1Xntnjm60gxR87jd8bFFuR8lE8ybPSNs4amt8qjGf
Xtl9Q+HHuA9tadGa2S9xN+ZWI9SnwCLz+o3oXc/Dv+ZBqmS7K/JHeYKJbiCFwikS4lI9i9bP2HJJ
RjrAivhy57Ot93s2X7UCr3CTFvecxvqB/Me39MJ8AiWP1l2w+HJRU+HDo5m06TJeFB40xRCixiF1
iy4PMQIqDp+jzZ1ukbIexUOpNvcAKByBlSIMb9MDiShn2pPxV9v94gNTf2Z2EGRf4+/0N7qeUb+f
7BwfamVwWdEboZnRydG4OEuwn2KhBOxI6PtNEiNGm2IeVrK38XRx6F1dLsJ8fMC3dyGIFoYnztsy
7DhNO9gek6+g0z9X2Az9dlGqwbR5xc7IOCXNwhMpVLIy4iFdiZmUUwrTBuvjl2HqBZPvp5srGEdH
z/OGg+3bC6dBuDQ1DZo0EHvI3YvepWWfKPUR4h7jNcO5eUrFcFajQ9xMz9Gikj+mq/G6K6k+nOH3
zTgO/W96ijsj2Y6XGSLTNfyeEeG9DauvuEZzX0J9xYZ7q3wjBqGCP6T/zUsChrfqiTs0J6K8t4eP
mcdH9lmE1FaBFOGFHS/Mz2bI/OzfE1ThUmH6U0ioAvNdfeaQ1eAbl1JziQBJmdb3ye8TZkFqttpe
GEo9Gbp8sVWzsT9sjaAUg3qWcGgPhFDLpkXAY7/yyhFlh88v/SH/s7pqktCLDpCQhhw2PKoRs877
xLLYT9BrEfIOzwHNkSIEoh/5PHhLd3Rs/yS/+dOmYspiO3snr2ZVUWPecINW3QRjf2V5mwzH3179
h5EGDldPxeM9D0gF0YGqgukEwuy3Bw0zXcM97Uf5AxsLPH/OBo+H1K9SN4es7F5R2uEgGFPwyIJ+
rdDa7jx234QVvfgJAIFPn9sOjQOAfCkyXzcwReY02vzDhNZHtS7/wYnn0pfuVGZJO4M9qPffVJit
RqSx4OiXFftXvNAes/i/j6ofEffvbPSHzji42SGyLXp2Wfjjla72cNZGYOVFCLlxUCo9SG5TwbfE
AiZVBzgQEQ+u+2BtsYjlA7JME0iXwAq6+vs7VcuQsezxit8bj7vAcHDb82hgVMCHxUzKy+AtEwok
QMWCM+tVdm/wj/pg8PuRIbh9g+gKuJJpoQSqY7tDpFejS4DvhaPqUA7i3L8SK+hA4b+Ub8ug8muT
PIZbk528VjH9j12tAHX0XFUe0CFKUtfkefDRrCR4oll+B6fufd8G1+AwPWytl0FvwsdGd3D4v97U
CNjGGVTnPh9BLyI5Xe/Xc1APbsgFXyr1qYbB2vko3K/0DVFlbsY9CD6aWifNj6qF/pcU1iXpdsKf
McjUuHeRMZGMgIKjEutrTPZL1zDlgGD10PQ3NH1h44OISlW/OOZ9vSXGKwpZXL48GaM1MTAdoDCt
2r9EbKR5Bi1uDmb5mIADEFxCjlmiQZlU0yNGV+Iatdwdp/uBv3nzYZSF3UZAgC1KlqEkbkI5SAKn
qh8A4cVHmOXIXhba/oLf4BDDofZewtG8J9+zfsw+diutmYJzLvWl4eLj65DC0Szb2kaQoT6uR2jl
xwKGL16E1d3DQabXmuMQBJL51Qot+kA4w+pMoqcMq734zMtj/6MNolHzro+k96uXXjOUzMKZb3jb
p+W8hZXq2thEGAJSFXSA7sZmjGFk1PVounT1UWcUoMGfSW38T+k4fgldYfk05bm9hh/8iwNqQ285
0WEtWkvxAvc5MFwSenQLf09aMsfFePY4WwWbHkup8kW1RbCvewvBSA3m/WePsZ5cKJfmaNJeB1P+
P+xNfvAO5H5cFakRJ5Rrm/Wj5MBNy3rgFe7EqYTjMhOmDGZYGIqZnczJjwlSa3YldrOw9A6WtyDB
r1hwbmfh6Vf0Y0pzDjaMv9cWQKOnMK9ejoTu40UE1LgYX5vOObJGCRK6jkImyYNy7EdXS+Ow1+si
O+zTFT0NOu97Mq3rKKqs1dYBcKX5VeFAoL3Mzri+b0m+p6qeiJYGMzw9dkCnqPh8fEO/w0I4kJP9
S5I8uNGxI+/oZa3C0+he+P1zZY2+kz+WkWDu41oNLyW16xeFeOp15eoHuShlDb/Wwo/mFt2xkPit
piQltJFAOPL+y7Dd3SUD3uD1rHVfa6NOPFLW3G2yyg9qR3G/uM6u8Cv3w279Ss917gy11YvG46S3
mrDnijnx7jcbgppoC3PjEXb+IdxZ+esZs3OolYKaDFmrp3183sxda+Kn1/yQ2WntERgAKj8z5l9m
JcFzQpgF/EyzXf0oQK+KNG6SXLEiznirqJGCAuiq7XqxW3JUuIci0VOKxa9VS9X8XP9ZhCXMHjp9
s0x/VB4eT0ZmxYIkRp6oCX2M/iL5dgCnKgRkmQIijJqpErdeRj7JpdHIOwtQf1AQFAkhm5oGMpro
PNzyCY6Gre5YXHuKNJaD1Kx9S6YXPyIuAkgvpr2phbnu1v0xpesa0UKVnX57uIYcPzmyT8f81XJW
pzqFolwuAOaJvn/TzdQdyD/pFUJFfDhA/VVFMH21AythIcU9jqhj/MqW7iGlU9W8k/1Oaa6tqT/Y
LKfi/mHWNugSmL3zBPbyIR8fUJfzWwOB8yEYIxACVuknvtkiuh5bmbgQJbMyBuULBPlCJh4RMSD5
uLI+Pyc9zh1/6WBTI9re96KAUM8si7tZnX7wLchgFCKF6KVMr1TH/7tIJe2/b6ujMaObGz6IN2QS
nvkaHuo4RdwbwD2Cm9g1/NPwZPt8lw0H3PzxIOh3OqvJbFKKXEvds6U80tvwulkRDTzwvyrGYCbi
kXwJR0FNsTGECd+ad17QwvomV5wCSTzfAzJfTqTunVE1upzdwtD13GgKfx8mMJteupV1Fv3pJ+jI
WdsJjGsQABTH5f8UFHTP/mgAcJYJG628P1Bek2KpUjRh2gdT8oEX/L0Kn7ilmuMXb9a6LWadO3pF
OBewpRo53fVDILYGDC4p5svriluHEc0SzX1NorbGf0CicDACMwaDKlX4cqOrv8+7nIzYQ1a5xcGl
AsGikZ0V3Al+9sEkbNKZ3b7arAKaUufdUMRnbLURfjhK6JRZv+s3aunFpkVysp1hkCL2ntB8WSvE
KR6z91NBWXAUhSy8X0uBJ2JXuFLPubkdlXvkmX/fAYKYa982yuCmV1c0NHpAzyeuwhkelqrsBtLf
4/OzF3Aeephg4WiI8mVDFPQ0kgTaF4eJ4amZuPES0YAaEfvasXhTFO/QBSVs5j5hGXDl53+3lFeO
YmeAuYwHsYXZIJlGG8Y6XpvL1YASfLhlbWeGxqGN7qrzKJJGe4OLxH4KasH4PLEDJlAqFnETyy0u
pBA0A1bT7b7PmyOFbyHufP9yfK5Yxwa4g5yJUyqr7fkJkHX9hL+2Cbx7eV32wfZNiQuy68l/q0yT
yDLatHThgapxr/q0NLcLYURBSSaVEzkvHSdXpOI1Eiwgx3fDhKVo/5jOgutPBDYHk77hVvu0hLC/
uolU2qZRdbLrVY+h2KKfKuPy8DqPqYnVJgetlhnliJRK2/aQ5InKF2t6GIoHYV8l7X4M/bXhWEEw
z2x2wH4GKDVXZy9Ddin6OaPDI7NESoHLaRQh/zFxRFSbxczYyMYO3mdt+AH6XIyOKPAqxNJxrXKG
tR6kLbxH24dyBLSLZ/UcQLRA1WULtATt3QDQ23d3Acj1gmQWPshSUqL5vvVx0uNoid9eQ68JA2ic
gMznAFG+CE4PSIX2sMz6Yv9Si+VoCTYl/sRKlERZSfFXEw2WL/UajCJEOwqG7KTTXoVcrhWa7+Ha
pM+J/G322sHu7lb19rCHhjmrL3BgZljjLUX4b6jCB+NG5oPNrFPgz8ehJPRRkHKGXxtlUi0iELhb
dfZRaoGosnZEAIJcS0hVSTEzwxkwUvpYWgXwcj6Ly1xQuK1d7XOeJQTs4/ZE3KzJKp1OEDc9mN0v
holFm9TKATnjS5JBEDHTf93UZDMokswrjpSUkmA7FmNzxV7UvseIEvGYqsa2VhXAo9nqu+i+KVt5
JQmCtetNHRdkBk2KpKF3RFsRSltBdwlwkRmQKLUDkVVhD+kLQgxO0Ie51121dRxSfbc0NAjNziFw
78hmD2hWaBE6S8HCPhdNalEukgso/Nt0zx1MRU27ncJvf8x9eYICpZr4+38j8gQaLXBX8JeTkhRX
fQhP7/aM2kA/3s0H/0NNSfilHyPlvKEZaxhHjrPkd1jLW4nuUPYMQ2qPOzozCK5a4czx2T0ixhMM
qijHCu6bgERWa7is8gvpnrivJpkaB4gRfsnoeyQ7Q6r4Wrc5YHTVDQdPearRwLem+VnAxfElY9Vm
xrumnkkBOHjdR5mt0Z3gyjEvFdrrNoWzpfrzr5oV5RkSljvUSlCYHVYFLKPAdmtoG1DlK4ExR08l
rnTI+vKjPDUs7+kkXsqhu0rww8FUduFOxsM9R6cP0IM58BcLY95SRhd5JXEQZI6dHmfbj8pxg5Ny
Jd15nvbjwzW+1leu2YxfblfubM28IE79a0PisFxmVidKO1JLfX666DG+9wfe3Ebd4ervwCSns4cd
uOYE0izBEleeoKV7/0Q34DBev6QG8xos3pdCu8pc0BpFHG2JDWykAlWdCMwFbuTlTCg36bsdX+vs
OquDgbVXnPZoh2cGthdTnXm6kj7zqg2XHiCbIo/CLKXlRJH6t8W8/8NK+hs3DYO9/GDJUPYnEwsM
EvpnzKJyeEXBRvkMaF0ES9HW7nuj1c8lgBFmJD5WLAKEznV5AYGNQM5oujh/R8iNIDJ17so9kv7o
34y15ScoFyhg5NGYTTeSmmk3Tgct1wR7rXOb1gGOst+BW7MGOrq8V05UmTrKp8rLKXd5w+fLVeYX
96G9XUtYIFKpUqghxXzUYr2SC8CRAV5LIEg8Vx+9tHq19IM75YRAfWJSawH00KzIturckz3wDxQR
kyUpZ0AuCY4Hf6DKTC9ISxQAeOELnnyPNSzdZrZlL61dNw2aHXFb5Y52nXWTW8nG6YoiIieQnmWt
tauSyDc6aC1RjYwtI+4VZy84CRcburBiYx3OuK8MTY4BYgEC+ny3ZNMGStXV8Ra7Ffp0rwXVp8CZ
ytHgj6qqzebfM4mqgPnbl9TDPWnhZNuW0lgK5N1jG1b6rv+pwFMqGhlK++JQLi/7mN61onePRj2V
FcBO5HV6zmgNCCVC80doCJGaCiyiDJKnP7O+bgcuvH7eaEJDUDdRYR8l6cWrEml+62vMvHQS8fQo
k1cKNCGqMhdaJX8U7FiiwZQcJux+syQaXbPMRPv8NfUjNAcNhz4IP1ht7pxCw2DFkXzOqOYdhNUy
lJqY3N8vrg0hxO748jlDlll6DgMruLa1mJmr2vUaev1H5zF3pNyMMCUwgw7k4iXubqIZYuOV8QMB
b/hjO/HIOWdyQg3HTHD1+VHYgUJZnx+SZEOxZXQ9TFyoSWk/8fVxUQPNAyZQZN57AKr3l/DgtOmQ
URpcmtvCwxavi56OuQaFoOBX7pPzLkwWX+I2lZqIlkFEGJ5NnUzvT3/5rnRFKE6qEIWTe5SSZYD3
kGT+M8n6LUe0aDyvLfbR/Ha0rno5/UaC8WVQKSd6pk+ByRWl3nJqIzBnVQKbdW2STMKLypamrwVr
ll+nefTjIu/nXujjwkxHn+N236DLThgwcdHbutv0+G7x1uKJjZCpbatDfva1i93dwPWra7/LzArM
RTmVgLt2rXbP4RwN8XUhABuponCrvJyZpebd/6aOLY3khEI/HvO6tk2qK5ma+Xn0sFddntuhGWWd
3OvCC+FxELt0Dns1Lh7FsFO5wluRBCHJ2jE7ZaU/9Z4OuDl6NvK8rZtGaAAF+6SkCP0c/aXcTewc
hmGI4p4YGEp/AQHCdfpvPwekW9So6hsWqrNGujx83F/h+Oxp5tdIVzSfqVZjNy2CPRcHBOi+eW+J
fQx6WOBLP/z4qjxRM08y6JTyR2HwgK0I28BKPmCnzDZoNFLZa3PEFfCviMYl6MzmirhUiXj7Y1Hz
nWQESlrCS8fsW0/sOs4U4NdhdJZBRtzPuDJAtF7Qk3HaWPOPg2l5JhbYbU4RdSJhsNaRXwfgR8Mm
Jmrja6oArOQyPBU1CmzBn1ErRQeV8zQ2+9E+jm9/10qC81WM/O5cxO5evAnuSFZTx7s3E3w61mqt
6vRAJ9KEOPVlEMEwuFCEj0o21uge4P4qGHgsstjyIMbvTRSJ6s1kb6YHJSd69h8BLw82CJIpgcp4
3FYmN8QONpePTlain3AyMgFCpklxJK0SsQRizIxyfQiy9Kf5A5FgrMk8uxLFGR7xL9GAZ84hfthW
Yy5F7BBCxJTFJALMUh1jnlSZyvmXHTjEzAIDt6ORziyHuZ2+LOq4HsnCanQBRg344UoiNC7dOWd4
ZlD8T9aCf+h7Ztj70sdc9LqNJ5wh5lwoz3jSWH/0Ja42yqUJjAnebJEfRIBw/fbLaHR8DmyQHVF3
mSHPsoaeI15/Q/ghbHQMDk3kRYLmWJSypvIpswB11UQ1949yZr94SBkff0hQch0w7crmC3Kh6tKc
+xAEOuoolgYeaRKJUkeifh/D3OldiCzrwJNFAx8isFew2hZMej65M3wS6t3j08KPJzOYLXlqeAGT
dHZsh3VPzCGnASjI5FuWsCA4Lb2akFTzPYVhLHHMpMCOrs1lYl6EsRBEw0O9mabO/7+O2NdSvMca
LPt2sv5njUm4lkUo7hL8bqlZEl27w3QLdlmrgoJ9Z4lUZktXuvT+hQKs7W9JsF/JcRPygEeflLBo
MMDFSoLZUqzqEOCEk1LfSUB8ZQbEI5+oNA2c+P6QYLg8VbtJlPBDE4M0PjDdlWT1Wnrqn11itK4w
pSxpMpFEtOBJVsggWftfvEBKqunDRPezFNnydveF0orkH+n/1AaDcLMWXLkFU1qDBet+29H52pdd
FI4QPbOvyyx5HJn523K0vazo/AbqYj3jTX3UYov8+TsoWO0btR0SuJLhCLlHS68sEKur8KrPInO/
6ENV9DU3lT0wwiIrKZtdEN58DEHB2B55TOT+Ru4C8gMTIE7Q3af27vh5qRqggVcnkqzDo64iYX7J
aAhLN7ns9JgfzLJK1/HpE04QToyJ7QkHmZjreTAPD5hiOZ06CXoC4ug5GgU9ZhkJM167dFhc0g5J
RzeI2ixT02BsvAyKi5MJbDl95Mg0NmnFAYU8lwinR6ST5Aag01d6adneBfLvh+UotMEd0+iWjAvh
6EdK6feTkPyg3IjdkW4bmV6VFEzlMfarVX7EdfJWj7VFZZ2TfF2uMNLa4dpHwmffUesVIO6K3dbS
9bfSF5hnq2poEyACYlXfufFiE45UF9CUXtqplXRPkt6gQyGMUt92usJgQvXpfbyjjFv29xK8FiNJ
lvnUKcw7hJexe1fkiP7+VQ5lKRwjkbQ03kGYRULk7Se5O/8UU/5i654Eoj3C2zo5sQ1G+IgKTZkX
XhoWga3k7hRdKfRtga86s1wx8aTxwLY+cOE4NkLa6NOBx+ltfKNgo7r0QiN4rIqamyPkunflpnUz
Ic2LBXxOVDKhjac/eeiTp65UP5zDJEpBR1OokYAynVwKSAXDE1NK7XmSG7iOF84C53YY4H3vS53+
aMYFgX18oyebmEdO+dQ0iKlgmpIo9QpEex4MkSDDctPDdRs649pOGrnEq7qCFLNteh3+LI2iGG/n
h3Io0C8CyilGsbyOYUFpUAPdxa/XwATIsbMqAN+7yX92E5UDtfegwizy3dk7+vSZi+nXf/XgMZUI
IfDEh5ZDQq3j84g1utxrL/fP2TCfzvfNAeVGluBD4hExjTz3LA9LYDfihVEUqCuLZX1KG3AD2Ri8
H12dbkLPBSQEXplGXwtJj9iehFTEZo1THcgwUIiRAeajie9dAQJabasEkd5XdVmcP+RoYNagIqVg
avviNNUMLvJFepgfZ6ARkQo7T/ubiuObgJVoDJ+ZyhBAvN76K2D+TNprXWQ3JCH2Mto1tZ3G6LeZ
Sw4wQrxARqufY2aYrmMQh69VOiu0SKzTvmUGRJ9/flZUJ8g/3XlVIEuVKGcyCydPQVJCUQ74DKTV
FeqK2/vz2B5LSvCLjyi3B7ub/ni703d9+lcRGjoVRjBGYueRLieuc3dnG1RJ1DNnels5mS/lvQwC
Ts7q88Gu2p8qvthyIrNp6E3gebrMreRcbkHZ68U6qCzVac5598PdCNmACyIKZLurUHni8hkr3KGD
PyWrKvXpAHUpUj8DlaBJ3OCTEPZBI4esj5SwI/wdHUkbjXG5QpK78139ACQv7d09Wo5y2ThZ4OZr
uSUyJ/m1vvXDbMIUd5HseoMHJlbTx8FjJIuFoxWinlkza2RI0+r0c4FJBzPQPGPJxZnG4fweDZhe
vhx840kJo+S1ndIBAT9gq90TLt/bCl/OydYQGsxGqfdYC1KC6OSVxeetCm1o2v/EZWhCXgCHQtWm
RMj5YA9/FgQJxd1cc7iWyNjXhCKkc5jhUjDHnYfKQSvAaMij6ijJooZvdmw/yzTVgRfhDE3I4M68
Y4H1M9FsCazW7dZTyONPWYn1CVi8DjtFa8yhHhq0YK+rVDytV228TQ+y35bvA7rWBXK4dUoh7Jcu
j2ylF7g8BcazHJ8EP1+GsjXlAYXtYtp48TNdDUHw9UHuBYbxyIAfqL4Au2mrr6bPx/OCRq0TAYCQ
prqccYhj80Y1KuecD2FOzV2wEBK1ubMT1XPGiPIIVrkhdeD3VCEgvsIiQmGGyrNoBI8Gge1lWztB
1SsfhFE7qtyigLXy50naoWv999pUl4UFJNZ85PHl7a6+0UFhytuIN2HnRJ0uHZFift38vGoTxsZh
5gea51ueKhGVKHFeGisNb3K+4hYTB39COTacxBluiG4YmhmYFuqXytqSq4hOYfGE9uynDjK9PsVT
svJLCKBLig+opJVNi6UIjqhy4LcRQelRr51HodKtZnDGWy0muXeW4a0U4QEIDxT4uCvYO65tp1ck
b0pW2nPJUbI7IfR6UaxtNz8kMfkSesecLObmc9ypKvFFSXWrFI5f+RGY9iH72pv/LEWNTdT0uoX6
pgjZ97COeQ0B9ZDhNh8zYGUdtDkCqg/ERV/6y3xRVScoF3NP38Q/pYZ3ndhBeSbByl97XomP/0F1
LHQwtizSIGqvnD/G+QRCUMf2pbtHU4PIE9QalKXsIasfFtYRXbfd3mVgRa3cSGdRTU5R+/SvbURm
0aYXKkflR/ev/DuOvhfPalpEkipKhpcyUEDRYBg5bWqBWbjEMlMXhebojaTJ4IL5tYU4cRKBVtna
Q/aviQjEOU/g2RC9tqx3HVixyfaFS9hQkoEvMEoaenqePhUDhoxVrxWK+UEn4pv5DHT3I56uk3E4
YdT2tdK4YYQ6gC6p7bfc8gEJpwtPACUnS00Gf2ouSHhvv1r/+7+hdVwfvGiuvjAEhiupEdwETx7C
DLW4eyQjYJekpM5Y5uLZW86M1FrHwxNSfQgXXei1avUYiZMrJUN+6eganQRYtLlNHJj6jxf2TkNF
0GyC4KUjVDDGVI03TP3otsqXcR3ulwXeb/Qa+8MO0xH+DUGO2GnOh9LfQEnYtxpsscFlNU8xnZOr
Tuw029GkFkHxKLYWnYomA8hAl8itCZo0rwrKcTKmXhb27rNcA8jHQIpQSF0ZXkGXUsbeWC2iwC5i
m+6ZrcqxqETb3oC8UNYvD6/3JRxmaedmmOfXcx0zSEZusNKuvs7nkLP+EhYzfkAddrG8c/vLMmZv
oz7+03Km8S1m9iFQ4HLMdUV4di0oS+LELeSkfiSaLUhHoUkPm+J7prVAwBV4sGE5ue+6vpFkvzyZ
Je4PjnsEddWsGSkTZgc8JNR0l9vZuQqv4TYpJ/5M5z4ZJHXPZt5dYpRk0gCrV+5LLE8mz78yKT+f
f72jvuK73e3m4AUiAXyJflTHwACWbEfF0gBGcWjZHWg7LUJYlJ0xIihBv5u8b4eLYf1TLFExJh1/
Nb9eb1LaoqsJiXcIrQYaz46k8mUd3RbkT2s+ffuGybIHiVJ5pk5BzLqde33yE/DvwkxHoDNtQPkZ
nV1MZv5YqrzShM7SfI19whtewOvBkklXshjcxGJw5+m0U4ZIgRIPtD5PtdJaw9vMVJPOUkXzJoi0
gWOrPsPVvSP+0m7cSJGHvDyidP2YhwGjTBVS9y7QCafLTUwDK46bw8f9rECR2RY/6Zq+DMZwaCej
XVgmbm1ITUg2TN5EwF41fCEmAm7zUYZY7t5hd9LmvwK+LuBxTpGi41SU9nYKnACUPZq+plor4A/e
r7daYatUjQhAaBfJxIpXwNQIArA2JBoil7/a4nnudwkbQSdmxbUVTVQdF7MWTAn1cZKp+5nwwY93
2l/rRZ+gcgHl2FwB60pca3rulVcBBL/6K3tXDwKlB9rCXpFz8qqN2JAo+8NK65kNMv3lKA8+z/vP
fEhy9IByE7ZvnVE1NZGyQ4HVzGP4STfhSsg0SIZCzfzyE78iXP485Abr56eNXy8WD8aKDeUiEWLO
LE+5Auw2PevPyZ2g/555gNcij1JUlEMdYL5XcJeneuXjQzc2JbWxvE6IHQ37m63cXftlxx/v+9rz
BDnsZ4OevS+AoHGemT0QPc1gHCYW/fS6KOQvLlk1jZ04vtul8GBOrPJnqfr/1xJug3+sb53wtvjA
UxbwikgYA0Rbv6B1G1P9DzPFyuWe3fRw2YPKGlVcQHUXUJ5g7YBiKbe7DyrvN3nTbs+xqIJTLz3p
PJSkCchVdRDUpEXi+2S9PgWEL/+CSZGXSQZhfurJVU+TupAuYJlt+qrQeWxMPWVqMIwXA0rLhj3P
EVmorzqTIQhPMFj7/8JEqZLLfMZnYzwSKHv3HdX/N1+OHccYOIjk7YIGb27DdUA8Hs36Ape5ZXEQ
e9i1qHMJQLd6Xq4aanLbhdO5dpGC/e5DgVHspKu3VLVoS6VvokdzpYK4/AydzWSilN3cxh5cmdoD
W9kbOJotS1JH9LhzANUmcQpOcdLc7i39+DT2sqnFotdO/vwZpcDfaZ8mK9cLDJO6yQprRCI78w84
QyoVRGThv0s0A5qQEbW1LZO1BgD4GoaVsdJD2zjvMvvAWSeuFyglxyyLi+r2yQLXUHYrWzuvjJnK
2rmPJ4LVkFGuj/WwqmZiZYfupdSUOwNWFC8TUzyngq61C2A1j6uqIu7QgOP2kQbkqentaWlGXeHV
1CFtaPjCdQ6HetGaOeEJi10uR+0GDwRb8H0GB5rsz3ZFcv0WTvWeD0sFcCKEAIcRLq1YLCpfZ5e9
DovDZEULw4ZdnXcnnu6CmYehZFG/6Wcot2x3HSCcgzslSPHJ8vWuGiamdJtpsYURDsDGAQcc7xoi
Wi57PyKMh3oNYIIT5WDg4bWvzvOxYw3Tibi170ZSR6BQZLrz+ZxgpTLzO63pNzfzILOi6wLBRWIb
QXo29Osihdi3nzryXqEIIwotLQnfVkbQZ0FAkow6+JSPZK+zSgdFZtdwm4+3JnwN86Wqt7Fb4B8+
oY535BVVMw5UBZh1HEAZ1NhrBSK2YuLEW37R1esbwTpDtQFH+QQvC8I6rn2dHq0TsGqPioLkGYXP
dQEHH642EOo++fgbtSCULAitgEKn9siuObCS5Rqo14x3D2Rw18Edl4DBo1YsuKc1STw1SkRnYGSD
wE56j0FOoPQDKzcvk1gEqmgF3giiycQpEgX3rp+9iiwQJbRbCe+d3cpjmkg/vsy3/o+7dO0IUzyU
ndVgwjBuPe/GGLWg2JGlpJXwnGsXoCZJb1eY87wjM7RwfErbHmqMZlExdRW4BTspzupHBHLbxFVG
s2unUMlJ2298uDP1ZnAptXuHcvxHLQlKeyv7+UL3CRbvqj2dExEoGArtrLNzC7CZKKT867kaIvmM
NUDId/PCQG+tXRxatYp8xzFe1bsscTB/IAM+2ux0m/HRemPjvqyCcLYXXiZfvWcNh4qvk7bJ6VEF
VuNvmGgKRsbbiw3d5Kzy8tuZa9AiPfYNfqttP6C7s9KEAKI8NCQrbx1J/LTZlYogAIo0HnfyT5BI
XKiZNqY3ExslTrsfqn9m/G+1EFrPEZzaZGWdm1OUdzmNXEpz9dD3hJteHS2k6glD3DdjqpHH9Xal
nSSitMBXkx3qpjjNHiqwZi6zE/uJi+YpT3wrhFQI6DpuGRhfHIOD4S3BtITMJ7871tfgL0PCA+NV
KALhBXQeF7f1Mt8EjH/OitkBf7jSsb6gDxNWiC3DyECudlEHA3CgHKdQm+/iOo7vfbKSKqpsuBFE
VANcOU9PLVw938y3eQJ1ivKb+FhAtF3rRjcinvOWiutjVjjryLIfe+eMkr97eX6RECyWuULBl+A4
VtIcMJ5/a6fVNP3mWfxAUcpv32Pe9XVCPiB89wPQrkED073THa8CebJBbpeYgiwiCor27lFk5eFQ
l7NWNd0hK4LND6nr/9Urs02P0gECd6zLEfq5YMJ6m1WL6eX0L+xJrT954n2rs18ZvsSJV1IsZhaa
UssF0u/ekireOJLBx9TXoN++++FZwhHHbOXLFj15D9TG0ajXihJiBFkv7pfH8vpb3z4vIJ6tY87f
Ct629uhg7v9Z0SPch7s+KiNixsWV+/vZ/divbyNhGz2JQN9MwrfPuU7A6OkKqwskdeDFgrkqCbcG
bqHDrchaE+BslU1HtbOu1ghyRlintWEhsUuCEfwTKcH+4QbB65oTEITP9b0Pt20B8tbXWCh3SJGB
9HORpumvRi9G8iPtJ+Pol+R+wQggEGSwolV8O+yxSyF7lxqb8/ycaxUdY8N7EHqtYHOLVwk+k2T6
2zi9igXwyZKgORHSCsigiiOkro+nKoqmJQBitMT8BfZwyCsNc1IWhuNA7X+3o3Dnsog3JSlOElN5
EQ11qw2xgLbXM7WClaNtP1pqCiNfir3DTJt4oBP2ec0Eod5tf/LbTJgI0ajELKOyu9HnI0+kYf36
nnOQbh3p+15mR8Q9YwhB6t6YnKPIJe0/kuVNGHoLgCKn9toMZAYDTRlPIXmTrngfRfq0DDsAs6nC
iFCqVpJ9JME+JFXAW5a31pQ6WPQoWZMzcXcvlGLhaBuh9dL35bZKQQTmTw8+J4GIMxbNqxGO4VDZ
+Rfy24j2jM9USZVAS7xKJda3LHRsXbhvcDSe2vGmqKOHpHYp/aMABM9DtFnz7nejSQUq5eAt09Zn
nt8bvrL19qKGXE9oeM4Wm4Br6yqxfZb/9Y9RfYmraFdFA4e3EBElCjP/yIT6cmZLuFMmTBH+DBA3
+yGdxAyQhhoW8aFbJixLJRBjf6sYwDAZgR2dDQUTkgo0YuT66QTyO3fmcXhxW9MDCQF38iX6N25L
RhQltuMT6DF0bRG2ya4Uvgzh70U1ZoXk3hPLLt+w91ebVflNmLUqwaFlpo29/6HDYR72g0M8rdDA
jM2xT1HWR91kosdwrE8YaWBmNbI90jU2htqC60OJRfsCkBPuI/n74StMwiyDFE2RPLMX0SIUBNRE
fLUMwGO4WRullAj0GKNIeXHM1Sub1LXMqi2WF3EeMYK6LQ7gboONVX+q/6SKyW1iuIwUNnhz1ZbT
uYzUdp1qxhStlHb99+NJWKN1U/p/ncUJI0/JWeDG5ZQOEAdY+kyNP7tFaIyBOBC2omXjMWhyd6cd
v4WfKHGmbTAVs2HTDK9VdVTExO5Ix+iDMi8NcqNYz2lIPbjGk9GgkOA/292JPcW0SGJBA4MbTUDl
Gg1pD0xF5mnX7Tvsb03U+HKJrCNfBY2qcIwABDoV65DGFvfdDjgfBfg8F5p8tbkrQujw/2boePrQ
WHM7AXZBTeYMn91Kip/WeIK6yrVsM0AnA1QdEkhNUnH8UG+YJDLXR7oebYIKQYYSaUxpGyqk9oBE
wY3odO2EVoHDVssKEpGMAQuSynvCZpzMNPT+NVjDbzBuadKUwJiz4cEASkxzNsIs3sFfyuT9xeiU
anPN/FZ421x8/4Uv7lUfneant04XE3knTkZXFUzKcrgh+vagy5X8FhpLc0nYjmeuxLiZcVxkqbMS
5QgwlOFpnNFDKktjopUVRjex6Nch0na3vmWmM5NB0zYQWVybWRWmZUlKe+KbpvqCEMwtXiMj/eBt
izb6PPLHl8LW57FjRZLGSPOGu2YUP09ohHq+Yd8g/1zhd0o5Br5sbDjTOdzVSjg2YPU/EH1IpmSg
2YrpdREUxT6B7kWCoeuxSi2SkEgR1S2kWZPEGC8LpX7pokeePsbEuxJW77q1hl762xzjBQcI5d5M
8vM98FUC8+ototUlRtLjpVCzD42qXfuhydZVpDVEultvLWXZ+oeIQY7xqNEi4qv2T2dMdUgilvie
9s64M6SA6k7TJ2sxx0Dr2Akm1FHlQFyR18GhzhXIK9gx783SfbB5duTsWRlVFI6sfUkw3ZODc1E5
g7El1knmEZtxK6XBngYvW6At6fPDQlVLKBZd/p3ps55HUdQRxglxZpUvhnKHbtAEeXc878mE1CvX
HWNo2KmLD2LQ3bCZ9sSDZpnPHo7kSd07WqqfF6yUdGToTtwqH9RlYSCAedKu19Moc/swQMSeTi/Z
WIwqgTaoEGaGLvpoFk/F2IxhHgipFnh9RMJMWZXrk9W107V4QDi03Es05A9Bb/G7HnfwF7GoebhJ
WzCqTd4CBlpdjsATgNteCdRGh1uczTW0kYRQXNyIHsoDbCjf+99MAiZH+CjvN2eeCMj867EVX4oC
zoS3PIythEwjrXXFe3UroegO9z5L1Nvi8tokvD2DNbX/LdMB9T0pWzxpAImGsru9q7f1UlYaPgg8
45aXIcyk6n3SMegs2fl6vBgsk61GMnq9PpP7PV9nI0TnWHKd9SnTiMqbhJraHWO9tH7vRCBQ2bMj
xrh0H2PrWKNrwocO0g6r0hGgblEsKcstIkYVXqTd6Ro7EUNNSZk2iFbZ4UTyWEbv8js1kMapBOUF
n5mH8Y6RLB+0ejKtBAVV2kze8pMUaFglvXQ2ZJ5wWlFXtYK2DbSUpY1FoIx5MtyDmBte7/WYGIMV
PpS2dq8EZvDOvWJUt31R+0yzJBfGWkc+Qct5PMWGgFamnahqVaIaDEpXD6k1trMa0IdX4+Im1oCq
OK7pKXElWb/0x3ZEsNc344juuN6ozuC2mKdkk6z5d76haZ+Ow3LBupqlFVzBf0ZzEStcUUr6fyZt
r08dKiW3Y5r54c6SwVEvRpbJyc1dBYZJLo1yIPlxJSSnERE1aX8eHaBwTILgtS45RPVsozHg+PWq
Dhomf45XfZ3e/JHYX//zuQrs1X9JAGkfee7iMeIpwEKzBXny4sk+9vJ/5YryCOcc3IInGj8qNEuW
VGSpKpkOHtR4vIeCz2WBaBl1kktSWPjW536lnnPsLRQVwi2nYo9/f//17uP99oB+1md5e+TbVU9M
AU51UJVrG4Ca8fzwQJIe6ITCGS/BUhM+Ovviq9lwDPafMokuRYF12yd+igpStIsaUYfI5BIHK2gM
jH5b4/dFgM4c4Hr/ooOomxn0Vgp08g9AJrVY2dtS6oaaMfTBZ51DJG7fzWETG7sXuhElvYtWJFBX
/w30JvT4ZqAqEy96xdRt8xvQ24tE7daUWWQZWLUMwqKcJ4pnkw1hadQ6tEzIASq9PY8+qVeOAx88
fS8N3BL3jpDjbgl5uVsSmBdSQ7a7PA28VU8wvnUAbYIWyJ7d9TQPmqM5VaiNvxcLsU744w9QhjZj
oszeNXNZWiYATrLrMf4IGT+31C6y7EE1h/QC/YrrIEEmTKv5YDZBlDYnesU+HkkRw2xABqlJHeDV
KpHeh4kqkUt2h6mvH2eJmM7CxP4PvecT/fJh62UhJqam/59HJB/jgVid/DN4R13u75fweTu9BdLk
HzoXznmb/iPg9/EoV/x2wJEHQfy3s5qbbwRCez27uSwL11mFlfzDO1Ustnxvs29b9ckssGOsvnkZ
bHVNRenc30YamhdqMMcBFCgWxReRxFPqn60420DHYdKNiLXG2CqsRo5xO2zFOJakpuwgt7iWgL8m
rHNcTrOaB+/fD9Fxk+4eO47b7xUvFcuviybDCtnuhoP40Hfh7wRYaynzVd8VgKNUzKQM6h5jMy8M
4V2bAUauZpQN2vY14+65aJ6zrF7ZPOPNYwTTmimUBM1ZSCNuObev2I0YOv4O5InRTbyiTlHd37SO
x7vWrc8X/O6IbQRbKQq4Nqyn/v3weA8s3+nZEC5oDZmQcIMpPmyMoQ9yYNGL2Ja86FJqX+Qh0/Tg
sBgGs+EQVOxwWiefuPKoGVDFOXj09tSmx4K6TEpmIs+2MVOScqPGBtNh4In1ROVCF87/z9JTvFw3
dop1jLkndA6Vf6O+kxSfitFyxcnPDuV80v76gZiFzVuV8Gj/UgOzMfJ/1roQfLthygkBz1eer3L9
MTSLRn0gP8XUfzpafMxRvqdMz4y4MMqNNC7i7bc2XiR9usyIephDjScbG7xlW67hKNmdlENzrj5m
cErmM/yabcc45+5NEs6926nVRKCko7Xo6dQIrcXscHEgXsKSoyGCvC4V6zeTC20MWxWOrVUn63fJ
14MMyQ5aOJfDRZYx0SZGqdWIwaQ3S4JyaCjUfygaWEf9010aLsRZwyDD+MBLoxF1ZVlHWcTY+qX/
ouYaDVr3BB1CTZFPkaPCjGHzdOJn+kJWg62Z4DNNq2G9Vj6UZ0ZSyNsQveHqZ+J5XWqsTTF4Q6SX
0nPGUvHpRvdjVej3m1nCTUFz9330z8o4/NMcr0z2aYV3uMtHcFt7vj5nxtraZdpgJ3U0c7Ji3rn2
6U8Q9u6NHiYohSB5oDAaOR96G3ZO1OMhLgMh1C6a5IFetmJA0vweDOfog0CRJ3L8+uL3oFiXnacS
zwwgHiriFDUDCyTJCScXjfFUyhE7hKYvcacgvfwyQM1GtJbq/s34cH+EO5zL+r3yfj0LDJBNhG8Y
ThfKX0JmAyHhk3F4ZRV9RJiM0IbMKZ/zZPDMf/QOlGp91QnA1VyQnDa8OieToRoP0j/UeYSSlgWt
VtZ75QdleFh6RkD6VA6BQ/AYg0Q4wILs/8+4IxbYvYrK9kCLNimuuRBHh4U3DGoRLIpobpGZUjyL
r0GSMjy1onSx7lPhaFt5JBxBZm8ru/VwJvjNz0oaXlLHZ9i+IaqjRvtox4i6TJp3T+GHZZrwZEG0
xjkXCET6sYvgOjA3gzF+qreINNEIEYpap0EGFkoC5z0LJSylK+ORuZliBaR0LIm0zEpR2CsJuu8t
i5Gg5dot2klLoqbZClZpfpcIAv4cVB/sMuMEaiACc5BwJ959nyWXYS2ckhaczq3Gcq2/XBBcuVK9
KCALDCpK2ntKWxt9EV7rFuOKfHMsX9x0nyKceoZ8CtC2OzPoScQLb2YOZvepvs5eEVWqtl1b9okK
NHt7ylPLrIdhLVkNK0UscxNeU/3NcU3vN32kavPWvKD8Bj2mkF6lOpboara0nQy/FM5NwMo6pijX
mBPma+y3EsUOiHSjPV2gh8cqqpGAfndMF1jXpHEbcbwar6AXlkQLQSLu4GzsESZ/SIafHNpF6cS3
bofY4CnI/NuhdCNb16FsgAdaht5xc3FjZ8HH4woGF/RxxGDF+yudiUltvFLBKAvwl11TedRjAlxF
b7g6qQ+io6tQJqb8UgGG3/c44WDuUgQlccw6Cz8g0yVPKDhbrPTMJyuprqDU4sRTg4pG0fDt8aOA
OhPMzvLmAGpR+iwtnUPF6mJNS+RY9oE4u54R8U2FF28xF/9i/0zNS5Qksog5R1fkXSSC4vAeT1/z
t9gvjrYiB5kISCkHvScxXS6lvPQapqPdD1Vgc3+qTAUTKOVufmR8zzx3NLjMuoXtc7fgeOg0Flr0
QLcZUyxSTlm1algbxao/CSXWzZLKRRrBgdIQT/WDhnguSievgD/I8tE5KBtwIcVbVVU5I2nkJWZi
regkZtthtqnTNjbcXDTrlqgMdOrIjdsydNma642ZaZ/XDiaIMm68MzdO9QQlMQMpdlCCEjOTE4uD
f2QMIFldYTxoCumaiTndS/Cl3nXOkbt+Xzym/E37aVIL/xWds1k+dzlZxX87tZEYPcgK/KUHA+U5
tdeOYrDi6rmhbv07MT/b8m1oeS1Jq/Y1/OGspzA3l1oD8hYuZGxR826v3SjTKdx30ta8iXq9yR2U
DRvWWqt7btTcUy3ELYAHxly4dsK0memw0WY8GFeKCSCPWJMUPrQmHIprlsvUDekKYnhM+mIimwFT
90OYodJJGXbMDP0h9s23NieRWysijgl/xFGqgTGVhmp7GnXqVcxNgm38xsO+g3hdUn0BJiMHenhT
W+N/sJAhoBxMngBnD9uB3jsSt1VoLsSQhafdeq3BjAq6M7K9uN9EAMYUupxHOo/iMnA0OU960eav
cFrmO6D44odFt8VsL+jK6yhKcfBnjiPVK2xuAmOaF1dAQwvucVYa3Muu8NPz0Noq5+vgAdYd5ozq
rogHmZi5he/usFTkoS1q66SMDi9MnogomO6uALmrB3g5SU2oBG5h1/lL/pWOjS8YsOj28mLHbQBo
UVi+xdMdhErFCXCw7OEV15vQ9ZaTCJOLOCnMLICfXC+hTEC06TvLoVWMKdeMdrMcj4/WYKPvP15O
LT98ehC1B0nKqGnj0pU39VT5RBbtv7Wl6l2qThYepeFkaU8SkGjbY54hUiiI6gmfJqm380IJeA+n
NO6juFb+kh2VVB+OR94F3nkykUn7LasMz+CAy34ZrqxJwFtMFtbYR9Sycp+Bi0YclLcBaQRLEUnL
1ZDUo+HYiORaIopnrRYg8Ivpwy3BNA/+SI1vxSr8EoTDfY3EFRGJuHafhoZ/lDv/dSM+n+YJAlc7
6AYtWwoEhmTmPrBxJsb1wt5sBJp+7ue/nVcJdvdiKS/a6akr9gDdutbAq0ffJn6YeQcorAwcR3Zv
pqSsjto8ZhJlfU1urU+sfu1ybay8igyxNItNShgY9DavcIL1Pf+TD5qKPX32whvvb2NXHzGv5rGr
o0lxBFGt4+jyxKz8EG5gFHJua6vTOvQH7ihqr71y1MvIfl/WRiuj6fO4GNykqHyegpK+jxRNVAWN
msnTkvjDAQ20RSKhqivNile3TiPKja6mdJnJBLo4Ofhxm1fjb6kUjD5OAxN2TTJTFd+WYdr6cVzP
BobydOYoW45TijMBNamGcFEwbbpQlFp0cNpzxdfx2GxmgpMcllFh7vOxcl9NMIh3QtpqXXvYKYLq
IlPQG46e6Ej/efbHQxChdM1lRy/0gtcL0LFEtM+dXCXJ1Te30o9613Y77iCETPvbvyOG4PnT61ga
L6MFkSHgygXNYjt1fh4TyS6xe819ssIBfLh3PEJLQKfV3pR7dQh/CT8ztGkU+G7beramrjU+QzgM
kZvGR2TMB5e2ZqrsCZSjTjulWtoRc7noHcO59OxBJYWYPwwB3cqkTzdZmZZzFVMX5bdJhVY+JGNe
OpZtuCQC0pE5N/+wJ2KHutb/s58bqy6eywyh8ESGYkZTPOKr1DRlX8jJcCEN1PXpvs7BHcS1NkiO
JLq/Nd+3dFwIS4JGwtRQnOjPwgE3nz05KQdxg1GynzYFtzlV0WASJPGFGtf5KJOJ3JQA4tUKPUl1
Y3IWzjphgyyv+JI7o+Xp0y5XLhq0HQ8hNe/cK5gzbq8FvELFy2riM8ZcS6yQZaSM3+nUPRfRNMre
a/jFRmh80h2BoH3wfeXx7luRusQA9lC7h9ObwmdP1ye8FzMBlPqd2H/5Jfq3WZnfGdq3pGwLCQXI
QZ8+Sg4D/phCS6zUQxFYLKfyB/8KYV19tNBRxeSmWdD5SXjQNMVVwq6kQeKMbXsXRJDMmwkE5dHo
Dkw4XGLc642f1WyQv+jNoLe+kRais93QQkhplQBhLt9994yReOt/EnKdLKk7f6BVR1vk39E5SFcv
D39/U/4LrxHLzBLBKRSILrxsS/AGSHtPt3F6VxuipRIG4+/M1akdMQ2A4JIxnX9uUxYmtcj/J/xt
LTCOBsedRBxFwimcSAz6H7e4Dkf4c6jGQMi2j5Nrf6nrvLjL8mFQk5kAnKuMNDg2wJ169CkdRVkw
VstgjvaeLz7Jll3XFlmMFltedeTA6JMUYemLrcqr5D/sIdN56cR/x3LSN9PiVOKyLvKxtBLAgO2u
MdMiq9AXU5cBoG+Dgrox2EvHzrYyxMKDvR2/QiflF+gtNaR3AgSGEiYnAejT7NWJr4iNcCvfUh84
2PJ+CVKWXKwhMdn9GOrQls+FxFTONZbT7X121UgACwQfmxKbfI4hPGFMkpP+afU3f8lAnSZQAfJc
jFopykWtBK9+xOZyD5DphEWr0moIERumqWZRfBGXnXBG+QUG9CmDiOPQw75bm+h2jzLfBUSgj6ca
L/wvToisGbFU7qlu0XMNnoravlX2jAAYdYd+8CMEIIHcfuEHjAjV5JUeJKq6z/yqnYULhxlFI32+
TKyGc1fo8rnEwqh3NS0tEstdIgXQwLnPjV5iywxGXPHaGbUl+OheVCNi0oZnlxaPa4yA9bDAfwa+
dH62ZU6wkiUdhoPpoYXhQFb/4exaN9hNVHzgmDM0luYEq/xivqs6khPVBHYRG6DBmkVV0MoNtuzt
HH54AuvcLWck1nIdk1pHB563SSqjOyuayXJv7Cxw1fjB+TMPZFVazvJqn+QYVKPtxVgjCYixn4Dh
AXh+SK8Kn+DfwBntTUMr9eUC0wqDPCTtt4n+oeYwpP47XG7Aece4Z0pRm+nQNyjeEDzsaNqqscPP
4MwZyusve1aJPLJiGp1goSQUR20knl4advacQg9PDBCas8tkviLVnfcJVninAXQMl1dOaZ9l5RuP
9F3V9nEfc2p2Ir6vCNc+IYW1WSRU3iwEtpSNK+iSNbVp75m+PUA14ScV7cSxcf2LFjydBnRW0Np7
BIdUVQUQxJz7MNRlvyMwk6AKb5evevLqu87KPFKG+ggLQ8WtDAjsn+z2PRrBTBIxCPDPwV2Nqwow
+HEQAKxzJ2Oe7jx64W7q8C3jKGkq/3PG3f1VXnBMPlxnSINzcOSKw6Jb0F3uqPMNDL58eGYt+gJk
s2fhhLBeAW0lT8cqApbT8JquU4t6vPtYn8lCCVJ+1BeK9AI/zCAZjIiyLJR45LDUwDtSAfv+OYKg
+BI6veQT8kpzG8s58cF31CpUZAYz+r3cIdGQRq7uUYcjKTd7DfDpHZpgiVWEs0m7NFDrZHpFBt3L
JcpCQC1kRJXhatPEyU2rIrBk1CWLvKnuB3fZ8Ooju8ml6gJQoG+u4f7JvjeJK+nkVhzo7Nb/xM9e
OqRq9rTUpmdhzyTLoBJijvtuw+mi7hh+JIes7ycBAVUXlT8My2THIoaSWS5bkE8swbD/KbKFC/1G
N4PFTqjNpZ74sL+JF9W5y88jRW1bmb/jJtcdFTMPdVamVaIeUIrEY/w/InBZdqNyz0SRlkmCMxqI
RXX047nhGwvHWSf41njcl3VY/49mEw5VYzVpq1A++LDgu1o3MuqIpTvSkvtYnKDW6TwyT2lG5yhp
56+fgHkrFosKgGhM2C8GUGnLHW1H7ozhcVJbkfAKkBxWUCRz2oBRZc/erNsROmbRgbd1DAcbHPo5
Tecj9l1IDs3BlnBWto8w3ZS9Dt1g/G5Vt5VJbC+auDYok93/aPgGgCBoNbfzKoIftpluKrGEX03V
I8FgkhQOAtDokZfUegKZS2SGvmE80DI9PZpsNKw9j+ASIMlyanX/e7jmGo2hGF3qk/0C+FE7uiOq
5DK5h//bnb+b+wUIkI1RkbTlrN22X4AwulKlR7moPSuIDanJQ74vX9zFxQ//7f3CjofmKdmqF8kO
5pvmcGm12yG8gTHjrp+Pl0yrC1AJXtURMvNi6Gs8vN7g4lxQ74+yZQ11tusMQyRrCC0MYl5sK4Zf
WnMrN/vLmtzwe+dq9cTIwsl9P60yACnq6TSOn1e+CA2unxkJG9tNH8VrAvYo8louO1UABw9obVdk
HD1wV62gvjdrna9U5tw5J1hvpQAgbWQBy2csTUX0xuPM8WIdeOQX0asCFarxGtQQEIKF+5Z+GYwc
iRiH+YBZtSRp/XJeR4kBIS/Xk38qJg4A80xnzuITeGdMxDZp4X0jUBp1vCY23rDm22x+54ZeUTo/
Jng8HfmUOWk6Mp+oUOXldsdvTujKe/HKNI4SCzTn/08/BLSIz3GivlEmZrjn+FlHY5aO2vLBRglL
ti/ULpY9KqHMUOtDcHogd7xyA2SDlKeauRdXm0iT1p6oOeyVPVzxgM49ug6Qt7rYlvQNdzeZtavi
NP42o6G8LSE46RH6/JfAEoRwdfqFDKkbCMuCe80deJM+1WvVVYFYx4ZGs5PjUyEZpL6BNoh0ZcIW
D5qNCNZ1VE5EYLWxx+aUBE+oDiTzBcl6TO1+peAChNvk2ZRL+ojisG+QoJlKAxmJMj4/Ub0ROwjO
wbnHOqXD9gSQj8b9+fq4zA6oQVpscXk3szGzqrvNl+p/345In9JqR4RbPl1Iy7T5rSWRAZZPPT3u
zJ3oIEGXw5ECCwQHTVVzWnBgvxPVkFUYHyUCm6687fWByw+lY4ulBtazwNDbqgLZ5Becr3slm0Yn
SinxsLHyrEylPvFlU9mMEe5Ohz28lRpquAktGmBQqY+Qk0dtrOVYWWi0FpRLhyCfVyGRKivwPBNK
rcXgjP/wwy0eG6yc2WSrj6UY3nQu0QtTuBKVN82mHSB+/hPdsCgTWGkXrD3Zaxx5GchAbGn13ej6
DAkijosesQmL4+IUcgmqp+w+Y8S8SZOJfywI9QeK3upQVCjDCrOTB09+Icn7q2HUtT4n3xWlVEbm
/Ihbb3oE9XP1W36LhFtAifABlrPjoUdjb3lLRC7BahfqK3fWeuh8yp7QbY1lmz0iztQ18jQlpsI/
qD5TfLNL+2kctNas3zTCDOwQnjx8OYSTu6pIZILvl6EpSkJeKhuRVltskB/xeyZEzfta5vb4qYKV
skr3AYhAatjRY361hUtQOf6c3KGTfWcTskzi3O3Z6iTIJr+S4H7nn2ixjDQe7WCvihUkQYIf6veJ
S9b0V7rXEqjKvw2tBWah96jECxNd+z/6a42NGQitOHvdR/hom3PTrqLO2ovo3J18WVx9yK24IJUa
3chRPvSYwJj2TT0FMx1Y1kqeo2QaQl+IQmkVbItWxT1oAmATL+De4DkBHIJqfRaz2lKYerqASpYG
d1Be0XrdGg1SFaX1TLm9p0Q2A1lS51warmNyQW2gVxTBpYSRx5jmLF2WJxO1hQ4PB8I2tLsnqsmJ
7UJP63ZHUI0Xzcv0LY8Jwa8u/T9ZBv4aD2Gag/kk9ywkEGlpFiZ8B8rTh8zDYgU5DpTQWyguYVpR
PDkwuq32ilXSboE3KAASHvD5GsfxaN0ru1gyYSpqGIaSe5EC3L4Hm99u6HC8qxiwD0RZL/lcFqly
oUG3aLQjs0+0BvLg7fpV6q5cn0zT/P6NF36O7UB3E/APV+YPS04K0H8nko9TJ1GBRlijHZaMZAfV
ZzrV1UgeVoQ/xiPMIdd+Rp4QmDxatAhLJ8rfdY9fMLH1QeuKTHcskgx7HR8oKO0rMIa5erv+guxw
nTPmRLOsJHqM8h5/L1z6+zGl3wG4Jr7L9poRKG5jYDXpbQ+ZaGFUpAhxGvpOZWyGZ47uvdTAjJRC
yN9w+N8ahxPFlPcaCBNTCrb+ziXZdHuVS+JNikk4hK9wbEUIQcGK0HklT4lE9d1tlb5QuF+a7zjs
mvx/eyXHpvBxGvr2RTfmbN8rIEuSXHNUz1G6Wp82pJX6fEXT0ADKvhfuTY53kfPxKR40sKecUHqb
fYW5KU7JB4245xrkuEQ/mA3J3RdexQWcbbvMs9MvvaeoKbK6Yhg/biFfKFtjtNnSFizfaSQsx6i+
lpDbkXc3XQ1NmpogJsF9oATlbTyNqyjEEG6W8GTYBooDUZK7Hgst/FTEh12SuGP6rvY9MMLNtdSC
ubnAtc6u7ihzBQYwXaEHhBYt48UFWd0/7mK0qf3l8PcAfkEGAwWJa8u4sDdhyGhT+LxVk4fROiHq
I8lYO0TfXReWWArpHJ/mmNu/PMf6cQNy2BPmEaSs9MqxFfCKbFufBSvdT/ADrz2Ridjq1OTgIzRT
obIdF5igKt6mvugt1FWcaUnXecyH7nF5mM8IxZtJuYuTgOvy/R2kqMewW1OdQSMzWrawlJSUYjWd
aSJDjEn6mpAi/ZAdWytOvMlRBrlrCP2UhJ3VjVr3JU8wJpFkFMpf1sbI5PPFEOlhdtzwv7o4/vJa
h/e30sZjbOPlOE5nb4OHjRUff4OAywgsjHYj8tFBYWdDm1uNfAMQh+bt68TjbIQ6QZ7ieHMjJvhc
kLFQaPvA0OLufyyWB0sV828WxC9ndqYA1TN9hwPBxg/X5COchOE4Q/2TWAbY6Svts+mWFiftMYOG
X95Gx0oneCrb3bk6gQqp8Q4arhVSdiLCFmfyOE1Owyq8Q3fu6faVv24siU+Nfog0oCAqwEmBYjHV
P5Kw17e9fisCPYA75V65EDT2Qw1FyDW9exNLgBxtfQPeJ/ohaxRY1e2h4YnxfftiZMHZJBb0h8Nu
NZGHC87cTlACX5AsUxCssZWYXpaizuOUQGr1X9xeUvokJbOV3dPCjF333VKSmmCN6y6AkSwqJJKL
pa+mge80e7jkSoQ2+G3O3i4IMRI2RutY8/actXJIqsG1iPBuGtXpcztLFlO0sxiKNrpxMp1/Fvd3
uBgucEK1VM/90CtWgtIkpf5etH0PJ7A6bcMcSrkNUdXmxqeumBYH59p3WB3NXgbshG+hTRhXtcq6
+1XzYgLZBtGJhCLtQEvYZLYbqNljJXpUzrXaIj+AHMznISf/CeyQ5M8HhJtQ7f44YA0rK9lN7v0T
+lTsoQYyb2Rnw1y7nbVaNPSnd45eFnEhJ35IR/0Mw+dKB1TV1yQgsypGvTUktF1t//kKAmX1Yin1
F9ZyZULbNjC7JXZG0oRY4jGNRRyp1h9kc6Uryg5CGR16ZawC/MwqzE4pKLVQAVu/rUnTeq7FTVju
gTHdXVTjbQEzIKmYzpo7UZzGSFS1iH9SDdMR+qCug/XErnIdXOoFjb8sr9ItMsYabGQh0qojm0CE
vcjDPQ5+QL513XuC0NPTf5Oi8VT287u1nf63CLL6Vpv8irjU/znGD6/OSEMbS6E8SU8nBVc4U396
dqgy1466uUAbGGMcW8fJhbmYWwNhM0NvDw5mj5EH1hWDxePRdLi9ir7aPWUXhDTvBJNSmz3sxDHG
fGWFTYys1m2P91EV1k0C8daclI/XAwqnUwq8FBYO++kEwUBj3wQ/lgw0Oggx8LuYDFavOoCBqKki
yEehWLlunpsKThSODsqRih4CSfzm0e4ee2d7YjmCBnwFzX7JYZYd7l56vR0y8wKfgbGTpYFM9nnS
lSUJyvXtt+NMyyxil00yllhblIvvtKGozH8mZ7X63jkOlWVfjuzkNDLsBT8720PyQNAlH6DA1L5e
IjwAU3dOoMwN9cvQCk5nSIxJZ7SrUIUSCK9FAYVOyeaOVlKmaQ8/uDsSvIJ3+mQ+E7GzDzGl5hgF
nINqswiQ9oY7hQ2WQhw9p5MIQDvaRcpIBnNJfae9xNxPoiWO2chX59TnLoD952irNM/SG6rHVVZX
WCfVN+8N9WY/V64QWy9nLmRa2260kHea1Kjr3ROuX3PeZfQgbVOjdUp6krnP3IWLaMwAdYDZb4ix
c9EU3sjqGqgPm+3J9SzZBsllKjvaqUto7WDsJSfSNxyMA60wQYAzGg43zBy7eGX39Y1jCWMagsqN
wcl8THoPSh9eMR7k7foZ5bx5yYLjS2r9ofPtM9jzJF4klYXD6x0Eld+MVyZBlV463OEVm1RPX5cU
jswAt4yTE0XJdKb4EqRdRe2axbyxKNtiRQlL6OpboIrM0G0P4VRNnms3Hxoiqk3yw4/G4yu+y3cB
exi1V30vRIcoxT3A+JGCJUaat0AQPRu6E0XU6kxo+EiSOESvBpdCIdSnhJw9+KKkNsSe3/pFNz75
ahr4dfyFJEebaqz2NbSKXf/lYD+IuxiahShYnjHtn3MhFHEsgJblq/n4KhqO4VQkRaC0B+8xHN4U
oPdyWQf0MOA8RWN/TWr7sKE6yBgPMSFEQSRcSgRREQb5/XNRx2HRVbOcO3qYHd0we8zoEAXNU5BD
639kvPq/204rfdrYbaIztY6/X6HUmGKt7WNI8t+XTNK6qklmOqNwBDU1+4/POZNEacWGphxE2l46
PDuXLkKM5WHtJhuZkjQBDgaW15XXJDZmfHgP78w79ALTKNAr/1SVM0bgG5P1WPNYcQwlETiy+0aM
ORrA1LH2mlqlWwRve6BomoIqyUI79HYeTLq1ac2PXSuaBehYXImwgDfenE32EaY/WYU2PPNTWT8R
uKJaQ2e+wdLqPvWXzebZres1XKVekGi3O4op37lWZWG4U21ucZB0jSuvPO8Fd+C0vqEeAxzlBSsc
v0Te7t2iOX9QXEGTzck6p7OMwKClXeGtDtG2LmKxQ5OQ5m1zaVRdextkEVZkKhQ/eYKvXtd+s8NZ
CJUPubNFeVSNUDqu4eucqNaVPgS8ykPri/tiPJSHCpz93hELRCRJCcQXOnC9KU1p2WSkNjI5XQPL
CBknvFbP9tGvNiEsLl1mg6/Z5QE94ml+UtVZDgeF10FzcXJ5KXai26lJ2Mbdsnf8BIsiKcTd/57b
LJgxvSOv4ptUP1dVn7XN7lIo1jjRJdlq6gwybZsVxqDT2oUK1n6AxuHcxeypwIKOh6UKf4NlIUf/
8ay+nGa7oNgAzG3Iu9pzPRm74zpvrS5Gf9bZ+bvJOIPt35mzTsdWu+PgLKilY9SBLvB5EMxNpF/K
nuK6CjQoU8qsomrRRgtG/28EtMVWVTVh1pJlhJm9Ll6yVGUJ1yjKK1wTZVRmW5EZqXHa8IWqrdzA
HQIMzugL9w1Sd6VlyYjIEZl8lSFBemV+bqaFQhXcSWt1LWFhpAYQD4Fpt6cOVGqAadejt0AZxcxh
jxwSwdKB/nuRNqwEFKrF5/u/1pJbdlRcz+w2m6fzNUkB4DoXz94Qr8uxMfNY9v1p2Qzd32u20uZY
YkBeLDNHX/Kajes4JH5LJet6JpSetFeB7zZ5XN5UDaop14ksQX0Xg5KvuMwkAcDoNrnSF8tPCP68
laAtlSU2GdjHRBiRwVFv9QSIz+uwZ10Je6JNHfIHVum2iAYEGbSuOXVOWCximAqMSVCssWiI8Zi7
RCp50EMVJ/VW4sLPYK/0/QzRZAuwwywheKpfJiinRMaqdy0U5ZPXRrMmVF4oL6BMTrro3UxEBaCR
ZD2kRDm0XamlWZKf9IrRukixIW4QHkziSGrE3pTqZNCVqrS8bMBHMyacUiqfniaS0a/K4XH5d/cw
5hJJYDzsPes3DIaO7LRyTS+rjWBHOCrpcG/UIyxx/QEuVXly/UlSu5IMgITjCMuKejdpWsVWmxq+
nMIaMS8unSM706ZFRqFRRHsADkSDp5Nf9/l/55RhB7zMzB53zSsCPuyfphLWoWN5EpqTtq1uwRcj
hZZeseTtkyHZDq6HtqBv/XCbeeVE8ZYcTvUi6fPG9DxdQvrBnVGWZi6z2q3nBP2UgRERBLvAJPc9
znWmMZnvBP8jOCYm0vU8tXKyB/FTNSTy7Htwf1cJRj16ObVEzToEyzIxsiUEhCqfl/OXRQFDNbIO
k+h33YpAqoBHzsn/IzcCAROduuYcevxLtO3axBqX3ucPF9E8v+7e32dBMhPAdwikjmafgGTObN9L
OcQ63BkLpC5IxPQT9rDOvQg/dGAKVNwPkHhnJSYyciVGtW9y673+xdRSc0vmlwmRF2Mo9hzLQW1d
l/0/Q5SUMDcPwEPvieiaIahGl807sImiSvnrBhyzmKk1qJOuT7rSCgzCxlmPvKCqO2c7LZEl+wWZ
3h2DVmeTTZIX01MyZaHQhnwoZoApX2vjg99mNZAWNIN8HTVZvIcgXAh4wnpSrdwwD/ThIkQIHQyB
XKUZijNNjwliNPrg3mJtS2X1I3zgEaUn7KEFzurcNewXKIjeiUdOpv8N8fxd9gFxdSBqjIe4mKFm
tC2de9Qyqh6oINWnk89QD0Qcj6JffCxtqKjr3Zp86HcKFl63IGIoJCvtTx3/NH+8QCQjEMQLV1PQ
yofefx2golBDNa65p5MFyjX6RdxbDQ4GlWHkZJhABWMlkp1z0kRFkOKBsLG/BNsVoYUO9VvjxkaM
6fHDN00rjk7qxoUOneyQxJGL99gmpuqhmQXQfLRK49jGIVAjw5sBMc2HlSNUAwdRQlLogu9DF5Ze
FxqpYFAk1kHNWYt0snDg6eOQ2X3H7htv5YuhK2JeUY4I+wxjCGG4sIxrYu2nl+RmDGQ86Wq5zAK/
6ZYa52OhpUqU/0YrPcY7wRF5SFtj6dXol9sNorUJopFDK0dT5e+wSVE47AmOikDidm7/GUAtKuLd
nRVZQIQgDQwyY6V69wDmqj6hsnRDPXooYg+WlTJvBkJu3q6eqqcg0aSMazqmf1pxsNMPz6dKzY8f
eNRXG/jA6LXxAv6t8R6F57stcl+/vVAFdbH2hYepPOxo7wtzpfBeuim4pSopdKY0K2gPC/iBH5VW
arleeS13vXAoRGJuvwyATuyYsbmE2ySuYgFTLt3aCSWY8cpvKGINpVD1EdjxJXKFM4cceIToSzTd
qoSE9m7CBZ7vK/3k6wSfqEoKH7w2eMVjhbCJTTTr8Qh/speIVMy7ZchPzdunqGSL9cXMQTt2aRWk
J22jFrHbNPQQJHCRodoAct/WdHJsRx4Qd4WeVoY2eqdV3X7jxGecoQuLEvihPSdewfINnwhpOfdy
PHjWZOnVZlCHnnPtGq4QcvxIcqKoS7vOYtkiRomfE5ZmU2tkplRSIcTknLcCrXxmk2g8zaQ1MgB/
AGivYA7olqWvkSZhwvh+UxbwRwSbiKj+GG97VgZSN15jkgqQ9w6frYd1Wyi7xlAwo60qKRHyYwzZ
GjLCOhAw6rlHViSUbnaWIOrh+IpRao2jPSGR45xe1wb44uwv7LbnR5Hf3e7x1PC/b70wmoSYPuH2
jMZSPe6H02nTV6qqSi2iKY+Ovl65k7AnV5QLt8CO79BmwQhfY4bSk363g5gzzzb2G5mq+xN04+lC
8xqX8CQGxGuPdNmu8l6feENwk/6isyNblrNXmTAzQJswN9qqUpWbfGgvqkC2gf7xl3tHdM9Jy6lP
FLV+ruIVgPGd4OEuPkKcSXX2ewapi5O3xgoTTtuLnnqGrazcYLvQ80nbYYL2suy5Nsld0YlUTi/5
B9J4IWm7rhKTh/dgNjKHJWJ1KBYN9/OKPrOyQN4VdbZSPPzwxSA3BqrtOHqGrRrd6ZuUKsg83Vkw
0m2bRd6w+UoBRsTLnDOB4UiWu28ufDRehLkpfcscSbvgVBxrYFdgVvidkWKEaIF1vpAy8YofrH3A
rv6dJ0fQ2xcfmRf7UDzxsxHdvzQfdOltzSNx3uzXXhxfh7l0Bg/Vw/t0fKteSjKQU1f59pCeUP/W
jLUU0w5AN6xQ+o6K9UPOOTmOH9sndwlPbcFCbpr55XjVZneM1Mbm9R9sge6N8mOcBQAbCj1mOfqa
CgN6jUW14Rwh7IBtzS90ca32bI6KEKq5pegkmoyastMqwVBKOeLYzD8eHZGZb/La4DfsB30sbm+2
HjpO6xGtCInEEr8s0sNCgktDyLUSLHwyxq5cicwtwY8JRZbW93JMMRo3NVEC4t3hiLPbPTK4sEKI
grcFGcKTKgOo+aSA7+RNyaYNX2lgy0Z7ztM2JvsM96e1imwNFnYV3XYy+6ckPyQBCON8sVWPD2rr
HSfNPe15E7woHgVez0rjpaf+eR7n066Hr5rZIBjZNrXKpNjjTy/3TI9Rblxy0yOeLBRa3z/T7a41
2snW3m13D5cMMZUfMcGQ+SqyLsPY1JhSe9sIbP7lEBF6XOh/VbINgdzVZFaHNBbaJE9u1PlLu3+r
6HCwzfc4bGjXf0PqqHTb2KyaicXyfX5h/PMfOToD00hdXCkWs/mf+/nbWtGMVKNujDlrsWqAGU5T
j6bpcN38IPPZ6hvyamHU0+3Yr+/tHJ5Xsfnb86r9EJDSVtYQBMsSlkPpUm0gfhqJfqNg1Vmo+vWZ
QnUxCx9KdRvsLUKEzfz+JrV1L1fKsxoCjM+IfjUQAPw73ey5Ms03Tq40BMNuYxBQpXMMKuiXWKL6
jAwvjcO1xYUDX7FtspAwwNXTfPG8mQDU9RU3aTpmNIbVNSUxf9XzHaxP4zBJj+8cOt7Fcrz/2EIU
ZD5wDzAQPoh6Og26GTklJnS4HqlmeeHQDXp7kuOZDsWlmAXv5n2tObl6xu0zgdgc12Wb89XgpQPY
GnY+IKZLHboJ4aAdo/qdD3G0yqfMzHpghQqMTsFZ7aNVC2YjtNaMsnTQ5X64Ed2plb14YYNFf9yK
kPxIQ+3e+lWGkmeTu6dUyh+lbJSvpW84FhAHcGLV06iwMJfbqOzxzAEn8B7IXkrLQMMheaOO85OO
b9CIsvKFxps8PiJmnrLWxtI3bMgzH7QnuDLWXmbEexOYXSF58vlOSbuB6aOXYCcFfqRnI28QsBZO
LNA1E1hX8ffNRdTdTmuOTCJlKgRFDTq4udQfu5TeA+PUnaoCO8oD1jDiN0MqhU/sHY5/PlxLuNTk
fYkvqu74O7Riv7H2t1LcA72ISfPYEzvYJrGpujOUqL9JD6gd625q8N/lcxMcd83FFfP9fZiPQWa6
/uuIS9Ka8qvXOspFT4cobU3YBWInBSOIdCmyAAbxYQ+pYzTb+XzEvpS7gs8Fu/mP1jOwTvN3WKTz
V+VtpunGoSKzU/yfQ3pBxDaAa3Sya3k8eKjGXfMKi7naDW1jWXUGGavWcRMpyUIMhakvbVfz7KVV
yM1/dKVI6Uvjuw4ivbP/M7dOecjgw3JErm2w7N3XLpLzQ5KB3sjTMgMaFfhwiobJu26eZBp8Mzzq
E/6TR5v410EI8IKjE3cPUncJO8xfaVSVnavvUYKXYf0MDHLhaWgutgRXZXXT9N30AAdgCaJ/d2w0
y/6+N5daiBe9Ezs0bXMrG6GydjbJ6sa9KjqdxcqxY3KLcZ1YzaK6YtlPhYt6QL29d7ZcQ9efsSIF
cfoFl+AV4yOWSvz510QTV35bObzYUuORhfc8Dwd5Q6Z/My56lvrqdVWvogqJqCrjjKG9KtIfJMXL
iQgB4cswnhVYEcmbCqJhfFOVXDMdfKpAqCKYa8hSbNfUrHuROcKoJBcRyUN09p1uT68tS1/H0BnP
S+krDqx8/VQ+4+O2xJNh+0BxKVEScjWvEK62REaRYe3waqYhKSXUv1ih/MsyIsmsf5CsrQd0s5JD
97jfyZ4JFwrdptOAjpqfnFCszWRnnWLCoXJtZHBTmLj39gxamSxNH2wr7vF1ylSAJ5jDmUkUoRN/
RuL0lRSYw4vsIKjU1MTosejyboXBHegpGeRfTuK6grJEjmDIyGBekiPbrG/Fb2LZbvtd0xVLnZ2X
nYiOrTBhEPvs6xNMvlqw/VXX42hOUVhJNaLfemMJfv1kKCmoFDnoT7WHDwcadit3hAt3Etvtkwn1
6lr2EyA49NCizqY26KsGjlMHEWv3HpmgM666m5okyF+JyePj597CKAVHV/YrqFP5sZ8iIZDzDI97
N7yQut2VQyqbi58Q6qGcPWxVR8HfFEFGtpLsjZJdg/DnqOODZNCO2cpjjUDM/PgfqzE4sjnnYce0
kB43PVN+PonZfMkdiqiMkelasknwsrEycpykh4lx1cgeAAW0Zxtk5E5+m2q/SMJcu12XvsNxTgBH
SkIwMwL182V/cxd9Opv3dUMSyuocU9RBGmf90bZKN0vkLIzZBXSsgrQ/zBGNHKx7WjSRmlTpFeMh
hYyXC0K4Ce8ODOAxHMLVa+EQFLc0pfA+SNcB9igNs3+uJj9Hfab6gFbNtoVgX3bTCq0LO4Hlj+dN
0cXn0ExAiOmA27/o43CEN2dReoYfMCHuvqClmQ5ZaGWmonpcwDpUciY0UpbKD1qqld7mrynSzdPk
SKxDMbh5i4HP22dx6fvIbnqz8DEvL96Cu5DFNJT7weKT0AYyFgFGR6LDgWHgtEzU3inZ2ApJ0J6s
qNtfEQ80lnWE/IR/KIc8vBV/jTYMltVvotrWdTMHsqML0q8TAIb03Fv9XuVeynJoH/ZADu39etjR
4v1axVtDHgbuLMMIGC34BGFxSzXNREwVkNLGu2rYhhuR3JWtF08d8EAHu3jKyJEGPPi4pY16aFpz
rrMDQzkJZEHtWkWczMf4YG7yrUY4pGRuEWWX1jn/zsLT9jmGTaYc70nmDvMuKqaSkTQ/LU48O+ts
cYm8KhJrSgWedqdmgL0SQsr8YN4miW+pPwvubO+z31UHUBam43DvawFM90TCDyn0c6UjBkNzqsOx
O3KMXboW/0Uk+Se8ywbctTHi/fZsSKtzCE4gmX1uVpV+edHy0AK/tadxiyADAvd6FMWyPOxpDyyz
6uztLrc3iPAJ4ZjVXlDenz/X8KVJNa0rNeOK4HWkp+mI5MeboqwhoXKtWv7BUq9BxuXPadOyoo54
QuHtcSZGuXdAXVMd91tzssJZP+cQbdkX12+rBN8IrqfWntZTo1MCKl7cMS2r85qe/ur3basZlf1F
fSBEuYdkwI3vDvQdeDC0Ud/Cvv7R+PLNsTrAujQvNqmzRz7YEU6Y5GohZNio+jGq3gdcJ4LYTlyV
H8TXqDwUalK4FTxmg4iC3MIK57JI5XxoClfTjGGjaQgaNaenl4rR0sxkitro5WIwPn2qvqJH6vQq
UPyo+q9I+qsp3mXQnnG7lwCPoXsn6ViQHvFuyzCIWLXSAQyM2L3V1DPylVq4y1pAyohEcNrkHlU4
WbU5hWQsSYFSsY9E7fTc9vJ05fJvdAvDdpN0efjMEDE8V0SYWi9z3eS0nLOloHAiX53yxD358zqf
gtGr8Q/3sEhRNt7bhxhgVxSlS9gyufVJORVDFZm+sgCqCneONL0x9vfdu5OLY/vpw23hrfPZ9jVZ
8xYU3w5rXnDXrNwqZicXzKIyMiX4bT3+guf5yAisHjQMc1gUCVMq4rb011/qE6tsvHDQM34ZR046
bYCsONE/mfwt1ByD4XQ4SDTnxu7f52mnJxr3QDSSaM70r1UQQukQWfNJSjyTVcfaxgw3WaBZftwQ
53OAxFOPwgWMu9TTsJHFAKGkihE1nCfKj4gvax7tYabtfdsYlJ7MmvrtLZ9abBhBD9EhkbhClCRL
yXqkrgdRZhFVSIdC+nMTWz5faEgdGofLZWDnkAbErHxX003Q/dKMyLugEx6E1XHFPjKkC8zzO4S6
u6N9NbbZU9JJmPdR0yzfBlNibcOizBUJC0ycB0FKHJXjAevFKStTWDsqgWHnTTNjjLhK4D2LLCRd
/n+QZSO359lYlA3IQydnfX4fngavccwZqhkyQ59yLgYXLMdMvBefDDFtc0ukUzRJlOvh9g5WgPD4
Dd/v+TDwhQm8DSgsZ4Y/mxA9q7mOz9Crj0FPz/MEZEEROSoorT8/V07McVsVXqk8q0sEK9b4YTRq
BYS91IAnGOLOIsPpMi1rsk/r3xRCYxdI2TpU5Rf73LfF/WQSCCaZN+auMLHEg2CCsPqW/Yjuspy8
tG/BGU1GdKvZEMFS0XahXUuNfVSty87RdQfMvV687SpDCQAIg65Yft34r3HNbuqce/UhcZqeX9um
5fq1wdDQ2we60KL/LH53nKlMaqK5s0c/2Z2cQinedIM30T1BUHfLCL02ZfxHTqry9RQg4AHWut2Q
SK14E6zvl/jHMtbxWaVkMp1WxZ2/J6FC3AmWi5whmXj0FbNsr66igazW6G6mgTz9p0EI7BvMjzWe
gdwa6B/9aTLjp8oiV+vSfSly5r3snaKsXgAmiLwR2TKebKR1sSOo2iNluTQ11arJSfY8IT2Lm6Ur
ENFQNll27O9J3+zqqT6go+UmWwIDzmg6zgma282UIGha73Gr0xYNklwIr6xneFbbWvfsmlOKXkWj
gx8Kk8HNCHXcAUJOhubXinOXkz84EZ34AJdG7PqAeLkjy+fCKdsj4ypgCL775EH/zy66efz7S3m8
Cnx55wb2kQ2I6J2aHMSWF4Bp0KjcgPacikbZiz7j88ZbsyPZYqCG0mv/jN5Ba/vtdGWdtSxN3JDf
afdEsI1E8NOgLO+B1Q03UmuNEmqghkSgTedw9gmVIkfDgxSpbnlynIP+wCgenooKClaeOzia9IH6
cC3NzmGyqk0hxpzTgHbfiqV2vf37Mn1ibyupOD4Mhe4IebSOvu9KLv3uxTKC6xc55LqtGOYyUdOS
vdWFlC/6af08RXL5EfOFUWRL4hGuTvbP2XCvMu35vUX78l4AXyESrtVO3UeIUbGLxkU3gJAR+boT
ub3pkQD2heiXp2qXc5Nr4r46QVrT+ZnShSX4pt7UJ7PnDEjVC+vFjLWymQAa8ZHFs7SGR+vPJTKJ
Cj2pQmSptD8JN1AudGaj8Suo0B1xBtUwWCjbbzARJHiDEzTPjDw35h7umIH8ky60IQFtmWMPG0CC
w+Bxy8rzOk5fKjOq4ZXAp5c0Yx5JYjYVpv4BWkZ2XVDUXLLpPuU0kaUT83xplbrujXhsh+AWaSp6
HLc2NYaldBkYrN2teWmHXmYT3VCii4MP6kRubZyR0rZ/x+3AuwbGTicE1p+0ecBZ8sOErPetnICD
yOfCtZpcWrjmbvfq8S4PKqGyAkBMRW+nScTLRsKvFrnE+i0A1DAbh6obNUArnFnnN+Q+dUC3gTYX
0MHrdSyGaBPy9PRlhjJXTp+lSKDguEr6ePKQFpT4hAV5rdVvGJcuD3mkU0UQa9bOQ1xkxwJkQnJV
H7BLZdIbZw+MLbXofoUygsmZJGZc/a7bIR99fTM4fKFJmEjEXe3N1fO3l01+QBUvv4WEhUz2qx5F
5WGXuc7fgGtfM8C2JaUL0N3L2JI/nsX6BcnN7pwWB/6m4SFSlk4o6GJ4FDrZWxYGKSs+lk+nuS+r
2qX1MGn/kDHe0vNQpROZp++/2WglQZqIo88qBDbEyEFeOxIFFQLlHbkaE2S9vjEuLUPi0AlskFQ6
9zCcjSTNa15D6K1dHS+ufIYciA/39iN6MZ3OeJeRWyfdEyrOJpB2fTPf4SJ6VrMKgfI+7yNdy93v
QwH8zxuOUosFpxsUPJX+2I+eQivoOY/+PeIdAK5QE+q5KrxXJvJVRexpjL3aK6xnTe78eUD66EY4
fCk05pFMMttufDz9YAgtdyl4PuN/5o5aCPfKkHJeLupdO5jLObOJ+3WpIi915YeVy9Wt6F9i7Jvg
KHnojD9Z4VycvhlXVA+1y3vJtgD1dGpOYuXVm9LwNHlRdfF73PUZwyLP9H49xNnlOBdprjABs09C
L3hyQGeonN2PTaX2LWEDuKdxd0SbyotFvWcQqe2T/aK5dhlMdidO4bDEOqp45q8EmKDaUpMa5Z88
2EAlmtr5DLXtjOrQnQMTNiwQU4fM8nrP7TtP+AFNvxv6Ipg6tc8eikuEzXWPZO+Sj8SjlcEh3ZNQ
7Y/hXN1kKjzD3ktiWKKef3bnW6XNfUrO9vjCY3wRUefdFi8xHk764ylDJEK9eNh3O+B8T0jJa2CY
QX6MKNdW22VyVXOTupRFcq1RnI6j4puw32Y8eXpYf9IWrAbw4StT15zIhkMD400VDWAL5b5mBgNl
E5daqIIOOB9YcwOLSkCpg6t41wI0WeS4JjrdmL9wT4Bj4SWE19b7IwO8ibt3X7Dg42QYXIv03QXl
FlsMHAsaVUUpXOX5maSO2aJGHlnMckccLVcpyCgiYpmQBA6L9ZrGUJCxH9yQVHdH5PYgb1g/3xfu
/RWotjkkJrx+f6YjobtLaAOZ4NIF87lZT0oqKInPoKk/1YtbALInZ2d0fllSbYvs0keJ7dh5SPhj
ggpuBGRxHIyzcQEL+LHBzxs16DDlEn2wy0eFmYe1QDqnC3iDfj6XTylSbNkbJw/sh1E2P9oXM5sL
k6ywFpU0cZd9CTtx29k9DQDkKdRZlfD0UR9BTywpM5foCfb/Qz5/W34p1zovQ28LO6YjT6SDp6UH
9vzZleiMK1d3+g7udyF50B8lXdqXVlWp4Y6meczgUzGzowcx6/YGo1qC3EjgC4GKX85wzNCahazk
+HcwVMSJxBP74QGrqjNcHEmyh+bCBX1188eNMuahkwv6CAbeuJYbtnqcqtzcVNrB/ILdVgCI4nSI
YyoGUTKmlYxfzzz2/LcajRGP6YvlBGKGHAQb6vUc4sxJTIuxAkG2BYU2BvZWluKJvqUX4tRcSPDw
mwP1rp37LjKYq1/pd+mcHQLjRbcUVG2xXDsU+Wt0/y1Zqw8bW4vG+NWzLXLyipcM55ZGgmHWbuP2
5w45JeNTSJT/I/MCd1EUstDeaXWkRMDverjcQlUYSzCBYJADmG2yxw9F2jN6xbBd+M/fu1ZZJBaH
EVwcOhV2lnUUAu2i48sH+esIn2o11cWlrhSzTB9OME8kLjcUt8DsyLmAsjcy9s1jxw8XvidD4Hn4
B6qE2/IKMlyDzSfLReU7bjZPs+Yy4RvIwhYlIr53bfVw0QSkexPQcPSdHC9TQvgv3JQfkIdJg4fi
Rm/M7cHgjzFg3TPCJ33nfJ+79WgzvOjUpg4p85gZYcUr6d1V/0UrFabBluE8Y2TtwImB/dfj1Cgv
1SaMKZ5iJJFdL668SRUMhvfDiHjrkBV9MVffJ1YIp50eWQLpTL1PQ8BvVfshrVjXeP9jYWsahH/x
/BY/cXgPu1UDAVYd6btvKtLA1jOS7veqlHAKEhWykgLG0DVE7kb3QLE2Bec8sAki1tBw5z7bYaEy
lhhKLBZbKPcZfHXSPJeIW+7RSQenwyz245jPiwVjb+ox0LGC2RNPSBCqvFRU0B0midBl+L87XpGb
q8KaUzRmklNfy0gg8b+PTLk/Cb/1NUf+yVYDazggcVUzxjrXWEiCJwx7vfxZPlsyt610LqOxk62Y
rmai7OMgigYxqVJbDFpVSK2aQ/MT7FJR8/v0f0CDxddNvpV+rJI2dMKGeiNOlouAPS6FW/B4vGRR
uOg6YNV6UZ9JGF0fUE4ULqZl9nUqUnPv264jEERf8pHee89D72tWrBIMB/QsRQjZS8N9Vz9+1sM9
/LorvxArkCJiGcU71KQmQdQiIxUuHfPxRngID4yZ/7p7KQykvm8kX42XAMeR+ENQYsHmEuWsx0IY
rhlpNTZ60EIILVknx9dLXEcKTUjlTc1iqnEMvk7ieoJX8qQGVQIPBiRhDYa7bzuwtLEPkRP8Frrg
uv3vJ0jk6eHoWUG877KOFvGd2tBT8ReZDkto3jrX+DyO78M1to5luSzAkL+oyp4WWWcyzXqUaJHp
mBAqcCs5yna/TGgxpEV6BEUrxdtVUbhKKK2uyhDNsS4Hu6BA/429sgtzzaAh5Ix/Txsw4/wOc5tO
QU0MObhOf902cNZaLhtbnunQHP7F8mOeoShRFVGmC+hekMO+NS8bS7Xp5GP4JPdNFILR71QSCer3
R0i60abWyGX/FN9unUN5g/lTEndB8C1lAgHpDWZXyfxqjPW9lqujtCt/k9vvd7m76BU5bL4tXM48
mNH9JuM78A86Zz+SGTv7JC1VFiC1KG9SqwmZL9E+Vwc06H3JNKLemtDy+8H1DmQlOaRNjaOVvhIn
4KK0FeoUNfr58VSoYjPKoA38q10/tsocby0WqZ2Hk3Q4OhI+5r2Htdq3o2Tw6pRoLzkOE9LX47rq
tCwuyOMgImInGDxORQLK55u6E02lwZO+yFb3LdgUXOeWc+tCs9BeL63IXa3FWlKns+MZoKCTK2Lw
EH5FSKSjVHaCrlByiiKQKn2ghdjDO9n6+UNBEVdQ2Kluj7WMBp/q0WX1HxCgXM/BBL/t6wnFNit7
eWZ74QmbOPrSxIM4yPLVo9iMRa67yOsSGNGTVvSrmSriguzxYoowW82+UuSGaExq0xU1gO71upCY
7A/jgFsY2XkxJkM3n5LagUdrWTOf/V6TH7NpSDzEwftmULK7TY4+kJY9KAResixYcd7WJpdcgW+A
P9Jq0kDkEzfgzpPMRx1/rnLrW3wp4p1Qi4i3rDRJXmhmmnw92RMGiZwx7qAEHkCa6rwvyFAeD5qE
k4zhwirtjiomEBWTnrc0rYMRyZv8uTNihMwmfmDdIg41T9xRnzB1+iLYjrX9EOZiyZ2T4yvJCS25
Tk5BCJePYlxwQDUVqHMmJWFQPMruCVPN8SfhuW8ioyj3C5QBqRu5Qsw+nw5HyNUlKtWlzY8fM67g
GipRLYbr4TeMWpKMaMTHkLSsaRVXHBBgoELpCZiDtu7sM2Xqy0rTnKTzXXZEw7v6aQzGMQN88H+6
zx/3IYVT+KDtmFRbQA/077+5TKm49bpYaz6b/wTrlR0Sk8ORJlbPccSid8j21Ymuk4/hk1TfhWKF
R4X9wpVKRQZMknHZQb57c42s8ybDsRzyCqnvtU7mgt/HB8Q5w/rtdvKq7QWB5cj20DSLo1B+2mjP
tbi7L81DN6rFDf3hnfqUuKG0eiky6g6xmTZfdkPacUJi5MdGlMJpR7licJPpOP+G36HE2xSTVmV0
7xS6XDv6JRyOAcPek8fI2NttZdZRKPEF5nc52Ppwq0zOkdTivHlAdx5tuybllk++4QSrAyruxggV
Cdq9QbQhnLhHI4BSA1CwhQAFK3oHHYU2H2vAokkIrI6GovpVmeLQ84Hh+EJdEl0v7EsodtgU3H5Z
JXYdRnaIAvTFpvDvNvuYBFcobe+6NihrQvwNYgG2qVJi/7dKjaB31MYllPUrshUJg7Md81WD6Y2+
KBzEMuqwtBgtiMSQYzby9ywEI/2ZnRZcDGltAaHB9wyJRK92dIhgSW9137DzySRXTT03e28j/O4X
rewTZBNNpLpIS9mo9f0SsrOBk3R45U5Tgin7wPdfqay3g1vaEPNFccOFiUYsWabH8XxwG2PfjHo6
E+i2YVEQUeddxXuDAYFCMn75C5s0K49qvdcgwBpZiTYgmWdlG3u5jjdSEoeMLP8EVlolvfBypvS9
vbGzKyErFoCRaO7GWGS/aK2rZO1GfW6jAqYOuxZYlck+QFXTQq2tq4Pas1nNrgojKIdx62jr44MD
LgXk44S4S0lrlp27Qdk/AcnepnPLAt7m09zVRAxKwgwRQ91MJ14+IGrxtwkZISyr+Md5wNn1vsmO
LeI6F3UGwzBuebAneFL4Zr8n5+PolVGrsWrvtWW21IhNP/Ybegu9fzuveorjNIf3lD/YyFgiezgn
XI+hj2XIR3NTTLKN3FqGrEQTh30NyuhCl0FAk+dkCt/O02YSG7hGeAi2hLnN5xCd9dic53EBWPkc
xdgtRYaN7WnXREKdv2pBFxT0LnhGbJkuKj/JGRasGp6mJ+nK3uIS2UhVbB0G6kxtzKhdqa66eGU7
JmWDjrNqE4c1QmoQnFbnKwe5uo0ICEVtpoo3XBr8KUvObYWr2gcHKKLwW3cj/fJB/psZpq2qPDfU
A3HlkeCGhaME4roq4kiyExQylOhy1jfGFqWeTB6SRbAraraEo14tUMZaOtuqAWynJdy4XCNPlc2N
jZAYs7ItAkZhr4sJKQJ1AN9jylz41u9BxPaWq1As+8NCqzKfCtCAoDxMmm7SAtg0kkSMUi/uyGRY
UKERGB2tgBYwd4m4DdJwAL44QUSuB1RatSjUXmTkN9AJAJdOdgzrByDCvWMm2WpM72uH7VSZeyG+
eocT/sRjMgn9Dtc5PjD59mkodVJDwRao+MBTAnSu1MGshiFK/NVNj8+AnMI20qphApXrfKtavSFz
4mIxpjCDfnxM9yoLdFDhYM44PnSrAHy1X62anDda74Im8wMK5hvOZRr6pN1yKlA5VI72al52/bZW
5Yz2BXYPrRHtkl9VqRd4WzHUCDnESR9f/7N2iLE55FoCH1g3AIY2r0YxVorXU1aUGKm/wCDM4mvn
Twe/zFabTYTH9YHFDmxU9cN1lpRgCU8NbqJwJLVOn9TMNXXex/f2U2gzejc0vf+/MaC/NRtQVItC
lgxC3oyfU209dJDKmj1q7bsfGs+msLy7XU9UZh/4T9Y5FVk2suJTEQC0pCu27BJWgaOtHXzTUuea
NjNzhQiSZIU7jV6zdWQK4nkuERPUCya5rptNNrZ4Ne1BkZ5edeKngBPSGFaIapL6i2k77adr4p1s
IP1dDLNAOomQvorxl8BR8FgpFWF9S/rBCg3KJwwzaw5iX7Pn9AEPcrFI+bZzIqdNauv137/9j6vH
HXg5BjEIlqiGTJWhlCSrIFNAH/O0lLTYrvzR8xSz0ZReWlzfeYCTRRpwW8xXQHVdHPJrXPzq7fnU
Wq0CmOg9ARyxm597rl/A2mZ8uEaZGuqIYHX/YEN10gpLQZW16rTKHCn6brFSYPsJ2XdGiz/dJy44
FESDOoRoY1VGSOgPbkTiBWSCQFHTrUWoTexnc/gcozrt1FsPugHPh8k5v/HMrq+h9L+jQFr53Qbx
8TJSbE4+k+tPE0M4q6wIPpyVmS9rn7GtLXgeQdWfk+Oy8/MULHKcZeBu5o7u7sYU37tKFKOgJlsd
pzr/z7PpKBHqfyKn5VDVNxdfhl7OWNI8qZuOzv/MbLm21aMaQPfgfqffzIwV3CcTncjGE4aKhDhM
rtK9c/358kYLcfnYQc0wWbA+4iqNcvk4eWyHYql/0hAcmHAqcoRXdAuGwypnEhAylwAYHeFSaF32
t2WVpprhTpLO0+2PgPVm/qagvnFg65aI4sQI2psqWuSJ+IQiHWAcuwrW7GdErGOQoiW3eLJgs5YN
6fCYjjxNz0p3pYcVnmM3C9kepEsC6wRBAVyNayy8cGPpTZWy/nzyDDBEf9wsBY5vtAoBsmh4/dgo
g2hmgTrds0TtgJWnAJOxyYJuPIRr5hNBomnX7/ws/1a1GxVGHtbulmSGs3zLMQKxTbso0xsoBLka
5ESmq1ul/+1Ne38256xQ6iwrKWh8ok0uVsK0q1bCtRG67mJsuWSo5C6fcP0GSCTsw/qDRd0ULJX6
g6UOiTG4lKGsh7oPdT1eWzISSM27iWT+1585aTDVzuqIVX9JQGJHaBcaqo+V+r5fRv1Szxg3+ttY
g1NFfz4kanVo3kvPMDaWBgNr113Y8U/QA0YKL3F17ueL8QKOXJO8zK89Mn6A3tKmAQHWAg1PgLhb
+JjZE6eFLBRK5sSBJe5frrPLm9D4PGQlH9WZ3j+xoVnwEQPskvTA4K9hfM9OmmorEVNhl/uHeERd
zkRDZRFKa5FbCEclSg0eQGM+yPhkwOfZ1gdQI8rAnI6qIvvZVtUBSVmasIpEEwoRbYm+CxYNkWnQ
hpxsTS1lZ66uOxIl/llRB6f6mqTcHKqnEIi5/IM/vCXLy0A8v0cMbuAamWtgWX4JuZgatjajQ68w
lhbCaNLa+EjgACOpk/V49TRRL0Np7JYNhH7nAnlnVkwxjxHUWXSnh1CyRM1I1xox6ZZtL052ySUC
kri/dVj3SYtp1OYrzzVKPF6LlhftaDyW8bMXHRg0o1UIC4rW0ZcBBtIW0WBlU6Ty1+SU5n95Ap4u
ZlROZMuY0ioKz9mOTlfi+6VxHlMdVYOq+UGksmFnW07+EiCVQ5J+ln1BROiDljShQffTmhHEl26L
pRWackhAnxPc3FM14V13DZ224LXn2BYxcyXyjFHUfXHhbAEC4BJJmEXeAFrsLIrisIbNCjVmk1SY
ps6NX8VxwziSdS/RRsU5IelfAs6LaixqkmC6RUBnG8qJoFuD1u1KH/9WyceqJIePdUIaSsYSW62D
wkTiFl8TCAzQu8T3kM1Bildcd+1pfhj6xzb2NMtoeBCmTShzv+vlkOUQJa/LDlhM0bX3pexLS7pD
NxFCnekwBLeHZPG0BeJj8g0qBS3Dp3MeftWS0SddtdVceQYdhG+TsYvHrQArC5K6I/s5IMbx9sQE
H8D4F8HFXEb6GpzfFcUuhWdyTNRQ69Kddu5wRaL5EVRGVJjYfQzNxDXinaKDLd+GdUdY7sI1idvY
HGwGm5EzKZFdn59RhhaFG2SPC1EBmSDyUAUzFkQ4NBEEZ0a9QGLgrKqY/MXl8OjAoNILpe6W2SRs
Z40TocEE2p3Ei2q55/XTsExJXA61fmWYfF9tEjWTT9GBYWfpbaVSiHPmEgQbGLYvyH7iU+8Uq7lZ
U7KzEJeWHzIzZBDEH4wdzDBTBlmvpIJLeO+T2TOjhe89upMH8uZedwBaYDpd5IxHYahla35ADQD7
a+RAzoX/AXPNzJxi86JJWwLu6LSm8niw/ulwUB8hnoAr02r/g9OIAkWYEZxgQ/2YwftlMUkXPt3A
f6VioXEuQINhRb40nHFl3oswRTHY3ky3DUdZvOo4KJgc6K+5sRgeaekTu8EVgtMovVZUD2T07tCb
XJj8vGb3JyYtx/mGZmIS+G/aWQ07fqQ4G07uDKwI6ADlPPSclJ35eifPIF+1Hobs9uFrUKLo+PWc
r+zs1zX3wSWKzrsy+tHJFKyHfxRqqcVLvOIW468Oth6phJzzjh1+yHjXzvhyWxfRF0mcXd0IMULT
4C2mexAbhhl58A6CR2wsRMvRgbMMR7OOZyJRecZWAP4x+tu35QVoKQbcMa4yIaJWyzFX0BD92jrr
HRx2zlSufn74zMMP3OTzLcFJPQVaKExFQMKfu/B0Th7yjicfqoGkFhcTuK9ssiJGsFvIiV25AqEO
jIhnnAzfKu+DQAyQH66glnoWTtBtsJYiLBFILgLqTwf08xyaCHBd7zdwcN7xn846F37okOnweeRi
6sPVc+4Mqj1kFp5RCm9EB9LoAHpPKgzLv2dJ3fpyjcMwQF/SBFW0CedPYmSc2mIQ2Y6gUKsM/68Q
PLo53gfjfCx8rI2Dl7S3SAdvo0VbdK38BkZM/xUbhLCQ05phZa5eN/++Egil1c3psIFaDEs6aIML
9gxBxdIdrBn/dG62JUrXKOUHiSLmaqlouervdw9LCz/g/wFLnK1rpsN+RUUZgadSstvr7CJSgco4
n3cOhbXMEzljNFbGTY7tTw2WBIUPpE0pyUwTT8S6G5uxxxAO5VJlB5M4Jf7AkOjUaJCtB2mCycRG
qYmQnfIoIyAaQ1ueMI23RDGZY533bDFmpLU2vMIs6KC2DQugiQoWene8JJ/ls8ab2XgBD6oyMOC2
97dbP9nOWatU2zuffDXfAAVfZw1+Ssb4QE8Y4hp+an587RKd9Sqp2MZ8ozsyD6qUTglE4iFbF6Ou
Lh0rxBPKQXcCKiPl2cYYXT7ZFQNiEv7J1tQd8CPhi/JBpUcVt/HcEYgo45l6WpH4T2vS3hLaTM18
wCru6SrOKXsM28D8djRJYwiMqvOT69shMoXRJ9p7PCqZzTejZ6XpR1QyzccC90EgNtrV878hJhv4
AZk1jPpSKhB6nnD7BfIjDNfnlTz97pd8NV2JBnJ2u6KjmFKimVfHaANR32MQw6wRX4zRx+iU+7nb
r8K0s5akpcEaspE/sPAob+XfLrdBM+5eN387LT8ZwBU/Yl9LqbsBxTznt7juBJd/TDJF/w+p61aw
LW7/TKnncdwKv0sX+099L/z9yTfot7GEx1BYXgUBZnetJxET+Ec0CU+/ohsYeKQg3G17g2sTE1i9
3Zx0sVaCg6tiw+HhZfadLoKP5v6jiKWCTM+AdfrD4cNwnIQGjuYGJWhryOPdxlUq7PkWNjJlvlNX
Ed0qONTD6N6sfRdkadv/rbKixLrPv98VErbAq1HYs9k7URYIvRjBPSpCOJs6vC5WfFPobXZO+tCD
9ke+Q6zkcEK4U+TH6VOMmEJZ2u+qGFDayqtMhXJSrDygEnNvVc85uMkuLTCQ/WeOprpsGu99a4tz
nOeir2jEIXeTOQyt1iIoofn2yip6MGfU7UmQ2KwImkpHv/LYu3wgJ/ovxlwd1hXppLMoJVubTwUU
xDxqNSNz0EspwwS5VCJhAXpU1mhZrEYPpDcePwCqD/61hhgJDJ6fYLyP2Z2/4DAqS0zlszST4N3V
d49mguP5Y8j4vPsx+NGHLzWAlQojqZo8ShVI3V0B+AvldsRoIx5C/1wTn9ezGm78AHiwbKCk4Pk9
LcgiMjgT5chbMNSPcCIk5gvqH3ebbV9aphaW/wb7LQRpG5p7U+/ERLRNUx8AUeUcykXAp8kRbI1l
J1zjP4uy46M72/rVxu+Dw9PPY6KRkUQ9ptBpnRUY+egucMxG3o5zU1bIU5fa5n3w83J6fcIFM6HI
vcZZPt9B3gJ3VC6HLraWfsVS1uQu5xJDq9qiHDlqkDJyy73qToji1pBwA5LbkWRlWBjGt2m7DOAM
Bry0e6prGdkiMud1yZqWl6KxZEpC2GXw4coWjzekpcbZqAJnr3nb/YMf8x+dtvc8OoE0jGeEyfrP
v2KdXhDYrV2J4if+3Nj90XoB4aeXbztqjB/6N+MlqBVZp3GMnz/orsFNGtOJ4uqQPxkp/dBSOH6h
hQ0YYOQX+D8B9/fE/tDP5CTkgmaWnqTF6p49b2gjDKtXzph9M5CNwPXppcATZaI3fMte+Rg2Qsr2
OlD8WglVawjKWi2Y4O16/D2IhjX9KI9HR/AetALUNwXbtQ64UDT2m8S0SbFHxovJIAQdh4ZonHYH
yuFuCcDcId88w39O5AgQYzc/Luecj7XePM4vwrzMgyPpUEUeJhBbacfe8BT2RqLboOKNdm5cL6qZ
nlQ17rGdZgd7SeZIV26860tS2Xc3+wXFnFPDE6RMp7m8U62st2LQlaucjPd+0tomUI8Q+a/oE6uf
ojtnH6cC/yqgU2L8UqQQDecdQmsqcthG9CGKWFeKOj8MLK1f9y1qkvA8W/pEKOXH0jiugxMUn1uN
yzej6oNogT6y8c5UOajSbc+WsVR20gu12p913DT6AqwQL/moNw07rn/Rf8FrofycDGQL6onkMnCu
HIruhfb/a341zmTj8woTBMD8gzC/ZPNuIog/YHbZnxtD3ZUrYZMNJT/zQPaPA4BjrVm8dJ+fzHrH
pvWRkOGepDChIVRR12KIN4jlShi1kamJXHDPJSz+kBwSU0ilwk4VGokND4mzxbYrCaGc1CNrBExh
B8PNpUv25POS9Brk4XWD6gyz4SSsrGl0oZ4ZVbtv9mIKrWoY55JXnWw4tlRYTAZye88kRT5nJ9uZ
6icmadKwRMCQx3VprRuhSo9nqT4XIQ5iOptxFqfrYHQ93K5QxIOhExdOH05e8q4ga5+JD8F/8l15
adnBN6EBtAQVf34bgOs049Z2v1kdPXXy7uouaSsHjR1tw9RUQADLHqSMUokbx765XXrS0ZW0LZFY
Y/ZP96biFkKUKdYOziYojhR0snhgC8GnG2k/fm3IuVmHzTfyK+7NC0kdYKhxjxJ1yVDk9NYURrpA
fw+bcMjk1VuSQNZeTqB4SMpybW87B30lIHU9ipseTJPC4Kv3gvYlRAOZsWZxS/lj83+wLcoQ4ZqG
rcB7S4qZVo0DXkycmGd4XMD/QkOMAhTLo37jSmNJfFyZzY6sIB97wwZDnsfz2ZLtOvKWAmF3b+jU
LyhMnDZUsnKCxAO8EB2KIxlS06U8i3UsizMrK5A3q8hhCuzb/Yt+9CE+IK160W51G+oaUcuvp8Po
gTjQh4zdLvH7ir2VUbFzKl3OroEKMGkO3J7/X7NPBeBdxTg5ppM32xlK68rxkDdngOq8r1IzFjXV
gAGClaog+o25px7kFCEs9ads5PC1eGXLPBUCiFchP9Eezn42LaAyg/aNrCennFAUTRSOp0UkrfFR
fc1dj0Y43mr3/PzpGvGujx8ISOUSEWMyoA8BExnt89UL6OPWLB78zcMX7bteDUQzEqzZyr6RBwGd
B8ghMc+JWnmhN5kRoO/HTOC/pEJ6rFZNPQmH94VhGoS36HS/kBwQYhRo/MYd2iZj+Bg0pZ4SYW3S
xeym9MeDafvhveODUcIyzy73pjRMV3qqdcPAdcB+OJNc31ZctWr4CndHqixJImcF53S11LkUcKGH
YyX3XCDemm5I+yt4fAvqUKB4WYOwCOLR6sduq89sGNot3JMmJAiVQIgXFOdhaBtEo+kwW3XpsxJJ
B77jDpQ/xBzFTvA34VjkcYIp067413CDFVjqvkx/kxXj972rrYkzWe2bSWhI3Pxzep1jYcpR6hez
RhTsBuhVtFlsWzIQbrBDyjib+1nYaZSfb4YVI/eQfqIHhXoip10v2Qq4juwuzLxc7lfwYPTZGiIf
qTkGohw/rKhzPpw10WCC3pCSJF3hTPCDob5etowIft3t0NOzCwWRBSULgwu1wfbYWvzVYiivhcWy
PE1MZKjJJXnaA8A91ZNZ1uFj/9LQXDh8WXlu1A52azCkGpWdNnD82/ejiq8M35xDDgOLbdidoKMG
uVRqQ/W84bvAOkpTYEhAwqTkbWaDyX4Y2f6rkZfCSn4TibRrM8IguOtRLiVwarvDNk6ouJoD25gf
4NP5JbZ02yja1DvgJ6wlAflz7SkcM082cJclHpVl62pTCg5hngD/TecegVqiH3DXLn9m9fKyx938
5TXbMJeKlannQ6r3ajruXGUkQjyxgPiJJC7bphnnVWjDIbE+jP1m9Vk9BRkn2vYufC0y5D9DQt8E
HJ18dQlHcndccYBIrmJPzJBxMIXF5Tjb3iAfSLNuEFsCVXVDIOqzJ1GbhmaFUV9wWK7MFtWLasxP
0BPlBxCDz+D8XX8cs0g5U9xU2gunGf/KM+pPW7gueOzbBqvzZBjHt0dVI93cDeDowV4PC313F28f
tIlBSCCCnsUoYZfcf0ydsH28EcIMx27o4q6yBdyQVPdGdjn8zGtn4G9kaWH6+aiuo+j5z0Ja2mNY
syk5wvqLYyVll/sevP+kD0ph7b8bIGeaUBTW5MgJ2n+oFW9vkgzIMG0dHLhf/8DwJEFdVpf4VO7I
yne6YkSLjH38hKdbWth5p1LPguJkbIJC/5fq/tYUzdUVduUhmDYbku8xKrCrNblSQDdLaUv4j6fE
pBCLcBdZee/zx2q6bf+zurwhPQrNUTjF+saTh+K7pBT6ndRJtjxtIvNtpfMOsAF3L543OlwLC6mI
eMkXMULfBdw38PP81M+z1ecbWLCnwVjld4lfOByNdMlTyxKrqfISgd5ECJT5cIg8dyecZAHkA6jD
S2QKmd1yAQQggI1ouqKlyarIJQFyK9JhfswYD+jyNCCd/3c1HrCJsipScgJjQppJHrHs1jTCIR2P
y4eaC9/c11hTBXEaost3t7mwP/8Strd7DjvZaHXTMeh5Q2dqZqzBN8VyWYo+P+VvRAH6dbJ/TEEf
1JNI+DC0AHC8CKDLkklZyhjl13aMXKTwgulfbyRBwVFFKgKAMYCCP5AYtbJfMBpEC6GJqogEtsD7
IltXpBs0v0XB6vOysemP2DP2O4DfJ0FpuhjmN121O8jlUaXwJPvxpfl0qhsFgZ7OFQuNTpIq0e4O
dXfmbJ5ZlnOGHhceRglYyUFjdfiHVlYs74rN/qgxYf0goeodP2/atfeIjT1yc2rB/Dx89mLHVLk/
sPDABXGaWH6LRm4usX27uTHE/zwuEYau1PQJCDS4Vvwz5tnzk61w9RTMpsenAfz4WNkUfQ0XaGU4
t4TqkoGY/eK1sOyMrLG0leBV8v/DTcivr5F8z640XCFeJ4UW/x/QQXowz4xHeXDRrd6oz5OUmhP7
nZ17DAyC6rfDCicEp4xkdez/nkT1FX5hYnB9XxMeaHtGphNYjuMfKSsyLXgSt6nGIgQq0ot/IB1U
5bwagrrQVZ2YUpIeSmwNPDpZ7HjNixltuUzwzbRHELqHohIh51RLyAxEU4ar+atn+SsQNI/zzc8c
bhKzjRaCn7v7+U0r/ihyAOA8Khct+9T4scDM0XW9CnsS5Vz0BFmjkdlODL+rZDyrfkvWrpK/gbYF
ffufKIroI9H6FErQdSKQmbSzCXufM47E5szwYPHa4FiF+q4kZSa91kHyGJ4Gm0Qani74rxN9eSqm
tMn+UrDVCUMqKXXgh4m7Kl7kjlVMqm22tdsTOGi1MlHUiRZ6cjfz1T5f+GYhzeZH04BM6seIE9fC
7xfSm5ZzneYqv7amiu2ViR7MQ3+wf57yv+lauhaLa288GzedXH1IJKzTbOeEoAfYbgKwqfhHWLW8
GBRL5BEHEzsRymp5omqxbk2lWs9Fv4j3UqKphySagQ3El2jIy3o7PrIk0pGjTRJB0lOLpGoMKkDx
xfPjbHo4p5MvJBCs/NV25AoyDGo9i6vaE4UiMvT1XeGnZfTo5V4rpLrvrc4bsGJDJ0NLJ0m8iv+x
hU8NTSoD62H5Dj2zDvEErZoqAALnmKn8A8edsqErHB+n8/A8UH85yMwWi332kPw1UHks1kc9O6zP
IiWPzMS9eQo8IjcajKVuuE/XDI7gpph2RLhEI5pMGCos2V7U+a53DfQTgOQlJjOgoFHgaRBnyUgv
/SisO/YfSRJFWzqkVQE9xONEV0W6u8WUk0RgU56kh/LRRyrEdqy6R6yPUR6hPypiKeGLsSMZl0FC
zef5oX/aplSp/GZ6vBmkkvjMgwYWAExT33XpnEGswF8VWXgyIwQ5JHvtUru/cF8B/bpw5aljl/qY
Mt9vY1ghSRTKAh73EupFXsfAk2FglcXhPencZnyHRA8/30la21pCoDxlUMnTXkQ09/J1vHdXdDNy
3iw8hcTVv8BnMhbzvGI7ZAyFciXrhTtzIHq8S6zljKKozT47/7f3yrVl5gkAkJZmUU5kSneanIOd
S+LbIPV5rgRdIzy7SX8eCYwcicBZRGspWgdEzApYt7Mji/OsDJnBeVPBHu+MGS1SZt3Tyj27zUzf
kUPO05rclhoSX5v3xFPxEuyb9h3heRIHvNTY4GoEJlYYGRSs69qe+RADpQN0ynfhFjtJidJ+Vtm7
c68VMAuqSV98gg6a6PfR9BZyCn2z2lGDMkR4EERfDxsV5VI7YkBJLGyqXdMvlgi+/zMHCnnLUmAB
zBYCzhbKC31l9p49sB+iNyCIN6qAiRpOdlBANY31OqkLXMbxQGQru2ekCKmLMLO0e1Zmbo+RFLsj
ABsxXuJRLn01Sp8VDvyg8IJ+tHZRl25V0+hnCpmFJ+scgHTluljVTB6yxTt3OahUdwnHE3qCXmRW
4W8YFJeGUlSNkC574Tf7r2suCHVXlvFWmotZwjh94j9Uzx7pEAhA4RqGyDp1UZzxnlQ8/1FkwEiY
QPnfIAL6hsAk1aBRCee57whREhJb5vgKd8zxfiYquZxH4gLhPtUPOH9XBrQvsdWnhCRcjndpt7ZI
IqjqDZBYSMFFlMmR2Rqxs/vAi1NgIaMAnXR584ClhiKEYRYZAK/9KCyrsk6WBEd/etlmC8wUbHhL
0glQ/wxOxjMCf61BFoC64cxUXt67y4Hx1mRvxkcCrMWxV3Iz0vlSCBssEMncuqyX10tUk1KNDsaP
wxfGEURF6f218sU5zZl+GbeXD7Fw0NOUXn+GifAuf5AtcsE6uPWT9laVjmVecfTbC3JCkURJME9N
aP1c2KYhz42zpGth+4Wnjx32Nid+nNkQh+NBZHW3yhLOUc0zabzpbnQ1pnshG3g2Hndj5s8ySH1A
QqJ7J3yskaUxgR3k5V9vnjNXSUa24A59WuSgETTpEo7vw7e6gAOUNmJc+gof0FRLSaa+n/xFPc4N
vE7SgG/dCQiZQzZ5o9kcsI9y81uQUeJJpsihmS4qS9MoyrakO3klZhJVFZmqrknt2b0WOGdnb1yG
MLe69fbQA6NgwI16uYYq+jFSLbEboy0tBnXF7ov4XfOy18V++cv+GkKRGZYRG9lQf7UPh0D+tUaD
flTRVa4ZcGYHtaN2q15y7cvTkpTe1t490OhHIeY7HrxxduKt4jqPC2wxVNJHkgc7wGGmhbvKHimU
STGUBlWWhkA2oOSQdOiMRq6apkuU+kK0wLJ4nwromXZ0MBubBQsCOBcokflaZTiKgxtLlu2Tl3zO
Jxgr1tIzHd5cUWyCeO073tUiluvnAIha30F52uRC9ZyAnjGlkycV7TUqS8iXkEbS61FlPmnP/X+l
0hzjYzPtnBzTmZ5v6p9AxspayzlNCZZN/DtlyBFSmvw9mX2PZdj/1CmJvZoBZzILa6dnGRz8EQSF
V1wwzZ+AJJirlsygLQm+/51be6wNOFQ4VpfRDTaRX/70+IQ4GLdHaL9b1zjvvGq2oQfTA6KriKYA
Gt3+7jbC/n4xY8Wd/SuWL5PC2nhhbZKi7gca07pnQDMWjyWxdVAfkmmDdRzc/G0MwYMYoFBSUvH3
K/tRMxYMxhyDzcGBTQCQsAevKM2rjaanppdc9aY5fL+90A3sypyOIGSxpq9xKrb5A/ynRNfbRU8b
T9RNxwf/i1WbRmv1KYfC65MqGSOMFJ4nhIE3IA93r0ceqrac983yrIrWXkcCIJyUTv3M3Ssw2r4w
1US6JUw3PJe6vFEGmqA6gyJmClRWlfDDOW3f0IVqbuSDa66U1SjCrTU+z381ikSuvGVwt2oiVh+U
G9WakvmvHY+dLKvv58OL2bvneA+roo6aLcIgHgxmKS6hp0E1K3Y2VnFwinVqPS/bpMCHLeDTH1Nt
JFjIU1VeOBSHWmOJoQFr4f7+vxAf+lMqCsUByU7I5xP2uSvZWFuFsu1Off39+9xRXPwv8WYOYmi6
TIZpSnImOt/FIQ2Fo1X2CQw9Klg5FLUcVK29DoSUT0tS/NRfgEBVPWnoXJ9k8oPfCq98syopq4m4
u3RbktvVhyzpvKhiN3X3KkHUzGKQL4YH8hrH5y9GmpWNamT2blvTiLbmSp4ORxMns/BgZUfiSYTM
PB1eLfOqRS3Hmnmdzhd8xkNYaPXA5S5oE+G+ZuVjpwkKR+CFsaUJIgSvXj+43yys/WtRmAsYVlHP
d5OE6UFTK8ACJhzG63p1WOkB6RwKuckZMxXVeF5iGdJMs6KcG5gyP8H+rdzOmcsz1VmWk+N/UtgJ
jrRnHXaxBSgTPRoSf6WJiFdrHWJZkj+iGBcrPYxsb/kXxQLFfjXuXxqpc7FcpmYcDiJvAKkDpLCv
rdwWgzMtencXnyjcXxGMJDj2y0pYjx1B/E1TiK12/1/g/tUMe6ZAF79CrAEQt+EO7CDoSm4e9q5W
cUmJZagoATd78j6rn+la488dlK1jB86Wm1VaCv9FElMQUSuagBEFpVvTrk0tTuc+i98H1t+QxDcC
WZpkOUHW1moUnLm2m1MwVmcxmKiWuG0qXOdHVKuQRt5c61uNwAt4IXiRtsi9HTn6GJl9WGkQnvYU
DUDhi+CezdKyHh5K4bmkby2tz4UhYtbUE66h9DAIUkqY0XT8ZRo+hNtS3ibiYZ/s6l6jED/d9dbp
FojWspvAutvOj0Dqf9+2RfC6XfV51s4r5NELJdkgW5Q/B60ioZSpL1FmuMuxGRouwV4EDTh4HrDl
vRFbc7WUUNgWl6EieAfiL8CVzGylCTxAzxtk9nj9fdalgwY+hQaCEIob9rZMxeFFTTJCiCgFhWNh
EAqGcO6DumKyxWFR4zPltEmRH64XYuVvyyhWk5wmrPWUGXcJ1joduGs85yvAR9LUvXKwIuO1rBHR
5X8vqoBEG/+s6BM3OE9UNvImBiiWsBTGtJM+Ouf5+uLn2+dfjPRrl+rO31oTKYgFUuAb0uIeTT+X
KT/+Oyfl3wfZUewIagsAimIePjE8Gt/SG0xi8+t/zr/6c3jbLOJglfhLgK7TMXI20qEv4f+yFAy+
tO/7ufp4hbV0oC3NloXU7cbCac3EmTUOTWvR9gLVuYq29dhKcHVOy33mPU2Mk0KNV/vzoiZgiC6f
dXJaoGbjR05jV+IJXMrMypve1FzSSxklrNVGBAdc6yz4FXTb5zE8OvIGGWd2a0iUmnsC1SegHukP
RznNfuQQK5sviAmF0cYwOAnha52IWD+sJLdV28iYAheu4PUjJXDAF/CdcdbB6QHq2/JEjHf57njq
gUj9purxb3o3iO+xKzz0/gE0zj9pam8CKXM6oD16hH9XSFNDu6+fj6QIpFa3ub2lZU2M+QeJ5Eka
N0Y2VfZltvbIAPGlnq2+P/XvT5SW+y/LZYOwc3Wr2qNnxWdqgCeHxbs6oEi8JC5K31RGaBhiY7o9
zgnmiN5Y+xIJGA3fcZ6sLuTAOXZ3fAKAK0gFEGnkAuETFoZgiiTiFl0w/tcVWqUb2hyxKbVt6dpL
nIAqIS9lZgNmBioLGGmf5dl1Pmv1NVU8Pf28PuUn4KaPaIWzTaRtrLJNCOL+n12mv/J6uL9EkiN/
Q+o2YVfDJjE/t0veklEZvSBz+RhJyK8lNdLQjL4K0v6VLKtSoqaGlFRU58b91/gR1Bx91mYDEuZ0
jceXxCHpky790liwQr1zhjIdTZ7nJtCRca+sPdaKpkOdKFwZ8AorwCxHWCJlGeeCcwDCg6pCQAVl
bGTJizynYgxOiEwyOGusxijW9R+gSZqOjG/sEcuff68fZuaGhSViXO/X/MHq8tMerdoWJY/InNLQ
aK6NzHBLVnvCdULr3Nq2O+67RdXaMT56W8B+qw9dtOZSGDX96hOJ23BP5OWcw06/L5Uft3EucqQ8
FpkMZL9yqs1Zf4wHzPYFpo2zTht+WNMTBk2ppovSv8jDNVz6xrsoPmpydWENre97X/y45k2ne2K1
27U/x0DIoyKXygs7B3L7s1qxJthXiTI9j3d5O+ZzMszegFKH1M4MnB/QGUpg4CLaaeZ6FZ9fJOHA
YkOrTJJGbo9JCLRBWyF31nGXxXTpHW7cVJMVqCN3u0MVLW8SD50b6F8T4voHym6JU73Co5yqbLo4
H2wsl4VcpHOUZMrAlE+mObyeXv4yFbQmUausI2hh4+bZH7ks5v32uQxgmzQSz850mgWysX+5Ijkh
X8ukXopjGzTE5JlGjIyBE538vPfsDcHPD4qhtWIAlUvpKIIqVgyQXJCWZYHHDbZKO4jp02zPapre
Pq3GW3oeVQr8ySL2W/6ZGrOemuAdmDz34tvu/h06eVn/NdJbDmh5U9Q9DuXYJi+eEWNfDNQemEPd
pw6nEaI2roAMX6PCuqkAbMxSSIoeLwkljaKNfa/e3RW3Ps+z7CrTxCpzoLAhilvUKC39gSVHYcjv
g+5Z7aWQmsL/7BYcWI5VwwCb4VNsmye6NTGcVFynnca6awU+LJC9u15KhggLIHxLWHUTW9trHsHU
wQ22UEaj7Prwnm/XLrz7ilerV/gRqOpMP2syHrkE+x5x42cHfWezgiOsqrjl9NEEddlzTp2dasx3
M0ZgTkw5Vy1Bgifxmencu3/lfpBccK0YNmUtyPEfpRt1pLtO+CXS/GrKKAJ3sHvCFK5fwirpgRZi
K8vtmRPjzQmshFnm3fz48KZZk1YNduSs1HFe2RunX8iDrSwO3rUuaRZSPwmspCg2u5BMWBEFTEsr
nO5LS4n9Ig9v4z21KmL0H3MNXowChjFc6Ql6yRGLIwtYtY/LdC6hUlgsrCZu9v7Jk8B0Pn0NFc+I
Ow4klstn2WirtJHAIEggnjq4HVcF7Vjk/GsGsKsfMK8ZWrzNMJIyDMEWvJPMqDdK89d9qDufvXwa
/gCW3SSGpdZrQM15VyuLRY1eLM2cNU5VGXL4sd+tpaQfr/93Jc2wRTnbr/L3nlPvAgs2STsRhQRd
lTZgiajpuTeVXjjSagzjL4oEKNjBurgXE5nBB3dYxnl7Pr6SOpN/EaGTOCTGboP3LlqB0lAKTPNa
Ug1VI+wwRa0EAxYmIie6GHRmEJn4ywXq6BTceXwCZ3jHQg5fTye/5FWaMCM7EXYDiZJC2pUUwxHa
gdXfxvOBMr5OPjjYOvrwuz0/moOdVZhSORTNMttrwsEXTO2ULJr4WXY45RibZ63vR8FywA7fB1BY
6qRoir1929O518mXyxpvYAq6Mbs8xIxTyscFpNPy8xSNNHqmFnG+eHhbq8tkJy6vG+8MB3Aajj5+
iUedYsMzJ9yv02+1isxsHqvBosEPZtz+3R769veqmj1YiofCvmwxu+antUXHPHyDRVQC2EADITlp
QtN41iy13z0937YiofX8zdKDnF0KZw6zCxpxleLXWz7tFnz7vkvfUJMrg5yZkWFNoSjiH/OhEJsn
bQ0Wdtz9WwZumP43tpyQ2vzzSFM+e/xx9bK/fEHN5glVyP9zkkkb8Xt8yWRraGnANO1mAYWlDtvC
zJq0eO7ow30jusZxkUjGcPDJ9EzGvhvMC6D3AeZKyB5Lp3HEW1Qz78YlzXJGA5cML2Z4lmHfO+I1
7DIC4xtRSH1MLevCWjm0MOFT/LY1uSxsNH/yC3HApKNdBx4KfuM1bDYkCx+a0TUd0DqUMbIkTaGF
ga+pWxzvq+NM/xTZRiMEwLBZeG3pc6Ehk8JrFoiFYXlgNxUaN2LAeBxd9km/mAcTRnaVDHVM99/Q
nyIzy/VXd4OKp36oJsd2vUoLcBDLfJMFXDX3sR/4yroyOjSnqffXdCDw7nQTTQRn/N2/0uS9/9e6
QfyEie+QTnWNEuM9Z/n+o0JAvcL/5vya9OrCBECrNz5oV4+hxsgEvzLnAefUWtKK9PyY/oJfoEDj
hQuCIKsaxgrjmihwadkBq2xHLM60pfw+i15r9nxjqGyi94NCuY8yb1ETOpnmntPnyw+SqkS9/LOr
GIUYgGm+c2ux6MGuKWFCrmNAjk7s4xUm3aG/dCTM9DQ9tLqNfqWNk4wLRL77O0KtM4BgFCYCAJVk
T+72OrC7/TsTq5RpmXXizhiHFCuoJRSn13sOTSr8+z8h4I+2Ba4MzU6e7mvJ5PrNCEgpHB/mm1Cx
AVdx+Knh058/32yRItZHcGfN0dlTm8tOtesfT4BvcM3tviSCXaGm2zHL9Py6WVe64N1a052Gopit
pdLlOVi2n+iLIms0DtEOkT0X60Ab+3ixFxePfco5G3Q3k7N2IMYjD7Dip75OctuDgDQ47MLlD3jB
ss4WH8AnvdGGqxyFH2nMAaywhEuZqbG8XBP12iP7T6qtjDN0d/bXje1naoGING7Sp2Sr4nDOA5bs
3D1EsV/sv/VsLHaQkyAOnqFgjOIgLKp4NL4ZygsPxk47OJKp9yB0jnWHEwquBfeVHe9RWJ6C+A35
OVSPl7ItO5TRi8vwPIfUGbifwCbPQRJovV3UqbHyoiFo/sOBhpkrZ0YXgnZ7WYqa2uZnHL/BVnZZ
5VeSFraE4K2grpfLvOTNGzU/PxtEN817neNjJsNUY3rlEaRz6/RqcFqI8WM/rIzAVQkrikJhtkWK
hvI0V02BLbkwPKkPPMiBqmD5/lEEHylx5KeRMJjbvXeuNsdJarbeXDhqfI1xZW3icoqDbgPCkz5p
2O040yLcc31Y1sSL9wzUaunEPpeS9HdyMrwiBFYCsQ+fMdlAxZDrzUVno4ODzxW33kyDlf5KxwL1
PerrBV8IQe425nHChMCo1Jg6/+uj6kUBSj1bfiZUXWC3J6IY4FPZCgbDl4/RziMpYF/Dr70fXZRa
urJ9I13Eml9jUGgXElNiIy4kwaUb5qvqSe6SFXxw4/o3/6wky4JP9KkYEPVlW/eoKYhnT/NXNSLD
YLQCQsq1BMl7sv/v0bsNmJhpbZJCuuI9CqTwGp0DkG5eEDLfDlPOUohNYvfTZY4tC648Dzfy9npG
SsqnsPw9n/wZCFyEe+sJkuC56G/66Y2kUZ3osmbg87kD/IF1sL4c4kHvwuOpa17Cqwg/DeLY4/8D
uBiXAFIFTpRIcrY46yBDtM4xC25iG0o/ECNe6ADUY9pWhe72YT9NZrfxdSBSSUHtXk5DJy+AP/NO
xNwsuzl1uV3BPRtdbbwiiMHuVmyvUmHlmKN7fs8d869GDJ6tAlcpHvlPTTUIeeVos2iY545YZCTr
/0t0hCBBPN05Mx5Gd9zBXSbqOIaEtK9O+tQDcQASN2HsgGZCNvgguTKYYQuz8P8hDQ+sfvw3urBH
A7BMZW6jMNj6xwBjlBdn5Ft+qG7u+V8U3yhAsYTTsT3T8kCQ9GT4wYT4yVI5W1fwIgUhdaGPGK8l
TcXNR9QMu8qtud6+Y5psNfIih4hbJPhFdkoqPGNvgiSErgWw8NUgwnDH6fTFJ9PgukP4TGlx2mJe
m1M1hiIXsf1CIQE+bxnJWXwdaLgkqpV6QRyy31CWgSIvDMqHJpyHOgOv6Ks0Ibr/660fLFtgZlW7
QYFNMT/WrKtZYc3VGJIsdbtc1stsKdVncyHhQIZ3pYX9U2o4lZQFxMTyhdeHW8A/JlMFkhYaxYuD
ElwGq8HGq7yOvOwb2cMToh1dLzZzYraH3mbBPp43d5VXPA1aG/05wtJ/RV+2ZKtJcOenmtB7cJul
wfAJuoIRy5Nidxl0ifcRIyeMx3WOa65+XkOmnko+a6H2IR+Rqdqvrq5fFxHbJf7Gsyars3VbfIhG
E8UtWeLAX2LamgGHROnlreoPFR7xMCTNITR2yJRSY6E6GvHG/AkEp1c99FPwM0rc29WAN1gbUGcz
p+xmrgDsV5soKztHjHcZwseWh3NHMfNp47DvCEk3PYVtbEe9h/lzoIlzBRbqZhO62ueX25+8L/mS
gRE6ud+JbPa9skNcnwrYdXLUuNlVTI/pamIy9fgAFozXsU6n45MrMWwrvCwGO5tRxrF1Bx5kk7lm
F6+t3f4MPJhJU39nzAjhy4+hn6o4gDWgNfZ5ASlstd+l22FXDLbq0KTIROjghJDk8XgoeJTFjl10
VD0gt3GxWkxKuEmqXSN+0Q3WT6i8PSnSYr8SD11tW4qQ4MivN9eAkArKCaf1Il5xXD4B/jNqM0Gn
LykNQ42tUCR1TK7X0aMrDzS2ILv4xhPqVleLXeuwPeDl6CqYBmdNdA0QSgFCHpv2p8O6KK3eI7hK
DWRpmP5rKDqoxDmLWIp1+9Zos84gDQrEGR5qfyoH2XJU+H0/9Ih7v6n0OrRPTUqEkn5fILfbEq+I
uWUe0lBOVXmkUywwGV/7PaDqpM5qgB6gPv8aaGxrzthBt17WWoOKggZlN1F1g1dGeYxoCFIl4A3B
UvGZ/a+R85Q56NxcVLXsoDjbXctmWs1Y5UMUau02s25blXdNVdgfGDso9LtnDY3VFWM9bJCwcIUQ
QDG99TWLDfIiBAHfqgfOeWaLaEDYX5K/Tl3Ytwc67IVELe1+UIDoXuL28o1puhCMFEJyqZPCfZb1
6MdRa5z4evZVT2DKSVZZhwhId8pemYmXMrRY1hawAORzqvll1UjnGDw0rY+X4XoeZLUsX9O+CdOb
/etFWxhcUhkQDCTFxgc6PPLYfb5IeN0N8Q7BhT2tE0b44deTjyK7nv0Kk5bJnaii2xkW7V0g1KX/
wJInUM7W//l7EdsonHz/N6klAP/HUFqZHVe7804ekVVP+JNEScI6zGS967q2y5h99OS7gp/kr2gq
U4N5Me+iz3oVXe98FzWjYaVgnBR1OhVuJ2s1Oim3PnO5Us296ytDkIloeiikFbuXnec5+ME7sepx
L9JQjX/2uP0RJoiYrD6AS0yiA1mIo8dHLZDEru4sbWpjfBzljpYG3yBz2/WntWmknvKZf9iOWvB7
WGzRytHB6dRKzod5j/ismWUckncyr3M3mUonbQWkky9EgRSy8c5uUaHiqEujrD5IADc/iligKrV2
DqeurH8F/UIlhtHoghlqaABl3zDKYCnAKnv6lJfphbCjiqZtYfqqVBve/HonobyWmi1U0VrWdRJX
hpzhfDyvBq6g8xePdVcDiXhIMtOXaKxXnc0/qqOnwo8W1dLFlzBiIoMaSQZzWVmqGUFYwG3vcyRq
nRei+c5+iiZtkCOsVEFWFPtsFr8FnqaKrvwGfMmTQbW3waOrS0F/zXojeNZL20hZF3bQEtDuYqSi
HDCsG5RuY/dCtGR/elSzz10z+uYCF1rXSRsEqtLxMvEQVtzJe01uHFmt93M1WMc5gNRA3VPbbc/N
vs3H3RRgqtmljNznf1WcISR18pR9/Qt2SYof1Wtb3zZyzSatlL4kEq3wVTGqwqjt3TIBf6keVDG+
PpZ4pxKhzFGRwbc9xprrbfdovNJUDQGL3R5UNlphH7KrpP1lKtLBIZx2oZnaCqGy337FB0QAjoYy
YxO5jVpUuk1gn55NaKg2BVdiC+E//NQyy5I0yo0qW+RViN6aN2SksKzPp3yFx8GlNmgneJX1i35w
0b5+6tOGFkgLiSL65Rb5N2tMCdw2dyetHhY4DzkO2XuOUzuCHsctKIS012HPD/ayb/6Deb+EhkT9
IhidqBfF89CLhUFUTdk69hROPygM0auw3BET+KyPl9NDuk3SpVU88I58fbb7yHFBQPaSTssiLYHM
5Ib8uOpbpQzaud1I1LojxR2s0dog36VF0tiNNIUS2u2WhMbEbZCimvD9Rxo858OTUfOezowm7dRc
HYgytv5DJsjPRYo2gz5vYug/ebwiwcMycFfkEbtfXeb2iCQ/A/0pWWCZSNebv88f0ZBE8hTGeEI9
7CpzcesqIRixGivxYzDrQWlnESD6s3pvUknJ/K2g116mUmwUVHIacuCs6A8lEMnrSvO7g2ZooAwE
GOulVaKF9FNxY1goAGaURAnCmkZGftauW4wRp3QXB7MGhX/5+drbcw6dNYfdmN5T/El2KdQsWDGB
QYtvBSYyk5msm+VinfOsagl202/ZTFVJx/X6qcAcKa2jlrdsUR/LgrQ6CgesLC+8umy2tBS95FCs
yKDxa5TmxOkZu34D5HAis4ID3Wb16plWrymxcMyKeelexn0uZw4KsJlDawvw2pku61bBGwepzwGn
18orfPsfd5SSsr8urNhZUjWt2e2eOE1HuAzc86iBdPXkXj+vrY/L1FLEngKdJUohJYREhcTDrKJf
u+VskXrMeS1QRyH9SgZIFK65uroDtSSr0ES0/nnRaJNQUqnPnKk+qfBZ+g6ysbWfPchrJzng9gh6
Vu9ifWysL/Zxu5WXDWL1e+G0BpOHl3IWQhXFIWugaygtpuv9Yt4YdvWvdlqdga0k3cmlgd18Xmh8
q4KAV7g9gviPi4mUGNgy3XZJHhIynDj4B7uacF6QOKMubMgSUrqOoJEKfOquX5OVWwTIlE1ULEd8
6wZl+fbQ8XvRhrOHsLmSg7o1XpT/diYGJAtmYoSc1lKYxxiLSkX/ffO896aeHXmp8NGqcfjszfyD
1MF8b1RkR5MHneZI5/4kDbpnG9MdzLqubO9CtpORRRJ/t6A/nCurL/3ymtlCxl57HuLpl011mEny
A5GwtlfRA0788x1PL/0wAMTxH1+yB2mWTXn3f1iEl23B6Ny5CTGSoUK6Bfb79w/aGPl5Q16R9Cxn
GMCSQ5IjxZX/bSAonydvzEihQPXAMStCgTSzPROWGhJDRK75yLVXyrKonLFGiGksDKGS/Jcpco+j
wI3ubDbOdyd3skhvzWFCD0hiCsLq2YAvxl314kGM/p4M4KCjR42FV/p1GmHI2p5u/cj7ttfB+xBC
Ip2OX50Riatw0ReJdfEDeZwrDaoYY2Ia7XZDJilDtU74q0E+6cuJN11GzqnAnyis3qRGq2S7NYKq
Jodp4KgiU+sKvm0uTYvjCmfgdNbeLx8bO4Q6miCfA868BvE6PQRDkUUAWXke15G0C6ebI7B2gdwO
2ZLXIZ/m/iLhZj+ARJQi7IDvALgNYjhRt8WWMU9y/7vwDs5RDera4UTBknpQSxTy4pVwHF5uaX4s
oOyICL/n1hYi63HBCpWZqBeSETesO5xih+XZZG/tLZrXc8BslAbNtJlKoR2qx6I4oUCh0qNupA+G
IJ+97xmJIfAh37rNahZqUTZYlaW9xbOmxB5+tgmt+MulYgwChETiMjbz5HLhYYQ03gFueXgRMvgc
qjbY6rB5x9X6LLjBAiv21lITLR2lIaa8N136txD1eS3D7Sl+X1Rl1XTuenmxVcSxZD/VKOFYn7pe
1dWAIlgDZhPX+y51uJqRp30cMYkdPtFc8Vb4lQihdViahUoeyEmf3L7JUGWRecwBoJEnoDzKj/Bf
twKDsZ3e0Lds7yZWZkKJrJwPZOmwP3WkbdoZiktC4J44IGuLIU8pMJXVnBVq4iqTQGBOxLI1GwDb
ZiI3l+KetDojtA3d5uP0cO3LwK8tYwXyFiiwl9Pj3JQ0l/5V2+RPxOTOXfHzQBMmk/AOIAy+pJpO
paRuf2yswk0To1rCBi2WywzDGMIcQOj3hfTUHzAW5JvYumMDI0L0Xb9XwdgenMKw+7yAnG3OWgCr
XSMhaipMpMww3iFRB/u4oTdf3T8mOIcTfGXyS88hNhvGDJeMpPSifAGd33DLi9MkbtkCw7PKvRQR
6JvMT3iPpcje8mKEv/h6dZI8cubUw8F7FsiDWRyp2cxFy2swPOMJOdtbbBAehK68muY5MctxfNGk
PdVpE+KPDZiwhdub4hJAwnzj+7NNTbBk1wRpcHI8ycXviVKUELekJk9U1BpAYWO+mVo2LzI1woGo
CtF10/34sUbOLhQqwoydGACSLMH9JucVcxiPT3m1p99bRDUEJY4bt+VX0/Qlxqv6CdfRFTJDpy0G
aO67D0W3ZLc5JNEOCcBayzIT89L/Fj5u4equFqorXhDrVQXQCy9ZOtIE2RorhjoUB3QHI9AmBv/8
w2x/dvNnb+gZLgP4FRjdRL8LCIDNdBXuocA/P9umY6iWqGxm44ZOt2UvszjHbLEhuJkbpcReQGnE
fq+RTe6kAAOyb0vbbL8N18iHnsTAWk5a72EQoXexJ++adUX2JkJhfZmyUEhN2x2SDKNVNUO05LCn
wXNOp8deHcwooHwLPCm2eZNa8LixDOUiOH4xYa+xN26cQLoBb65d59IBpunBsaEzPo8xhgo6jfVg
AlKRVKPi6PwYSAYjWuyjEjfi1HLF7g4sT5vVdfRQ8reiAq2+65DIIPI+QprqpU311w0smXBrCPnL
HPBUCb3I4oUx07noj5ualRBG7SWawr/pnaUtSA/mPX107U2qYUb+wkxDzrJpSuXUJF3st/2SI8bL
EdL0Hj4yxDeMvvnlnJG+j5G36VKXELShsdX3KsnaaAwHu0hSddQ/2/72GaiolcmyScmZnvj2+LE6
MJKUK5+LLePJY8MIA/i402sA+WEHZfdDCqVQVITzzSErhof8QZOSVNYY9e65BfPhw6uFSc5EdYs5
0e4KqprsLngi6febdYPW4uUJ4ULpDRal82/YD5dkygaN3X4zFux9RHRZh1ZD7dt3Hc/bFXNHgE26
Zn3IxDgG6HgKDCLqyOJbcK8EDYZjZYdu7+CEzmpC5nlbbJhyGFgpRbwmpr0pao6oR4h28dXvAS+T
0tKKyNi7/qnEru2pbplRuht130F8VKX+LJtdA1LrQ+J3msNtS5uFiKmc5US+djtrvG2mjtK8z9M3
XZFf0JRmLRpHr247P/agB9ZzRnqnmPSsL3dQpyQVIaiOxDzgE6AH0oynVvhf0rUFhOy9ecjKpHyw
NAfs/Q7+LCrew0CioAyMOpJJvmqflBYyrVz8KmMTqZR/mSMDy+QbVqeM6OXVH5gF3CILnw4ezp08
k0saw4ZlEF6uRQv68TfxDSp3XEYAwrWnjkrpccCVbAqcbQT8ee7xSazg15+9Jh9vGA0y/EejFB5I
uyGUNmQ8oK0uypoInAXqZywupJm2gpSuh5glRGyadFRYpd/k+hSZ+RFclZkEmkrQcrbBBG1gjUkw
nycPVr3LootKq9Kc+ie9/N4GuLFxJ0+e6eAaKiMegQuJVBmH1Ymk4KfFxAjSJ7itABEduikIKW3P
ZLwIqZRwbU7ZLXX/gdjI9MDDP1+PS09Ac5bzvvdOr1zjGF4iGZUOAgEfJuo0ttGjTmc6Fv5plf9B
C9DWCrRfANwlPQhZHG2qkyAHbqfK/JzUQJrh2w61me1EcFSxLCXMOrKP6e0UqyMhPSUTBlpYUZZr
4Rs1apFARpbWnkrigl2FhL425VzNYt2ILkJ31QIXAz8u8JrWQ5vUB6QJ1kkCD7HhgoJwPbkcZQET
vTgIAxpYwmKGoFMI3HbOOCGVHqjnZ+7xKXyR1pyMCbas6mnbMD/PgtPDZ/fOeqWkSkTGrLg23GiW
IiS++Ui3Iilt/qpIiWIEnCUoe4fIIzmat8cLvTWeNdgpCeZjGyixWR/95qE1wsNxR8OrKotFTwJd
+zQnnmJRSjMvViC3q/fCza/n8dhYranZnWfJlGl5RreoTf+9cEgWEo4loG3fo5Hc4xXpCTsDUZep
PErugohsq5dEFApzRLClfA4lMKtlHLpKyKMHlDvTpd6DutBEVngMAsTuqqp61MosugXbHYz7EfLV
3IpZBh8KgK2GNnGisZvuVVLySW4X1u09wdd2sb5+xsIq3UcJfSh7XhFMsm3ojaSdsidnB7iFkyL9
fMt0E/UlOsll28RCS0U2kjQhx3IVpl7wKcKPKVs5HYVelCbkggAM3aHJ4RopaMQGiBGvnTzebaZf
nxKdm7HWknKXfEuum3sYeuJaIpKCI34HAiI0H0Zs4zXc7BQPpIoRnbAIsPsGTgdPO9CNHrY0bM6s
H+Lc1ehagNvBTsLmFt83O+MWvyZAz92+ptElzBrveZA1R4Qnze5Tw5uQubY2oGThmeSRhjJwXht+
jAvO7gdK/prRhGj1DYakhw026hAid2FoU3V0JpUZZP/BRUAWlvyzkBGXw1bLGgbtpE8SglwA8pCj
0K+er8fc9ziFlHCmI3n3Fac08bpTIBVFtkvJnxFLIF5tHQMc/KVjmqPJPUfkgQh9GpdHnJFM6KHl
i6iKEjOHELoRl7HD64uDPtYxJstuOes28kGDgST18w8DY7EfPsxqDBrh86O4j7v0t5JibhlLhwW7
hmv2TNnf0MxtPSk1X90ZLxdIZAu7/aZIU0dVpRkmYCNaoBKG4Pp7/wQL36jq1DHXdyNlFdlcXNsr
7jVwNDhBzzx33MN1CVzBE6chHoWVMOLWKtATUS3wBgZy2EmjfuJxJK1KU56bOyaspMXjaPECGvSP
OBhq6z10CCTW3HPtKHq2LA0LqLC+l6BT6vEhVTQpuA8Z1874nxtXpSPm24FwLbAM1i1W5GQr4AVZ
f+edKvwgTK2GyZkxhCL6QuuwVsdAMdbVdNnZ+Gepy0iXvwNruRDuDXH9aChcvHgdgcnYekZFMm/4
CLcpNJU8EhH3HL2e0FYy+9aWuqGwhnzH+T4VJ3oRYjF0xfmq83BF2p0bTW6LderW3v5edEXfXjK8
eCfShTwtVBuj2J8TCX3WrSeUc9pf7Je33CeTSlrs0FPfDy/+wluVTrd9uhmLs+EsU/yu36KsXzIO
pEbqmWHp0YmzrA4ZQ/JA6lFuP8j373yvjZHrDsk+DcTwrCjoUPRsrvJ2ZVIqu6lRYqHolQxIY0Wu
3e+NgNcQrX2Nuk/M1azhyETRwFyepv3LD369SpsGjOetdakWoQRDWByRnXrSkTMkpsfO9r0X5KBK
9yAmzaUsAXSwD8E9k27fcbe/ku2Il92D7dQW0/+1C8HAUR9lTWvwA7di/XuPRIUYCO2fCvFgC0Rb
RMGgdXzS2GMTjNBiMGNmRvIXmxFzh8QYOLx7lc3jpJovDQcT7r4t6YitCie5Eb3L58HPuttdKDgV
NmbKvoKXxjCxknq8RVXi8CL3SWsNcn2TyzTIL1GngMk/eCTy0tFZ6jiLi/pl/g6W7rrW2MK9PK/n
FnrZc6kQnJOIdxzqIAikIP8Vd2VBGKDqktnvSo/WAG6wVX4dBp8403FkvY6LlhldoEiSGeEI7jd2
PpxbhZAzM7f7Crj//jVy7rp04x6a+SqblAWEGrABdea8TyV7CtowW0/nd6dxF1/VQncoMthjcAgY
H80J93ZTQdNOJBol6UxVjXBYZh1wBWr0Rna43s/O9IEG91alpXs/LG/EqP7eCoXajG1LRNXvrWaO
z+aK3ALWZtYR5onNES5updgK3blzTaGeEklp0S21gTq4s0tjOEQhoxWOSo3QWPXnyLn/d9EYVxpu
U0qlO/YPoEXqzTj4lQAFsfmzIxVfTysoqlUU5u6qUaPfnl+kO5/aebGnhOUajQZZabXLPeJdN6MS
+zv/VoFioq8eht9JPypyOnMVRUtCJZcDy4ToP2InBzB46J8BsOr0FiZic80TuEE3ep9h+mE8a89J
AS1Sg+h993RFPyG5rMo9k+QZezatyyT/c3zL5KkBDYUl5rQVd4JXrRg9BnF0ZPcLJQMKPYBnYATj
xyyJw0+ezL+DsTQTqMGIZqmFE+6OpKxOn6XhtetHtr9OmVz01osoNt5HBlxUPsGYvP8U2GqN70IO
F7Fx/dEF6N2KsW8RtGwvY0MCHSm0TsaI64XRycvBsfye84EVwdb0KlOnI7ogrrcRT3tC0FPMNvZh
TN6lkYeISTH3Spk/lY4JBSFeynCUOsj5qGZgo4dff6hGkFHTe8Gz0HBMKA1gWfd+/0m5Kes/eT/q
JiAPoqbyl6FcMm06PNJaK9FpKtoMCi1cUhnWdgiiN4aSk+RlvysJtWbxhz2IEzkgHBRfivb7Z2JK
wOpRiGkFl0EHwdLSBCWCGIp0GEGpmZdon8CHdvI/KM7UonVw36NLMhq7deMILxVbb+S3m6bpIBkm
P+LKWHtf4IX6FI70hMGogBHE9wwkcUZ24ny1+jK+7H6R1R3stQtsxkg/4O/BCNkIJCC5UsXVILlC
PyKtbJI5SENpqMzy06V4j4KVhDk460bSePfQAV5XDUubwPK/HKpPm6dDX8tL+x8ecM2t8DIGDo6B
agH0Ac90suEdTsF8iPex3hxCZFS/mKbxqXS0P1up6uMC4FfVIIRXeHCxeqpkphRIecoOXrcqyeaE
MOE9uFcJryG2qz/44IFW7D5o+lBCZzMQTIks/SzSHiw3J6MG/X+6m6X4A8Dla1FVUPjMfrbjnyLj
gpy++h1RU/y6ffIr833Qj/l2GcKCRY+dxWI9moofSwU+eYbD3Vv70QPzcT9smmVVEO+l0UO4vlgs
g3XrPj23PKkwLzvJOw4fPk5CID/bKRutw1bp5U1hJ+zhEkrwLhBC+EEOofAE4D35DQgWyNZtJAjr
mHZxALGK9DSgoiEfhGThlGmNNt3GNVHCzu4FsJy+rqUus+3KGvBpdbhsZF/PCcZFSqHf4mB8rVDE
liacE3w0ZyKb2nFZf6Q9wDLqw5vOELYXJE8yp+6g+fPVMy+IEdOVcSv0bRtbYvyLkYFGfMpqFgnV
yrxKvEv10jlOceuPtw92ndF8UXtBdMdnp6uRe/b5bXrov2IkQaju8z7rR6N/We37EAkQcaCBtD2A
dyIKBqWsFSXvg/4oamLNWkhbR7sZMNTnCDa+FrMqfpMaNXACAAhMsn+8MwYNgPaLeP6ZtTbrBz++
0ffbJSEmw9S/kt5zQIizruIc50SlxjFfTbB6GqS01wH3ZwJcim4EZQvNfpwKe0uUf9EO9AGBXCpj
12cjMJNcH1D0v1vjgTODVNpVYYMg91eCdX+q1lZ3TUByIsOOT0LGJmFXDNn0rBbCrcR9A9UyVTNm
4p20VklJ7XExYB7C/cgxtxqOhwHH/j7X/nwEWGRGShdXcck5JMN7UsVN5RHM4VkYp9cksZtwGE9u
cmfQoQ67w6ISM7py2acGuAkqyT6k/w7w2MsI5d2SuYGaw1CW3fwM7S6kCyJeISr0ckxlXdP5dZrN
Tuy1dJYd4SNMz0wnjR9/utjzmm0UUsj4GM+abW9XybomN4B0de6Ou7RVsNoUosLF3uFmL3NxRZC2
uihb2enMluZMBpC1984nMml6vCs+XkBDLFeKXZtK/Br7jye2exl+lWJzhQD5Eh/xrflMc+wSBv+w
5aGzhPGjEIHF1pAyN0K/A4lBAxyVatK2BdQY/1u1bmgQStc5eLILdNhPYtCqdLqw9IUCITw2PdTT
jh5wU7OlnRjvHArOl3cjgmZ7cvZ3VaqfmgMlTCRZPCmbwNSn6htHei+BqM9vAy8l4BlajphuMX9R
MN+gmpUrCnxlcwQwFUbq6JnNGwnWRe9W2C1RsSb06Ns3ItgM3ZtZLTgRxrt4m6xr2mebHViSCew6
bpByMv9XATj+mkZlmv05fszIGlfQHPWsgK6Hdv5t5SXxlyo529TpCU8/vSgstEOWjB8vT5n9uxzr
d35I8JQKDbiDmZooyv26HhTmRDXLvCwDFulrPIcUSXzojw/cj95Nleiz8cNFeiN2rv2dxpgN1oWv
gpPBWqrI1KPdAdUtYksOTPZVvDVPkqrz9/qwP8/KlDYf1jyeOLn2RRU4mpJp/0j4ZeImQhqVPqPs
jncj7UhZ+QpgZdN+Pug4oGi8OfdRPVa9KiTEhTiRvVcmohQNPvajM2hP5OD5umOEgF0I30yZRWhU
xUmsxExwRDRFLQy6nJR0rx6sU08llRPBDnzXPWu+kQoFEu0iMdVikn70et2OQECuLud7xHeMA5jw
rk1AmE0u9vhNv//p3qjgTc0bQfRX8xcacwcPQqNb23FxnKka4TAeSYATS1TCsGmpi/qP3/dDl/vz
IQxoRBCRUbVROxFJURHwAdHfWjzWLwoxmc3+/f1uSa0aDfwliFpTbdzwfgpgB8lIM9cAtFoX7zU+
QezVLJy1a6zG0lpLieHyfBfnJbnHPiLJrXEC5HnEmcNyB4+XMqfy8rpKLBFnPyC9opuk6bjribTB
Nr2aLJc1ackgUkOkedYKWr7sjQP4JMt4rwCtqTq6VQW/caOwYx6gfFr5VCLE543EeKQWs3TouIQu
RWlzNZddjG3VMgkfqTvXwoDiFPzN4L0FZDW6ejTx3j3XxP+Nfrd4mPanvakSV0NZK4V3iO4T1JXM
deVus2+o8RcG1PoCXtIuA5MCQh7nt1J4J8eldrnFuHN5x/TMdbFKH0T753CHIHlTb9yZbCJIt9j6
mQ60+V18U5tUSl3sLrA8xC3mqfbjyzXw4Ksz6BAWHKsFvdaEdttWD7hArDUK4VYvGZcEqHW2fru7
iW1Dxiql2K8ohl9QOT2Wn1eyJBdyDjXoFi6jwyUr5qM8nSkzB3XeB4nskpVN2febVZmiNE/Up1wU
/payUxmObeywf5fngelK+CayJtB0xZfeoZTtpLirgIc+uKN0Ayn3v/b0dNx+T8+oy+tZS8zQj8OV
6Qm7yJgmdgUris4Z/ndXSWrgAt5k2qeCBj1wkchz1bq5S0fW3bB7l615MnEozQdAAMp3L8meCz8t
nX18fhCUptMbEfG4N5pSspTYLhggwzqMpYNcSiHlNLKFCE/Q6Vz83phkmYMm0Yjpn08GqB1batbW
Td1MwDmW2Tj4P2atWAOOB9e03IiIaqdOZ/Cfkmrmn16tvcWbF5sijzj0WtddQJS27vPZkH62Bc7j
mMgeRvp9H1rCRAeJuRy4MJGH5J/w8Wn3/13arYmxWlXgzyGbyllklkQUAViRhFehLHedOuRAmn14
WCWPjszBPnm3N+4C/IKUJmpOLSrRZmUeF+eJc107LPQ9A15c1ZL7BfltYuQNHmc9PUBV/Pg6U41e
TeqVkue92JZ/9GJjxiPjuphMZA7dCN/F4x0fu0vI68C5tt3Y37skCUTZjLFr0+2KyKzDELsSQU1k
F032Hkp4UVzuVfSVO6FFo2LwyEa+LdaucL6HmREOiHrzhEN4mqzMepsZyTPs92bikzaECop06F90
DAbT8EfIvbabaTBRTKkGq16eIGkSW2Udjijsc6zGwONCt731MozRb7rRgQ6y50q21icaSYrgeHI6
FjsGNHDi3rwODfCkbNy91ZqbpWGZeaCgn01kJKUMDTYLQ96HihhChKL9jxgNPnBan3vWpKwIemiV
Oe6G4Hm7KnRuhBGU8ZrKqMOegsM6wqeasTy51gNWQ6R1eyJIUaN/0Xpf+wqzgHnYJbPV2illlxFE
E8tkts7JJszetWvoSnr6tc9FIrqx3fxfC4UyH266J28QdR/O9HcubENQ7oF77ojdthGdlQ7ALN5A
CWtUQIF2Q5kVJwbloK+Gnh/ZGQ81AGp8XGMUUJGE4O8yqZyqNez9LBajAqIRHp5hMTvT9x0Hy+k+
2njwurDXdD04VE7BP1Jsa04sKEwEQQlQGVnM7cxMfSHUkttXAVBfp7RQlgQtFMQSrY7G+fuFnGCm
kmLdtXO7NaaAJ6n8Ne8ZwVw8YeEs5EZUe7028guuUN7391RlJaoLjMgCJsAJCT/R1Wtz8VkshV+S
1NZhAMG9Cr6n+90Q55tp/XSAPAwAi4ayuqM3wpNVg3OcsqTvwz+Kg6oBYH/PCqML7iH5R9sxWj3x
EOW53QqvgrzAsM42ePwq5Ojqlf10tCZCP+HGcnu5n1tBw0QElYTKgid31MdvkQ92IUQBjUO4mH4W
sBwc0h1J+q4Qpz0RMW7o/iecEbJC7qHjI1nj+IpSyQZQryg5Pj15T7l4QyS5YTupB7EGJ/IRaBpQ
B1Ynw4HX5f0CLi5T2krXTrsX7GC9Z9jqF64RvbcERnIgXzkDNCaD9xRQt2ezEBCDE/Ro51WQJ2fW
kntG1BWG2bWLefnRT8F4R+RunGlzgYemIrLhjH+LeZ1jMQH5NBcRtXh9oBkdL5Hs2n97OTIrJ8Z1
ZXrYnjOT6CMb8u56qGWfNHn368ifw2rZMtUXZ6NOG5UiWdh8HTEj3BsEiiCvN0NpJbMCO+S7LOty
4iRDstUnhfhImF+AExNkXTi9SkngqffdbYs32PEZ8EEQVsYzC25GWxX3groqDYgTcAomCnjyMHJR
Dxbny0VFsA/4WDCA9d5sTyckq8/gAnjkLMmlCAh4/Qycp5RIcQwnlAjKQujr2W88YQ9kKHnLJid0
RW5YGBOcaqU+zb/Y2LcBGoeP++8/QwLCFM9Hwk6Ai4oG9SF35hm9cbKKL2Fq+GKiVY3XrlgB++hz
PQ/kcyD5rpeVUapLPeTLnYgSWz1IelF0ih7LaG3yhxFshcTyCyQAX3d5xsF6uL7O6dsKWGlsFSCB
UtP/sPjQHEFfwyy9BVdNLkyE4uwrwyh+E5ps7W4LqJjMP1GqdriGtUa/+/dvBvCcp9mkA/kT7soe
l+A2fb1hcm082lw5+k5qHGsecfuKRQ31L0K8yOTps8ZJULcjGnSXey6+LK9PS9Qf/bQWe0DQcU/L
D0wab0f29jfZ2ECnXjrTLmMT+Dfm+aY5r6hvYeMYABUFh9B57iUaP8XLgVLUHsYh9IBJmxnfqFg+
JMKXySdTDfNUsQWBhSOQDJjmceNzV/GCDAlMePcgXPzIG2E9iAEyNVmPg8bTA6MKYx2xjDlOYcvh
5dwxyOTUtmzIEcBxIAvTPxu/q1Xlrp8jLmkK+8zedGweCMc8txyGS7PsamnI2HtEf27vGYCmi+H0
iPABjCnCTlXVvOZdnAuSuBCqvSM/EiRVOnPibRfh5eC5gqFg2pb+jvinkXsA55ZzABA54mUHuimw
Iot0cENeRYk99fTToBkXOoPrOUyp0cWcgkVA60miS7ov5aCMYzyY3d9Hn9KH8x2A4S2XYRoKgqSz
dXTOiO5qpv4e8Ft7EoKal5G+iMdiDRaBdsd8NXUeO9S9vnA1Zq2yHeGJzt8KRru2jMy5e8sfY2a5
Gpt2RdSxeUIgoByRQ/ePXCPvF1xAiurV8QwKfJMTdVpdBLsLsXCHTmkRK6QSxMLnALKEuTekyDQh
/NoUtR2Kr9PSPvvhYbvcT+C47hPG7ybF33mmNH/EX3eWOrmWN+vY0c8JxgYPSoc94bvBRZV6j6BS
/4Vdwja32sbDHsTTKTP7kRa4Zl9FlqUHlNLdK3go3DTDVuLvzPNpcYJUDdf21bP2u2SupHG3BNVm
P7yXLZe35jFb0feTgVc/HM0brLjD4czrNBcIKr7f0tFFSDgYn/QslRvuhMD6baernoZiVjmSbpDt
8zBC3tRgTleJsnolQnJB4GZQhCG0Q9Zxeut+ZXv51dCPBEQPifizJN1QbiNjtBHed38lfUGDU53W
mxnpIb/qvt47/96A678o0p1pflLzQ9y0EgXt8wW9taV8t+v+7Ou4kljJXMOoGINSkXmwuGxQv67j
dstsxE85CoCt+eIe6KphNEJVX7bJUnQM7UJZrF+0r9jRCO6PGXaNfkjOHky3qX54l93H20GtdCqJ
HcJPkjKlnSJAOdiMigDf7K24JCl5tqljjRKny7bjoRqXiN35rULg+eemcnnFS72jhmOab7/w7Nv7
/TEaChJDgYGo0G1+ypyb2bRyyI94eh4YoRP7Jmo9NovNPO/AkMDRlE1uZ5ZiyaWsluXijPcRsoSO
zYEydA3eVMWe16DOKA7saVhfTcL+NEEhPwQSyAQbC6a85Ka9Wmz82DGjLw35xxHDAxjk51wEoHnE
ulYqhYQAeqHfw8kvEsq2DpUpRKSHov6QbBnof2B4fprGfkzcWv0gpvm+tLtDWo4S0fBYtdxNyP8V
sGCvvAkoLFjLdvi8zSaQowAcFSR2fZ+y5jhUA78yAPF/KkKaVG0qhAOTl9wD3wx8H7zVldmt6Nzf
j5QzeSFvcbv2RlbKMBJdCnIo8MHo+eoW4tLb2CI38aNCTYrs7g85NYtDwu6Lt7/+Wx0Rvi5QI1BW
CLzVQ9lyARnHepPECgNtDBDBb0ASEV/p17rrv75RqPICkGrVPrg6FYurBeZdRMwk7nTC2Xl+jJ1x
dTW6vDYzxU2Z89o8opIqkS0VMDx/3n4K3uHoMAhUczes1BE8g5WNezRJQXoZrIZ0WqF8HIJJJBQe
10wEVUoZsJR8BTZ+0PvQwf9hYY0IkvAXiZPZwCsqcFeUFbG3Deyt1iib87/AdjCq3UXE9UjsRarh
hS9FWEWOjueKnwZHXkw2yLzpAHfeacw44lPWE9JspP/NpBjsq2o5e3MpqRYuQlfP2Bf4gRY/to9J
6leUOQoOCGSXGdsWdKgnhpPir03L5l81AJVBAWnXVLfFEu0dHQ5HBJkzx1OinKAc4e9eHc+8AU3s
LhPFfuDnoeOJVSqrAVLAPrnG9Bnhv53omhAY5ToVnIRNYJM2gU2NO8v50ZRbtXuaKAposQmpBJpy
GKPOiXBee7bScv/CQvvlMGNBIAFENzEECkoRbu/YVKKWBCaEBZbvPfPJWb2A1jQfPhUNol6micNO
kmocZCXN6iFfpmNvgKX6q7hB7ixvDxy5xUAZ4i7viMjZXLm23AwpgwhEdSE51Wl+g4omiVKSlcx8
FaU6LcinEwwWY0U4kzbSnHVjNyXRWK9MVgpACBsN+OEHvKRD7kLL8lgmx49c/BOZlMoQdkejCYU8
ioq6WqvlBw1wWTwCsBrqq17LgJtnxZwVE4LcWmsPsxzSnvebeBvFv7cK/tNFBl+vwgEbB2Fv4V+e
BgsoJwmjcUT2l/xvoyIn4OIj8sJqDyHbAIh/1qxEApBlOsb1+648Rq4zPb70qlrUIKfraYWoDv5H
MLr6PjgewSvAbTd8olCRNIvgu7JguuBT3pLVXCjkiKxs+KmnvvJC184hEIVoVim7f3EqmDwrY8sR
zErkjzWXGTsz1MebnXUUOTkuS2m7IcfFJepZl3+EtXjKOfM5mndvGz3d8fbwzBd+n55LY/CgTJjX
VQK9dNYkCGZykGHtNsvcTXTNRrXrGdw+BlbXpYdJElT7zi/HdeHjeOEutCubQxC9ODfQDN0GIfXA
4rvLQ9u+6xfu/nbx0mQpJ3bH+nw/Sq+89/9tD1j8B/FGFpn46QfYDwx3jKkyycbcT/uElDQlfDAn
rZOEre1OIDYw3L9k4qIx317osBUdXNkOm3CQU16aEuSSYooU2kmdXInp9B2d0ak24syvQN21jsbT
baNn9BfrSJfeHsZLZMarXYZBfHUj7I9CYuta39MdqrQUFEcpCmbtZb1kRZLFRX4OzPO1M9BHOxgg
gUOoBD64jxbeq/444bnchhgAopdc3WGkOni4d3AqciDs6atFCyU/mGOvJIbwxYYEt1uTNVqmgYKk
h3RtGTnv7iJHZwMWo0mlxT2Iq2t53osPxUSnhMxDLy4gvflnsFh4WlnhbdH7yopGfvtQ8vdiumpo
Z2fjyeZZgZ4a2+ohxrHRLQuXVy+n46/eX372AhBwcz+xEzVnUe5pVyfHegFFPOQWn4SqZhgskNrK
LV7q88RF+5nBPx68DlzpoJ5pHHy2fGzli3bdrZmCGd6s4GRJ215GSs2YGTArxQe1TN31Y4iyLwJx
aCLwhvPMRgIS+pUjDbBGW3S/QjMCRErqwYhPw5uo85ykX5xGnG4LJUDRmbNklwT5O8E7/X9N+Wzi
g+kR9i1rW7UMm7FgFvXDigf8ErhsXpI5u1KOctfMCzQPJCQue6ZXXxsEVRy2m+ID5jFGtO3bZ/uy
vBmWLkd3FiRcV8bTLGFBD2N3F+DgNsaHyf0kk1J2RwWuc3sL+TCNgQNRvQNsPObTjDmUD3G+fYyI
wS7as7AcWSmtX61blwHAJkiNEr8Hbx3acSpupszT0oCwp8I3genkYsTwmJjLOyUi3LP0K3+Wzy6B
jkSSnXWn339ROIwM62KTeTFQkghvX3YCKlPKocVqqpu0xr2y8YXHlOKgYqCdwBR+tcCWMp3tkyRN
GeL5+ny47fGYboWA0eo7Cn3WgppusW08VxVDSOfpi9Mhl1PlCWosZLSGZQWAZ+HkYTQl3ue1jrCw
E+EFzlP+YpX16/AprEtMo7Qye17ocdLxpNW2QJcW2E/zyZb14sWucHYWzW9lus30zB3x5ksg2MJo
uta+NmqOZVQwVSFcY4D3KMbGYL3n+2oDDv7fO2R+QLdUJSikUcnUcu0A6A/+S46Hxuc/P00Hrv1w
qHIEpKB/YxCAXtEXUxo+luYC8emN1YZoAXWLxeyR52BVWWGvnM0gO+i06U60EGu12immeKDRmFbr
wN+uiOpFNs0iR85u1gzaOsgCxT8mSU59zztayWB8IQN/pKTDSv2ngx55jyav7WJBMWZ/cKWMnwpl
MLKW08dLEmOeD0LjTcBRc6qqAbcRrIWByEqdUk1ycZlgcYip+k1eaMFAjrenagUfREvqJMadPGoD
SC2Q+UBroxwv0SGm8k57a6k3GtTbUDW1XvzmCsndxhH0FB7pQ7Zaxbrr75wDU1tG9Xvh5T6KYp3w
m//rNBRRvhh7c+zWKoH9KUpjDmf2DWynWM+AhwHmxeP4Ooc9INcMQote/EWwTLOTjofQvv2xHgxy
UFThFxra9R4yx70CfOpFZ/hZHJ4uHfNkCAS85JwWl6YCTTfLQTrnd4pKv3VU9FWKz1MtbWfoWvCH
2OQmuC1adaUZN+amltRN1DvSW+ornoK5JbSKIE4yiVYLKnrVLf+52/uqG8+2C81AhjCdQvnO3Wu7
nazFY2mqKD2BOO7Jdeh2okYZgnpXgqFIjAeVjKcqYm/O9+EO6Kqzf44v5Gv02w/VAS6t16lGjK8x
FBB9jyUCt6u3se5KZlQLQ9zbVFEc1WDp0tnj4QMgZr2N/voHdmCJ4s7E/+vjV+iDnTzac6FOLnYN
S5gnQ7kauOmkaA2EdwFKZuTE1OsD5wfDgSPHpei2jqEB7GOuzFfyyntUezVkkmApiJPBljd9ObfI
eyh7oCzlsurzEkj/hnUcCyW5LFChvlcwuGMt9quX6zBKZTbdPaiICzJI1mg9uV4aD/ORUeVOBesN
62yBvPMMgMzNdWuEvOuNTkgHVSKRqp8VyEKm7leoRZeHZ0s/O7C0tHDx5AswI3QYWlGfg1boSu0J
CvT/Wi31kzXn8MA3PAAt0xOFe2RyFPjM++RCjTf4e3Kp8R607R9CoTbSzlYrEiHgXbEE6OrIpS78
AGr7DrqMUl+LbvUk5R49q6MHDgIMQWPxf8YaL5ydJvHgeMXWWH315xWfG92UxcqsdafUibvguqTV
R+sQbyRLbfyJZ2vCic3kk2p47M48Ap2dHbvImW4SuJYZ28hcbwgNRj17vCAf3bzdjA4EWprxIqsS
NYgPKa+elJLqQ4kO1U5Kja5DjZasmf9uTyUppiwqmiEyqO9s0QszWdcV9c1fbbq1K7/9NcUiHsay
jbVmeEBW4fL+uCVgTeliWXl1E/hlYtiq/uz1AWdGWs9JNQ5CbZ91PK1rsgItuRFeju4MY5w6bKiW
82CiETN02ykvcrCgjSFvqla42D96nBGKId4EGSHtqtx2xfxF5MNWqRzjMA5GuSYfDju7dnx40M6n
l2jXKJDDvi5UciMxZjXbM6cAbNML6y/zokvMh82WfUIVGf0uIwh1+8Drsj4zD4iDAABH1LyMJloo
YDJ5omUhjC5LbuHwAZy8P5GFMzTk7T30LlZV6aZUzXP36k1bLrMyxg2thX/Xwi/sk7Fdzuq8j/7S
zYip7AqIk94OSh831yyhvATym3T0M6D46e9MNaOP9mrIEdXqTz5/5sdSx8Gl4TroZhsUFUMT4Xy5
pizSn+npPX7pz832KmmvInAgxgFWppisT5ck6XRAxX0CpJQt/5wFVpu5V3Aa5erZzt7i4MY6HCjr
gYkSmCeVsZM8mtnRVbyPpfRvsZsiqoLEZ1DMXdwZ1aD2tvS+8/2z/mUXj2xWbAS+uR1l52pWMoAB
RfCCx5Wwn4TJMRudXcyOwPBNio1B3xl05L08SBpbcQ67GrTIfX0Tg4tjSOtJkyacIzCLJGXNbE7O
m5LNxjTc4DK7K946Qfhr3p/EGngHmyFpxMoSdcDSioCcTnp+wS5/Ou7q+hIxATa8g3Ah8iSE8bCd
3nMa0eI/BHN+6xcLiH0M7hPWpZ5E1GU2z15Sn/rCKZ83xS1DQqr+oMlKfdIEyuWCEyA8jUDvHlq7
pCLLjBQEUiJwWhTPnIchRtqKc2kYqxKLI/+ptULSL/wOhZekGgTKTy6jIE9Nehx3Z603tzhOfrG0
DUIKnGwcL7p7XsVf70JhQ9jXHcG84/bHISyrSsonmZXLhgM8wnDzs++uqBUfRkUdkBQ+vu7kSyWz
SGxUVN7l2sFlU6PhO/S3fKMKgnT4uryt8khUs96W2+/xVs5/rJtYi+gQLXVkwcwH0eUUDDitcmTK
N4Iqhh0l2ckB5F8Q8RfynxjndVwKPfYxmAfnCCvya4E20JYTMFNp937NBguBoovqf50DwkHZUsNC
I+VT0GHw/mGyd/01UbEUImgjNEmME87iV9jeI1QjaCMyZiE+WU+Z9bXekeLzxlkEgOZI50T54WGP
aeuhb4J7D947s/GzuEsjwgN9NYfmnFrCwu65WEtpQ4oGulVVGhMYJn24Z9+VeNlU4emshzi1cD41
XTpLIvhFCihm/mYyADALa/rkeDEk9HPeeXk6QZeAwXhzDME98+kyoAcmtciw74XAHbO9wzPYZWPJ
t3aKq/aSL/GE2/TwXz6J5h0SFvDHahwzP7k8ytPs1LFB0C8T33EVESrpHB0befFs1L9IuPrXN1In
gPNguSReuTEdffSwGhj+QZ9ikWFEFGyZVnN/O5pWR4nUOJK/S0VAd+OvV+UKh6/rZmueP+ZU6QHq
rTiyTBcZ6om6pBGKCOrKkarHfs9ul5tVoOFS1Rr47DnCts/6PL8AKkiGddHgzpIFFnGPp60psJQT
n7mfkm40+Hq8etwn6N4mCRGHCoKggGymxNvSMbP+pwg6wCwsEJ3MXlXDrOA5LMCJbJK8JPoQvLbc
ZPDwQvVKjFsPrfI+1QNaEh1YeIDfmdYCSxiN4606+BPf3B7v//jKRO6bFWaJaXGvW7IZSnZ4svoX
S7/lGXES8YwcjQvxoY6TSf9K32BBdkA+UVX4kM3hM4hozRBJRDpWka5mfslRPNEe18DkN/MJqAsk
cERFtqYC9FQjbrZk3cvWyUtzq/agwdht423+IN1xCHb4lfK9qaPKTKeLTJ5sgQlbNM/huxMctq76
JLGvACwNeNwnukCJTFu0yOMIJ2n6dfZxu3Y2AkDVUV+9E97B8Xk1WMM4fnqwE+GubgceetjnYa+a
wCpMHOwMsmzUDBuv2yDCXSNv3PsnmpUelkDfhskpnG3YuMHBE3txFA/1Djl/DeEqixGkpfi3UvP8
FzXp7dbQVmarYHDZIA8p3wUwjTUdhCRdiYXkldXrn6c+LLHRxPQCg8bfiLYEUYtIFkCDwlW9OzTn
4ylYvBboUGmHDVtSiiwiFhkRjFvul+B63CIQC/EtAi87l0wt4tIm0Wvk1vnH4h4MUg8By50zgCEA
ihT28fGlOyQVBYaOPol9w7yxpKWz2RfgiRO4fIdAmjJcZe60X77Ws/xvvKActeRPn85HiHnFJGi/
cUQ7L6ChJ1WvTOdlpKnOn78tfkrqD+HAoky8CncGYPBZzFI52dq5/yWCrhBgKjdyi+e+OG4+W3eV
/BR+8dvQxtN3aj/pzQI5+YaWIjnvdQI+NLQ+tZ6iAC/iYiAtCp1IM6u4HfMGhVxNkEM9s0ZHycOP
DdI9HNrAjCzLVkeTyvkkql1Wynx0BAsJF0j6+e3hutOHXozWfGVFmGusU4pLnCsehWBBqeGbeNVg
GD2+kiAZxN5pA5B3Ja139ukIgbe37myCoV5ARpKT0q5/eIoNjaZ22LzdP2NktbEcM9IItlUFXbEm
WjXQFEigJHd021/7qxUXQ/LTqmNXdMO+Ci400o4vUUCEfv+S6S9fj1e0w13nkv1xBAEZJWaYuBfi
iyNz7IQubZ7xJ4o2e9JZ0bjiporAyH0kctadwD4sORwEEkQ7h+N/4KJpdrLQmyJomh5zQ5wcbwQb
P9jZWwW0/FgC80LqJgaKTEF2hcHQsW8sQYi5ZJFmT2t1e5XWA8nB64Qo2C158+3Lkju9BxrZjOZ7
aC7MQWl7yswKgfe9JHTwoi1pvlIIPjIyawHkoMgkPLcgbjykRPih3+/qRhnG9bh15Cez02Ht1XpM
wLr5QIJ09gZPtJqGS4mMjbBNaAPXJ0y3VcLuLO8KnjMUZubwEzKjYDUrL3ZTPsnnxijaAS+GI/7O
ObUB2AQdgVA0jPcNHJFz5wOiUnMskRLTkwahfoWhGEa2oAqvROEVzjIijm0RaUnFxX57GCpU3hrx
piE5kTAcR/4kQUAbLOs8BBMiGUQNMJZN9IzwslLJDEgN5O0+HwfISZRmispAssktA7EtMqtnc1Dw
JbzXj/f8quv1X8z2q2jLAblPBZSqogiUVo7Jzi15TNbOpqFVl0cQtjyJGKB484QClemE0Du4eO83
gES+fs5rdd7jH0EUOc6/AGEzP28k+bYg99VViw/ol5xaSw6MLHuJt4UQ6nA2mBxWQw2rwH6hzDfO
20WOaPEVHKipXeKi0B8+3odYeAn+dsY/NF/I3jU2TJEKK/IPMugqs4QLpAuUVMGnt37UsymzO7Cc
EgSfiqy0phcu8Lz4ETtTFzdZFAzIhXu7rwY5NYkLWMZVC7aKQew9VdK02ex9YknGz+zK+gwwzyTf
QwpKRn1+ghcIIUZWr9V7Ls3agi0SYXqaa/1O2yg0Veg/2XBKOzlJc3gjlBAl80mxI0BBC+x3xz+y
ZTadN/JZcTCpySK49sc+skSgy7VyX0uKufd6z/QKbgbWhgNG+BskeBx3sFz15HSyMlUEoOPg92HC
I0tc9ySAuC5kj9C1XjStykkNlKcMX576QW/ELuyAJTh5+tr2Hr4p9b0gFAO8o61pu4uomKzKK18N
108hTp8xrmb7su9cgVEyC1foSoDX+FOJpR6CQ4Z3nkdm5BNZz9t9lLVt9J+6I0D5FT8SWmu79hnu
8lk62OyN7Fu9+EoEc2x/gVmQITl1zwVYTPbJWVNLYDQcmTuK/BmHUOheflo/UKkor6MAkQCoiSAi
P4zRILTnSpypvEs0B0HwkTWQjnELyF+ybM0+7sU585RfFR1omlWnBLzTJ2nHNlnBp9QowZa41ivF
kShZnPRv5bvf99Y55wvTrVQVIieV/SdCBHHO4fSIsZax79ihKgc8B3mHEOZOWHvY/hdav4RfQEWE
f1mkPoRaTx8m/0aNE7MmUyf33p5MYB8DunHTTpx03gG0MwzSX/HchsW1A/Sjhyvptg7zJFia5LMF
kq7d8I14FFVICkltd2s74NoFIOkx+AMgFTIiFwI+OUTK/8RRMGBb5j9qYOku4bBEZs22And5mkvU
NJYq+jSJcx+LjV0aMIkfDfzzgqYU2M2pbbRVZeMO9ZUZjSqsMJq4iPYKA4hgwXe71Qh4ERY4Od/E
T0AabvebZFoQjDaTR323nnYieaBNQHw9f4Rr4Jaw6e+ITydgyz2RFc5O0Q0oYXzzfIZgmtln2XTt
Ni/23qlrUE8vmo9nkzHQA84JHtCI6TRUvg2J4uMJZ6wbMj/icT3S4QrFSwMKeLsE6N7OvZ/9Kff3
73FeqeZiDMp3qSA1li6r68qJFKgGyo5iNQ80S74GRc6dh7rNFTosZcF5dZkJBGmSut9gFcZ4gAUX
f+z1PpgHJy3wcpRzkODMY3FMqjNPn/1df/vZmeA9M+MX13Fm30VttRan330LkIfMUI7kXaz+pkW8
HgClbQscjJf4XVn+H69rfooGeYVhZiEUIxk7PhqKYVp2DfRqitNSWSE07UVCMS2HSdXcmrGMjzF+
mWdF3hcAPXKqPlibweRc7bi8t22Gpt6+tZCyIOrXfzgbIoRvw8Rj6nwxtbFZgv67HAYnzKpOB+wC
Polf18/dD+PtcIDtwKNYEidKaLdMA0HA1Qs8AkbV5USUz2Pai7F+OpviWZVFQ/cgNmOL08XFmG2X
zaNTd00xtdIAqrQzmiXqM33YAKjtpOXrY3QUHq3HrhG7oUifIG0L1IqEteMaQyGTk81yuZpyNfU/
CDE75wgckP7I/tW2jiL4+rocy6IPALfqgnB2/PBPeC8axXUobrykfxREASj0kgAl4I+mbO0KWIPs
l3GM3WmfByLXGo82YdriSUVA1YgBr/nfY4U3KnPsgivO8wal1knYjSWbqPszg2TXUr1CZ0d2INHF
KXkVhbzG/4S6A/jfogHOqdMglw/nDg5zTa356k0eoM78jlJw5X8QJFtdatCDlDd0iVbUGwCtDI4s
L+MpmO8RtFqHGL6Es0y5foogiS9AQpi9NveBXoUQLed9kTQL9vP5FuBFyQBg8u/mypaUEwlGl9Df
UUQonEpteYfEVeVdrrr+akifqWdGqRcp3vt5FxCl46HRnEoR/hYzsBbw9UTEH5Uq5iZ4xk4bwhFV
SORIp8CqKXBRzfLxC4yYIaElncwG1YTLNnie7pVPQIvY2tqBqZumgt+Wbut1e9o6qPvgET9RjXwy
jdbe5DYsIRsypaLl8EFTmGAOQ/BuvUsGPKgG7sWYrUQm1YpaU4BmAz//da7wC9CzuasEHGmq6u0v
aX2fECBr/JoXT72FTC6riOajBA35CyhKy5XCKPWH9/NRta2jLkDCFFMsrCQQ4XQqfJn1RiUFUmbM
X/PfwfBkCks2uu9N8AlCk6R4hbpx3J+PJOopF1C6qkcyX591gyS27dCBL9U0dNCC6TYD27+LxwNA
UHqXEm6OTnZspMORS7IJdm4jMe4HoGhh52iulfwFz2nfrFN74M5b3Azmn8rFwNqlVJv1yGgiFTna
Ruj6YHSABvzKwV1uX0MirnXPY+IGfTKka6feGOTVlciYsa6avv7v8A6/VgNRa7FdvuW54/JAZxaL
6oYO5IXXypBxExzvVADXkZ4DKRWtf70FIJu7RTYpRBs9SGqea8a3FdPMIsbwTofMEMq5BJEtMNfC
EGdikMa91oaXIfzLgGv6BZBnSLFKlqM9D1a2ybKoXUATcvsFxjA9QvzPVhre99MbGnlq0cyWtYsi
19U+E7OxT9NHhg6CK9tiHIVQ9nCEStC7x+8yBTBYUGPHjES+R7HC64gT3pi+ii9dqoIyhuahOP6V
dU1YzFosHkb41UtjHxBE/TDin5kEYIgbKbxIYf04NGLy0NzTrAqYmGSpR5g9MT8dpHoDHb2iIeLP
qz/wGEWX4x7uvfihtYSeBFor0Zzzh5IEnF/Dh1ojTqgPoaYK6AsZjGWyt0VYuaokLjsT/6HMRTVW
RLQMQZGHFLAnKPyMZ1+/oiiO9nWrf0LW/SMkZRqNyX6ARrEdB/tJ+IzMMRI2XLBO5IjMyZg/ykUD
QG+viAcmxzKcpDAPvKu8jwWiX1Rx13/BTFu9l8G5Hgf09gbDQNowmGmFru3MNbklazJTe12hv5Br
+f83gRf1fwCO9GXoXyX4WPNevsHAn8E1jniX91PVnyeaDTOE8OvRoqmPQTRfjwZh0NQodaaAdi5r
hZ3qFZ+/qr0HJ/AnshYvF2V1pwnq/+w17Z+CE92irky/ulHjgV4awj4ahh3t3kXM926vqWD5f+v0
f+1Hlsb2AKPujdoRTWTQ4GaQ3W1qtvgPskZpZOlMzyxO0tI+yJoudzOAK06mzPil7pfkLDiqio0D
kmdLBpMGdMEqh3E3yrE4xIqrhYoKQYhaKVt9OdD3Gzt+CoeBoTFMQjuoHV0Acysg4Jc0qGCFWx8k
+a8olyqKRRI++69FmWd9q2BpImZbaM6h9T4wSvnfqEF42YrdC01OTV/dJqIogyjWpuFUaSy8K3dp
ZIkOHpR0hVjc4rsh67XiDYjQwjOjDTIHfFZ182EijkUCipcn+x7THOEMNCnOYx19uaCdSMrlvwlu
vjUZoKUYZtL10i+zs2C91q0XunODgBzJs/4yjlgndfsSvrXJ9Yb29zNVv6MjEFiSwLgalPxjj554
5CQRC5I5SLRRqcPLFJXwge7XPf5H4l0JkdY6KNvMHDoDQnBydupBGAgzdwejYif1fn41LPSrpzIx
t64ODbuxHythNVR+xSWVBwGh0i6aIeVmMjHpMCEY6BAuqXZgff9mHys6IyXAcUqeu10W838oCfzI
ra+5moEUSYRsqmZkvRjh4sAphdD9Y9RaNpZag/FeRHKSDGqZrpvOP+MaoM83BrcqFWzpB9Be+viQ
oGkLzsLYxzIxfS4XPrC4mVGZ/tEwm/GI3dtJCQo/zE9yWzumpGVaz/rbb4WNdwfd3Opme8d9iOCU
1c7rSFzYTY0N5KpcxqIDWGXWY940Z+oACaAZgwkbHyJCX5vWdQtpTiL7E00WQlO6FTS+/vzZh88b
5UL1pCiu05Pj0DeaeKStEnzsm0CAsnfKJBeBtUndr5JfOP/IkT3OUwlGW8xvvy3GoNgRyCeSadSs
9PYTkz/yOC2kNKyga8X/gSCGf2OQDW0/ubgO9fzgru3598LbmJLmNFUtzABShsMpDUMzngi5KcWh
FOKjTACXklSRj0Wv8bnL75GTz58a83PEsxxgum/7MRSfKtfO18v6X55cCuFdvHqN7nsXaKVEm6g1
7Zz8mN4yTJZ9X0YrZP1s3w6Ozx5N+PIAencauO5HJoXRy0FZdmLatfq0xUdQFBCd1VMcCJacTcTl
yrEGGeE30kEdP20nSpkgbWUTiIpcs895gaRzyU84Cg6P/l7P+tV7EKpYDCXD3MZv6AASj2vOLZ/M
68UtcubxZERhYhK/1BFEsi+HuBVLhhv1yPCTZId2GpV+IbeZta5qutrjK+pSyUwlCe5sLnVsG7Al
gJWGP7tu2qe1PH70XPK+1raylH2WB64d4B6eCzCUC1BdjzG1V0PQnxjJ3heUQR+8rgI4KXz2zS4c
j5Ym7YVY3NWYAIGOISyTvhOHtp95+NHhEj6tlsHqDo7rWUEZLFmIFddRMFzJvNlR8umi2OP9gahK
M3FsAvPnaCcAHsl/vpsyAZpJn+GSjDhNvfdNEGXXyjW43yjdemra1kbjWdZ3HMnycvU+gxlVOSdz
wAFoSsjLzfXOXH7ULqfkPmJrfMn4jyqVwN3YbtppmEzt7hggqTLk3gt/g1u9KRUpDGWTonMVoB6d
L4ilDaLx+QWCLQnUMH5uJj6JhoF+SAuOaoiYX+azY362AU5qmrCskvQkpIPu5TulNz6/zqzA7Kx/
CBk24bBeTYHSEY/9uYZnTDVTmM2RAVX6/F2O3xFGztzCOirxn9iZ/2t0A+zVIsD6zKCuEP5BRsgG
Ob1jAt4eMebDNfOcsqYamRfEYMQDLObuwwp0kFmdDNyEi/0YK8tVeYq4wmb3UZr/k0842xYS4+mX
1jc4QW9IMjG+mkAj9XkHlerHajD3NzfY/YZN1E/+CWt9oG4pzjPJ1bFToy5YdrvLWbDmCEOMhfAZ
cZLRVK80H4g8vhYwkXrAg4lUiBiwxBBeD0Ox3l0z5gHUFWD00Br1Ns86kEo1Curk2FjNC1h0pBAN
VDdIKyppM/VlQtOovYDfpZHYHWH4MEOq/YuxjeKQq1QK+YcBsyAm8mK5WKILmfRs8DeDQn9CN07Z
jl+f3W+6EGOgN6XKdsFkTo/sZu88U/au0676OseErM5gk9C1clqeVAEGexcc0Lv38i8n3O39j951
55ctpK+haY4ZGxs5RsgWpaawTFFJaO1S6OgSwIguHXC/7GlCUwwzpmCstxBq5dYur8xt16AdQVdr
IxoGaYtg2QFGYOIZoGPHXqmFv4isBqcU10Nfw/xmQkeWizzpjnWcfKZFMnsWOIDAvHn/JwY4xHNf
JiKXYCOmxtstSLvUv4oy+9MIH7vUt+trY4ynUFnRKQ9ih+3a7RZXqoKDReqNHUwgYdeUa1SD6qhE
Cx9SK0lmdRo9cJNZ/VXRB3lf3fyXPj9Zu8RjpJRTgt+bWuTqX6JIUt0H9K2C7XPYuqTtpqesFDbv
RDfkhLOzhwje5cZRNfgAXHmgbPkgDHrQHobYGa2aSHF7dlgIBTEYI8Trk/GcCfwlIYIkOkStsYlt
dCon0DgALLIM2KbWmqdBUZdObIyUYMzCfWVWS8bRP5dftGUwk++RlLXgFEXMw7wJQTAttwTq1e+C
Cwh0gPu7U+ofw2reY/DFmzf4b+OSCzyaCys6eB2aWeJCU9PEOLo4owMSQhdEMLeq9gBKpfSt1VDB
KddL2p/zjP5xmJrhsABlvM8dRUAUQw3IJ+vuEw5V8frTmSzhO0U8AKHE8+ozlQgM4mLCcZDZzU06
4NMWSx9e/6Tl4ci46q0sRRg7Wt2aOLiKdq+wnunsVAsTp7DN3YTLnXagqiKDlRt5FPrjruknmP8L
+oWfaIavQSNPK/+BAfXaBgODznt+iEe4A0QPn7lX5KfkvYNZzK/D7gyyPCAbeHE2Vv61zgrt58Jp
5jaLaO9wpf9TOCphvbl+NZcTwV7gnoVIqk/FKYe27GlqFJaRxCPvVfp6Y+Dmhka/Jgn4K9CyfGJn
ELgrymzW398Y8YdJ6ykmjk13RfH31goAcFnqQNNoiQfamcDMj0//o/CpgBiSLxjzjKSU6NOzfzAf
rNf9Rq60KzRRNkk0RGy8a9tLZgsYEcybHeIzdp867WZ5k1uvN3o86dkPKZdsPhqC3srPr0fj7m60
fieV3vWGtTkE4CXXsobi/6WIJttp2O8GRXTPwGx9KFGGpeuZfNtusT28+zc/wvEJ91zfDaSHWjb1
Cc0i7A5sXMvbLUSA3YuoXJiVeqDQZgFSAgHi6rsYqRnaaknnTo/xVR6aJRm9Xdr6ft6u2Ioks4py
/xrXQjt4XBw4awqO3sSTAI6rYoAZcW6RI3iOmR8dMfrFaL0Gc+lxqL/ElsQlt6P4blqF4lf29IIZ
4g/TLhA6KBIia0xlzsEXTUM/b7Ec7NIURvKi5objq3rGQ+sWDnZj05/vC0abPXv3BnUyYffXu0c0
Duxnvo8IbX4KGvJQy6wQdb0uDKgiGdJKLtLBMqw068LNjYKGdXO/o8PZjImHBhxFntQAx7N8w0Bs
4ucsbEsFR3zMdnlpEbhHLgMRu8upID7l/2xiGFpXomSJD3Kccld8CjRXz2D8g7WkZf0AJVjcC3dg
XxrW7Z8StqESwksjxGisVeALcPtXRLcWPp+HFmLvjPFmqr5TxuPl667ZUldgYJ3ezJkuKvdDNPxV
W/TzWRleWK4l1H8HpShV4PvHBIx/zA07V8mcLoJZYcDkEdia349Iz6x2OmlGOds7bf49DJPpqPPb
bnBapePo2W61OwQ+mR9uNGhKXNuYgYU+clL0H7LmGabsgzDITpl9nF4WmhHmNZ0SXPUmAtyazyH1
ANVBd0DuhXonK518wHRqTn0eDFNN+aU4ybgduVnD8AymYhAUSg6b/WjTPwUu6Ar8c4V6y008IhQX
QmsoAVF0IT8LK+2WNtvh2EL59ZwPlwgrnBuaM9y4NnUbCK06fiJOGiegHVXCmEr0ui8RcO5zo9S1
R3Ld/0rVtMUI/fGyMCLfsjla4ELLmSSE27v6dLFb6yzXtIeDsiviDGoiYyUKNL1n1VMyqMj+QyQr
IUAwRYgLZh2mvBnY0nXD5HCPuFEDVYzyVzrrHwvpK61qxqnTL9KvCK2/sE5Qv+Ca1f7ZFCnvzPi1
5KhzbiyWtcdKQY9FHBkmz3PHPg9VU7MIeG1BZ9PE65vpL7rpwYK8bTiZAEloeSDD27COMXVWlHZw
5QIB5gfdIA8bs0/YTC9SbM3mlCWsxGaL8GP+V0tTEQli040nW2kTw4oAzzwOWBayyg/jTE6k5WI+
oL64I1TeA9G3uzg0V53Yua82Z6JDMqVXXbT6ao7Kll5f7vKg45MP+cl5/sX873zJ/v1GibmgnDEJ
6TZfYJ5Z7DbJ20K+rruiaucVFuPLbQ/4jAVpFoTb/I6nLgee9xX4QkcWoAhXoQf4gwdtgUIfymWm
YrH6a2JJ6wo7gX21CyywVGepJLX4EIiKjfK+TvQ3S5H/42kTaEk9YZqYHKiPo3wrZ3F4P1yzx3pc
OYp66s48T7V4qbeci5X3jyxrVLoPW62gQ8vBDyUG59VbpajMViRi/f+/4Zadq/kYRWkGvPlgikgT
QUsjLp6pnsmTsknAEDvmFe7Pt0QQyyAAI4IJByECFdzXejmqtQNPKBIeCdBrUBAW70ZckW3ozke2
rMFPZmleywECQbTJRqJD0JkhGRfSkFX2yrIU/5OTf3kYxMu+9hsINz/Itvyh0strusi0r2SM0Th5
cRp1U96FeiOlFLlclCuFJbo1a6f6kVO+PaaNwRwC1ONv8iomtayNqfiDjk2Sas46riJ0IytSJwNm
eDaJZFQ8ocp4O30WWUMJc9iDSwKFcrgFTSCAGoiktTUWhbpW69ml2IWSxqthXq6BpkeVKM/p1a6i
s5jStXmcVp3ado29uicxbyUiz4WFRfVHbqyJUlpgbRyY2wqzRDi2iS+IFrUW5sTcwNSb34Vtbj5j
l7FRrwNhd5xLHrUFw1xEh1iIPwlytPkwqZt+k0zzh6n7wbm0D+lzEtfmkCue+VQ1ZmxaFFc+adOr
m/duModDXY6ruJhY4Y6O+bZwJW9pWWYrzr4RD0qzaDbIT4n/LDidMIbKdbzWMJYA99DFeiPDQ4cg
egLIOwUmyImaJcOR7qAcHQjnZAT5cI7fxErXOqy4hKojXtX0o40z6nwaPBmOnAfywTMtHbVp3Fn6
WlalMnAJeizCHMA4SOAw5PIWxuc964tn3S1hADOfEGCiJHbW3nC8NyF/kgVpcegpVwESlSQlH7Ri
NVj4jXrn9QlajLoT9P3HfAP4+BIXW61u0H0C6uq1JZDjbPSwRXLR/XqEf0Rm9OuviyIGnCyTAotv
/ZNkMxaBECrof8A3DgJn44sQwL5kvJb813N8Mia8fWWymrg2JmwpQpFi75BegDaJ1oWghwDanudj
S/7KONx05quKMl/7eweruIrX9w50lnxslDcg0jCRS17oeTtoH/CxXuC+fkOxo+0906SBABrbbxOS
5Uul7n7R8Zb8iyud/1bAoxKapCvIfw743NN34+9CnUqYML3hr/uAcp19lnSdBM/DElv434RRTixo
TmbfaLK6fA3Huk/IsWF0vvweoXVkEFnydznrwKL+MeCJNU+wU1pNEfVjzwW7JBf96Egvr2/zEqas
drHFNg7Zwc0WXF7pRie07dTEAKw0DJwbZ/HqSHRKCUgQIcBS0qhk3EROSlOH50/yVp+HAhPdDaYH
aiRBlzq8hrD4ruUsvPOU0rJ9rrVnYT/aDcRLCMxcJyhmPpMhtktPNWJ+JN2K+ceujC+gxsQCNtWu
9YOc/ipoVf6DfpFvrHBakyUL5aQVQ+U9hZI7XD2tVD3C8SCuNdgGvt/yrrsdzErRRVa6HKhkKYLX
Ey/u3v//lbAUMKkVPIBWkNRmYkoaHxsefzH4tTe/fZfNdvu/ZogkGvQwRe64RIcnm0omyrNvxmbG
hpwTgNQjjbKjOBvMT1CSw3xVnZ5kXcAUQg7GzQCC6oAk5kQAw5f9NQRsnYL9/FpZLS2EOhNpwo5d
rkvtJOMFCpxIc9irxGLVPs21BkCiATT3tnxSMgSCYrs/gw+zuQdPJx8tXJZQRH2RfPCnrP0X9B1w
bFX7By2jtLYaRASBbfjGjWyztfMoa0gbmeU5+9svTWRNQkrWIIbJBY8w3tl8eFUH4SC9uENLrKQR
OTV6guX9kQaqU1Oa8A7tMoECWlZocBbPdCr2C0cg2b8LIw//DaQJSMrYUdl7+mpNLvEgRXCEmVwP
jtv7AcOUnUsgi7VvrUVsD5l7FV+WhfCXIqTEyLVDdqkogkcF66CEfWvEfHkesaWltF7w6EWzj0h+
5qs5MH/Ux80vbN812taj40f5cfcmgMk4TlI/172jaiwh98Lt0nAzCQjIVT5IHJP91LVJB+614SfQ
+W/7PwI8SyDLjpUcYTb213jLBjopQNQ7EF672AoTEJA/NWI9FwIUPe1IEgDNqt3YfXCxW6E0GABl
zVx3AFsuTYwJE7m7EOmwnLncACYMaxp6yL4RThR5idw7D+3G80bPq3V2JtufCAXI1F4Q0oFb02JY
PGx7jOn/E22xnyzxtpjMCYz6Q7iMyujTckt406eduWU0VeictHoPwjLnmBk2WsBaXTPJZ7v4ODq9
7PB5+LAITUTzdFaLS8PvSyT/a4RK0Kpno3gsJKodo5XX0qtbXEyFq05yrYfseNLl3zw0GfUfPpfh
9R2tWQydNKGT+D58SL6ROXM9UW/AAJszNU5PihEzkL/74wxGgXTWOjSajMr1FF2OIrd4ZliB0G8W
TIjB3NkkwWqelnY0Hn0onjmbVsIMMLjTCYRaHo6qi4TSCTsuI7V05N4SEVvi+zGz1wIEXnoR5hT9
+S8FziWCRMPsWQSL3jaMBo5mbl0eycate5NVjla2ujW6uSt4n4oDTYaFZGEu0cG2+U3y0kTG9CwD
Fefe5SP5Jd3Dqdh22YkKLiAx+arXHNnJvSI/69+vn+xAgIueOiK1C3k6LKFHx5b+v4CU7oAsEqfU
iQ1lvJYi3kKFrtFlDHhOFFDaLWqpa/L6PzCI7CCDcx4mbGIxHB7flqMPcvg/CA7Dgai+/hoRZ3Yn
E9jeXKLsyksA2CogAogi14dwZrU1DY6ApqxkKabclTI1FmFP1BtEB4gGgKD3+yIk7SwEd/VppN86
qhz1FfKQn8c6hyW7UqF0jojhThJxNZBSiMI5tdxbVaH5vFnvxeKPL1B8/6yg4F+r1FMNi5DHohBf
ZYH/5Rl4ESsFaFeNGo2D6+as8c2sx42La42+MBbjLdGJSqleSdBNIVJSM0Kbn/a/IDGzJlvomjRY
HQjXgaOVDniaQFS3ijiBSx03ETF5ZNLfkMnDoUjoY2buFGFp+WWrQK2yuQZZqky/zvTthS5gMQzA
k8T6nCrL8OzRNj2NeQxi7zzhHAlT+OT1Zlc7uppPa3S+vb8S81Vr7X/CiXtuyvxAWvPEDni5dwLc
VN3dmDfym8Gb/r2ypniI+levareqB0RQcIuklnshWzA17dzXEQu/L7h3sGIVTvp68WasWe+5VAhS
ZKhb/+ghlu2J/CgSFOujEr81x5nZfDNfoNNIzD3VIOWPUH41zO1SbHtcHBqY1KUdXSwSbqN049iI
uWHs7YIIK+4WY463HdJ/WO27DXNrrdvJw9Os61tRrEjtuUlLndVzeH5zOD660O73Qj0RKDtSnej7
Zl4nLMhsbRkm8kzuTaFJa/TGKcpJbAaBJ2TgKNFnSGtNjyC5ps34A1GNDv65BSx3bZ+9KE+5KTHL
a/5Il1P6ZSZF6HxFn7yKaRroz1aLhPyA0ueh6/v3gu74JDsumRPdzA98xLacUYMjmLYTNdTqOCQI
xD09l92FcoF4sukloJJmGw9iwkAz1ZD8K/STYnCt8cX1ekrypx+FahNaZzXuKJ3ghskiUSR5Gw+b
0a9yQUUSH3En1BLmy7PvL6cKd59gvSPO3lsoy543A59xpV5/tPWht/RrTzK9wjWoNzxOshygq5+6
tUtpDQ7oZagWHvZSocJ8DY3KrF5jR4zGkT6MxICBRtEPIjgBycd+lnoEC/WLsM9NGe3OomugSSNr
1B67nAp/AC0WvCMQpUFO0/HiJ/rxJZ4+Na9SqCc+8INN9/nrn8YsyHXqaMQaIaA3f+ugjTYhqbu1
qWqzA8W910MfLTaI45B71680YjiiLxY6SDamMLG7myBwtpkICBc1BnHB4I9qsaCum00ZF3ocbpDP
YtSfZWIBEngeBE3VIihSOoAYBK0m47yhLfTS9GV1fa1bDRXR8VX1Y7p+fkMWpyC1CUTHC6C/xlAE
FKZbwjUFG4ZGFh4QdZv90bXMPzFQYvvXycpB06G/oLiWQ0OOwCpFNRGYjwQLsWNMY7MId8MToKW9
fkqf9tk9I4u5qkktkl0gS9ii+aJ8vh4n54D9XiafftN8U7z8e+0A95mHqCjK0qvML7GRBKdFVQcl
Se7UvgmIu9F5Lp3IWFWFhndfEoAak1GgHEQ5UEYaFHQ+Nu330Ea9tT5Q9DlL7nSRVnqC1XbNnjL6
VRsMnYOhikQAB0pIqEumH35jmnGe8/zLHDIZaISMvhmo1/2VsGBzoakU9UIYjilBAyge/A67Jxe+
GKbOa17amoJt5T0cCAQeQSxDA/fegx0OwPbS/ULPI4EEaNcbT4QGobibbP9fZmVUhccGGYbw/igH
9Zx7hoBv4weqzmTapCCOReRmV3uADG/60npz0owZ44maBQvMUOzweEQHFGDcBNv5IIO6uYOffEW6
8IQpKlJUortAMEngItkBvgKsjLj2LSXrJ2HoWf+LqPkM2pIfExLcVS82TvImy0Xqv0HCP3AZJFFj
Ki+TT0LQ7wRFuYFN+oz5rrGYJxwLsrVdNZGA/zZqJdqO71ZGA7W0RwM7DyuSuhrQKgqPs7c/UFZp
OeSxbxuBp+of2eG8jMkLpLtXecOQ1EkTgnusw4uYg5yp7Qj+MP2rN5GK93SloCNVKA02Y8sZkHvx
S6Yc/32HEl6rgbP5uTPlh0GxWu1sfRMxlDR6Glm/9CiRd42+iev+5Qzj/jiDs/cmwbM44ot80/e8
zM8+fvCOaDIzvE9aCEmSglnxcFlC81yjeq1OKxGKL/WAbe/zU0rR1qdrwhDk3c4x0hP/zWS895eW
Dv4Fk5u4r1pFLWLymw+dcZFJ1CuXTnoSdZC1iXdFlIC+b7ts15nEHk23wScA5cTI1LDhEWcSI04n
17PkZ9ovDKe6SSq+ti9WoBKrcpK5l+5LqqafOt1Ttq/FWc/TGrSBsQxkOW15DzsVpdE6q2cnN6Av
Pef1JRzdz7e6K9+K8WjvEmbcXClGZ+XVKM3uwN/qEpL5kuwhCZvYX6tqUrgZjguOo4aGgah5rn1B
3jOEj+cYqQ/nDrSls9OiKIcPQ7WUj3VYM8ikaglYCm226y84FXInDFJDsr6Eyco75iEEEMr28sqr
L9mjQQPJyyieHG0DOazqOgxs/2gV/DSmoV9HK6dTCJBnvg2pEdWHoSqRsU3kWXhu0at2MWh1NzP0
n2zRTYS6LLnxyQXn2w4DZ+aCdJPdbf5MjFsOOL1Quo4m5gj+LuhmfqoNtH0bmAsime2MB/3YrM/x
8b6kPVrju1OrrSH+c4QzTDPHP0B4Kdtoma5GusCwbzwINl3La2DR+1e59dQqB38SrwKMYqYUj5/N
nIYomjj7pGe+3aZrHYAbwKObHBeZY45Asv9JwxxwcLJx3rKxDHdxZ+hvVTbFwBZ11VOGSarb/HGh
VrKA1iS7z/vXWxirbcVG2nK+4elqJ/VvnzKz93SZUmumCsmSzgosgu78kIapZaAViQVELQzvNyh2
ChxoQlJus6L8SF+pjtCoczzoMEsxyCetMz95jro+Yl37sXaK1CuCd52gtLezfidTNuVh4LsInley
/VPs8jTqFIk65Bo4f+ki3XB9VsuKtDLTP4TbIR1QgYLTlMrH3nzAgpeKtsBfQwgq4uajcazkRoHS
1HOOtZG0C9U5GC3zhWiIVpJN6eK60Ozi2IWmDE/EWVydmZte/rz5xk6EBhrZYtMIW5JJEQjVmsOc
+aMVKdWlB6RTs3QRPX5OWPn1LmpXddau9tp1B3rpVZ0CX50hahLSC1ESx0kiYGXtfyqf8qBu5IP3
wbOOOlDP9Py65w3R5yDFjGnduk85dX97s9jz0+3oByW0OXrqLjd1NuZp86wtMbAVAbVQV9Sm6T2w
9EMoGNphlATIBoHdH6ESHGo6o5Om9KgeL+VUK3iv1jiqax2QKvnvCq/pn+muYgYJm6JPQYy7ZmzW
q9rb0/s6zWomyKCf61R6Czvz3DqL6ybk1ERIwBGqQIAHQXaVqdM5W4cWIhfITF+2oYH8AiC3IW/k
VrIW4PssmQzgBKIB9Wl/vzx1gOGEZHrbQGz2tN4Qf0tG3Eo3tgoMnkEEBS9FMBiFcPDR9hfCbNvn
UB6IIUa4X+RHHLvfCZcpFcF5wcSQPdeKd8hFuBBwcGm1WjoEeo8044f/PWRGfpijVyQopaxM3dQK
7/NMXSLu+CxmaXbbpsGzvpDFPw/qv2zlcJY9RwtOTNohIn8dA1C3KmzzNRcSYxYSDfOMn9EFQ6G3
4u1d9zGjQ7mtyTFwr8zZyhuQQKvqvhdExloZ8XMp7zTdaXSpdWnDwxCXYjNotnTPXP23lx3Eh6PZ
cg9U3gEfgHvlLF4fc0K6NETHVWWdpQlm2XCAnso30tjD5/c0nfLtlUbFuBEpgZWEx4GJe3aqLwNf
lo8RCAgBVo6xVg2z/MDgNSO7/0oVU4LsWqi8f3R4wJs27LQD2PbZEX6LUmi4ibmOGbqB4HPQi14v
ehYgltzbcYk3kj3R+USTU9g4U/KWB6J0fAJoimo0yqZjXYykGyWNKFbNVb/deE/oRbV/Wziu8Uu0
vTKeYzpeKECknVJJFRHFMNfvBxC+s47aX+udbCb9WCCBpQgn1CO0dKS5FyYBq06lwLPHDPjrODI9
vRpYQg++fl4tnIcK4Ba21xS38btw6OzowYtFmREjDLV5JuSNViHR81l3PnqwmhUensDXGD5BUi0m
m2Q9fbykksm3v5m+wmi1w/zHaFdNWMyQjuAERTx19ZwoLVVYg/sc6hQHWTKwjSlLwrYgAbOiRt1z
lCY17P4AI8Ua22mnxJUl4wxOc4Ya7Kp3wJxdBwSm/6aRV6Q4K6INAPE6kznfBABAgdjgU5eM8tXB
TEKmIezEu85qv7npKw/YzGSOHSv3JTTxp/DeQQaUcR8qjxRWQRXWnOf7pHpXXjOwGZEsfu6JKCEG
mlK6IbsqL+IfZR1X8Q4IRmhjMpvomg5hDm1HX4ajV/6GtyWdk1Qxc4Xq0hDfaJEQv0OaJKd5TIwQ
dqUP2yde7KL0QPB1cjTVAWAWvSXN6U2rzCxj2hS6AJZj87//fMe2mf6BTVai//C+vE5djfXbvdNt
ICMyM1K+IkmLUxjz5V2bHVPdWnW8ykbTpnQ49D6CIMyp8geXE4XMQhWgvduKy/BewlTItagp4+WQ
4YZMk5WXGEmVKS7fY9QAa85XRjWhTsB0s24U4jmlq94IAv0EVpVF3YH9uUt/GxN3vwMbzAAZe0+7
PaYM2TfWcGVprOhvlBbGL6+DkD8nCGVJRxdJafIafz1RPqjUMpdUt5mxqVrpssSsUSQwZqbqye91
0MlJzFyKUuHCMnVtBPBydPAR3ZNyZ5R7J+53g9zmV1JIQLuYp1Khaz8mRsPmTMb0BwLGwGEtNPQA
Qtpyxq6h40XIZkuARYn99qGf13dTHJaVePH5M4fGjmMbI+1WgETsOoaQUpK7dHuJsSe+n6I/PNg6
fHK2G1UrjjL7YrkEESRKnObDpw2uStD5bjB1erGfcK0dBkXYR7/v45c9MGXSCUZ9YD/H8AXP8ZuE
ydTc1sbRPGw/pik8eodc2KuyIeYEVKa/meQfecZDUJ64t0rAwEeA8ToliCMsHA/ywk5OMEObL9TH
hx7hXyCVSl1kOlS9Ag+b1I/BJksDP02h9bmQKaLHsg2pece611tmp81lbFGqWZUGpXpJaHM+wRtP
hlr7O7uaqA0uxWj6pbsyM98c8ZzLRkVJw3nkoZIJpjCWmlEqNQl9kNBNuQu/OcPBp/bI83zKyfeD
qdPa/M/ctMVtyPQ90mzcj/DfAhTFWqVGR1FrDR/Ki184xyXTWpJwie9U5MN6cxsGGTI5fzYvjK5H
58489oRoyx+Gubv9x/vHevzaQaRyJWz5f77aWJ0/wMlf717s/7SwqlDvR5XfkUnxK/tFfxPEwQ9y
DnecJKDfhtCJpIz90gsPXZvUvlWbNlTNmdrDGi9Qgo4J/AL6eYAhHyJ/oD+L3+VPf511tJvvQ8QR
ZGvm4FlsxbP6cb9xFRuG9MTk+Z8FI0u3wtTe7N04xCPrubzW8rd7JiyvwWMFAwD02ecPloHXziaV
buedOi1vvQ75/nY3xGumFvP0l2dNERomO2YFJ50EMvRRJxv9/2jLTRtf/8aubcfWVi4tDW/pCiA5
jsEaJO8hYINiZhnrlhz9HhFHPE3wKBNCGvD/uEBgJFPdca7Z1nbLMWhHS70zQaCUsBlwsiwbeRN6
NO5w1P3tqkEwIAhEBDTmk4NwRvhlxMJiWzbKR9c3Eq/WWga8OG1xWvMeFOrBCPF7RGx7tf4SO52k
sMFUTKk7Ey9n7v/wGjtGquhzMUtnjqlUCVfuLU7af2Yo0Ytj7RX+TN46jD5cWJHar8FCFHwgIOZ0
9H79SHZJPLzQi9G6DVBI3OjeX/egZhvoQwj5QzI+48wbz6ydRAQ9ca8OsaQPh6XlpBTxvzi/3w7p
L9yM+dAsc77vDVZRvSvLZYfRn4fEKzLJAbHcxDTgbeepK1nackGLIWJpxn4quRw+PR2IkkE+lGKs
HLweQGgpTLp+P7JchcTnJy8QAv+MSV9yW+RSHaPUtt+ByBiE+hL3QLGmkwr+m2T8bi/jl7ZpJWWj
5Ec+QN4aPp6YB5xhBT2Bqw2+UNMpXWhjnJwnMBEDebRodJXkawEvnvbmz/CUL1uHQlIshYiSWKGO
1713j2QaM8QctYpA1f10OJsPuSPi3bqjsJHg4Rv+CwLA/5BSir9+bczrfwB0GVRpLkDuiOLQSRfZ
1wcXYIJvLlT0FPYYo2gcZLB0I1v9udCL9i3w2azzmVhJnDROvZ8ar5J3Lds0kQ6dlM7HatFYHD/o
WYSSAe2zK/t6ejab2al1s9W0FhOs2vKkPidEPq1bvVb4zaqzW6k8AcFCsW7MOZr6JS0w5CimCe4Y
+dmjC41f4ZKkSKL1j1/jxqXx1a2UOUt3lInF5O8pADOa3FstxzBeJt8ARV7w6OG6ogv3d0A7tkLb
GjEN6jgJ36YwbbDQKQWKrIYMfWndOdrG2qN9QGhOYf/P581wb8NZjDOVO9ncK4cpjHv+3gA9aVoO
d0z99zkk1+d9YQmTieSuaUZfLP+1yhBP6pQ0YiPKTSZKVmuD9CR5kUkkBJrzqd+9zvxiEn2MXEvT
18fEXyV7/vb1FNcVl/6DQ0m22oLrU4ezxb5ugd/89YaqgFK5NHTNChN0YhrwBl9o2qhkAxlOU9dg
RhJuLAX7XnLVXv63fVpPP9e3/velTcyQLT4lrMzGBLsW/kDvExtQEpOVrPKsXAeotH8ztzNI8QZZ
gsLcMYbb0ar7j1cwv6VMWXBHxG5mYqnk6XQ2FWMs7zOOBv/E9IsGJv/X+amtWqXi6rYCwPsm+JRe
dkD0BEkNtv0vCLLiQhmWXr6r5qQCT0mCR8xRFlSnlq1ksOmM6jLfJV4GKAn+03WjX++ZjyMvHs8/
nbO59ttPYcL9QDOIldOHpF8I2jYcH3vX1+8n4Q25FG/hRMcxJi/4vBpIxbBzZjZsUaZ+MCMVlrTa
LaytvVH6Sjh5oAn+M7+xXGdG+7Y27pR8GwtXdH72eFHigSjpBT+us9jh+ZCj/y5cc8ANzC8sqSAc
niuURrVpqP/e2Sg58nKx6UEwAVxusJM04hy8n80L8IxCPDS7TdBHCG04ugeIUJHSBrDJqA8ngYWv
YIpHamISWqRihu3qYk14JxAoG+980DunyaKaeXUhjm7RSdv0XIFOhJw/jjmwpyvsZOMOQVnkIK+O
lJ9IKIonMbkiVVotcoKif9Q0sBZUgyV82UF53f43DSmJxf2zWzXy0NOb6rR1G7PT7ofAMVTL5v+q
8G9Ztji/3pQldRwbc1uv1bYdFiFsEBnJL6/KYn96GFSLrZ1dvMdBzMz9+3jGWIQfz09mzFOySdmc
hu5ibFrAzdj5J01x7dz4xZrVQeuk4fCbKGxH+CQ5WMWe2azoaZzuQm1HtESymo2BYdbObBqBj4Qp
oHFzvk8AGVPsQweNw4UpiGkuEwt6DUs7k5KP2witU8+P6s7r1Xln0QmEHKzb8Bq6Gr8yeWjk9ma0
bup7WhM9wRQ/VwaLZi3ECliz1PnVBACTuLg9MjtW4qc1hceQZ22Dm6nUMpXrs32PLMdn4Uo5yvxm
FRiZpUVPv3hstLp0QpXx+TaYvBGTOgUU/GEDhz784pRUuXEOxUlMByZct1FckaHw+LoLje3TJHI3
Gqdv4AkgMC0UU0LmiE+guZVAJ0H17+34MO53tbsS+8f0bV6XCKIjEzrHRWXM90iefAEG9DKgGijL
Jdz1S8Gnb8uNRMO7zN3EwfRiKRTxHnTtt3uorpMLkYIn5z31AGXO8Kq6dL2m9DC+FDsW88cCH594
GQB4VeShbGvw9EuR86lls/z6o+k2oUEVbArwYK6znwCtO+3XyhgSxq8VG/CiTboe4/UewfX97u0J
XzM1TWxIQS0w/SOrAR+BeDBEYvRBtdFgZd9kWKObh9tKoeP0V70a6+VRcozv4EanI+2sw9k89erF
UzHkUtOkv8yF4xyoqEwwwD7I/YRtBAJJRZLq4nGB2sbga1rqkGm4z44jeBX9A7XbZrbIwYtZlf8F
/+vG/Uy02t6fCjEFvdLgC8S/H7Dj1IxVgoaRXsqoiQSIMQJ/x12Uk8jKlv7Wx55ygAuw5KT1x+rM
J1I1gLQXrPTHzEh5795hV7e6rSHiul5Sw4Rw06SmjDRcA9mtyJF19++F5iFmtIHXzny8oZicDmvq
ACnNBav8bHDqI60xtX+t8eZsEh4ccEIhls6s0KH7xuIe5amDqd5lyobpXQ4JuVe5tgO5Rxkqap0P
MFudxGhiVeYAYyF6RcR3pfZHovGkTK9gBPrmN2CXnyGsnca4LnKZYMg5SxntmMXriYiAYmbQHzjh
yH75pV3DklRZ9EWKBvnlMWB1zvTDl7ApRMQx8UoBPWLfa832IjPQ56Fckb7FeQpLS3qa7Z/V5T8D
9k3gsAKI65cmVCD0yikFIM+xTvYp+sxlyVRUcIhw1Q8l8Mv1+64y+OdX+oAK7xfod8BRI4d7bdlO
l7836j9U4xbaxKazV32IqWcodr5QkBITcx3kjqXRpMGExzZgCq8oEvj4wcPDZp+MzDz4mJodhr0g
zHKifgaPk2Bcb0y67I68o+2HBOafb08WeZYAMWxbRjxGWZFUrUEq/ohGShcXzWb4++8t46/KhIoq
rDhSKtk54IjirRj4MBUnwsjsR3gkrPBj80G3Y5kMdDG4qEw0GeqSmaNn6857UlPtXivpViDuwYJg
sguHhtOfRTDEdDwX2HqVhxzKpSoLiK3KAGrMcw+U2cMgKIi0Ii0gVhs4YvqfpX6AJd8qN1H7/LDJ
qMhIIO7tOX0VTMAwgYambpqnRpvpuTDRX6bLrhIdIR8WG8yb6PG5cANlP8WhdeflgUK6+zx9iUJW
wXDNMQQKoaaOv/6gFwW/5cLWU56ashvolQGCD6TLNe7SU7ETZyMKJqJRk8t+NSnHnlig2L0pbEoL
ChVYHp3W9Ult9g9+VfL61/7q+iZh1UUPuVACxBZ1SmVkNkTWTQgGlz8mUO0IcAOJwI5VBdr8PlS9
EozU3QfIY1NewF3RRA3FGYdoHc0F0DaC5RqFm7/6dhpVaKAgnqQP3likzTBEs/Rk7xL4rtLhf1vi
Efm+zjWPqpExP4jAXzeSWV/l91F3qa3052L74MI0kJJobI0g+c+0g5CfZO4+gT/Dmk2no/sjRXEw
qY7tNHH9N52PZMqp6V6Q8wx+Ct+xqTQpPdLRSySW4qhzEbZweY48nkV9fDk5etCEEbEPqut2PVOm
zn5CqpJKo/aXrPwVqslW8yEPrZ2Gzl8a4xzGM+JordeSRRMKjYkCYdutEOaryj/dyfh7mHmBYWrd
RktTrORBAV+dlY1AtBlmG0xoyczMbF4LSOvjjA5HFSHe3fN5PtekUAdSzcec53xtKK5TbKTZoCeU
Xm1d8J5/v/MeqoGkFAe/Dn6s0aEahuxRJZp3j9O0apfGp7/aH/ClOuwnSARMR+xn7Y/0sMG8HJr9
0M7j+ZA3FXOM7i7VRhe2QB7rfFJjxyCixMRomULAazIzTkoBMwS1hdr6AUnTxfJorAPTKI1C4rP/
aUzIHK8tAQwD88UTK9WkWlpIyWMRNz6o9gH+Tl79jMgI7AeeaJzv35gHsFToAAkJ174l1eH7ByV8
i3f0QOAtqd4SY6JvBHLFxkWLoK3bvMybHL5PbRA+wyfKiF+AVkQxCBpXl1wBylDuau0sliP0d3U+
Ue97NSZtu+s1b6Uh4vU60bWxsXeL/BVcipNPhCJAkHo1LlfC4DqXKrm/sVg2F1EXQENpkZspdSEB
c2g4vVfTnoGodMCZFqat1TVJNXsPbN5SnJ1Seua6JG16PFpaLZ5Yvd3lcywHaO6fZ3NCfYIOAg1Q
XnJF/MJqai3LrCFz+DHI5qsC//6538WqrB/FqN5Eg/H9ehDVZT8hPmwFzGuAB2gCbS00LA0HUBPU
miupdg6LLB8yBnbX/CFNLnANMVhj2Wt3sohTT3/2fMEyWAL/EiodNDRKyi/5ZH9vvLG7k4FyJy4g
k33E9X5iZyLJaV3x2QcXbdIimUVJy3B1lYbsFhwLqn6SYFIqdvBIzTAWZhRmC04wAIbLqmu/fGn6
d+JsjrAlYoD5a/Hrye/2+FbOyVlUqnYcPtqRsvb9ZZNC+yUR4yQHNUYNyYCvMWjY2V/JMtJ1FJjB
ZnH52K/gSe3itIEchu87RR59JlflM0yngw3w0woXBEX9wGINHK36bmYLkPc0+IkQjac/tkdW8NSS
bFRCfG9H67hr7IdCpODnv4VaN69+iIj01qGBOSR618f231Ly2Day/y8zro0F1sntER7dd7nIvSSQ
UQH70EPNzW8AX/P8HKFfV5/BbvM3nV06L8gu07xjR4yLAECu9WL+t8CpKIspCy64B1TugIJyr++O
ldyY1j/nIlSQTl4jatD5qHj/L0bR8iSrITKC4OxUmsEOJ4PLgT1Gk5Aow+oNJEm+52+SPTqlkvNq
YdksBnWiOfhtB2EIYYr9MWYE6ivpWHfhF8OMBXNdylt5IaJxuol9S+sMW7Y3z9HTfCp4Fhup4+jT
+LaF1AKBTY+dBp+eRtBulh5PDDFG90AV34MlGLf/x32KhvH+lJ0iZQnPfrRWqcwbtmJkhlMBKuyI
BUPUrUWsYVDSyf0VLN0M/rJvrN2kEwxPu/uFp/CxPLGPDMIrPvMtrx7g78wCyuIo09O5FhOUKJ56
7C4DJFPH4Lf4oJI7SGVzRFWw5zRwzR0uaetyPsytS4oHgG9RsK8BHqoZGR2HRItTJuvLE1VQ7jS7
Q4O94e5pxWRqSsj1jD3o55bzbDua7QlgEM3QgHFhVzsMXftr5I3EHA0odnKNzA7XrJnKZIPPdZ6z
fvkLWnF71Ba9/v71MAsjRGGqT5m/y4KZ55qajaCmQV2/T56g3YEREP2MJGWgsnLio8mqblkDt/vl
ERlYKOT/7SR9MZpHxXdYzCUjzFCOuxff+OHGCjX3CDEQP3CJiBigjQqqOYhBQPI4AyH2TXpZ3Q/a
kctayf9B/GeGKITnxYQXbOdsE4qV5Wb+86U2eoy7MLlxy5px5vUUSyYhTd0t4nNDpplz6dxO8K5G
eNt8GxpmfDJePQrG5IieOufCIT438APzmeyZbDCGKs3AqfvNsp9omDkFZjv2408e9AB1jDkC5R2/
u0c44mAJM6Ca2rEr4HIHrIZH4rzk0FvePP1TIxfHLtim0c+a19Npj8+w7WAfkglCPtoBSFZMyRrm
tGEKWXEECh2DvjzKMnOZgTX57mOnBsKm7dn0wNlcHACV1CD2nC4w2uKFw+/+azvqWF6GyPL8XRyN
khH5mIJ2eSRv9/872oPJl5GGa7/xdSNr9XkEqtojHsp55aUIebB0NUzN9V2/dtZ69wfgojxCqP4e
dIzEyHkhXCYoN8tmj/eo9HZYZNCsHoyO1wx1dgc9FbHrmSoc/YotMpUFRh5akTBiwczuyI/hCr8B
QLHRt9nErQInJyUPeWHqvOZ8i+3qm+RMUwGzL+4Dg7+ysk7x1lddqCT0yJdryLGMsKV1rqfGvUFP
FFlImV5N7KoLrbP3DZ8hmKO/RPNMe4Gw3a5iVLDROfNzmX8x0yKZ+tlbVkKxuCKS6hh5fmzmQjS3
IsSuQD5Uv2mzoW/9iy1ZUjR4MNRq4oRpOcwCA2mITenXM0L7aaz/4WeCtYEU2+ohEQ6STZOatH1e
DroopfF0cIOF+8aJzUcUFMG/at7HiC2ibzEz7tlRxreY68gD7se2Swx0jrFulfCAR2KMm0cyG1dE
0Zzx6mP2QDlPJrwcPXu5mhGl43LrDYmi/Hsn1183TXadd09/yBqz1i9ij4TF9JmlBGsSy1sndVWx
9DQw7Rax6e7feFdnU4RquRWqdmT2Uyw9TYtvV6WgRcuJxfGOSPI1X9xhlonrgbmXJQBg3cMBIqMW
2SmpJeDgxAV7UroIpVqRDTIC+nCsvrdMxlC2ecvltkN2XarZD9YEgeiFnmKr9D9dPLi921qOOlgR
fyW5DqOz7lWAzGYasuTwf1CA/fvsFnikGEvz+SArO9u+Xi/lgX1QM/tpal1vbDoh5eCkywiOvlXL
hfYlFVAsdNSzOtzxSTE/iNwy/mw94D4Uw/dSitGolBubx+WvfKwJdJkHIbw8MJq5q5ihQK3+ITFq
1Lrbj+nmx2QJ1MRZIp+8mI+Lh3g2rlxf2NDK5yybydtqYMV/FCP9HY4zsfke7wE0KlT+BXdCfrJC
9tXb/LSnWDV5/DvhS0gIwvGvl2QRzCsbU/41PRN0le1rmiDYaOib9Rpv9hWZ15E4ZivSJ4GNdc+6
fLj9r/hNfc2p9F5PE0e9tJerkDJSUYHdlnIrPuJSa7vRAAkaZK1UrYaU2d60xG1dbRYX04c+/LU4
1NUk01r1l/Hcjiz5cXsUu99qLfz1Da6SywPj3e0eUiEyA6NyalOrESjDvoWRe2Tp2z2eyQzjeO15
i+MPtOEvN0p3m8a5ktloRP/Jd2LKYtfjQrU+ZLXWrWbm8LZzfDKvJ9lY95i6vDmxG8SghXP2KqNM
XGc3lhjhvxi6OSPbvyJN72wNsILZXuzG1uhIR722q2HRA/Ks5097pkDhGM0wqvaxgP/2R/Faao0H
UCRzLxU7OX6sQ8gikaDp1uQVVokIx6WOlvHmNt1R2y0JcDmR9afUsqfjqnvM6BKjaxxFezRHE/VO
wMpEGnMYmAR0PC+Jffhql65/no+cZRrDIbEUJRJELm+xFPscuLdA+CkWqXC6oKY0FhxAxU+GqZyx
VTjec2r9arJb+tm3N1M0tZdCPK/pQ/PDrLqUdXoKpO1KCYUH3d6Vm1Y/ky9oASKFUYCm+gy8sdBE
HVR5VSkHMGGpKfwdWUb2I8I4ncuQH4HZ7PIO63lfMovaSahXnIB7cV1bKZPvILHS9Cn/ahOzSMfd
m4BGVJKfZmuTEFzdjtlCYvvc91ptFE8hXJMM/tCROpJqmZbIOWtm2MImCz7u6PZqpcxVJVT//4FJ
YBzm4fol38U7MuFr3tigG/T0msmxLNtekA0bv9Iz85/PSKZ/mshBhzDHiWqL2a7yDjm2n98evX5k
XfD3j7Ly/zap1E2LlgHCGSrLLY2okMwSY5W4HV0+IK3Qb/8mQVDX2VNnPnKDaIuE2o6rLw4DbTsJ
fe+kyUeEjEQFZPWUgAzjDbwC0mp0b3Ed7kl60gWigdIGGv37HU/zNkjr+lJpwoie6P2ZWvd3DksR
4ru1bUAB8gvHRmkdBPBJqeojyTlUdrgAPh3Vl0stxd6U1OpQRGaSBruuW9PR6wkpsmceYfph7LVq
cosWnVzlaG3M1tMdKb1cr0EtvV6H9KgMDEm2IAW6o4ui46oFUd+5gRfUonfNNv3TTLIJbJGG3UC9
rF7z7KfAQPOagc+cVPHW8TUPlZa0uYowyhZRskTXMZdLKhR7OJJBktVl2Qsv8DabcaI2w2cC0yqu
gH2dKvdmS1k6K1FwfA79h+ueKdceRSeFx7+TMRZJCGb0Vlc01ZuidB+PZqCZOAePam1QWu7RlIej
yyu9EpfJYkSI7wojJ0mIbqZpRxA/xbOBaIbxSzYSGDfOzYmic5nP5pRg6o/HYdWcTq697eBrRX/q
INiJcT5hd0qUHM9INqO8GKj9axCzIyC2Dl557ypn0EywS2zP6dxCsstGn5MuABa1Kw8QcUrfzTlt
RixYiqOo6HYHFWjt/NYt9vDLI1AdnCIJBlenTc9+Wbs0iLpWhEHrZG0BQ3HxNSFWa0p8fSo8EskJ
41h79RU50rWu5wpmUukXSHDvPwkXGJfUR7imaWJDzSisgor0CWqaaOIwRmWym8K3SDaDM9IIgy5P
h5rkTB2OcaO9ARm27wgCBzYWiJXEQixef0IPv2X+Ge5Ym7pO/GeFci+7diSEMJCz7Cku30n9nk+N
PYOz0At3H1/xP/q79tIp0vZr7ktIx8/44/cNHAJLPjojIYM6ipDTjpmk7BMt0CfDW0TvzjojSUkI
xTSai/VuzE3DJ7CwjkwTSqCFZUPaT1xqgxMK0tsfFlOPcjymPcTDnqwb3Y6V7g8ZQWmqSJcFIzLP
nuiDgqnQ1byUekQi3IpumPgWxjK8xNFYw/U9wGf4yARTqBfJ+J7JZrWVpWZB9UlCEKknQPsiFSQe
xqglONxCC7PksO5pALNA82ksH0QD5C+WvQv8aUALdgYzvYtjiOHH8qPgesA/E22oJND2ORue/6pp
f2YVgnxO7g5Ly9dnK4Cx1sfb/a8SgyotNDPXzIBeE7KcYisbwyMKwsFyzVmZBTLgVLOQQ2MY+shl
XGW7o91cFT3C1O3VilRv4rZxvSMmJe2LngLSu2iPeDfITMqdt0uD4u0eWlqIk/wtwj99eP0m3ITw
q5TpGqrP2NSJpec7E7d6hT6JWq1dZ8pzulZv5HGW9/fSs8faTPvZp0wq0kSj5oB54P2KccKSqYxo
132AFLi7eFDsoZuMJLufy/qrF9l4vaL69rRWevXvsVoG30kDlCQP+Jjh9lhxGfcuq8OgNflgKDlK
7dv5vqX/44uHxYFB2OEena/Uj57NRTo1kMv0rx/XQ3oK68+kzjwGj0zEOVjYtShADdAp30X8qWqy
2hNrSameW9Ak8/5JJeChwsFXW6Sf7QwASO9B4JJMWK7blKGRW3aoLKbV+vMPrI9r1+RB9Uok9xve
ncZ5megVbXBhlngWmhcZowte7FlsooWWjGkgrggsRDtQnb94CEvtLVc/AQoN02UrO3uq1XTWgFPW
9n8FCAydPl4tptUYBLl+FuMswNX55RTLyx/+VXJW0rdK9NDkZbWGR6/QVpUiFqrt92diF6kjkIT0
tCbrUcsiONUBxrPzUPXRKHfujxjuYC5hJYI4iMQW5WjzmeuvGw1i5LytyU3vCQDPWOkAXd+gRDVe
4gzDoLonDRXNFuu+avl2ek/NST6Q/g+syVfQcQgliWW2FaSZOu5UM6cb3xeQ4PkjaIlTmNR099L5
ESDkUBfy0b+Hdv5loYYnkdy/LBi49POLv9qinsbFemINQNn5uToOYCeKbhANeL1LH7B8irTjIW8J
fFHco+ZfyRcrYsTSZ81Yv2sozu9wjeTx3fl5eILBgJeH5KlnE433IjuRmeoI956uTrf6dLMNZq0I
F5NZUDByUMq5plryEfPjJ6mM5Wtv0U8fnPBaJvpTGF/WEiX41uKWwRGTjI3PbG36Y+gdgCIq194Q
RZnzGV3qeO4c06uHG0NblzjCCFEOini4Z2HdYFr/uh8EQSwJKE0kQGIJLr9UXFbn6dzs7PTKxwaj
5U8l3/2m5i13a3olep/KNiiRMJIW5DS6HNCuhnrxPxp4+1X0z4RXNwtsll1TlexXlsUqwJQhqZiM
7/QT+Ii+AFQk+yeMNQweTQW8lQz1RFbsrvuBTvDY21uazs3NAMvVNzx65p6Wg6gw5AXP/6qdNI2O
gKm3o6vt9jeBuyzpNXxVMGoi7uy0ZDB7cDhyday6y84w+3b/n2cQyX+1MQQgrpzHBwp8qXQzERCw
whC2zSUPb5yBjHPBKnItCQ2qeLZIWpZD/4GgAHmibqWRBrt5lMrMCYPluJsJt8rNA5EwnM37/Aij
VXXRhBudBKXZlfhcf4sItLcXHjiIXuWM1VGecdaRMz/3VWxlSo81w6u88tUfnHMQ3QWd++XtjXmK
ixo0igrlbBs6biHerlhWysjdnFuNYq+ik6unUcaAyqcp8ezZefCixdfO9VLNxADpONgtCK9RY+7t
096VpaiXz2s7Zv2MmjLTLdlUxv+dqPaWX0b9ejETvE/bTciLEVHBT8Z1v3dBMS4bl4YgSb9UC2u/
K92WolNlnbGzAmrxiAuUbcbs4L3asL77Vo9edKH1T9oifc+YldBiOCav0o8q1Cd+J+8psD6qYCTp
1DcvHHflNeYpR4HF9zo9ugAyZGxbMvSZjqnhYuGlkj52EWmnV2AqTxEiyjoXyPVgal4qprwxIPVT
/dvbcd24rwLHZTty5l/9UIIQ1lKCIXvR93Co/GsTriB0+3YJjgavqIlkH5Nel7mx/4j/4p3mwkc2
S6Q4JrX0HwvyPyAAvBeGjrDy5iowr4zfIzJy6BFL4JODUZwvaAqBgp4TJQf2e42vTl990iSUQ8gT
CgcCiCqcTB0Oc0P5eCgHoVLkJ6aqHE5kbR2U4IcNv13IvniB8W0YrVU9pCAUc9ydGN7WfTa64VQR
wiDqXXFNnFmC/7JM8TSHQcLnn39OsmAOvs+LUqgbXSyZ+Wbex65wylRYbruetUlQDsL2KN3Hu64o
uWRiL1y7L1Vc+lm5GlepiyNkWRyj6y1uS2sgP+06vMSasSnVyRLfBSscdzFo2VK1iqu2p5s0NftH
bLFMi6XFZoQ0ekJ25JhY3r+gyKRyG2MYBVEYwHHonndaEQZUUIzMl75IKLA31DvDic2sPs/IGAlh
GqhnLYtCx0Y9ZGSPA0WgNliHsJi9AFpekDuLSSAyZWF5jRpAR54iHrsO7A2212nJrMwuuvKkmDFT
9M8WLlLxKzuv3vIvg7onocIGieAX9kMGpVrxvWUT8Ml7va6xjUu1qJZY0PGg80Sofs0l8VHisB2/
p4YCuHZ0MpD8VlT80tcLkSvjc/C4kHIvFYPKIvYzhdeufF6gdqFRbmsDJHtZ00ZQHkxpkkM+alqw
mmr5plVipFYmSki5nCL5wJtGXh8KSaXZD68ZJpq6nomQ5ks8eccUOP/2/s5yn3P5t8UXnkwzQCPn
08Wbsw7QnGdxnODEkMm7ERlqTvDRqrg6YQsHU2OLG4GueYuWO6kxvWzvsA5IsLFbbUYObm41RM4t
4Hd8XrC6WZpNxhe7q4/HhAOhOl9LChzaGsnPgkmcY4hXtxDM2exEGbj2X3aZIxYDa0EvYQfjQRzL
P0oEwZrM8JKkzfONnCfFC0iDnxk1bCaZfZysgV10afntq96LEybB6K5XgAWlEw2nM3anxPW+83BJ
lctRh7xfBP79GN43bhFAZdFSUNkORcK+UpSQHwxywZWDeCOK6mTBKLK7Q7rgvlC1QePv+iNEAQUV
6pzkGgRhWP8ddQmAUcM2f1MWtSv1H//D1cySweqFMeXhOoomNBoV/kVGURiwbSq9pbjBUkaP/cdM
Pfh+B3E6w+0B2j86tCW49U+B+8i/VLza1WA95DBzdLvuoVz3VM2S8DfQHz+JOmrTDFM+Qn6sygNl
5HH28+rEvANiCkdqnMEZ1BzkbuGg4Gr04jzH5XT+7G3F7ZqICJSYXw5aMIUjGVbC7FjuGivoCjCw
NAKEICYWZmkfhA3Lgqtf9njUpk/9K/ed2jyFuDNjGvqm7iPcudk3aDdb3vbrABGI9tsTyaBJGjeo
aCp6SAdKG5P8hkgoK2rkSkDXATsXCl8P472thIhTNQHV/LOKoq4tl5h3awYuEtJbRDeiVMAtyHPN
dqLXwVYdRFzUm1OSXAKHfP1P1ME+j8zPdR91Kw6BGxjnyoqIniXgaZUOh0B9RLWsB5vzPuLdYUDV
/SUQ8s9kP2+I3SeYvT6+HU95M11QCSJxTQqpUTWPO8TIagAYyc3EUFcA4ynZ8WwnrD8L5kFPWK7+
SUiRStt7DbduegOw6Ze3+yEGBnBzcnYzlsDr+lwcddzXpaqzRBzMbIqmC3oudmkWkZGy7CDUOaFJ
hxFdXlA7IGkWEC6cIm754GuUtQxZRvObYjiCEGF8eCL0n0WeZlBv+ryNzWiL7jq09qAPE1Y0kQHG
akhrcYOt0vtol0G4rJNv6cTp7kAFkQf9S2yVh3Sr3/t4PxeYCOFTp0oA7KaPamO0hoBkh+xTqCeR
lVdbQRMgmL1LwVfBU9RfcUNWHqH02ZY1kfrgdla5TKLZBeZH001g1XLgeqETNkc3pGw1tTkRMBVq
Q/IwEJgHvPBR1rpPP2JmjsOUZH5wWFc+AH4xi0esiRgOIg0Hw+houQlZtpxnlKmDArbhOrttheI/
94Vw+kZiRQGPig4/hUgDjZB+tBv3OrEhAxqYhKNQJETzZqs+pOPlselQgyKFvkls0AT5qxl4oWqm
3lT/xoAlJbm3fCNDyzwxL0qaEsP9X4ZrRO7ErRLbX+KpCPAwsqZFkZooRNBAV1G+8taCv+FvxRro
un0ZvzbFFtutgxWf5DZZKWEnmZOSShzvXt+GgdP+bAL4ArM7DGiR/xcenGyh3E66yaSn4hywft4k
I0K3fi2txwfmPX9baj5rdXSYcDyS04g563Qj1AFcOvr/uhba+KtLxw0i1Qd00oP2rLlXDUXSblX3
3pou/2Lo/NvaWqd3tVqI+fz0A4SD1Ahb0MM+OZs0KzKphQlfcq97b5eafJ5eiWr75yoVTIsfU+W5
qyPrggeVWgIfkGPRz3Eqssh2Oc4lLFV5n0SzhXwf7zqYSCOzekg0DJfQXfPT+A8YFrkFUQu6IjyB
sjkDnyrMdhISHPX6m3WjaSb9IwF65eaOUPIl6OxgUjEBClUc4Zn0xxpxKvpLHGIjPUsa3u0dmCje
+lN9Zhtf4gG5c15ztgV+Rw4Bcaw9fNap8Tow5UGvW52zxSNhy0z67w7btOelX8jB7aYXMK5wUth6
6Mzgb7hOuD8TPtgjcZVjwxOOVBgMUOQQbgPI5IXZSmCUlVinpjSDhXQsVgCnCklZlEGnHCgHe0kg
dV19RiotGi4/5yDE66gO/CKsLmSulCNAiJ/BYaWgPlOad0d3ZCnWvufRQlpaM9nIoN6IMtAsJ6+6
gw0rPxqqird3GS14EaY0ACliMmVJyiH39U/nassAWFsHEjfmvG/LBV0tX6wPM+s8plBOrZGcGrVk
24dTFIvXAAydxZD0hV9xcI8vcM3DWCCUuTh0hsURRr22Nr5BY/Bb0Qe5fflmlCXyNefdvOdYmu/m
rwi8eRGMJScX4+J8vQi8mlNM0GGR8BsipQdyjKbaHE/zgnpOw2jKRmFOxBDdxZOGVe7Cyg4uwozi
jG5x6Kl+16zSfVR1SnnNfEgSoAaDOIK3/iuaTUTjaefIvY5mEzpoH7g08JeRKPi0Po8oS/f+A/CX
YkYaK8a2KVDBZ9SQK1t2WRCpFtyw97X3hZ3PH1ELc3r4vy0Ncc0pIx9rAc1Lu4gOAzhFdqtK3U/8
wUFgZxtYKfRsONVsq+LRDreXEXy5XdL1KQbqYr5ziuvGEfB9/xVTfaNiuCaj2ayLosS9O4L3YhzY
Tjb+7V3EzcbvWwChNJjYfOjB3gTAX/Su74v3geMM/r3i1EbQ7w/7TicIFfXeUy/h2wtyfTqljoRF
UX3LuldnSHuV/89LLuQ/VMwdU+3fbwYfu3c87fibJ9gzjF8cZSgB/CFBhlyxVI3xKtgJcsmHsEUC
RJS9sTSX0579NX95aDL6IuVd/7ls4n/kE12grmNXpfBzm/z5xVG+35uDWvb0cxA1q8JdQE7zRtNj
PRwhxjEfFMrp3SL5a2VJlTzrMdF7HjeV86+ME9IAgBLk8xQF4l6c3RbJI5HTzfwgYbF0FA8eK2TN
4BjOxuz69q1nZNwB/73I4sKTJ7l5v8uJhP4LFAwHpk71ETLo2MouI24mvQ9ANFElRjj1QWq9lZ9q
FDL5RCKxJ6R7W2WUTSSCFlt5exnKL/Uk2cD1qiBcJzWyX8Fy3c9j5PmG8u0e5IlQYwYdDdqu99Yv
NnTOi1tyrwdNF2r8hhf8YFUrwgfk95xcKYdNVziYQou0mtiZSG4rO8bz8TgEQODbTxDfTDBUl8vz
Op7Mp47Bc6pZRt+dDsw9Isb3ubOq2ZVRjanLt4hBqy4FUjQGVPwxikC7sgrI8/9WEjf9WXzXXso3
3oZGwEewPs1j33n0muA2pYbU8CPjYoM+Egw5zfBBrjzc1py+DG9P07zKp7hjon2lGzXT/48RkjU8
ZGDcsEzv5zacajgb0O/+ZYMhtgM08izye+3hHnCSX6PKp1iK7nEFqDHYR0KZYoX4z19GbcPEdY1a
Yq+HLHXSlY9fatE9stfGQ5WXjZSHu2T2zzQX4+rVGDSPajXO7ie+nkKfHfX1qztbrl/eTU/Cmqwx
NaLtKykxQnNc9+JZ1FUyJiwccy5b9E+hGPmlyQ1JxAkqBV+h4GLFLPsuGFQOKMFUlPMRaNkxfS+b
JVR7dAtR34Oodv0Mx+teqP2n+SJJbqbmoxAwguHXD630upeE47ITDs+zy5eFRb3hyrPZoXeW6p5C
fl61NPSWrhT4C5DU7s3XwZ291mXGYv2v4W1YQ1XmLM3gsrA/esYekd0EEgEuoOn8O3h3SMUXY4wE
1bFMDUkgfX/U5zWRwqSl9tXZ//s1N4DuNSuCIjbk39WQS9UnIaYJhHwUxY1FXlTSPgn45uDLOQ6o
YxLKrLAxvRo0G3HuvfxtL7hsAMSlKTLb9Pi/OYwBTQ9GluJYAja/kDokwNST0FWuRVQWEZVIpfzc
hzSzth3NgVzadZvtXngjsWQcXNZO39KeX2r1Xuv16UaZqfDxqLV5MhEz6XuEZ7l0t4cahnPSeBZ5
gTJTR6jt1yq8IxKk7uYLv8uRLy/4l8518L/WOC3TiZhqq1CnZ6DIX6/+jNOMIJB4jW81ecc75x61
/y7Pkw1KKblZn2v2DyShTlX7mV69zrbKAkOSg9ttGOpo2SZvm6ZHjZx+1WyY/lKDA3b9pCqi4Aa7
fKlUrdXqUrkqrhatA+KX5PkLP16Xx4ZMhDsW8dA/X8Imr+XNuShcLsoJlR5A1H7AC7MmWw6avvMI
fmATN81za6YzJAGhRfLIVuhVvtQUFByMLife0pcoFnL4D4XHQ3Bx8JvJE9O/Q29/q2apwGmRzA+d
DcSQ0u850dTwzS2/hY+D5iXdOdCuXwto+vTXGI4if6Pw3WyR8dBu3/cEUS+6qjAs1f6eMnArJUfz
32LQNgUiIAAubtE6kjlQr1PyqxHuf1zspcJVeNHOPU0K7hJWsTuTzgOZ127dOW4eyf0TAHX20WfF
eMbMmOY7VVU2aCEZcw3mDjZI4YNaWJ4NbJxg7q6zctThvpVmSPaPgLOQ5fTYApaAAOxu4DqoDzmS
7GutwzPDbAN1FtR9cfVagNPLTKBpn3gRpJGkLFryrVy8KkzwRIaEb8TD8q0q5WnJeDbpZMVwA1iR
Gn25uFfH1XJd7VrB5V4fTA9ReH5UA05Qfq+HSISSsl5XUh/dymTOdUE/OYCllSUIAO94+4LWFtd+
hCOxdR8Om5rW0pdB8sta9oWMpE62F7yhHB7h4iNtmtbJUni82tHcv7p0/Vy1ySGSkl+1XOfqtu9C
D9StbBygCvMGji9CatkBl05rwM1hGRmJgI77cr0SGKiEo7nfM07urI9gTD4ME+EA92ejieGeDT34
JLONc2266FzHGHu9tdbqgsoMBa3XS6HxpdStvIOk6PLJ96ALaPrCWtzMEpAgiDFS445t9rjgDiAb
nrQ8YR6uUyr/b6205tdH1e75MdZ6jQyuvOiWGAjm2ZhTTltBGAqmBKghscnvA/TDO4s+A+y6r1eW
Nx8Gt+o3b11bX64jJ4bU5RRsZAF/q3X1NMzQNc4+WTcQ7kXxqBlgNLNr0DzTbc9uC59pWWgQEcMJ
19HmYzkYe5AUkH+ranTEORG63krr0HSnLrHjGxpbUSBnDYfado/dJyTpBeqasvFHBxcCnr+W81GK
jwRA4IyixqwcSM8eb/cgTLiJWfXWud3DPcKseVXESfpQxCj2wRlbgCwmneyM9MYP9nornbFkUh6g
Wm/RxQ94YBuBrBFjVfDyXaGDHDxAnpmyFHG7PYEq1zv/JpzPtk9dsCt+H6sGpaOhMaets9xqqUHk
CzOLYE/dkoE8j4HmNeiA0WInhETW6eB6D4xKVIHR8TjSdVCjGuIjQjeVOBX9v3gPR5D1WXUu4y+X
kUoXWHKfRVw0Ks+cDX/AajF7ANEFF9XBeoi3ZhMvA922zEgrufU7i9wU6BbSTRdY+bXnDQdlQ/es
ngX5yfVQVFgx5R1NY/gGPenS7K1cbJD/7/Pc7cdUntrhiGXxr8XBVzHp0P2z/+LcYnPnH6sluL06
sIYiGAXNpv59fOFKoRj/Ch9kr11HYP/QDndaF57f36/2tEZt3v66LWw4Y/pxqCwiUjeRROusffD/
CG4LhyT5HDxH0qiyVm3B9odscatvTv9SuVFgKMi/o9Kf5xeN7tGIAKo4oiGD6jWBGLutbFdI0SAm
yqTh13+IV9jqFzhULl5P/tUdwXr8ikz7OcXJ9M5l6uGg4IIYK1PGlLC2sVb9/0BdkmDILEhD1yd9
fcLKOKKwHkkWE7K1N7FRg/rNLOwz8gVcZQborqP8sfi+YWDJBREaXP0DelGz3x/eRjV51E1FOvgb
bslZ/EVabD0y3ekjpW294pBWGcir+mAB/NMN9EWyrgFDB1JmE4xOFtRRd4iXOqPSta2KS3mlZXCG
g8LpblVuAgqqFIol6RsifQfi1BfvbtMRIrRlXe5abb9fbrlyf5lSM9qob5EAyd1mrbyPe4p5DhsE
ufU0CskoLnZLQzo6IYZSSq9G4QNNEdmFdrWN6R2Sjd4ANa5E+HONJzUmEGiE9ULIInO23TK+LMoj
XPrBAgUtFN9UKjhydtVJbNHcqTWqNYYBK8fp3OMnSw8qfkqXXJ0R8SJoTudVdLdtNHeB3xxdcHgv
Bzxb5d006OMDDa2S955s6RJPxtGt36BbTI/z75mdsYBtdr13mFTWqkfZRPY77dnZGWN72ah3OtoJ
izZGF2PNV3adVgxqsAL7mSEcP17OJiHq/510b838KO3tJA/QKAkLKR3yegFmBCDk8iXaAvBViP4i
oZfixps2l0oCTEEeSFX/CoJJVAU/lxOC68qp76ErAJXiSuztXP0fTrH0xkoEeFfD0EAZYVoDKC0a
4zxN5Bj44UDwdhHTGpZuJwbVgutQmvR6krrchmE+K8gNPK1M97sgpBXFBZV3Mp2Ic0okyRXn8aAM
ishoygdEQxcDVzsVedqqQrNEYNvW9uJ+p2H9y5myTtxJ55qxUuYO1XMc34eIxPMMOO03E2H2f2M0
Sfz7fFhMKPLwFohhAIfmG0gC27OUr8cjuSDMDNO/OO9jKl5FvCf/2H/49/q/80cYk0PMbFCFVpMs
KEQcsarlqZGJtOQMMRcRCrzwZuKgaeREiPyxnm6Y25N8ewQkQVJ5b1cPfaHupTfiNcJQMwUEtbVY
y/kegg+7qz36B9xdNMtQo08XY+rkhVj1wxQ6AcM6I+hwYwnwxGDTfZHGtwJVLtPi99tPGc+HLyxG
K89M/mAuJLY8UQ7NvqciNaTYoV/vfazd1klozoHVSMQq/S40y3kUcxPj/7m6MnW2fHupvXcBT0Bq
A2S4/KsyOHmzq2ba/MNKLEam56BCZMpViipO7r8GGf4l7/PI3+9lS39vo6CkEoRjalcIj83WnGH6
WlXxYnunn33M7nUwYylR0HNrowZVCJIYGIf6OdWhC05nQEDQ/xQgXW36VGy1mmDoH/RVNoAwAnzg
dpDkCgyHZCofD0acLsgyHgYs77edUg04YXmTZO9lGcweUdU3rgF3XVvFWhEsmbv5ZUT+WPq8zghS
bVgPh+PhS2kNeKwvn8+V08Mkw89uJCjApbv3srzyJtuubnPOD22/FLMzY3HEOvpPMCKSsNhCK4/7
Lzrcq+DVH4DWnbLjuYX0vkDtYnoSeoA9wO/juUulqeCpOehgsSBFsklssc+VIWkZisSPMDqUOT0u
wzuCUNqAyK6Dta6FWLqXCiJ04vcz+2kiXvttw6Lns1S4PPrY/RGSPcfN8O0Vnr4kDSFmqSAijOx1
FMWo4J/1u5vajRATAIDoiEi2HBxfjdrT6I64x4HYdko8FzpDANOGcVIxsDpJxWW1iGoi/K253dC+
+ZXszlAokNQcZUOKArzFEd9bZrkvqjgusD3o2CUOTl8VzAX/8mEMLiF9R0M3JSY4gIaW3gzykZGE
Hn16WE+F4Hb087I647Crsi0ymcy17QC2gvUglWLAehAFVnezjIdqQ7GCih0vJwHQE+zuuPC6645a
1yADd/L/9lWA6cQmlhw7Q47eYdNPMdPwwtFcxb7Gq2FoKmZP/5BYIk2AXQ3k/KC/V8U+XUd4Rr80
OQbcpp7Itw3cQHfa2wjyVnEqKB4k/kGiv4RjeL0XIZHPuuiGacFKlSSW7M1blG2SsCjYBRsWfnOw
tPHILKbm+aFTQ0nk+ayPLr2BdStdUlBzAZAEgSUOiqGae1lhZwMwBNmFbokaj9jpaVK9qTlpQ3CI
+H0HIcDyxr4o7WmmAOXHUbcTjTHI824Gwyfmv/IAN6KvN0Hp8GNi7lgrrpKAG2S53of6UCd0rYkN
rzZsX0jCuWzPySB/WqSryhXtxYpnq0O6lrGRUlYLHZ4orepAA5mndmGTLjDbswisQ7QWFxbRtv2P
plIUq1WrEDO8bbbBNDn94sGRGsnYYgKPUjKqvyYWixVQCM0MnWhqgWnpWRlwKQU1u5dr9aPfT8Uj
SVuHYlXhnVM+XJMPmR0cByUA7Y6bVkBdlWSNAj2/gqzJo0jTltHSSkxGyAYTLv7qHyQQoPm+UO1b
lxrsD6SRzxc3vmgk2C2esfp7dkPxA/wJGgCGxcSraOw/y+cNv/qBfJUJ8TNlFAMSeGJtaNcZrOxb
/r/wjcmPPuVOnLkG8P8fH0BVCR9p1zzmEWVYZnS+KNC+5VTfv4wZFmXOSyrTHmArSqT6jFSPTxuy
bvIUi+k/Wsuu4ARbDQT0V5iqy7+udr93IzdEzdvIsGxQ8KAxxv2QPePP5a946fdbWDZQ+ZyDJGWp
aaSOfNhadxNLkB/7o7HGPdZCff7VYv85DoBV/0CG89uAjAYDeWWGbEkNPh68QSmC7riNOOwR7+k4
ewuzo8/NsEAi180Kko3HUCO2aQNKy1KP5AYT4SfWnE3AS58PmATbuIFjDBArJTJFUZsvdPVpQFtX
99R0z+c4HzPTYCLzHR+D1HJtkpptXIuEVF6l+CUv8f9UIWXB4dhnrcJQNsKNDL7PKvgB8F/XzS8h
thrywm3kkEezuq7DK1IFRT0/RLlDCfNXEHXeqTz0nr3SHGa828NR9XRYF7ZQdcZc8s5JTKzCwa4d
I9kfeUu0unqg9Lh/motXRJ2XCMHHZjCPsCifo52SjNBczCZ83DZiQrePwOBreLTfDr4LdW+BM0kB
OY52kd+VAnFETqgPKjjqMFAMg1uP7Uln8kKszcT8xApat4Hr6wTjwFxbVaxPPa4fSumsEMQcDUsQ
6MdyorkRcxHhnZT61YHy+9IDJ7SDA9H6dZm7y3772/OFOpkBxLg4c5I5jf4aa+KFHCO5tp9sc/U3
qhFZoJfFlgUa5g0+E54uIRcSTalkSfUsUW7/Wm6Bw3dFSCCz74v9lk/dWmvTLz0w/FwioQPJTZ5O
g7pNvPRmilKb1O0kYsMnEeCnTTzuYO/wDZp7c7/Bn8mdVVw0+YDRdv7d+qFpzBjk9sIuNcFxeA/X
ZyAOYuI5nCVSlU/OdathVGMRBVFqFzT63GbgBK5qrSW8DK3rit+8Qdd4H5Uabxck9mU0KsXb5WsX
aSZ7RCmv+rY1tpuUGIjSoRGHTWXGHPKW3nGvB5Lmrek5KI+TUJtSA694Az54LdSeuhHr7DJ1PIbD
ftEZgLExISdwoWIUQX47idUqbqb9xWzTTt7//nRPgnZCRieRldAQ6BtlBBtb2aoPSw6Eh1IggaSq
+XyKRPQYqjHCRs+xn9Kx0HaDolzG5pZB11JoQHx5sA5YWXvFilh7cqupXP2BGBbIMY/OpVYwewvX
csKzN9KDWVceR2b5C+caOh2WRIJBUxsOoXrLI/vVQsQAOsJXoSPlZlq3i8FctMHHkPt7feEfIlTb
JLKJ3b4kVyXDJEl40gtJveHkj/IkAQXDH8mrbwGbPNywLMV9bHpTvRtCkEBC4OxZO3Key4d5soDr
Yqn2GvfPsqiiCb78HJDxprbW27bUD+TA1/N9mr/P07CaXYtYIdesjjJdTGE/3cbObsu2+EpXEncX
wmoa2+zLs7WJLCYO1PWZtPpS4KLB9weyL9cyblBCGedy+tVYU3xh8CR0wI7cjAL+XEd8KCRp3Zqu
RHjnYmAQz7SjIcb8e+dxNMoZHum+HaXdZjsC3iHHdjWwBTSi3S9oOzVG5dM1IL8RNWFKtew6jpqc
qsjsSaI/Jju/pDdv2eevKR9exdAdJqBtIy4AIEtDKGW0TNVR2hooTfeRKqA9nhdIxnb1l3YYUJge
RLBkc0us/4nyPLpY8RjGswJ37qLHu01bFGGS1fO4hyHtq9l1ztbgjHEbDp8i+TawHOt7YS3A4EmU
Qn6xELkiKiFMMijZnylXPxbxCwCZmwPTm7PsJDQdKdQvWpvysXHabzhD2lybCjtWM/YnQzYeR/Ym
CSZV5mMRsQZ09VDNjrjX9kDN4UEQ9IVpt7kZQ55Fg0AWf+Y1HROWjbRwdeKVUmFZ5V6Ih+IkpdCp
mMMAjCFcV+k9Bebz5zKQZUrerW4JaF/7hLh/A8GuwaX4ZXCvG6da2pvseqgApN4cpGa43PXZFfXj
OPpUmdgKWFEMU2I7Jpvkq8oYq5gVUPeT4NQQwf4LBvqoL3hl5gzKc+fZYYDBVcwy/5kqjXUPZLGx
XdKQJ1vEVSMoVywOtLWH7UROrwmnb448Oz8dKjpVRwaHibTwRNX5zwXRZspipYduJEiWO20x0WfO
da7s6zaLbjG9U8A9NjX/kRrEXT0NGCuIfQoptQYIh3GiBnOd681dO+TdvCBGkt0c1Duhm7JLelr+
K2tdLioX9WdFwsgg8GRn/XPe9fIivAu38nJGUW77KiaClSdCpd3z6Vp8wYAEESHSpMXCQhLA5CuB
w3a5KjTX3nLP8awFyvBcg6m6sqByoQ6/zQw9i72pW7+pfMwis2e5A4udV/xqUzu4UKSS7r1rGrBS
DtIs0CBdCuIk1Qmmnuky08SPWLBPs3lGRrYs1937pR3yaBSn5t21u9l6m1p6hMf7Hnyv2g68MjEQ
NxgJ6EUjulLEVVeX+ZaIWnaaLbHHv+Hp9fFU65ZrNtms0gqgiFmcRlljrVup87/Asv5d8dDXShtZ
ZpozruNg4Yx6Lzd0gQprP/89TvtC0xEPTCvSTqJRyYNuT7l9CL08em2S+XwcYSRs9T+Tc0aAqvW1
bxxjE9KW/lr/jn5rtP4qFOVWTFPA1sKGD1C9K9lYBvv9kaoWse4sMkb6V6hfy3RGdRId8PLYIMwB
82u10L+/geuQXSYS9F8m4clqc+1FPxmcHMPleuzee+CFiwjZdy38fx4oCWbSXeEd+3DKcvVjS30P
3WX7yrwFytRrv/ojMdUBuO16Cp1UKYwb6j+W8DX/QlmybyHDDIH0Z+HTKbCbPewW2MJ24s+iElZg
DvoTQxdbOOiXIEoOtWRlwF6RJi9D4SLqP4dGgNpArdTg+582rDNceUfHn61SR9OU36xkJWKV4lzx
PT40usRgeMofRcnHWkOzEuRjWlr9rYaWoAm0GqkFIBOG1JQ25BefZ7/MH1I/X05psnoLmhq/oMlL
Bwc7s9bvssWIhCUcEAjGSIqMRtPs0u6kV+YIb4LsldF/qkjui574j2VpjvWidMbt371viWUXhN9S
E9B2UEPm2WfVZmydsjzAUPAzc/7H81OhJ5OTuZ24GapMRz3yjFF4HjtkZWxOa42O+EjkWjhlos17
cpJjQw7wOxdY7UAnJlHmMZReQW7TBLSJ1+p4BbL/VEoE2BPbrAYqJd6ik5er33xSRpCUiZZwKFMc
RBrUErNp6nuzLiPKZ8szAImCF8keNjQZ1kA0SzTCwTUsoi1+WMpkG9d87ooIThL+3iNSSoxH0J3f
cgZsI/bko+71Ol7QaANQYctk4fK1xbwzBGGoF21yPRdNaPLJ7AY837mw3/KnWtON2CUJn9dXS7RH
sIjGcqMOAjvKckVvrFg+O0+ijnhWFXPGsSZ3onYhNg5YoaEi5xk2KCEBxW0ahhDYZHkajvZW+7zj
QCPf5aTQK4YOhidz0sS/4wwW64X5/58ovdt309eTGmo/elXdJaHuHncG3tRHvfNfd7cbJaiqpFAj
fwhkDGNsxSUC+eftZLIMQEencpg//jDjxj8pOSMBvXhVz0k9CCq6iblhsh+sCR3NKfDEcxbC0mtr
ULslG4SMnwyFkNmM+a1OZky1eidtM07PGuWY1tSh83YFPSQafkaxVUg3/wZLdip4SFLJ6F1fXGUc
NOcroOgG/v3meU1U7CbAFhXMZj+2zJgXJumfRnnzI7Vbg8/EBTeTajLAFTPF+iuZKoYZleEUXIGw
9MnvXigbKglkNHp/O7irTtHD8HA9Ze8wvvmkk9p0Fuz2Oo4cjtN7ujn8o09N8s4GBR0HJXjxScmR
gdPwJ2rZRPnYK9WNNjWwk2ZcLC06tDaHP0eUMcy15kzHjfbP7Ujhb6UC5GO4mMagD05tQ7VVWoiS
RW+sTMjs5sAWn1b2O1pC+eIgYdzZpe3kW23mimyha1XTEaTNuqut9BNzO71JpYMeH+Cgs0aE8Cig
ZsSoJuiVThfVhNHr7f4KRWZ9inP3EcWlgY1tTAbhmOx/ba3CFUExhxg3TPVeIGjpuuNYnrPFQ9Ry
O3UKpUx0INBfyM4dsDeKNQTgOE1CsQg+VnlFLoJWXFs0zOs9eZEM8zEnRFuexvRweeDoHfREQGTk
d5xG3aIlmzgtmhqQHbtV9HilQl3hdsBvFMxmnsP101qyu00jWIAG6xUaVnSRY9oDFFiiEIAUeehx
5KfOCNdc4zFgct3fdJO0Wjxb5Ck+uc1pWAePQq5hk4sAKKbC+6Rt3Sn+luLtxkKUz7oEzSJ5OXMq
uhAG9QdyNa3JT5g0xa8r2oVXLtMeSFrjg2hQTcBKcZUiXS0K5nn6rHKuMRt9OXb8fcOVMzzNtY40
aihjCQjupTOEWZRWWXqYHty5mCAMo/I76PtPv2hYfTYUb0qugz/+VKeuknl+cITvd4Bu9FqDuRfq
wj2sepYr+s99ClNTz27BBk0aAl2PBh5W4wLzvJ+Qj1H5Bzz+eWXtbSR7Sw92TxeRc8FO+GR5Rt/x
Kq4fSV9xPgFKwG5GCDq3LzYr4WMxZZaHVTUKVPKuH/8d2eZGKefkvb/46zvC7VG4lqWZNt+mQYSu
EPK3asyWVWldUdGp8Xyp/0i3Wt+auEw6shP4pkkS1XGIPnD1sP8ROHFeBCgbOcFxrNa8kMO/k8Oa
88mF4mIxPtCdFKH0rn8BtdfY3KBnBfuJGmrqUshE7jnSQgvoJ/ZGURaVHffMwYzHqAxuVgs6rlgT
pFY6GckXv0/g79ZK1+4tdOtMWhiEoua1W8jXxsnwitFOP9vITb1CkRwVvaUUQU413mLKDGr+4zQv
F53VTPUrr39B/sEVWPTsbj6y63vXeA765VG8dVYWLGeWpUHgmS4MGPsVPJFc5nf1SA5MYX5hOsjw
HiRaYoExpOEwzKLpk6Cb5NbF85WRh736fsn9Tvy5qt9ePMcqml94WZnwp79kG9+Umpco+cIR3G/7
hLYnKZNp0xa3ogIyGkpmnporN7Qu9k0Myhr0tg1zxHvD/9CCB3z8RThfoh7gMQagSooHvb8eu/oW
aL8hpjAH8dqHKasosHnJKU1LTXBYuj0q9YUnzWqMtPDPQposck9bZPhPcwfaihy6fvy/zWfkuZ0D
FPEOlyiJf00jfNeaWUVvAR5BJtXQtnYzdQu4bNbeQ1dqhZTQ814MVGPXZl92spEIq3xIoZn0j6ee
MV7RhnYH+J0jB/+2n7Es51EFcWp4x0qGoVnkblrnmbNNuBcSnNskCGH+Vgfn4ieLdj+fqp6pGJ4O
tYMoRbVIzXcm5YkXhz+ablnpkWIgH5+heoi/jBA/Lj6+3fxU0IjJgZ4YqGHLBJPfGtBCyB82vYtu
1RJHOBQKBAtgzRG9KCu6HPxO8CXocurvx/hqhau1gDJoen6ZKrvAjYDUkGSABvj34q17+hLMyX5f
SnTfFMtYTluY9bDzZZ7pk19fKuOVy5X2Jatuf9HN/9w3CeNqLvNPZqiPwcU4BP0APc5amwvIJk6E
d1ROr4tEzY4k1gfV39E9Bf7XRQgCQCrNxVPI9jGzgifxvHBQ6yDMXyZKCzHtTrHmTy+vfxhDV9Ht
zd8eNbBqMBvpEq7XuOA98THsawS+4UFtH4DpjK8Fyd9oHyU4zARPG8K9FLZpS2JVE7KxFbejaDrK
+MgEmGCTxLQLBTMXc3kQMxyleFFpk8YVti90tzI/7WmrYAcMydzHqUEUsCb38phzF5npRuJmf7/G
4Uge/0uiKNM5pYHFoNYVHKIMVrQwCCAzSJYiGPsNOE3Ysu0WE0RT78Rh0IPdV2XJFnL9WixU95D6
MYNhrkI58Dkt0urHzeReZYVjmgT1PPXVVf5ckDag5x6mNi0TUl0iBd0Ya5eLlBt/+w4CQTZUF5aO
WqC7vH7qELDYrWAwOEF8eW5LlYigF3z6G0VvHYVF2fhLJApcQHtA41CkoFZVGhlc034Z1XaKGngg
tqglU1N6dwO+aQ17tsrYWJ7RYa+mcUtbUdXwoFWnqHW3iNGk62+UbwgXon8pI5hhMzh/ZFbMiBZU
UpcW66TBgdSLbuqPU6bjwr+flZJZeRq5TKHZhtHsl9F4PL029INVDAUj+TBgzSjsxqzppV8bDfCm
DN3rJx3TVKy2Vb8nVkqHaOIr/rl7+At39J9oCKR8gs0vE0yFpsl+bZSMMEjbSNubTuuDEaQIvkyn
VzmDH0+mrpBcce7l3Ts8LC8BVKV6N6Hunk+B+BNa/H29+yOwzrhYfHfqJj3/YNntIVIcjgjeGqg6
7f6FQ/oVONzAaTxIo8qS1zm2NjzgAc8h23Ai63xshpETo1qv4vb6j1P244AeLGP/2ASc0jbvisNw
scATPrCfhulwI6CtzINDiiu/zZRA95M5IF2XzoDIMXEfIyAyJHo7g/RTcni0/G0l8x17QJk5aeV3
H5U5ZkePQPVspmGsUN6L28FXfekAE64oGU0XCHUgmFIWgq2HOpkXuSuLE5rIeehZS93zDfSQFQAZ
X/MQKZgyXwWNiCpR9Ps5Z7bq5lq0gzOacZyCenojnAt0sMmx3wM5STaMgh21qExBn8z8fe44zMJ8
uqbttnhK9CemnBNtEyiFbZsE1OKmwaWvkjLqiKQLxHqnZg0U/RpxUQt0k8Sn+3ek18jNFsjAtalS
Z3o52erDTJRFITOzYynD2vdrQFvv9aJYwE74q3Y/BNfH3v9gr92TkzALFALzsc5e7k7CIL1/5M/H
CL7z1xAYfWd6XwzK/bBSC9RAyS+UlkyOORU7hZHc5R8+oMINOm3Xpnwo/ekJGK9dWZCNiCyvoc7M
JsPcaTRtRR0v3FIA6HrhxCA6zN0Gc6IDexNFlyas9qoxK/Uj0rejjikZNcuZft0RyYvipe8tXAR6
S/PzY0CyDUgIHuku1F+j4nzGJIbj8lPQZ/psuKXLRJWwb4wLGvwjPfYbOaYMdbJWO+GljAtvXpCa
IjBboDXxwukXjzvE8ETVmS2bSEngL9rJ9lChKsQ0oBxh7Jbj9Ct6FDecoF44bAKukvCz/FR80ctv
ZrTYtZcEoFFjQFcg2b+0NVQNOgfZ32OEyWQbHgVTGbpMw45ublpJWEUVScXw9+Tmbwp06XukDtok
C/t8VJngL41WoLqGrb5fp173sgOid0KilUAUP1wnlGNWnBVCiAk7gF6Ucqccs5s7NUOzt2Loma3y
V+vywekCbQndnRhc2tQMs2Hkag09HTSoMO/h7mCQVEboyhx7WuLd3Uo7B83iTO9t0VZRo+3jHhn0
MARNgnyzxreSr3Cj/8h/4vsvGep4S022BIqDtclWenBRuiHKv9rQkUz3Y4ilM1exf+3Gw2NyeyvZ
F5B1cLn1U2SuzeNBgonxdGQ3id5ppOUQ9CP8t/QMw9fJQ2/WIzgTvGKrcTWxYewEwEnlqeVHjS8a
/smxg7KTE1gcVQEaUKmA8XwXCEe2P8Z9z0vcv9pr10vCR63PJj8iio0TxJK87FnWjeqX3zqhuoHW
Qq7Mt86XoE5HxtyOfdQBTKybm+g2vP6I5pcDQ1I1oEzwuYaINqbXPzazFGpGKjgTaOmTRqeJQfDf
i02Ht46dxd44oXzxUuzGqovSIr8kpWkgcdc+Zb/v2lP4/5Wk38ZiUhjlRf852IAgLXMuON1PBEFn
HJTeTKxxOCZOg+Np+MgIdLHhQLpRSq5QutP1j8lOHyRmg07XdkSQT8TbEdgal2eLe8PrxeGjdivL
QP7KfvZiAfXcVgx4VbrL31TgVXx4EwakXjCcEfnO4m0GWmK/JPx7zTOpe8XRC5vl5B8c/73huv0A
jhq1LN/+/a5fVpnrg4tUJQWEdrxDbC1NtI3EcLqmTNXzvp6jjSu/B0xNWZFpefk/c1gsPeQzaS1Y
qjyFKEKz4B6QrNbfomatvGWFs1038NixDiQb21p3j0sVJO+RHr/BKWmtZHJjYFC3DLM2jTE3AZWR
W8v43d3RKmy7ia8Ej6CtAHl5/leNcvlaVGDWLd53byEsCoxmMiHatIbbJ09AUFxY43s0mU4ZjNy7
FvJXAT90SjMpjUWfZBkI0SxFVx5eYRTnLbZ95g07OTjx14wrdiiif/gQJUo8FDaKSUOsjpYXr6p6
Q0KFJ/Sh+DZj4BQpgsIQc8BCKE1l6NNWcLsA5E773Flu0wVVhveYvAtnB+IAxRx5/YTSXPO8Sysl
VjZU+Vx2MXfXRVU50/V7D18p5BoJTKakZE6VLYXLOcqDVovZLXfSqw7hc6T78KjdyXNOE9lRZeXZ
U56TznYeJDfAVoHeNNGPX1xEDMpk20KSX4ddAgzri72PEQUSuqLa1tyfOHcHsSxjXZ8BrRJ7ar/L
EbiNBfI8MrUWrTD4z8q89zQeSR18PlKP/L9uhozV1BpsXgmUcBVM1Nc7sFqk9v4mc2Rpfkgfg7Q9
vYXesM1JuCnPIdYO3dCU9Ug0NTVZNsnxmbUD9InXWBxUQR7mZoQ6JMwoOnZWsijuLX9RT9mz1JgO
h2rCYmHWmXfoI2BVYf6+yGAAZCEGCfRldeOTkZBQT/MPaaxJKGMWCI45LldTBzawYeFMWHVLfsfO
o3OlgIM6qh4ktMH9wZIFgR3eI5vYkXVY2SOZOSic92Xyor2IomseIPV1ZHXv3XGSyU+lwJsVJuFT
NofRcHh7U+Ba5UvHzKVYsdHbcDsacpLOiPCiivDoyS+K8gFABI5B3FKG0YdnQCF8FymEKPbgr/w8
lV76PLS3bD64NSGKdRSu04rnPAk5/XG3f2cky/hkUHBb7e+X/7TAlC2fjM2vNGymW3k8W41goHvg
f472m1XSs1OTu48clBIrh3mbH0SroZC5TeJfnBV10xjzbiWm5XOzEsYfpSxwcS2CMF3pplIb39hM
JnWgeErF+doEj/eFxqEtj7CqaaGfY4Ek4TRwA9Vyt76REhM+hHKKtTst5kYTF7q8paeSzpa5Y84a
4tGFJzZ1+FcV8kzjKLjA1CsysxWTmm+1UPcutMVJOys5CRFm9ZpiqUvO2aTc2MtJYiXbTJ/3oZe0
Ph7Q7I7GLZ5UNI4V+qVQoiHORjgih3dRoRSKLpx/NCn5mJdrCO5fTar88HlFqEuvjlVfaM7haDfM
YHPi1tDEpB5twTSFMDheOaIgDiSLBkup9OyRqnvuZf8Zo8Ol9z4qJEsO51VFMD8WWIoaOj55WPIF
wLoN8JDRuUqPKzO2rqHgy5TD7dDRax/xpG/Nh2dpkXIEhH6m0IRzZ0JgnWWt8Pb1+pvlruqKaqAM
gEU++8f/2hWgKGnI9WbpYvQeLg5/geAG+YeWJTK27OD/INfxW5dFxh1IeqCxN/ksUplsi8YN3Ev8
l/80zeTDXvRnMnxyrdhbpjnb6xyla4ygSya/uQpGbJbfs4Mt6gfeB1w9AKBDgs5j4EwMRLQbonoh
5qBifbN1OTSzNWkVAbq5Vr7jjtHKUvxVQMgZpg5ThfwI9WkJmu06zad0azBbmvdsC4mCDExdqT0J
c3KDHge/FAudvzbj1k4KCWFRL1vJm+nybYo1NWKCbs4w6kcOl39V782TLCQnl1dVvg75o6Z+fBCA
NvKdeoO+eRRu1czKo/RsjSlfWHmz661yLmmzRXWXFB5XvPI9LGxEdUvJVOparanKZ4al/x+YdBd3
Vzz/5YLZA50Dvi5+wAlpNjg5RMbq+7ZwtZLvJPJq2SnZ7R6KfMDdk6bDuHzerMNl2u1HhO76Ai3X
I6NJ0/STt48sr/imWaY0/lqQm7rAUBqgA/lbGWpJUspmc2W2mwn7QDklsMKklRJPawe6rAl7IRAG
+tBhAROlRZNR7vn/u7hJkrYePasCN13daPWlR9Qgcd1KM8jTXnaZROwb/v6T+HsdcTSXLo9PhqF+
OH6m1G4679G3wfb9W9ay/yjmEFZw4EOGb7o5b4Gt6/FZVp/aEX5GhVM4mZ8KcT+mUJrO1KCwZeeL
61Q4wd8x4ALSjM/0f2ahcs/tTxqityna0O416ImgNtHkuldOzJVAr7vNcFCi43SIEQWlNdgl9g6J
LCColk1uuHJ3V0NXYK2JS+j5i69J88XcMmqM37CVNNkxT/FGEso6SBa5DQ2V0TNUg22Z0i5XcK4M
OA4ZQciSQe/wJDOBNVGi6VtUfnmdE96/RtoPVn99RQ9NkVGlZkPuUKWVuCjHFElQ9SMM9w8HAHZq
thQEcsbNlQ7dCmFsozgPPlMMupp4uUpAcajLER/BIH/gNC5E6qRpcMAZrxTBZOChWfHWddEUVJX7
GSstI+RzBnFMc6lWNRjCTe16Thd8INaNdWesADv5+yOAes3OwRjzb8eDs79g5FAchKo5GytxahW0
Q95EFHW7nTGffRBBK6Xd2emshczujl4L+4HGbjYc4itnOx4xItovMODYAT3YJmDkYPFtCFJ/F1xM
GnZkre07hHfHFIjrQGRC24DzTB7aw/AeewuK9EA0sAemuZaBFv6aYDG2jkYZJulg5siWlNZLoyNO
FM590OnmQRwGzGaNvW8zqbOVla6vASFv+TNn12hEVDzBYhgC7jfWIHbqJcT4AXFIDNv8P4BeSXAW
Ejz+pYQplMaotLNaRvWnK+iTn145JWQwsjJnEb0Draw/r8mBFN+dRqYy28vpIoud69+VcfDbykF3
mD0VdtrmibahL5nJ9Wp+jn/oKuMRIm7dJJ6wmbyDh7hvAajUE2KalUdXj5i+9Q38hMluLh8+0R5G
5Cl2HhegkQ1MgK+POSzvFSsGxLAbdTYo0iiu9vr9fgX2da3/U8vnWEidM7fC03VQQJhBvdG/Miyi
JnxZW5GeXNcK8oGwaAfsd7VYMr/2AjD1OTyyzYJEZLiXKXUITZ1742DbH8m2W8dtjhpiUNaq7IcS
DS/h6eKmoTIz4y1bnpQBtWHWQfpuSXj5GxuHp+5eP6e8f9O2o6GLP0v7XeovQHN1s5abBHEAPLr0
CsSwzy9Kc/NaLz/mGRQHVpo4CVOtOhx0fjyo97/NTVvwoiIal/GLu8RQIGS2FeklJJKFhCx6xFAL
ioT4qdBlxMOmk1R28KM+VLhFya49h3R1mOp21qIK0XfPJlge+OBsPmMMK4Y3jUC8duDQ9ukfpGXq
knY8pSUmA+yoJSATHngmLKuNEDEWCgLfqULqrE15WIStAVriHlELHREppbn7G6Hpjniw0pLGPsni
caeU4snZGZ0Dbx1RafSaMwZfA5RP/56MxiqOS8REUXSSzMjXuCAnl1C55J3lnNDpMaGdF2UJdyR5
rbZVfS8DrpCl2a7xIicn/4fRBw7e9MHhx/5jNHPgjLu8go9O7ttXeNrNZGtCynGrOioOVb9kYiAV
RKGoyHmfr+d3dQFxEQhfoKrNA+6vXjOJKlBr6EZ4nQGS9p6G0d2rtvbFiu1pocz/Z+rQA6hjTEDZ
B8wo5jrZAkrSJjLlAnOwcShaoCno3A7C2pQrzHmMv8NgT/AuVRi8YLB4ZfdexL8IoSmHIs+qdh6r
/TMOYpkr6RyprE426C4wVCM=
`protect end_protected
