-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iSDGvjoRrRf4LwE16oL1LvZIsWvS6vVIhApeF6v2SZ4iBoSpTzfvy0JViH7aI8Ri59NQmDqFnxnh
JfH6jRi9JrKVfoaMsD/3en7JwfwDlPVzHdrL8Y/c7xXDbJweZI712FvkMgwK2iRqMbddURXsn9uu
RO8zfdbAjJXaJeOuqracGRfMg+ZgDy8BHC+i1aWDOHD+iGLbll4sBgl8btietR3+8gks2pghb3Kr
eHczcje51VCdP7TSXwkTYuN8MLOdZ2xd9XwM7wd0VJyFrkfb5VsIy3W9nawjLECcWF7yM6HDV6uH
g4UYrFyiK/KxA3u+/WoLH5ePKmm5O5N1i+1PQg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
pHr0udFkrDUyZSjxxh+Vyy2M2py+rxutm1pK3AZkfqcs9mIZ9Vl7EfV8PsNpBDZdfr2cSHMg/CY1
OFBHdGC8P3fPlfiqUPNjvwaHzlG1TaE4lZc7bsmDtSuKAdpjso+vrvtH8o3eWNFdUkMQsF/03Dno
llJROrfP6+2iP24waU4nvCzxH/pRdOEcJnuOrI5vcuQB9wVWPyixqAkGc9bhkGOpUEjjYQ941vGu
w/nznIOlGKc3Wgk5a1WdQC7HChfUc4XBBdizT5C06qb3SGWlFn+UMp5UStW7kI484WvT1pgEK/re
lOMGRWKLnER3ST4Euz3iApJkz8hfSoMY09Z1rPZi3a8Yk8Dip4COM6SLQcB4D5HfKuworadDEbvh
Gc4f+EF55mGQ1gPxqwjs3c4EHlOS/lrsfZyfZ8U8K8TmKL94ano6CdWYIU5s6xECyHHPNCkyMZWm
SFKWsd6WEzp//dHe9x5QsNW2mneyp0ym3gpcEPGO23Rsp68+7sAY7pKZaPh79MH0trSU8T8HUcTQ
IUE5elGOkN6v0XMCGx/Ol7qfO+YMFug12PWn65gUVHFL5V0rnulmoTKiz0nqoFPLByHXzhsfZpQu
FLXLhHd3ImYZCiNbknSpERYtnGGNm5ngCy1hCJFGZnL4OAznYR3Oma3S7iJROLMWx5EDyO6Gc6gA
yRG4xS+Z9ADvWhcy6tota8O+ErQxmJsxgPUMiGvcPbaxrLlBcqoR6/vZHi4R03Rcxf81D+ybYh0S
7kzbo7Y0jzE4jsIV7YkrW3izr4l6xRjfXLtzI7/q0rw7boUHzmOHydy668E0UGTce3EXyEy4XC4j
6QHkdt9Qv/fVYhmKARx4s+yDim7Gg4uR3KdwWxnevzlmuTXQKPBO7Ita1lHbGjlG1P1PzM88zioC
xYNWLJeVkwTKbgopK8bB71j2QNsKntVXSxbYXO2CkKKRiGxP0xYNrCv2BxEj4hQC3Tc3RjZt4KcI
nBLaFciY7ZaJv9pCxU9htVvLGKvgl7gRsrsC6j7iitacF+kk9ZiXdtL8ZCAP3KZ3ycI8dIKn3c+J
MngLWtEqyyEPFvRtLiH66DSleWQ8H/c1sGIxSg6AjgFutsGn5Xgrz+ZewEIFEwFdI8MvZ6D3XSLj
HrcMQRZQDBjUgKYrP0AbwNUAj1qR3m6uFVJPaqXATIpuG5gJwZYdjmcwtKSG5ZlYOlKTfMwESktc
xQUjYkzQjFMlVNsc+Gl5yJk1104r2UAK0tpSymJgbPjlpZsH++t31H5i1ODvQLc5agrako3huNVg
OD9GrIufFE1mSTwHZ1UUaozZb4Jyj7CpEjhyY/ZGqsDwzfKTWTwjQ24Kj0BrTR5pr0Hc2e4jyrUY
y4PlvB4rQ00s25fZ0QxPhaqOWuRiVwPgD4x02AAQcME9lCfytEXUbs/Mu5+KT2PlK/6RNWzlvxxx
sYy6fVnRPfRJlEweUEcZXxWQK7wopYg2Yc7QMyr2Ydi6oF3QMhc6F9GLCJuDwPf7Sjmmau/hxhbp
BGUz5ByKgnKbg0uO9G5d7ROJNcNm26CxEWTyw/T/dOgO6fpDjlZNaKOSXGs9u+ELv8y1Os0dOeEs
HLJr2ax8wZMSKzikaJLLb17UmQCDx0GnCO19i311iK0AeFDx2xpN9YWVe57+L2PRsVTMXH0e+icF
YR5lhRRGtEzj/uzOzG1VYwBk4Dzt/its9of0yMWULPAwgBP68vWgHQbo6yevzC7hQkFe28QWmznh
tmloG54zK3+iSpK01Xm37JKfvu4CxxBj+0RNF0Dk4vfEHj7seygszaBHBJZM7BhtzqILHHf0eYE3
pEOr5vraBHbVmXpRDWWP+v42vEkMzywpLkszO5KIjHyNI4k62VHm/NW7cYOrhcCIqVUMYocOK+sE
JG0laZRS8UEAnhc7AnqA7eJoyTc8i+wwWlPiiRswdiz4TB452gBCu8K/yXJsgnJftNTJ/tDz9vCV
He7GQ45DYZ16Q8ngtM6B7P7hO46jLCGa+vLOGA9FOlbhBV0lGiBcQ84v7NdJVlGDOpEl0KXCuoCT
dwAJJ7HY6XDSiAihVs3mqBGMVFKG/fxnH/80R6LsMWyOW3L9pit/988ConOFqrKdtdCEz6KJoyUI
FHz6DgPiKpttpMYEtV0fOBjRFBlzlpYyB63IWxPHdZY1upYrlyo2HAiBJch236AFHvaHPWRGIOi7
1FZH5mhfgNzSa4pDAJKPtT/IQPe39qJaI38PCT0Qm0jRsuUgzjg+s9cxC2JP6hcJNI9BclY5vatC
JBuN6iSZih3lBiHkAr7H2DuPBE4lqr/RTYCmd4z4cR35RCFg6ZFW4IzqY3UbX1+Qb+hNfVXfuptu
v1FzFjzrpWy8psfB5RQe7M0pb1/7k+c4VcKjEf4/2hN6/1LOyUHP6BOIy2wt6/YvhTtZZxwnAJqh
FlMuMFSGzwJsdroQLje/U+w3hzYFwNcySMIvFWINwA+SAr89BfA8oP3vTEZz30gfDUioX6/vpp8I
B+Frs7zQURAZJIT6zUUzh2+PbSckOtVukaalPdGZtpQoUA1B+KRhLm74LtGOlPwX2ftvXolV9vJ9
hASVDhi336KK71RBLE0/2DjKFicUt0D2IEIXcq5VTxPugPoZ9+EOh9+9i1h9nSquRxARS/0WPBR5
7swLcCG8vsnXnPkVKOlimjQFgNmWP+QVlS3202r5hWIpoMN4/C2whKLl9Xrp6Whg+pPMJhVfXJws
0dbKpRC/YzErvgQtgQgFJLnH2FduWPE/RFAfsPM+yD5VXeCh2c8PUnG++VfJROIE4xEWmi35hAAS
WmTcM9KZNaX89pWk/gaW2QuxHvvorwPIint68qX0uB1sEJNTlYVYgkg6XNVzroFrcwEpnnnmfW39
QZJwYOMmiLKjZrEFWEYydkn2bMSnhZkbT8Ge17zP7XeyMrc+KUwB6u2aTSrXwt6MQAzsmHPfdZmA
aO1MbNMXhuM1sh6EOInNA5fxouphpaRkzKPF+NumkefIZYvixXtuJT/0F12TBSYccmcGCIhtNAdc
4W1EYs3JQQjZdcSNHEmwkMCkxaFyzn0u2Gq76cFdHByQnzSDgBQtp0vADnLROmgjewmVsMrWbMAj
xVLouTIfS2n2UaBLm8V4kZfbpCC6mRpz5dBxw8hSxil7VTwr4juoJManL7PLQRw16aKb5SSpDFhE
IcjkoHIojHyjdrXC8cColFHwyK53Qk3ABlOjvEI2cZsvdlgjneAX3NhiINaJMDuM8e7FblW95H4c
/eMlx8/IYfOsC6vEU+qye50Is/YO9/Mxez56I7LvlltSq6U2c3wjIWV/4yWDiI2v13COxaHq3Hea
83dFrVtvVcX2LsvBPqTssBPh4bHUpZbMXhwsk7Fuy/8lT4Oukp1LRwQHHvaUwcN+j4yB9ZmbMe9F
2S+mrUR0gpfP4zQi0H3OIvgzU3n1q/bBE86HeMLIhZJ5KLLmiXJzc3ObDRVMO2nOqbplo/EKPCKw
p0h5CuP14m7JrSfvsRL4FgSjMiB+Umfa7JgmHOHWozXRzjnu73HuvjbDgpDn9vnJ6nfWFSU4N2Gt
kiPeXJEked7SgavEtTHYktTbErg2en161j9D40hKP2i9k57qnUsInrw2X6N3trrrk8hKoEeDX4YQ
f9434DZ8ZUxd7DbeDg5Av9P7e3WQQAl0wY1iyJfjwI/5xHm+u2t9hW7iLJoQPHwiPFGPEgqXxC3E
xbpGdn+D8BrX+i9aylC3pcjB7VrY0YeYiArJ/7quieVp7SU0u2Q80hvzO+u3dbCWe7hmYSUjU2gQ
KkhLZGO2z68XMW/OL/ZAMg/mb20G0YxKY1bRWw0hUsOeR8ZbDmC83NEqJZf8b940DF1R2rO1IOTh
bTmRLKdbbC4AvJDVjMEObeuWlisSMlaSMNZb6SCNcD7xQh633oGmHU5hit6jfIO8EWLjQKqxZjnA
zlrRvAGisc/onSUoFxBaZw82rRSVTsFvY/uiKOgEnhnb1Ex447rdVo9aXpJv41EVB7/fRUUBARG5
KlF8ck5+yEbMRaXkZ+2fr6SIOhfLhDQbOESFiy6yegntN9Yw4b4FOq9//VzxISsJsCZF0o5HxXSp
8Jj0BJo0W8JUB0saXD1Khjai53EFLyYpKFCPz6wE7+0E/DMTmCpRX0VCgnfNNcBk7u5+KKwGREsW
3wnxxU2QvsSpSv2VZjOBxuu+h8GClr5ruzwDsXhmn7llKqGCHT0umML7+rtqkh2Dns5q0oGQnIPj
68KK6Q7N63wH0WKi7LEWd516+vckFlcP9z+Zu4XfshFory9Og+svQsuLzcB7KM6Twom+B7XvImPk
4TLUIzIFSNXEKnEzdLclHWG4dPKrrmmN8LX77dJu9JbWFpolG8aW8dXfOSsoHn26qoaElGcOC5xM
4F3OWExRh41I8RoZ6XT2tcz7h4U8s7KyoniF+q79rUa/jZ2jdnSvLx526p/iYMpeHbz8kskO6j5n
snGmNbIkcZ3qdOwbu10He6+xHrFwyHtDuuhJ0MOH4Idc8RA8sUGeBRIhvh22tcfkOhbE5Q8WLjiJ
3e1N5PAVPh8j+iEPfir/eqpiW2oJvjHZkZDVXwoFR83QU81Bll4CBRtOFXczjdssIcb9+de04lD6
+00sNziNz/Q7x/HVwNkundrk+ELvjn1aPbLbWtFVVC1/TJVUsETQATL1qS3J9x/4K86EV2t1RaUN
OgFW/1mzUEoLcEhjw+qrrKznk7GUxsJZc/IZ8F/joji3vbH1vAMHOT8LSX5tjCpbuYotWGhBrYoN
sSConEDtd/DbrlXwaTDDppqyBLsP0YbEtCyVCcv+zQLYNiHpw6dsX/TntyZVBkhVvmVx32chFfLH
lbIuDAnCNFMJrTGkGcsvAf3AM1FoEmpakuBfChLNvDiBJQnQktaD1tzgCtq6ifqg50n+nhInNYTY
pvLXs3LNe5aokuZ9jbcfxzE0X0TzBsZpSfXDM4pJOXplvnwIeGnsmZggHn8KkxPvatqckDausHYh
7k/yaz8q2jiL9Sl+vnUrbOFnDeW/gsKQeEc1Lc5bOAPRsEARLl2ogAJ8XkoPb9rH66atMLCeKxxr
FzuHXMm5050MLnGTAR0HwOxeDpPV319K7oBxyampzWGo2OIQAq4Rjwa82W3yDtbqVdv9RClUB1ee
G9jT38zWtDE/IHrh6r0nhOMtg+Kqk/Shoc7kgvU4TbjdryQNlMZsxE91dccHSbcJwKJImAnNvgBz
/r1278U0Ik7gF8PYYBdmPvev0b5En0RyjPVMshMpGPrYjSGj0dP1HGVRdKmehynSs1XrIcdDi4yv
RwjObF4BS7z7eZ1DBSXHtsQ1sqbrFeyjKlcrj0TyY4RbmWaPB7z2A9jb0auAZa7EpJLeoSqDqC7Y
yTiqWmM6+htz7S1K2Gf1VxWKzlL48Oj1tx0ada30DOxCe36muyeS+TnxNQ3a943AdqO0AdFttG+m
cngfALAhaOtZ9WvGdhLgqyK0f4URelv1oMoE/Yyr7weIta+Hn3j9HdOH5qbdmutPMJd11c0HwVke
fY+1CL1qRSz+2lZo1E6ivzFsl/xuiW5ANwxHTlg5OCrMAF1M7B7Y/POED8L0UACZD1CQa6IqGeZw
DXyngs5NMWiJcRJ0jmUvXCJEWO1I5FhoKbVgx22nD45arfhrhyYTcY7T1MENXK5U0MQr/Xelg4X0
pLDG48BLrLDxpfywQV6X6xYU+3IFFhuFz3BPL/x+UXi7otVretTvwpSJkmglUrf7wXOipoYBk4Nz
EY0R45zN83GzkZ4ount5pI4TMUH43dAn63pVP05Unq0iSFJoeH0ToXuia4szG2HBzojHKs04KINj
5q3lKNl+ARbBrtUoy/c+UrLxOA6rGK4VB9cm2mM/OAZMtZGOEFttOmrVQJPyZmFJOX8TunJvC7R2
yV2N+Iyu5vEnTkr2ISYAMXrd1dcobrJvAeGz5cGISLtYwbW6YPh1u+FoJw0d+5+jmPTKXCYko0iE
YRHDCjMSkH8EmYT1OFny7gRhejv6H559Cjkplbe82XdBgxwBIFK6DRxkDc1pY5YkF9lBuzC8lHrx
dxuQxCTTEY9U4jw8iVJ9tLGcXfvOXDnbaH0qudlHOSnjYCUiflU9yZhxHYGrLkIcYPhFiF8GqqhU
fNS3+IBSTHRAG3MMWYRbGlTXkCpzm9rui8N3pLu3unLpifsyqORE9/TFtFeJHQybPDrQRmOo5STM
TUa2BWROub00cElOCltL8MUNmeD0bwnBxiZI5PlK6NAyFSWYZQ38fr9XflY+XZz0XtM/Rvt6VijL
6iugobc2twS9jDz+K2S/Yz4xbxJis1UJ5wMOn7EwMGAf/dvvxjzEvChFoWDgX4E3lCukNoMNwaSc
QCK7f5H4i1E+84veqxw4TZal859lVbxUQkNos2D+ofY466qT5VVeAKwqfguZ7RqEYfAS/9e+7xKN
kBqqvPnvmv4GoZMBhSWw+ntH0p2p1fU6MDEerfo4BYniCSWBayEww27SDtmEraihZ2fmo4d6kJHb
Bc/rQxh9YDcO2mAGew4KhFGdebStZftWqGwuQAKgy47IinsF0WcViB0c60g7HDFKSNOkw5wPPw04
Fio9hjZyJMHyntOYWFYJB3UYz2cIt1cfdMF5d+Zl5fGhUXonAIte9hwx5c62Ls5LrnJi3oNRW4AW
J7NhetnUN0Q+dnVwskyprypn7syiSHjeSlssGtsmEQbk9jNALkcb8IxQj6t1e0gXH+nzISba0aqe
yYwZ5LQr8jEIu4Sq4Kxr92PEjqNIpMNymsIJ+tIlabNlF3YtXVqRTzqA9VvttrOdK++LlDDO3Ryn
YlOmoegSLv6MCPRdeAb8cBtVtBVWkh6oEotLnu/xDvwrA1OqFXzmcRS7DY3VCa1Xkgws4ccXC99q
urk5VpeD5x7Xv0NAutDOCvma8b+T/DBboFTKkP97FKblVuAWv4i1OWUIS4rG2PWDhvdRBi1NhmdZ
cmb2urV5D21nlA/SSg4UotG935titCzxRfLzdQxQ9qQcYqWSaEBMih8Y8YQSVEC5uhhajc6Cs0IU
jhapIMYVxxvSmqPolU3tPg8Ij9iZimnUNNS591hVE44PudQlO+/Uza3sO3RILZcU3EQylvuTMzmo
my9fvEHRJi2VK0LfCIowySmB7YccB6MObuLEqW+LaJGK3tJ8nGDr3ln+bRHg9U0Dbz870aguDp3f
gcdZB0JECcgz7NQcWkSLxcrYip0Avi1BVFKtRkTZR7DgnWc3gnIlYQGgruvT5Z8pHBpUu50hb56K
RwhyrEVc2uV16iknhhX25Q4AZ5VqBm+tafkWlE7QtgKXjVQuPiRFiiil3q9pXlv9ZVe3ZnWgK36a
pI0uLFGKcOh9r6Hrob1AvYvXAWWaUi9/FMPaiQisbmi8m3hSIZpcEfDzUnEal1iaM0gV2yPDS0Mq
ybNQvN0zwOX/SBS2zr2b1D8p/7J7rRRz7RYOido3Umsm5LYPWciaohdoFUfH56VRIIkto6e0cnk+
cfP8d/7LTHaeD5xx2jUPoOiOgtbYnCYwODjhvtSbB2g0PEf4lq7QFaIkwhVRCqwnUMQkAb1Z58uS
nEiTYjgvRPlvXg+Ycr3/Mtc0vBKPnF5bLwdtHrmcZ/S6A79apGw2sGemFVSDuAkwP/3X9gGZV0Ea
rK5NpGxOQgpu/MgJL5YL0UtftFO5Biuvn4S6Ij3Z8XHmB9PaDbTlyeeRDA+mT+skSiqMFh4TOkAQ
rDlvKm+7azJjP8q2mAu2dv94SwGsQiPwToQ8RXq5Qn2hpBJhxoNusVeMxhBV6dXuLcHBAm361R5q
OZr0k7D6Y7twp5RloKiZSOar4Mjkm9lAY8+HHR0+pppxjocK+otPKQmYtW/pu9MKEZIiUS/l5zV4
FLSVAxepv49l65Xtld5zjc5ZeMyIfffJ8x+tX5CbOql6M+6UE8znC81waKi20aNV04lycksnNqjh
il8YbkSmnH/7Tere18qQWiTyyGHgtsKQsvIUcazTzBD32VOiu2asXgxTmoifQkT+QoaneQDghhNk
8vx54Ie8n4m04c2rZlnFBcjyvTNMKCxQdPOn9aMUGGvkeWc+zHlIVCKzStz1pTm1E+lm+rXFHoni
m4S1dIi2H4wD6paS/5gpqCe7hnBEmYYzJ6TRB6WmYnqjCdwxoBPV+hCL2epQs4pzsfXCGjzoI5Ml
iN2a/NBeOgEzPTjIGNSKzJMyBtqUNnItd/QhodttfN/zaAlxmkeFWCP/grMj1BpcEFa/AG9LbmFK
wkqVHrPTXnXY9AOrXlSNxUhgOcc2K0IGvJaxYSYjCc386cdEGjo3RylLaPSdq2qYeO0HQ3cdv+7F
AexuluWs5oSvCE3BqgxfTo3FidmSaXHkCDEnNHyFiWcHcsu4hRbkgL5QRlBupUpVoFMdSyuNgQb3
ejve5N5VN8Aep/C4LveY+5lhUOsCpihUPXd7Iqjn3p5lUZ9fwnpxazB5Pi4tTq9LXkXfaadXeYTe
crcxPaNo/YiPxM+iYSj2wtIQfUGcE3WUR8rxsic90ILyrPkmuvmb6VyRILXgZ+BUKnsbP/5d8qOv
I10XGeIr6CyqoYMCA+E21w4zx71zZ+cGoWQkJ+/MZgpDrGAT2Usfc680IvQax/RCDgSrsGpGM1TN
UUGY90nhvHkrlzlBg5/0EpP2+vHvMmRfT4WUZcC2htaYYhiqzFdBIk/sxSFoFPKQZBc3+Ih7WgFN
OSJd/rFGognejY/doY+exDtS10BVSnCb6Cn8OyL3+JgK0EQnVlf+gw8vQY6VECUAPUaTUN525bx4
VN03g+GPhzD7k9hKwhkiNOw+jSDsUxvLcZmt5BlyLXKKdmW4Py17+FR4zHc+iHdzomrW+oZ8AUbb
cjvvvkPnsqhJPH+UL86WyxfkOZFkI+3qytaJKvOShh4tKnnpaioQolGngpcGazRkqo7eqb+RxAfX
dQuhGQFpHHn54FKKq185tdRrZ2yqdRrX+muPyrWSRz68fblLfWJP4NgZifX7SpeQhI5gsPYAi6NY
2HmmPdIfVTs8ZLFOgJduN1uOzvfX0og8+0gDPaJjtVa23l3AgpXbZIDqfF5JcAhvd7tEwUhU+jQH
6lu1CsZlmCdxGtplSpNf9RV0YFAlUsQbVrKuX129ax4aDuho8rKgmA7vkgyMTnSelCDvU7Yi8VYS
F3ABaxAvxwjZ/LGli98dzrFhV9aUCU7pBTtgFDFOCkL2+0+FxH4SKsu5vrABSSLJWeigmRStMj3b
A13M3QK4RYZAdpkABIg6fIMvG3UewvBgCtSRb6CDuXVc+CXRp3qt7nFuTl2XSfDSMdN98jslRZbT
rogI9M6tNPnsMw3xDzOkcYGK4zK7sJagrXBohzXMQy3K4gkxclOaLKVELfkW7m2WN+58YWl+Wc0m
As7kvbqmkvs/mtOfQ/cCx1XNYSvFrXTcbg4GG3TRwgXIJjd0jK/uO5A9Eheeu4JDeUU5oTMFtj7M
14uGHdmo6yzojZAch8KUQT9gP4QwHPOBFN9unPVr/T/oW1baBdSZfXZ6+51XYYbYKJ4K/bTmbyQS
OOkUoLcLGxyrLKhT2vMlV4xuI4nVjSdGEsRFVAW7i5Lawx2IS01YYBJu9l8Cb7zwB9g4AL0sMGWu
AvWnadab1KECS0KUF+tJc3U7Ak5Qu4ZYBrBMEI73v+C0eFcn2pztTW6mQE2i54/Ig6c5GaNpYN0P
h3XuOCECwuAWRgTo2YM5hNpPMhGELMSUX3MyqiOlr9+OjExA6CblwUl/ekNHD2u0xOnYMDBO0Fr9
naP+kP12rqIwTi2bBYNym9/p0hyyk+5X7iD0qrpJVG0fw5tXUPhSWyBWpaMur5BuuloptFoUFpyd
CZNeM/5hP5mm85I3/iWMsu91cjdBtmgRfXVIKKtnI8YT3sDXKpwiFsLRMsJYJEW6qi31umL+oNpH
pvhO82whpptfWeqYo8wBeUXOhBp56ywnuv88ncmhIE3g2pMM4vsLLPMk2gYgKTkMpnSBj+cVNbPA
cctJpgmW08wilClX7wjw+xl9nB5fI+lA8nuMemO1cinf0tY54aS2m0SQ47XXXT84r7rCiJTvW82+
WGPO8zkVMr2XLA4ohsYCQadg7WuyKsE8hd0dtPu8v+i0Gf7mYmfL6i/1vCQQZ1RHRTV+qE/iGn5D
BeJvBorxuoodRnUZhQdgDVBPrn+11n9r21OvPXWC0ALTF5gDCl3fI5PdiBj4YrnQ1QXPNK6K1DMx
hEWnQ5YC8h+JtQgYHqRgWtPXA9SneU68momwizbiCfS802xgWbL8+AMOL9MSH5C/c1/BHfL5fevj
P3VI/zSTWmwL6yjhkYmJx42qq1uhiZshSL/czzmhEvZp4LttMs0+U2b5M9hC0FVAgx/mGGL63WOE
rn0uaX+AEjQuroFb5rpKaz7ZHc8IniYzk7C+GU4EVRyjg3hXlHRTFzCfRr//mtVl/9cnO/Ff6B3H
3e1s9Pn5ReXzQgbQgipm2KQdVV2ppzUVVyghBGIAwDK5CDth9OxGsIELvZXHNtFZcMqvqE7SAQ3c
rAxKCVaT6VtU9im3SlQwYIRY+bhtN1CPHGt1WUy1lgFSz27+Vs3vkVRyb5pn0K0wdcWGp0Z7EzZj
Jvt8stH5pdRNfo5XIdUVT1U8WtUMoZkIKY3AMjrMXtyqPATC6hlj8NAMBOSv5dn3Q7UEtvE2yIiF
/xI0cEIxXgOBMPIoJJiw0JQvRPJRWarLOdi1HA3gtDLr2lfU/Vbs+NTKvvc/0bw4cIzrVyG4CSef
SZV8W+0yKSVtsj9BYZqSCfpuqrcgoSSncH/51fmdpj/P5lSXqG9nAgVBj/vC0lZU29hPvuKWGc9u
uYRhL2Ct7AOGMDamhHURgE4pROCreGaBxtgTpGozfxlQc0htB424XqGK3GHJ1TXhJsyrJnuBTP5X
OzgeinbsjncuOPVsjqbRNNgBwS4fFj1gtT7mVQLgD7TuaYPCw8vNOGAwRwAjiwrp0F/LEeDolZfl
6v1sUDooYHjG/4IppaLtN//1IJEt6NxeiwNfSPubJLKsJdMt/nJJqhfTMZ7iwcswNl8lvTycwAh7
ehqO0U5x/NyjEj7oCVcp2Ao8LKuo1f3AsTOjmrzSfuqc1lBANQ8GhXGGzH4+46BH4EpJcdn02sdZ
cRhzvDu0VOQsqgmmk77iF+xv3mzQnA5ojY2gZt+gGD0VaZB1Ksg4PcdEt39e/eiMXOtduxLuKWBK
JtB28L82fZGHCkn1iXu97tbw/xx1G0CmHXgaNgOMsVWBu9wWlQAO5kKpZAKXnXcI6H2CitziqLOH
Wpx13VBC/pqx+ujn0GRD4lVLKcC7TE3kc21+YH+iYb2K1YlArtECHzI75sIPClP07tzee4q7kRzE
GYAtfWegfR0v6OEV1aMAI892mhrlNp/w9LH+BuD/AXTWMrviv9d/bxSTM+bCZ+uG/pB4JJEpJ6Ud
iYAZJiUFARtZK9uIBOVGLeY/b8JLzTZdXCneMCH3f3l0PJDriciTY11+53McLB95HwafpHt5Dw1H
orXJFnt5T5iMXrREs5tpa8EpXOB1sA2iDukLjnv6KUFhSzKNs4kfGKN5J9a1c9cCpnKWer633t1f
XZMWBssZnk3NrayMgy+NoDVJdlunT0Mdtn6fCAh/bGXYx4I+yUjIr4RDi9kYUx3TkBDgjzrya6hA
fAHNHuSxruIuAem/6F4SoN0Z4NcsUVCaI4ev3sAixGuLAMtwooNJBdqGGT1+ewTGP+fMIsfS+7kv
o3md6+rTfGJcFqx49j2yEkaIiXSaHtztbl4gpM+F+HVY1e5huH9LWt4yDJQB+2nR9buQokV5LF1b
0CYKDlREwSz4VMIm5OkyzHNbda8SOuY9Qa2A1y16snspgfPNaKiBaR+GF10mAQAcl6dgDyKXaVDb
kW/UxA1HbErZRxHj1OqV3L94/Ftffhu4egisVEkjGOvg7amjmLuej4fpD66CWEXwjs7ly6GY3baD
WdjiEJglg4UCXBcdi+AAhiJgE2/8u3nUWHtEMEQfAstj0tUpqY9T6ukOCtQ+k9yrNynwFpVr6TnM
cghWVlsmBpBd6QXck5jiieKW5TE1ysb18b6A57a01kXQy9S8LzSEnYD3XCdkX/jdgk4CWb2v7X9B
ny0atz1e4Po9NrGgvX02tybODAhYcU0Wkoim/yJoIGLkcgZpa9WyVjwJdeZHogYIK3sayZH/Wcrm
IStoZpYtHFXoDV7lr3CXbfOsGu8WoA5YPSYxS9XytRwNshjyXzLWaKBVbV72Jfa6WJ9D679I8AI7
Ihc2iqV0e3emljmXTSBWMb1dQJwAmZzGWxp9sOMmjwYE5Zr7y+nY8XhTADCC1jnYMkoNoH8YBmEC
GWu/Jp4WDeHeytZj4DeWWTjZL2LWRjkOwWZFX/LD3AaV2yMExrbpnZItp6mIjFOXHe3cRtDeNkxK
kgw3gdxNcTvGbHa9S4cl0lvN7pOZXTRK+KOje8AupAVx9AQsG40VwxH9W+TNKTHEVrNMyasEhw/j
UHkGbLz6sAyDPOcBSHH/msl322hAkOpHIjfB4zFwgowP/jO9AsoGASiBq9thArfjLdKZ6446PR3I
DeXqm4Y8B2j/abaZGTcMz3D8X8PtLRu9uV+WTMilJxnxoNQG6zOZvsSZ+l1orY4+AbcLgmAdppvu
147fLS7rZiHhyosq0GQeljgXRyUWJ8eoVeaorl0EMMEANUUBFNFT+JGg8XLzd6THU8P07/9PYTjw
zYQPxCM2INkHKjozuwVDglLqaCpOXsLXlwOFwhZ5r89R28Hd4Qo2TsAOLCwq4Y64wmS7W9is2kmc
rUcS9ZbLWxFwLO5dWTV4ALwu+14oqfKzv1KL+ZBgnZHaMJvOEEh/8SHD6cuUpT0UCibK0q/5zK7S
pEsvlbYPnhxKWLqIEqLy9k6/A6CdxgSP8+GLEtx93k7JcNQ6chnkmsWHb00vMO4ozO1D0Fi4HofT
wzLCyq+zL4VO52SnyWAJcDvzwoUhRWo4pEc33n5MUrFqsTc4Q/WC8Fbzg5ZH5kkw0hmjbj8GwgmH
wmuNyPAwA/DTx7MF75R8uFIvmGBKlOzNOxCD0h1LRGw2k6zhvYzyytbf4IvHG6b8esvl4BEJj4dy
gvFyFPTcdKzKp7E1tQpmC45zz/XO73urVSEhxNF+WTnNNBp12iQtDjMo6DyFWA90v00epaVwuzGM
R8hRk6lX0e2xIzkswO8d4PlEkAEh4rTjjyQR+LscKk/Rv+nq1X6Vmbv4M15z39nZsAK0l5TWaNmo
qMdyD+LUu4m8FIhCHiVewvDB7+1G9WrBmzgFNYJV99Ir0fTlh87Q91W61i92Wre1q18sp5BZ6mmA
zNgL8dYFKex+f0m9DG6FfV3WKserLGd674nCfKEKKoOah/MPEVl5YQUtTVeYfXn2MKuLHyEx7FrH
QqeAZy8JL60TwtgqvPZiEJ2XuVZ2SlEBwND7m7A1pP6KQcIRAvidmaWWTft1Wum4WnBQRiXHb2jq
3m/QI9jNDRxUALIw5QC7PD2WzFA6Zjyh/8YebmqEZN2S7Lo/We08heHtD98wu9CrpNztLLgaA/Yp
ppATVAijLNyMSv3CqZHF38wj3B+YIrbsrScSPGgLtgcn3S+9i/UCoKt1k465eHUSiH1RA01rk0TV
CIO/q4YphRadQtm3lGesz7Mga+6o21DYAZKYlMl6EI3joGHqyIyyDBkv5Iz6no4r7olLXVlEAs17
VSvKkqRWs2ym2ArmMC8oNY8hHq9lyXkLftSjykchfDP2yhsL3DnXMeaCfpSKVcY2zgRFYFpssvU0
9jGDLy3oYr0zDPq7faZ7etHtRII9iw1c0jV8UuIgF4aI59iOdUXLCqLxO3dhkBTdI2DqJCYRcPU8
VCj/z7ny6I+Ly45avcndJgzWU5c5WWUK2MOJSh4/cjnuQ1xzWQmC4+AcpuIJrDCwb3LwxC1LE30B
6XtiDMHXKOJY234R57JlnykMIW3uOsPZnu4PdLiDeHI+MfSJk51SrQiF3F/qlQcf5fnILTmbalFP
hNnbVNdDquBMrMRNxp7bY5wW3J/hfv3hsG1n/eaBeKltWVMA/x/KmuV8mcbmVds55pnvgNVzC8Jf
sTFWRE6aRyFH59Dl7hMq8GKsw6uUGc7LtHITQLBAs3gEjY9TUyj1acL0cwt6rMTYKlwRx+iTDqgk
rT53TZL9YLcNvynyalrEo8c2Ca3mOiqba8W5upL7fUe+PgYZZmtpm68uvK01X+hBO04Q0mLz2acq
gX6cw2r3AR9eHOxioTrUH6gBY8akg3LKAq8FaqEsPMssxjNz87XLgvlv8IIgniFf6eKleLL8FG3z
oMcsKaTzG0NLkPny3/xlRoe7QxVxINPvxHc5gzgcyN3QysY22biymRR895RBrdtsWZGMLOBYabdA
UOLqViApMndoIXFeLMLypqSWGLUxU5P1/dzRmgeqjhp00pSnWqmHkfhgjrYny/SD6mNLZKErGDGb
zI0GuqVSHtGXysSWOtWCDfqqrUH5t7xqjZZNtP4Cq78g7TNjMiVujbkhW5hb4JrhxsXYb8nzgE50
iq/jsIqMlGxeVDY4EufERYcRpK8W4vgSQNQNDe+QVIviJrtjdxTBlE25z89AVroYuhdSvBntcjbm
98ocnPQTDmUh8P/O/WuKSkvywgOQqFmb44YHzGMu4ZexNIjO3shtij/yGYGo+qXFF4xW4glAYKs2
gK3wsyzXCV8/njeqjDV+FsBaHf13FvDuvSXgUdvI6AtvsLcWJ+P3K76wAKUMutBkcNCakTfnscxV
O7EP+D/rY3Ii3KvW49LV6FUeY7dyqo1Eh8D1XOBlZy6nuW82G6zcpenSdL8rxnTrradi4Plv3jUc
+IhHJ54D3V8+WWFCV6RGjlw+qZdbSRgV9rzC8oy5d0QwJK1qk+YXGoWM//j9aiAZeLvM94pAAjtp
xykNi4sImQlv/ZuIcbYJSAIyIzR4WjwsINyVk8mc5/0xVRdulnhGmgiguRBvCzTl3oVpVM7qMX/t
WjRq97g9cYy8IwE4se5TgcSDmanL0g6vPZyaGAuL8BDZFxPKHAjGxEPdVV/Z98zI+u8u4bkrl9M9
Rbc9fPriVMoSlLZzLdm3M+naCo68pZvJYeNxm2mjphlu/UV7Fh9vL/eG92raM1EI8OoAMDJae+ZC
0/WrC1lj95N2ZAwD1SAMesauLoGpLS4n84pG5bFvhXz2GkEOQXkXpqlYI6IpWU6Gd3LfB6R2BvOU
lMZklDxSyPN5NLKwEAwWEpXnl0NaLfBvYtDms00xFXCVDPZFFYNBxDs5NrdSDpfsEPjsRtZgthn2
2xo6VAHHxGKBErAStLzgdA4qkv6fB0hp6qfvEu+uXhWsbT1zhGumKCgs5lbY0jL00WdurdW5oKtb
PHOqeV9B7qzvWniVRrjHR/V/dUqgpUdiFoCrxMTuGL5gJTRJkXwdFIrO95TpmGMxG5YG4ssyhO7Y
P2v+xngXyUdFNzfhqQUEkkkhcck+WBdBIheq04AIlJzwpCcCR9dNnSvgv2JQ7vm+E8SVeNmNxhOi
Kecif1nlgYBpwcre9NC/nPHiPpHuieCD1P407Y6+1dzqr+q6pdRMo9ozIPicW0FpEvsj39GlEUSE
5VXBWAxQwyC7GSv2gFW2lE1sL9o2qtpbunGjhSm4CQ4/6WmX7kKjhD0zsDYkQqP6tDyZvwOAYnk0
gqeEGHwgJVsvzVBjuK4/9Cbb0f/XIm1y4VOQK+gs0e2GnUa6is0CcvbEDjRQoOXyQMJqdNw9ihrq
k2JcU7tKZlnvNBD8cAkIIOSJD7OxzRWZdBH285n+WdDTn+IxmuMQ8tleoR/3JgyRmq8e0Io5OAZC
zrrQvwJnkBtQMwxDv+r7+K9AUk6M0+nBH+j9hbzqd4EqXZJDR0jnNivfNJ+7KR2VFSyHgNoXjT2a
lTBUASpJTTXg/qq4hzFDXEjzSXAPszsAwaChQ16YzTfRw3v1ZQuTALdMHFLglVLIlcQ4hcdcLrko
rnVjhWcRuMbCSGnsC4GUdquE+/J3kjL785O3N1Fm08pUUyHqZ42a2hdeA/1JgU5bL/sij5/YZelF
fGyVoD8b0IbGmoCwwC/M7YnhYG13+SmbXFFG1FrmL+OqkrBGq3Ifkx0RwhbSGjRFe9M1D6bzc6TH
0ROAlRmF0RaK3XqwnYOkFQLbjgbWTiwvM3of+lGXI97xRIlh1LzGS9S198Dx8uTq5+oCKz0IJspS
aOd/Yo0mnxxHZhquW7gj8BDIiMUhPFQ+CCcMaHzt6EHK3Xa9VNMpktktE4ZbYFN5I7JWjN9q9dm3
4kJgv7h645gFTdaJ2reSBsWJ4dSjOTl8Is+xrZKcC6+Lcq75nW4vSFafcJsc2u8SaEYBewHLAgp9
K8e0UyQHcuhnQiskN3IoGMkxMh6KH29qPDkvAeyXU5sWlqA3+mxQpgBMhbRk+vh6BVwAtes5OQ95
DnGglk4z7eXKd01B883gHekVu+0fM9s2Rby3rpHbmPfpD0wcIMVrd5MK1ukpvVXBpvpbfc1BdXdI
cKnCFyE4VZQEUOmPuiwCl78qVKsJ3EpC0sPs72JXNJcOe0n0cRrIbKRC5yUVLKhkTwghPuVv3VDJ
I0sgDi6Y31RKBrnZcVhlY/WdeTPkZeYNiAUdOLSmufR9EcEAMEEuVOdLqXB+pNW5pF5FE7Bbiw0R
DUVnZi+GExAd3C6MT3B2zGlWpiRF6W63Im13a8o3jM8yTE46I+9uMD71+ARG3k3bv6TS5Ao+hx4f
GToDm2yX1S7f9TBRJMSCj3/86N5vfTseod45McQ53j3eZrz/kg6oexXkaSpEXOg9qMd50Zetckqi
7LW2sk1/4OVChN5hU7NC+hvgbjqzCC/z3JOkWSlTF/hQNJkXEmOV+6rWbWVV5QzWJzq20WzSvI83
FngPhAUCpCJfVDRhpws/l1xJcS/XADTXTXFNwVy1RbJ/KZZEaaDUxRtPBg9WQWVH+L58wYvcMFYo
H3a4cau7AuY+Vj3EE2+z6n+42nJxS2yCMitFrRdpGQZ6FdgwW1eYrSxsc2pgeq18bImshcKZTwFt
o2VCwUrD3DWPYzSSzFs2l4ZrqekwCR9aKdowlsBHaVpDd7ZuS42DEo/pCJ9sScB1srykEOk83Zzm
n0RMBoAYXKXwQNIJGZqOjTCEZo90iq/efsUFyyYXwYm96H/pMi/gbtEBzMQI2PDyMCVBS2hJ38/b
kO/72J3n7b5fe7853upmuoU3jkZIwZqzaY2suE04xfokoS9ZMhQnykY9E9cTnEW9dajLVAsuBCyT
+9+wgnwdUSbusOxztlT3sFSng2LPK6dJEbWjgEtLuUhrE/zI9LT/A5ONDopXviOAJYWlSbtcOUjG
clzEVf6Q2caRQjwzvy9CRS0Z23cGWayMlRaZGKrBn/lQ38uvaIZ0mNw9cfwvVmyL1cks9KUp4X5j
T7YBCFk+YWdS61nj6RsJQzvfpLx77+fn8w+5vhK/ahNY5jmtFh8jfbx6fkxKIANZbXBdNzkeb6Ln
Kft8VtDBuytDjkb0NH97rXvm5vxyaInkF+h4z4RBzKp+mc4gpaME/KOb96FaLqmRA7r9hDczUvY6
bXEL1WFU34HyclECQl/eXcbWNy4H+2ajL1u3c7dX/eIKX9eFtUv981ssD5hPgASeOuZ35oshEAS4
av1a6RUOXUpVAq3ZWB23YnMj/Soxu+5WTao76vxWuMz4b+NEgrE3OmhvgxkaR7FBaXRV8k/b19qb
Dh+BAFHl7VW3r8rWhhzKekXiHbLKT12EZytCEqd+fkZRT8A36UKw5WgnPfKpXqQ69UMZ00R9Vzo1
p15X6pes4nXjnO5s4MScXqsU+r77gw07OI6ms1evGpWegpChAXAK5prgS8V3rJ4CE1AjQrpS2HET
MQA8umooD+SH3O/r2xRw7hx1hakJ/krdbybKN1xWhFQzm5goINiZBK9uCtjBcPzLFGMsFzi84npq
gtOw8ibS8laq6ZBldszvQWigoBhVAJGNb4AwkBdkqr0lUibdCEfLK0Zgu4YO5t+OkWJ6Ozq5vuDW
MWlmCudEs6MmJlv7xOsmzkIwVuRiO7g30whzoobW+R30Um7EpPuk6PGd4xwh5+XjBUtYe950r4xi
wDHnEskDIIlwH5l653/TFGstpBs2r3L3ZUQGtp0G3xDMdefWU1kRCmPD3CqPhOGHyLTr6gI8dwAu
Jpc/kewGFXewnneGpWzUusEOg2xiXSxEiFpWVDqEeLoF/8c7rnSm3K+vOATxB3S8kiAHvbckw79C
rONmgZg38XbVtCjdECEKLClvX2e+nrVyg4q85h6xlsAxiriYI3m6D+9NnX+uO5e4nNSPjZmL94Ta
AAsyEsetZmKoX/WPw7QcUvs46Pz2c4lHW/L/XKaqxRJ8EFrFNIFfAMLqgpDf3Xws28YO3OJbgfFc
tJKbzPv7XEQzIBhefSaq3TV1Kw42+8FLXRp214gspXcajWDYfgv06L5X60cI+OT8nMkvrVQgJpT9
POYrJyFeBabixILaFRYWdnHOPyFoYz3zzRgSE8dQF7aDj4BoKgs6D1LgYQppXaxC6YOvzEMX2Uvq
Jfpbs/vZv7kCkL+qX2WdsO6JGDNLpVNuePCh2E/kN4dubVqIplZia/syz7/b8je6K8B4r/3qOXKZ
qaX7167ulbuk+MgOigLyBLXuONYlgzrPi4ndgc9R24aR2zP/DfIfhqv4SxqBozSI9uovPe/6UhZM
Z+ZEokWBW0JFa8kFpxc0NdRhQ9/9xWxuYASzkjZ6y4WIoIV+BDsceZYVisqIDm8/+Bh2e96bzVqj
qWbaXUe8U8APzZMmIFhmDzGLcW3+gOZafgWhrW7n/AGVQ10/sxxegpUt3ehf7IBxrchdJaLYT/Xl
3k/KAMP2hFSJbFKekWHP/9kn4iqNwzffE3TmjF5dNdat6Gx6Z3ssmL1INvi3mDjN9trj54ooEqsV
Y6/pIqv/4P4u/XNHYZQnmvmnGorH1bvq0y/l8IUL1S7PBZXsBkW/YQBrhyrZe9RekhOIBDpz3nQ2
ESpU7PJ2jxrlRX4Ac9ZKluCfinw74PvgGM/P0P31iqtgQB7Rvri4hatC7fa6QVXJzI7wUH++ztQh
yBX/qQhgInu/lGXjl61BZ8A9n07jGThCYXTWQxEsnvUgFNYwRQkH7HXG9kqhZaCyz18OEHs0nIPZ
IIwliOORNVDSa1X8VUPBImEETJmlGg3X3l4FBCAtf+Nh+H0eSnQFikEDb1WB5RAy5UGWvrMSWfKm
4WWWHpYItPATF8hSpne1jIakEs01l93KhycONMIwyrosCFes18vDEvI0Kl9NuZb+8G4rlEyXaxE8
SIer6A0DURbMKzV/LAqMx4/VA3j8xJsRkftsfLJ8tyl23Rl6fCvMgVGFdSrnwWBdEub1vm9E+36I
oKx1R0dlgtLVGXsNzw1CVLczEoyYDAt2r6M6FTZc3MZyDdA0kcTJodfkUvvxQC5NPsxouq9Igrbw
sdBrnJrQr61Q5+XJJrwyDh+kwtT7U4uU/5onfb3US8TSNlBXnicf193FtiD1stSRzj8NzUEW6y7Z
1SKpO7iezvx9qyplvOdBlweejv+Mi/5Ol2EQa7uPcUwgrdzBcXk0wxGt3DHQZO5IG0KqRbSlWIkX
Zve/RAqNfyExzb6Zl0SRLJL4l273gn92WIxtb71F7ghyE+lV0RMvtUi/ftWDla3XzW6D0en6CyP5
e/It7EZelFA8HCSCFuWOxzn73IZFCZ+ax9X5ILcryYEuRkRy9u6F/w4MNuMgzF5E5URhPoGR+Jci
FagXeiXfbcEJQyfLenJOUjWCfcvpTy49Z8kKQCB02vGznJcuQuqVOyuI7MiCE5eJ1BrUSluNr5jq
r5VG+YSCKfYV9OAHcGLTOIL0H/B4rbNLn/ow3DUQApfkVvFOUckMZoZVOM9G4GJDnEaQsEapgEj+
mvg6v2072MrrAYeONuNsSN26YnyRK35J6fI36hZNdJX7Up2HzPVJGprx/K3PTZnk11rDYtgxdK+Z
SjgKklaNSH/P7H4YARTUwB8XTjMHhfK4t5pFVJAfqkh1rALv7NE1z40ENGU+l9rs1zfF95MEzA+H
VLoeFdw/cITPPNT5cI75lGzXjpR1Xv7mi/tiXQcqd3jB2F+xvc9DynbSSNY714tmyWPpxMehKXCo
0Hpilm8mUMwxTsw2qWXyo/v12A8YIpD5dow9Jm18MRAg40b8OOGLvMPF3aWq4eKkAXRd5fACxFaF
M4zptOSIpj0+yMZfFNIPYtJlSVKt/KEwf7emu01ZkaMtjjQeTv3gVN78VzM5wz5a+DXeUg1iQzcG
4rCiZ47ccVv0tG9ZBgTt0+N2Bu9R6QuVRzvz5wnPofluKUsbRASFy1T6hwynSQmQZUwGOQpjJlEt
RBzL+hGPlhh/S0IuWUChNwUNdOYfb2NVH7s1orNTQt4Zse3Wme0Aroy20dpnOISHIE9botqBUpGU
5ljQUp35vHmbGkTFu2i6RMYet+OU72MAt2g1spUJ0EDBI3G6AREHtPQ+QHevWeZ7PGFSI81K4ZJk
pw7Wov+mQGrLhnKiVhx14rhZu28hfuVd+jYaiJQZMqvikS5EPmmqdp5R1WrxaoIc1apxDDxVpP4i
KVqcEXLzgpyVstj9p+Wt3BBRZ04HM7DedmqI8kQZT9XgGkWu82LrT+sI6q8HtKWt2f3HHLPdspYc
PiDLB1dDU0kFcoVcuQo8TOcSEc8Bg1x3Lb54cuPArpC7RU9hhb4dCnWE3h6ualA7kcnE6MnQQ+vW
vZwNKwvUzO92Ps8USekMaa88PQWreOTrnmbXRTSme9mIJ2lxJGdUM8DxJREUg3rd6A4GojN3igIN
Velsp5GmqP59mPEX0orfyYFsqlkcpfiE9cyu4ryG9BGnAmJVFgdviuxjMcp+lAhlsfTbJgjrHFWm
iIBxD93m3Y91FDF0l7HAaoHYPDUc3HC74IHaaRQeUByVEb7AJxCjIyh2ch3zTzq48SgDkhicEPoB
GFlHXk8nSL0R+lVaDdxcPlFiLD9iX4J4ctQOS0yQJm0A/4nJvua3IJsZqB70ap+DA4LFUg8+4qhA
V33mUk9r+M/w7JVRs/T61bxcC9b1guf3uCmU33xiZJLEN+n+6JxeRP6nWJxE6wAKiVy7mL3lOUru
u/IEcfcxjOwwO7eI3fs9+3hbJMfJmny5HFeIPyGsfBwgsRGm9RZGSj7pGo11cga4Z5jzfQ9A7I5a
3eW87FFAfU3a+SQkXin9MqbEQXjXl0vVnNM8VTmDqA/1TOJmQeTe1W+SxhtmF/mj3fvXHhLTZcEg
1BuRFgCcWThSwl26HqDCKTWylV0tvQJUMl4GY2PtejRZu0OJmk1UytZrc1kNpxJ/xvzHndt4vDI2
094KK1rZJ2gS1/MgRUsJu5I8xqmaqYx/ybYBWrpfY6jZGevc61g1Tk2go2vIcWZIlBtS6rOxnyNJ
kckEKWL4TBgNR94Mhas4kKunbsxg6upiQOCVQ1lApq5Nv8QRK7KyKB7qPl2vNT90JbzKmr4PbJy7
JzP41OwsXmvjXlFcDZnmNbPpTVEvS9QjFHH/WHkbc2V+EUnkc/4ZhuR9Bodx129OFgCQJ2IS0dhL
Nh0J517j5mmOflxxgyMB8BY2ApivAfS5pBbrTWMkYpelnr0/7BB9BazRh0duMzqWhwe9c6ylN/VI
7kMCFGvAaSesGN2XCs1li+of8o4jTTEgZPw6LxIh5HIV6ABLEf6LBy7fFl9JEBy9nR5rtu4kg0n+
Yon8k6nxN1t36hdrzEOMH84zUcJLwspQ2rJ+0cCGMTyHth1W4BksnYEMuCYkcJYyJsqWPZhZazFA
pwO/NZ8886u9hGnJd95KO9uBLaMT5VoK6O+2UNFKu7XH1WuBkFyJzCHO9p/6UHBjYrJHG71I3ZwG
M2OpeEnctR6Dg15TroG6wLo7ZstbUe05+Y/zz6RiWInclK25vba3aXrSI4kOfRoattj4h+D5z0hX
xZHjOpAiZF9BXFUMkSrk5F6ei/0bXQ1qllfMAsQKkxHQnJ2KeBn3BiNLKQD7bpA9Tw963M9ftn7C
EFJMG2rBpLG/MS5yHn2eYw65uFnKqVgEhNwKniTLwFE1i6Utfay93U9w8JfxouGexBTEb9FjfrcD
i0zEK2monfppoPLshFthKwmDIVZgpRUDvMjUyHNG9pyvkhdMu4+w5bG1I82wdwbpZIMpeRB6HdcP
j0zLQIpaWoAtxDEcrUK+RDQYxJRJ9aZQJxMviTGZUxg0xTAhxEG4xCcajZTl65jlwsVs6innBNWy
B27dweGfdakWqsh7Jf8e60QjAbwWrKkD80t/eRAIFLC3+5XHFeYubaZNhI4K/QoSkSka+LHFO+FE
B2BWdYGVvc/+25gSGGoxIOfSGouHakd8FVoyr1Vq3qTLKbZ3PrlzqqIl91NpMJI7J435+9shkkgo
g226nsV4LBHZL8+x0fq6ihQLeHZJ5QKNK+UO0pfTaZRMHmFUqM0KwbIagmisKI+qKaxlDyrCy9GC
phJP77EfqwPiZ6ErG0EeOAeUvD5/SvABv57/f+zoq3mAHhRaqYx4t8DeHna+MffqRANhThcOKyP/
CCMOuepnRj92wnzKoCnhMorCneSC43o6IQrE3vAu2y9GVpb/c61XrAoCNq3RrjPUmANEWFlKlO9W
o2ItS9XEnhPAGG7Rf/kutisewQ9FtQWVydm5zW4t0lxTfeBAf66hTbWp9Y8iLO4bXJgoweYwnN5H
WS2kZoqq0RnQbaHc2licY4jfcdRYqEal3U9xwzpPKwKZDKJZYZNjDPTE5liGl9DLUlRR5pczY/ZG
BbQsHZlVwlVIzy2AfXZJwtQeSQ7mfpZr2qADiKql3caQlIh+hJrwv/ezohb8ViIy8+IzxU7m+/i8
NqIsjUjDXU372YFfDC8vSeoCeERXrLSsCaZXTfc7YN1i7tkt+efZ35L6ewPtXHWrVbo9vxrt5xyC
ZxfVsM1WWwJlp4wNqaK3/rAQg3a0bCV4TJpVKaElhUCpq1PL+0J1AoZEsAScuV5SXOmBCFHAsihB
UqdlAX6Wdx7/H8cIQiix9207HWF1LeLixszj1unm6E+I7fLPf7VL97dHqlTwLWv7n5Kpa8MYeoZ5
UJhBBdD5wH4qhcyuFxw3XvZNZEEAk9TZlgcP3BaiPtdOGFf/o3Zq04NRONa3rnVUlbXYqFBNlkOR
s0rrbnnEHJPbW7h0QZn9q6Mc1jJs7BktAQfR5nCH7A91o8eRgawL2o6yze0eDGk5EUHW5xJ43kLG
AXtdQqZkgrgpKW5egFQKV37WWTPOCMGaAzoPoW49vuUMyEJB8XJu9sjnsYfX79D8f2b+uOzQWW64
TPZU+rS7b8NbjbjlyKPAvEgcDmNMuK+VCXg2K0LgWAM9/Z3jkrcxDeCDs89TdoMD0Vqld8h1ThAm
s4dJG4Ctyt78idL8vN5gSF1w3fEAYF64hwA03BhLIL4+aWBOWJWpi6UiD57fElgwy5zbj/MvYzZB
QM/JoVyDpVuPuD+oV7tC7NzNUQMeXcsiog/+YI+G7vGkKzSeyBBIT5UKahV66UDVwCxnBmMdEZfV
e/uuB2olnA0zNgB5e/tFuzGxffD6/9NQzmGCH0BW1/lPELfDU/0GPcCDVuKcrb/yp8vW1t8YS3/U
swnqFwBw5vE+MV7Dfz3GO4pXoAu6yzJlFhkKXrO7SAWJwXZ2k8NQn9QcUNfbhAjz/6FtXLKcfA6K
M1sTLUJYIL7N8jMQm3Pr8Q5NA+GwH65+Bg0vD37bruL4exv1Rx5lHWbFS8s3zsFtjgZexUafWGzt
jMmM+38MBxo+narhYUeylr6AcRthiwQNVgAHQfdB17OBasuAVTqE7SuGS+uARhCzcWl2SIpQcjm/
bXKoZwBM0/tWHqgiJdPAupZimRfzwaYXyv5D7jhCnLaGYW0TIZCHC0V/NCgx8rtMmg337+8zG2q3
BjqFy3HEj8UF3nGNHeUm/DNzeoNI3VXPABSlKVguDAwsyeYIJDNNqPLQ1cKjx3zuz6ClxwJt735a
aptIkc3jS5ggryoeoVF0rb46WjFGVzD9oGOezEWu8DR6nZNHzTdzXDxxKlpZrC8k/GVz2w2vEVcT
m30g5m8KwUO/vYF+Ik/ipTqX8zSkqWtvwtD7cea3DGEAew8iK4d6nsLAbyn9j/YCro5feQMa0KiG
o0LEzIJfy/5GR3ihYb27idZm8bZ+zDkiRZR7fO77Q/zWz6eTbP0r0dFSXvuZvdg7uy9xnqRdWq06
ikPVSvOx8Iv3q8q0q9k4ZVVDLa9/cm+9DMInnU/rhKZiOWgX7ht92AEpGb5EVtLwpdXNGnFyuPrS
aV5rs+CtKYHGcOuV4kLaeWwoIGsmFQb+gfLxhcN9bxLU1MaYOB2BNg3VK63A6sqhvo0EZQXPM008
Oucy2+hLi5Lz7u9CWAiYfl2938hMUeKNQ4mGU5pwxXDocNRWDgcra+D2DOTF/vWSRHBwxenZjNTg
HZEybaRA1jlKioD6JCw70XZ2i9tbRugKgItYRFMoRekN8b4oK1cheh4ZapHrxS3jrAlXdRVOMhgh
pw8m1ld3XzMwbSknAWkNyVIRVFbt/taebUb8CBhbt0qHWFOQPPbKuqNYkYQmrG0ABnA7KuPsJfv1
36mA0refz9GSkbM1toD1B/ZIv2313cgi4vzm6YElsZ6ucvxfJ/PMsjUlX/lzP50bW/s861s7/zhj
IiBTjcnrg/9UF7FisPZpoxWE7Mwrc6BN+MuNoxxC0Fqx1awEBcTqdHgE9lzkAWD4q2/77ah3TE2/
dOb8knjmd7kboOzA9tHO2VXUBDXvF3mouzUa+D5PKWpNC6+NL3Iocvgct9A5c0tIPg60geO7hE1W
oislt866yW6qEf7SIfxKnchBhN4cBNienxRp/1PIR7/iZmAI3newl20t8ZC2c1etwQqtIi98DC+O
GdzUT9QhZirqPtBSXoFaKojv+C5x2D3/fPgAv1zW2UU+vjcyg9LE7qxNf7ojOUkulD8VkTxM19G7
vP1xa2KrVoKmQKRHg2hE64sqdbUKyBRdiuIqqKQGuSFJB4ph4/yL3SYmnjcGoxg9mgt3zBy9zBbO
y8WcOxMRSjHal0COLdBfP4GX01SkykAiB20Y6zOOobbf22mQRH/2L0GzsZUemWgLVf4i6+P+5iF9
L3y2akVoniUmN/v+1E7XAkju9lLmyLNDmF3NsXV+d6fvKxcdtcg6dNM2/tXkPVZLPv9xYu9SVqZz
26zIw0T+3PSMw8FkoGeyQROx8cfBIyR9JZf5PhGINBGxPTqVm28ADTXrV84E9NfLFFTW3r7SvD8u
NM+hNXe43AYXALTfvBsQ87HmycRIyBYCkdChWEEUF54eXeDWurdCKspoig1kiDrd51rgXLzKEBdX
pibVd0O388yM3oZkxuIl7fdm1Ksh93jaZHFceoN7MMI9nW/CGbTc4SuHiTYjD/0BQQlFM4KNTWnT
K1a+hiYSaAMdYKpaDEH/cwlTrYtDxky5CpE+1CxCUlErFb3bD6n2mbQ267qM94fOvWwybqphR9Du
aQnjrZ+WKWWqMYV6CYz74/naZJhBPUhpT6fv1VgaPfaoJ06WZ9PTJRtijRZPqvEabB0IJuSzMXZM
rF7Yo+IliD6+RqqoHeBOjLss6xMV1N8U1uDyHy5Avtxf/rBI4CB5E8naEoN9qYAl4T7mQqEknYTU
3RE75JmFfMy2wkl61v9W6z2l0xPE9SzZrPKDcJ3NX8PXlPOnRNvnKbf8xDDrhMmRt/oNODg/lYi0
49D44bQxmHFBeQgW5gPqbhdyanw2KbH/9ilvt0oPN+RCRyMpRVW4wSzjXsKhCJN6446P7+3UpOFa
sJentPVOtzh6dkPXAS5OPxD5ABEGFLdt3yiIbVQ/ERqOjhhQ3ooMnPsZAH7r5Fzwsdm63ePUEWwK
S85DUrcoZg2TPq/AbRCer5ZqdkLJsGw/t/XAC86HwrQ5ZsB1yOj4SxsaciJ5M1nHQroMmH0xT9cE
+b5MtK0JG8z5PCX0lbB64m/HLgUbh1snlidyOULm21XjT/Zdd1U+7mD9Za1FzE1wG7ZrPgII+wfM
hNhFfjaWx6/Pq8ZVWA+5AVSTo5XVT7iM3dwg9YhRWJMXaFHXXY70imtFtdnnPl4If8MrMcSm/9n4
H4F5IdRpTNVf82A9Xi3umNnIXMzg0sqOJz2nm7Vjvl6zSr75Al+Yc+Q/jmcKLzsYDzh6vrDEPs3q
KFmq0arWOW1xSOxvAZWZCusi1FrW+fIhrCz6fsPd3sNk4tGW5dWgWkGxVFhUup9mBczgOy0A7ZyS
iwAhBkwM3G3FSThUiz28PPMOA0eWdrzN+5AMUL+xzkdgeReMmDEusCOElGsUEBK14mOrCeIU/yJT
XDOmvpWnON8uNV7lCOCrmk2WWxqRHK0qkVBiouLhJa0V8cjkO7hfHW9wPYSjZzhWxx4bb3DUv1fl
9kNYFu6rwZ6ixMPCytZH9uVWnf60JTGyfTh0ZST525dw9VrFpuHbec83HQmDGWul91Sez7DV83mr
AaYjitcXGV8ZaPZTYPTLnspAFkYGv2sKG5ucUbR9b6sB4qDwFXPy2KfcQDBu1gc4ph58Z+ntmY6W
0TR20paz4yC+tYKrvKZPCfmWE56yqq+FrNVYHI+LrQK20t47IVBmOvwjA48KhS46vE3pAbGw27N/
vizRu7YnYp5U/YjpkjANxfy6XKaTy7l/3qRtDZfM/UBnCVyKHoIG9D/0+rypK3l6QGrXfjZs0FTR
zPIKvkGFR6xSoIhMIM66MZVWU+vqJUwriM4g73D/kPqJU7iiMcPuvhqpicfu1z2dAknNxO4Zh+Gx
EKQ7VOFFcQvuhjxr3PFaFVPEVPS7h4dUIFdZgBqXRKU6dFbrZkfV3Kp5lBCzFcb4rtAYMnpfFanb
O+cMPO5WyYUOfK4/oxNyLEvh4nu5nzDvkN8GE7ptT7nFsHuA++fUwc5yu+Tv5Q6GkeW3KkVA1PAO
KyhlZwlCst6l9ZSYvMayFluL5YRI7wZpr1925j3fOrZshpWdESaaU7sp2+Nqe4EcZK5OtaQmfh09
EYD9nKGMGoIM2+JxYQ+0BtyNKWISEoRhA0RubC/iP0QXYcRzHV/0uGMyFowHI1cKd7gW9jBkN5yW
iZdakDZTqhDxhyFEBUVE2k2DaOdC6BEsvbmoQ7ipZyPWs/ZiuRK1fiihOOS50J2ij8BRDgcVYyWL
MLONS0IcfbCfd/8Td5atVsmc7BSDXEIpS2H6S5o9FcIFm+2UURkotpwR20qGZQqUnorbZQX3QIqS
ERLfbMBA5yE2N7iZ3ks1t18s8WDmm08KViFH91jHQRMbDFLAL2+pCaMVtnKv8Z3/zg7NCfTIBI6S
eMkCRRQS8Zu1tKHLRbiBK9XsQXMqql+Hnh1l6ej7q5eOeeTReQU/fZbbQIN/qXLlw2I3ClQbJBdv
q/RtBaooeMsyExiZPy0YLYkI+xbMA7dErhzReuwlCpPLHYV8h8c6/jkxgFUMQ7Y8fF2twCuSA+wQ
xfhvJgEy12Vus+eETew4zWrF+EucHqXCgzW2wuQe7v3nWMFgLTtNsa7jDKynAZ67FbB/qXWUVsfo
7KRFZsfw2dlX3FDoV25rmgmQKUbxh6uNR7QEd2URfrv4JFEisiui/fW3xcgkpuHlNSGIm5spaLjr
QTZ7NXaoKoVoaJdrnr5plWVFsZGmk3glm9pDP6PzsUPLJq/fIz3fKzwOhPk5oy7z3fitBC9u9K9d
IGZhDlHjZm1qqLt5G4/iJhuZ36UhNWGqzGOcKzETAFl3503YUL01rmwWeA/Ozqj8bWeUxnIyWxFV
/KZGWYMn+LwOuFIEmIegWE9YaSGLzhHAtBmVlq8fIby9jjOKVHNYKxGSqApwQJcP+Fi5LxttruhZ
GJnkGo40IHN93ZCL7eqEG9LfG9dttadSmzcT6DDearBUR7TzmhuFs2vnherp+UsODDZduxC28fXl
Aed/TFgN2+kD1jAVPix12Gx5Mcytw7UYzb9VaLhYsaVCo2l6MkjsfCBLvQJCmVtG9UbTA2v42L0S
gxnIV1K99oSBAm9w1wXD53kYxRnHHAiAoaVCWCiwWhcMRAXLVvm5fgrEBWaCz9pSR4ofpUKm8Btm
T8OTnnUXUSI6GYRYi+pS4J8S6a7Q0jC3th1aCWtI8azczc1YMZ8k6Gedk9hJHI9pjGYoPfgHdvaS
KhOjJwetqPSytOcQuBkCvsP/g7GXzwSFAIRcWEmf54JVB+vzDkCsIQkP4EeHY6JSG74ShOn2FGJg
YbTNmZtiE09lPIVagdXLSCyfHN1+aOZ/3WfMmoovvKHZ+icOcjff+LpDjZfEMKhYQNX7J39DtGaE
7aMXWJBjY0YCvFy49jz2ssQtzgT4l596ih8LND3N+QXMvS6D786PvholViTwrmav72B7znfysuL1
BO7GC354KALRX1uHQgkopjZwYT82z61cXodF8M5e+zqty7V+uGSKWIuaNh1Mh/PmJ57dC6BEgcnH
Xf4UArlrFQmogl7VJFyb9NJJ1KfPd6fMsyQr4L62KULRFhvDwqek0RsAYTABr79ioF+zD8w/ktnT
EPE4obuqrQ8+D+l+mzjvJIeGN/ukCCee0OqlJYVWx5hd/xDvgjJ/lmrhw8B+oj799QtpIhuu1M5I
oBy/ZjJ8jghSIZKrZx6w4GvxRkeVd/djJc4fhcQFbUIfBEnLkSToIpEmk0u+CPrffVjCAdFM1Wba
4sMOb8t/6RiqxeU2320+hUKW8ge/xEYH5r+SV+NNkoFaU7FaDuOlSwVBVKIR2YZ4H3LLYX7wDOYC
apaiTxvy2pcZSBtRTOa6F7EnEWhySToIApBLV1KILqnozNf0WodFNpMtouZhEUcj6MN16X2u/c+9
l+YQZENokezHFPgxv9Ti+jecCOePQHm8/nUTOCboBeLIyejfeaLp4wvUBZZviHbLAPrFhzC56YxG
eTURfsP3NoooYRf0p5L7TL7BQu3dLnY52TXRidgkmnxSvjBWKUvn7oUMlF3/l7Nhj+z4p4BqFGTm
1qx9x1oHBdNc2L5sUV9WmDjkJUrkSrQ48WqbI+bTDbGZJZ59J1NA5QPlHCZ1tuO5ErEcn7nySA2r
BeBX+CkVOmqiEinLXPRS57Jl6ey4qeJd2pBW+eC6/G3ubK6gujYCokCDaLWDfX8b7ZszMeZykVbD
Tq5GBwgELhbHWmI1J1AEeX8o76sJ/kFLxKPDIKIAQayDnnfdxfN08U44G2+fR6KKkSwGH1SWKPkd
qAsQo5vcQKTUtgyQpfSkLGbvJiH1EoHop581DC+1xVKmRVNJ9GTxIgsbwx+5JxrdrhlD1wb2lHr2
aNTRu8O64l2mXTaUc0Jt18worb5G8ODztXSuP3JYuIu+89jbsNNWBJMEi4nPjFGcAgqHJzbxZ3xN
6GTf8mwSAlXgJd2IV9o0ayph15KHTber1q6MFmIRXm/wjkFTqUBTo5xiK+HrQFqvftF4qO4qx14V
fRNNiDBXFCnnJrnF+GqenZgwK7uzoXxJEKipPq5601xW+yCw0S3HGokdqwmB+MReRa3AA/iUVQQS
urqTKaMi7rPccohcv0Y9GIxJyVfsjJaZXNChbjzcaH+OOjpVEAQcOBO65iU1pHcUDhckkj/7/+Gp
cEGMZZCl3dzNBnaoX2cDHdOyRW86jyiaZRF7zhEZncK08HpywVi89dg5Qa6swMD3kYMcmxlYlgUh
g2AASZc1XazZIPHGGT+7LTmkK6PLaVr3TI3lRu0Zww2uYq2LvNwAojlvbPcOdeFQgSvL+9Z2Ln3p
XI9cQni1pHat8JpFizTcPwI0CdNUCwkMTiSudX2c26UGDgsfCOxVrpZyseJLET4dvF8K3W54sShG
ghErzX0ErgiajfaLO4qNZOarJ74x+m/dy6VQ/dTPezXF1Tc1NyX5m8jcMggRDRLqfh+JsDihYCDj
XD2oWyDFqVPJNelSvQAD61+1o/sq+opAIy3NdNZUNAX/HN42CitGoY5oCeLegIwelB9K9grHysBO
rML6XKbmtGqQ0yp829XZoLXdAnXggZshvD0F/fSflECQXN5kkM2iBsnuhUYxye1TIqQLlIudMCOC
rJ8VGCkE25jgNAXucZXjN94F3d3WcNCo/WUWVNfYvlZRKlmgXoUYyfe0t+elQbui4ZXintvRbGjK
oE5pBg63Bpj9CYv1OjUjTWIOsqg2GcpayMqiKza9NytQFH6FzTNH/WUwbrUVJAGaj3hWL1R9iezQ
BecVr9G5I11gUaVU10yfOrFWEDqHzFUnBSZSqPqjyyvyBNMUJ/eJtt6yeRTHOTvOicHjO+5qwyVO
W6H1XP1R3JYUKRtmltdhTcru2pJU4D4+CUinfB63/oYZ2fHUJjISMR6Upi71GOipgmfK3efJ2LSt
l5hkRB0lqZzmX0mblPle8gEh9P5abx+SH9IcvF1YYXS5e2/wybxtKIVA0MIak0PlvFA1ZiX0RKPu
+PgPTwY9E/OfSY8FG3ZhdICm/0h8AwIs+UtUTe0ZDXtidoHPoSvh/d9tNbg1MWO0psuFP9ES+j7e
Mxeroumk52vAa2GNAVtA4IWnPe0205Z/DSOwg7bcNaIo0AmFhNZN76K4f+RRPtRbTxpEj8Z2qdaB
ktKuvthPwCgikCjhXW8yXBAb9OhrSfgxVcd0Xog7Lfbir7IQyW7oI/BcRbsdTHdGUpSchScnNqaa
sbM6HBrr2Pu9ZV8L4YmansiM7FyHwUhmYQUGz4AkqkvpCfhuuK8qI8VWrmDPzHWMnoibCf/2TS3Z
M5otvF2+6WeKK1xQ66Sya6FidUDsN3x4yBz0O5ZXj+o0d7rUWR/BeAz3f5lS8Vo4qxxfPxcYZFBk
5yPl7E3+z3mqxjf+gAgcxNj+EumVEioR9fOWBH402/UjxgUIZZ6K3gZh6MPprR+qaC/zP8HZQPM5
rpvv6K+yRt5uZkjXKaFaRU5m8o/0Qnkj82bejgDSyGj0b07d2JiYwGV7EGH0lMGrSLw2j43zAI3G
AXWjHHTNV4hmwQyW8Jes7ZfvK0wZHcvgWGFH/sGYKdXlxr+PVM/JsJbohfeF9efnY9JblRn+Izlo
p4tFm9FhR3cmKJ8FEIHJ9va4pxxER12rYm9it6rsEjQWozpv8xdgD3Lm9NSIyl5GK6qXlt2PUWC/
mDgbyPr1iTx8wuJCcySxmKvcNp7xLg73XOix+5p3T2npJBIBMPHLkfiFQ5/lywnox/PYCS0SOmqy
6plUlmk5FZO8n5LSwck3+vANo59l7wwIqbI0sdYB2mkGT6rtj3aFqEyQ7g+qG1DwUncg320+2bM9
rFiTmVGIfuLn5qpMNmOUMFD5dHrB3oglBZz0DNl3uoCEfXIhaVtDYQillEjMI6jeTgB4FJlTrIgZ
REEVfRirxp60xVVdf+uV2SZwoBcvbtPOSNAFZePfryL46QxptcszISIy9PEGc0glHdto9LshYJbe
htyi/qCvQ6Hon/DL3GjtF1l99ND8N7mTbD+wohXOGoGGF5eqGhUP0QUAe8R3bU2jt1S57RjyhgoM
Z5ZqXhfxPjiGSKpZv7Y9lP4sUawex+O/fvm1aCuhCvoDmndeU9e25oGVrwTPTbsoiXHWrksLpvoD
FoUCVTEKWiAu+Svyh4aeSzYolbO9FF23f/bs82ftkkow0AQk+ddCeSkCSDGSRD+TVFcx4Qv/2WFi
iE1JnSBcLdkJSbt6h4IxLkdroshWX7G5gXtSsvUtzRqrMjIs60l/ooemxmmhrTTe1f9KNUhNohig
dmeNfsNEKvZYPXAOP/GWJlxsHjY8yzA4g5A9qBEAK17knBxswB8/KfhdmOgWJr7cemavakO5MyyM
FB62e1rt/kbzTtegHTqK3KR1SLXgHoMBFitibcKdIVeXDC0ygu0FfWvuPlsg5hWlX3dXi1Q/G1QN
idJD5FYuVPsd8IRKpUDzCcwIyOPcLsWuMKPpKbR043JsU3kAQx1R50lElCAsZyZh0DOYcwaKYlRa
5SIzeR6NCwI1NQyKfFqCliqBnDTy+w+F/sWF5zBd/o9PicQBY1OFk2/8OxO7vyORBbspTDSHFTJH
bW2Il8htkifvjRYub9UnbPqB0g/0najOPUkTP7D1zQzlQWAwq8qo/tZpFCnKm/Bte4vqr0YS8aSd
Yl12HyE89akzOzMWt2WYmwehbAFFy2ZU4Ym6LJCwgmvSIZlJZPUDt8Y3psR0C9YBm6lt4SZLOxqQ
UFuZrCmLaisbKdYHJ/GPQHtkJvXWvfOvJI8kLnu4JGAlf5PPFUMJdRhf4EJSI5eo1NGel6vnGtHZ
VpR4z5Lpp1q73pc+2ByczJMAsDE66XrW7kIzUsAMm7US8O/ZIR/K3KocbYMdyH1o6Cz5XHWQxYKY
UhqtX5yCQzYdAMo4EFMSXkwl1pOnjGtuUL83wPea30zazUoU3qjgFCvMS0qb/HIUBg4iw3u5WHkE
Frbg99dD/sFMhDTZ5JZX5k3Tx5EzFGyFxTIC+eC0cb4lHzz2VrcjIGPSWd+z8y98Gyc7ZXziiP9K
cs7OD/AB8fZ0VaHiI10OMwCmGMngd691Nvv06+hRzYhCdf3uM2IlgJzHX+0/5ToXJNlK88q8EfFj
I+iVFvoynhi3Dpf3iKAXB7kMZ0BsJ+hGib1jUJkJOY3f8UkWba19OC8qeRub9XDIGKJKXkfuOrXa
N7ioJE7HLvs3KwR3eyeESHEAHTNtLTQjeOXpM0lOYzFClMsI2l74SdDJ/IXDXo/jnwpp6nM3WGoh
XPc0eHzkpMghLapqtEu6xM26YixCtidVCWe3qwtkXkrPvNmH55MHOwKKmf2RhqtPljnPiu/Fym3F
Nv64Jv3e7LNSaQZho6Qucv4VS3/ev3BQQT8WmU9EZdGKOra0b2IZi5Pgoapzl2a/Fv6c9yTgtRxA
J9GxTipojCz9U95SZyFdxTTBwFq45LptUngNQETYNohi5nbci2kfzScpNtcLMZEUj08lYfmN6DWY
JURw2LvvI+iMlmiVsFfMdaNRlgbI3BdGkVnjAIzGlaYsQaZwjgWAv7BIhDiS758fV67bkbBjWjo+
TkNsf7m0PHo6XtGT6RxV1uD8eiLJhhbBN3XkMeJaJeIqgsGpwFfX0LzV0PhrDlZAvaB9nFT2RKvS
A7TrS2FeXAGq49/Ro0OkkenPFHhhf4OA4YY5S5OsLNRYaYoIrAit4cEi98jvLCmBT4VUf1+MFggs
1KIbJ4F/fmKknQH35LWMjWqNa5ZiboAYI7zmpvc954u/JntTgB33b3aykJHyCM0VMftT1fYmDPbo
MRjqsdweIfJCsi5P+/DvacS1ELQN7GSihzYMx0JZnGNEzADndvy5+XudvYy/eUrMFXJPV9OczD+Y
LpvXkogtT50EYzP+nety9ga6nbF1Yw5aqW6cuAEV8mvdGfg2GBOYQr4XogCfV9HJaWxKOW1rHIEX
2FzwmINbXuCo1Q3z4xlh9XDnT0GbCyvoPX/hQk2aCZfmZukOMsUFbfG0EB9+Bw96SfPgSO0V5JqX
qrNN8PlJtR331Av0A3EIMO4Y6Uhw5vGmA/rTlw3hXBAz4Nw0GjtKs+Iq57d/qCkU56S4m7kaoYAO
glIGc+dbbhCTYLa1p6XRqKJdqtZH9VCrpmIhN/J0IhaKt09OG25JMRKYXDLug5qkPNWaQ5e5F1El
kg2+beEwsNcJu+ifoGZZlvUcfD8OqLoPNIyzM98e5kXedB7XiyCyEwBbuIyMD2l+xQQukO4FMr9+
pWzqNjJDD1tyNj5wGMNgwcgKCIVB4FERENSw9F0HNEXOaOnXzOIOgVjBnxEyYTEzy6CqUzDzW9Df
H97Bl47Hzh67DZg4WSI7ZLWcNC+k6f9dYusbysy5wHKekjENQ7pW1jXr/flJzYH37gAy43vfb0LQ
QWv0TbmBp50/wDSsuTatUc5b8idPhjKQWrDLIlGwWwgdc20+h/BGFlCWXBeptNW6E7y+JdJKHt/R
6IDdTurPlTuRdSYrhWwkekubyKPkw3/hGuZyzxp/pIr39BB9OVo1S2ljF1zGRhMjfnpLt9+DoMK8
ZaS0klaPf12wUHtbIWTly2rdckmVejffaOx4YHRPoC0s5Bfx53LuVmFuoCF/06AVakPR1twAEGbz
4/crowAd6e6nlMmMyh4JEUwydSwXv32l48focZOWQNWynC5BW9fQlDapGEUcWSvIlf8xKnEUguYD
3qVaYIqC4kPAdJk0Eat1gXZmwgL5h2cuEODvmG7tz3ei27VDhRySamxxkDNdSo1tVkrD1ui4/dKQ
veQ0XaAcVp195TI3/ZmJgjs0dFL8RDJWQK1k3dWSIf4uDQQLU/qJ9ERVUmltkLJnoSJMZT6mwAuP
ZxicmLer9otMLRZQ4qtg02ULLN+Pa74vaCmf4QmRfFOktQWOtS9zPhhi5pLPr7FXukzUEuts9Zub
wisAFIqYC8dFmL7NciIiVOXFoH9y5BSR4sjON5Wg3ltFJmWc2HPxgDkVr6quf+taUx+NsFkpiwLJ
Eu5pZCkK2wgs23WGC1ainpd6a1suFfHpvh/L/XQpmJDcePmYdewYU4FktEHcBi0y2hiGhA0qkaC7
9pqTdabIcWaadFo+oQm/79tyOnAmJsuiI3IwW2KL9FSJ9c+ykMPGiJWxUHyy32msL7TOcmotRIR0
op5ssaCgwp11VvVIqTzJPzEqWOLz3OAjnSNgdHxy6SV6V3s9hhWcbVD5OfNviLVTI0jMUIRR/4kO
U0f97T+tZ+UmSRdnrR50BunI3cWqlxZJGikZNLpuH9xXj7ZTUsFnfeAJSYqrOhun5XBxLhAiU5Vc
LbKye5cbL6ZZDmwBl6oC1NPWZZHKs3hvMwY+7njI6g3WLy39k0yYZfTjxqzDlGKJNCDrK+jrYnQb
/E+tFn+b7zs64nysMAsDkCkAvJsonvyEXZTqDLB1BAwX6FhOaM35V9YE1cWHBfCljFXDhjDdTFaG
4O7TWzk2h7rOrSaOyda2JHZ2bSBXbKr7MF1skS2D1cpKPYuLg4PbCgKhru4BPUCZwXLRxF3hwi/3
W3m1eTUUiFx3vtVPMWw7+J6MvTZpw0ijuhcgawAKI3T9oo/26BtT0nmwjgmnsR8FF5rcuoApQKlv
ahtgjmmJqxU4ooh2NLngcRoXBddvIwmjiols/VPbxXS5fL5qnjh/lHTmg1DsSkscZOA7G0knNvsp
8JEKru1vX3Oar2bB6YrA0c1uZpX4wM3C6yr4jkRU1kS5zAd4MUPoTMghS83/9oC96grUwE+vgM5i
V5lUfOZ08e78OWgGLN6hqgqr4RJTkIpITZt1IKH0+8jPtnEaZ4R1jSSFmtcSrF/shukj4IFJ0H7K
h2X/UHV+yp1mMRpaNw3FaGAg+HfICtxp/nTPt/rJJCmWq5oURNBg9yzKE7jtm43RmhSDHKB4BrdJ
BnTHL+9EHjY50bkqcdM6AKBgNm8FxNJjJERUT51SL/UZHLJeERzxKLYOuGv5f56Dz8uKLG1kJ3Dx
4cdTe/r4Tn81YgfePPNRfdWOkcuCGXnIgrQkWtEmq6QzyBwdjk3i4OB4Yq7tyIXQT8CWB5Ac79UP
5wuyPclUVnxAffKjZEd2jqsuKeWfmQavhUijaXx57bN7SClUt8Oy1+DpeH3tkh3D5iAsv5HzgyxE
GRgAlWRD075KRbpiZBmisRxYvVo4RAAkEuic4C2qA//MeAhbxu1t0LQE9qCPW9HGemIxG3hqzKMn
Ua8apn9XdghAJRzIyD7tgitFlecDNvC+qO5iH0C5twcF74e757oXxUSu3tKoJ6OEhom/U2P9C5j8
KOWM//U2giDwsIiyGo8ATqC28itF44YOLg7AdY3QlJqdZGxhxS04Sxz/JQPv1FHqLqmV1JKK/NgD
Rs6ECPM7LodejvkP51X/Uvfk4Oz5a5b0RSl03zLsBpEKK7jSVN9gRRaW0u8CS5Q36JW7eYVdTp2L
Nqy7E+TqJNpjq8Ql0ZeQlmIOBaybK+ZNRfG0P9vCjbAQYc54JSLR6lESihNf6QVVcriDK2Yid6WO
3uE8omgkxekXzr9tIhwFqmGbDeNkmLc8zYchTGB0Wkeekv6JbA8fH6Lg8IZJWZ2YpJdm9QSX9bTx
jKpo036TCWuUFBaYZ7FdWp7vAwbLFgJZablZlRME14xyECB7Vx7e/BnennQw0eHTG5sRsHjZYlkD
4D5YZ9Fvxt7g9/SwxlEGx5hqyhInXbdKGEED5Ov89zGtt++iQ5ELXNK6Chx0kiUJGZKv1ErmHOUd
0wpDNQjVy5iDWu6/wRdzXGtOUjqaufV3OsAzs8UV7D+6WwmLxZfssBlLjLb/qLH8Tc1v/uBQqSAa
g9vEtBBxXF2Gfze0NQA10caAzdlOD+7vNQhbXPZ5VWjM3XM0VUs7OwzkP4RPzwNsTVOeS6Z1Uamg
IPYehMwOsYpxkuk8iHq4xHrmUpoBrShlUd/lf9gh2edGmQUqOL77A77fkVhPGkp5ADJtRvsR1WB4
PWuj5h2mGqibts/O5o8xIYBxIzc7RHVeNsRMPsOuF99Bf27+IsONmhlgLj5bkiu2XWUR5plqLVzS
ppoDswlSWlLhHLYPYLal9Sa223mHRem46H0zPtvw0bKKAuL6DwnliE01Rfvv/klX6NJ+KGgiZZ5E
C3CZ2gwMupAPZKoEXknEesen9OltiHEp7UrQSz25SqTFf1TGtVfJfIeQ9YUoiGLTwxasAAG4/oXV
p2/n33TS4+5euBvWzXsUfo853kwr5BUklBLHoh41xJI/YPKTburobFsC8nstPHtCK3tPUbT9xJkE
Zxo6WpjsFnfA2W/AaWMVXF6OhlXAW9IAhQaGCA+UDb/WYjj2d03Pf8Yjd99HT5nQtdi/VI1dH16L
WsvJiCGERzq3LLT0PKR4Wk1VsgmrEWjBzYTue8gc49eTY34Yd/D2y9skpy2/zSpuUgmt0REv6QxC
ZEYv6YbaCQNVeBHzkGub9LYjrljgOx2BBjpzORODk9hk+9MDtEq7qSy+q2yD82P1Tz4R/WC5fKM3
akpECvhEFpEJuul/m9pYnrned+9CGCkls9jipvnZODqCvSs9mLXSJxC0UyuATT4+kIJNy+vYRJT6
4ETUutkJdpuTLvCHqNySUTZLyYwBE9ORcqnUI6VZOQjsIAy1bk5L/dxX101HbuFbuCjWn/OaUTZ9
XeI3Pvt5zVJLA1GRCII0ltsA+NnRRe6wc4qZqUG29dmHAlIyQ1Xx1gu6/E3yAKbR/ZK1EJsGxAAO
iDAZv3+xzdWDGGN2M/qV/7JminDjUm0nSshhNjpkpDGz3EItIuROrKwdBv5T8oCUW57woZgu2vqp
6VXs5M1mppuPl71py3sVRjx3D3Uyfc4gfjAM8u6AiGnvIc3qp3hwN4B2JHrnitLHPRwjDMhlAhUv
X13O+ts9ZFMuIH98KL+aCkO4TriMPzq3GG7TzF4Wn5x6Lj+UI4VapKZZvd9wl1BIOmPjA1C4lLQS
Fyw5HlZilAxml2HHYf9BAXwEMq5nRHRHeLpzKyIAiFEhP8DMKJAhZMCxQ1G3MWK6E1bG3uEKxpdw
vejJNJ0UmQbYI3ZmB1Hx8Tl0ChLF+EQnqSzdIn+iVPLzzH9cvXptTP1oaBYPFUliFLebOqpYkbO3
elxyTqBcdRx0x2BEzUiC+ONVXJT7/tU8JNCK7Jke1NGVGK5PcKOd7AqKDSnB9gFewwxDoeX+/NrY
RE7T2Wj8QBMetqCQjMT8yr0tH+XQaKuSapCoEPc35x4m3KD3fteoEqUGo1ZXFsyOABFWzs/JTb5H
2pkoFVqzqf8VyL5pxE/kMvXncapWgv85yjmj8p5DmHqd2QNASy7U9kB87tTM4e94TdrxH2LHtCy2
vNTkMs+V/eYE/YdMEWaOJXEw/9s9ZkGYSJoxfreKP5Qtf3cNlxaS56NoD1qUwwEWuYqA61TK7wpz
X7XX8lhRdPRzzU76+FwWiIHlcJYSjkk1Jummj9EcySij+FKo1EUwGoG2gyZSvNUytQqBeAslBPIY
W2Cit+e8aLuwV9fAuCnH50CFx0RyZieTM/R60RC4IeHsEUM1IPWcY/C0VVl+/LosDklyfn3NuMY4
6RVFi9NOWLJSsaIu/FXIzLASKN/AJLRAnNdB/bj2t4cnLD43x2Rq4uLmQCaPApSUZePGUpO2sG56
d/CperbRqpgE5VkChT/Lef1onSkUkWNAUyJvMkhhA3L2FiYFHCcp1nBRt45gj5UeFHCpAWJKxR4F
F3HySHTo7aD4d0daI578nftLN2LJBfSuEcH5GvXh71reu+lb5JzydjE09rB/J2+/31+MP97jkRdG
6ivjunCSsm7i1WXq3aYzh1PNQ808V65ZYr076N+fkoBj77paZWgDt/wMxZ/lRTw5aDL0n/ttLnlu
YwD27lQ4/JOS4Rg6w8LWsP0zom7brldGWsMKZgEJMaSayv4uGB7wFuxZY9OoB5HepJEF6x1vIR2k
sogqhfs7qWBjB3zUgHO6c2or7Ggx63iEEhzYBF5b7vr+9BtdphZouPXF9zs9cGUYjbea07oeWE7I
CEljVcqQAu/p4pJ8lWdQ7+c5bfmMQEsPTP1CDxA+76BGIQPBwbD08FX+A5ke1lhyIsq8c1WTZoLd
Q7RcjmAvOXfhj4ST0JMDR1W/YvlkVuakPdc0bWK9IYHPjvl2cPg9potRVmKg0QO9v7oGRFdN2PNo
/e9jTJgG8bb7ZxcqGuS/I/YgWvy7a6ZweG6l11T2GPXBQhRLgril7VJg8ybawehaRjDGWb16Xpdm
qZlc+DPDExM+an6XVD1QomQZm22pkBVnfdNlLNgM2nbK+GIP76Dvv7Ddi2fwrm2D9V5NCT+B8lqT
7oUY1HZWuDZRKQSzEo4z3NwDMBu1cMyaw+Sv+KabcbXuzDm0NLrsHWOSxBowcKJkUzulBlhAfE1B
tCcJg13aF3wXvRbAuhyCCY8wE8FoKCPmQvTzXXHSQ7lqid3laajHVesbxMOaqo31ySew2iqdyYoi
+mvIUjYgHwevKwDO4vUe9hDomYhTl95FpGOsczCLYpa86LJU673jlt+reSONzRE0cnojDQ5UeQpw
RgobcuNoF4thk54PecZ7N9s1aa1IAjknuERvKZx8tiBSnSMn7ER7fF3VLJ+pOVTQ9Jh+9DvRPMjr
ABjlQINFpnxvmL7p4euWVtOMPd40qE4e4G4XPP+Qnl90zchsSuhsrPJ0nmrtyKdS2MknWRf4fIMA
h4B5+NFVD9GbzG1HbziiaDdPXqoDbndpuzlmnniMMvEj1CikL6J3ceEN5Qg19k+hBCmGh+kE1grr
ROKzO1HnbPPo/xBadwRd2ZidGJ99W0QEAwlRtXFpZhG1JzYBGJf47YOTGub0eLTc8Dvz7A/XZXIM
M8lN1P1lqn8kDozfAs49iUPdINK7kUaxsHZ1vZQ+3clAkS8ThsjLBWBvaGaffcLn5B+UWQyknQX2
8ZUrR0qsIlILrLDVprOHMz7hshZ4Lun1wIO8zoUDNAxSOvrf2oa64pIJdueb5DK+Uk3VVyNkHR+H
m8Mn3p1EkaMUoiawbBxhtF7pLX8HsXKJVMp4d3iQgHzdRH2wVfSt5WfFel5P07VcFVhj6uPmoei+
BE8H8y8Z8i2NIC3Nhe5U43VbzQps6xqcPSLLmobRv3bypbjEr5aghNzhCSe1qW5L7n1QNmw+OjIZ
51/4ziWzvQfIni2Zh9uTnLvKxGxLxG4VAV5G574FRA+RMVFCrJKdOycJ3CTSh5/GN5FcksEV2vzc
PpT0D4mUasoLpJDxjBlczVqK3Ey7Wx3HcuuIYhjzQU9lHOmOB9s6A3pCXjtKH2IzmNJl82W48eUl
F/b4HaOBmgOoIoMk07CliOtDmK+hg+pjZMxmAO+G2EUuaWPHPdmc+TG0EmJI0hp9OlqpcduVIx63
WuW72NBjly+pJj+p7F3IdvxYsRbmxwTDXd8J/n2Gqc0mGjYTrD+1L0c5ox2UFeZ2mpv9s1z0sPi7
DHdgRIVuIFdUi76wwRapiVDeLpTC/WciRNRkHukateJr3HbJKe2el3m5/0J69iGigPQZPg5p+nPM
`protect end_protected
