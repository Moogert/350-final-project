-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OPD+nZGyf2SM8NdhibnvcX6dqqtpMbOqIvjmZbb5Bxu/gl1MmyHE6GlMJ44BTLVEI1vZ0KYxAAcZ
pbMbdu9TnWAns30ku7cRUmwkPfpd8OrkBKx5lBqAvYE1HSCDv1ErEY52kB8dWAUUcY03wIjZirON
Ai2KGOXrU9aUtNi0nSbIE23ROCwbX2V6x/Xpjw9HCrHerH46fMsLVC0Ho9HIFvK31xtLo7TcNU8h
M1HjS+K07gDgVcB1GhWGJ5y663SKoK+w6jWHwQb3RDyiEfJC4sKcXWf6EkDDzMf4ikTlTrKymvJJ
1W+forFvu0DU3EL+7dyTuZPx6jm87jxM0c9LXw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
/zsAQSIcBkBPtr/X2qtoZPC0ZMkAIBT9WSgQHaKSMRaxK27hgSo7j0kKhKg7W7HrwpqpW8npc5KB
IYksPIcxP/aKee4syxdXbq/XGQdSQ6RuLbJHw1fRr2DIj3TXFoVWRkEZHEf1OcVW4VNOMltujFk1
MyCnMfbPB8AAZSK5ckhKamqX1evnGnqpem5M3yTbsf5xTXCknKDNxIIyunx2aQBwUwBadOFvwezB
nl6qPdHdVR/bv+6j9oosdJoVA1vy9/ag9FuZjCnVFepF9Zwx4pfliXODzXvMGIR5gDxyZNEVXZ50
0eKhcrtGWUkOo/ADVh9T0B/Cp4H1Jn8diz9LeKL4gQnP0omej4iDsZr5WdsF1Ron32iIE+UZyudR
pKWZ2Zcv3D3NgsiFNhMeGzL8yG0QKeESsm6VnldHcVRxVcJY0C7Cv2QAEW6r9ZkHm0duVvzA6pnV
w1p2OzA/F28JoXn6+yNve2V8Ce8Ya46LLAkaFPQyFjHWUiXSNMpavymLxOAIEVxzFf36Y88jiVOW
QMEJg3EHtPTC8iXlaIZcs1KpmDUtimHVv5os6bR+2u27nA7SwDvMaEsjMnc25aoj/PMZ+TuW8PNh
yMtMiVhv8LiUQ88CE2yVWPeBvO5EyMyWnxXUUVs+jX+VFRLmKHT7BXzpCK4M+JOy7WwliGfXGJh3
Z6Gu56BGYCP7FnGJ1XQ2We6gJwAUhYmCJqFqJaSDAzAVEZcGbldA8F5Cl99OKR6o8IdWx6jeEZAf
l8KADAXCoL801nGOBrmzUEs54SZ7wxhvuDE4FlxCOo4M4fgidlEz/fLMNFOgKz2rdK7PIAi2UrE7
nGBXFC7ABtFZ/nVXgyabDY35aGnYqV61HeHYfa7ZDCfdl/YoTZa82LRnoKrjsSVz2cvNHKhU4RjF
qU5a5JYoaI/xDLbIfzexp7rc+68+ACG2lUAvef+Y3s6JsU061VPSJiF3Xz//0viC5lZ614YVyKE2
rLBiq9uv/9rW2PjFu5bxdYrJQT3kDu0Nx/LpV75qwuKEzNeG2LwirDFv3s+dMKlzI6sorLm/b0q0
XIMEjbmVYjsc2KoKUJ6sPv+lEXzAHWj/QwJqpyKgRDq/oxmxMX2MY3+zrs7mYbTRgy44HlHu7vdi
bh6TM9a2Jj1Ao+zWs2R+Imggqowk7DtlTtqnWibI1AUhYmbBwggJfwgbSFCv10EtBCBi390d6EK0
oTElyZ+XPUpEvKXMjH3XdZl77VkPdJAFp1kaFaYdNBumkZFa9Bahw1NPTSdHF5/B7DpBcSMevSj9
oWKHgoZ76P7XOY/9GRdXtjeqYaVcL3TtcSF5OnMOj2kb8oGaspvLWTpNp545v2zPOTNHfokue2Dc
d86Tvrb8dbStwtcf8o48dyOGUd35nwHbtoKkAiHHkLv0vYSaSMmsS6TTJh0whqfpA0rpauM15owJ
2G7FVd+hc4UkPc6zkY0pGE0saALSJARail/pTkB4sJxPa/2h6C5/rJyfYjgvWXZqo973dCr12rls
kRlHAnd1Uc1H/gpQ2Q7GMyLX4wmV9cWAykLDKlwcC+9NdffSNymODKEPzLWQh3Re7maNztVmP3T9
UTTUoGUx9Ky24vA8X8DOeebjdovz/wwoTc+RqpV5nZ4HaavnsXmIkVVXz4+uHsXYIOp5db2PqdeW
+4NHIRFiW+GskS+UcZb9niGXtCsK629nSaaHfZ9g687d2cukakEZSL7uq3YUYuTmA4AVpiZsrh1C
uH3plHEdceVd3IKHLkQr89mZiIdmdtzY5LO7iSiiqm9G1T5H8c1SBjN37P5qaz1lICOxgfnz05Ab
8P/ACUqz4LCfFYFyHPPjyMc44kWEoPcIGCLI1d7PXQwU01FkPh2pesPMbFMPQXQc0lNktvVEFOff
sfw6iF7T9xZQm8bR7PmNSY1SOFm12ltq63z5t37AqWrBNT52qiz6ZswpgaqXQtlTBrBiJBfQWhtn
PtQQ24gHnq2gfftWS7XI8pD2pdo3E7WkwMbSVlT3FUX2PgHnNzfg3um2Wquev8D3uukcYAygjbKh
Eym13GcgchQIy7j0B+tvZSaifkKQ+7vtCB7OR5fVse6S5erCKY+mj0kMO1N4QKRVqCVLA3vWgLgf
6qDI1r/FSPH4s4PRUIui6zXB8V6ybN33lUC44w/6S+F/HfEV5yJ/c5aHKf5RGYQqWogrgP9oK0pC
V6UJgQzpbjSHHl8N4kCBxAY7T1ZP+3roK60FYqZHZKXNuBY5fId/zDinszFjKwgLqNkUx4My8B8V
n7jqC3FAmN5un/NS6ExeBCNX3BLDlOysnlgogJbj2hvFQL5IkPczDND0A5FZ454pAtKpF1d7WDK9
ovN9dwM6AxkViCbFn5eznNuDkyVs7L/IGvFiEOP3BbLS7UCJb1i0cloV2cv04GrGNShTomcGs57Z
KaVSeFhyeou5/Wizu/qn6hbMhh/o8SALn6WGpEnR4ZF6uzZHfEXmYYWbcXd0yxtgWwR7vCupHhrG
9K6sleoMFiQo9kuQSXOxyrGp7m6oexQKtNkVv2o6VThK4VbbJxGhEXJhLhFvDnMffKV0zPLNRVvN
D94MDlWw7RVjxnJCzsYQ21Mv39cN2UP8x73pA9BHU9BKi1E3sIAaQMO2wYvlyF7bfFQcxuy9zfqs
oWOeFXXVT409W0zOUedWE+K6BNRCycwh8xKcmqoWhGMJx970mCnF70A8pSwyuM8cgg8tAhpnLsAH
DApzDtfPVqY9+nVmvhC7BjnO6ihUjjoiHd7SApDjrvE/T9kFttF9oz1or40toV+bEzUJx/MmrQi3
zknhRcAtV3O6TuIVtqY7OsJlUE/4Yg6QVeFjxojnOS92kXhBKJSrLRJVSfjw97GMqPKihub1IkrO
DRAao5SALMAWfMM4YBulYySj23xofv/l5uRn8GDaPVeR6okCYuND9/9T/9lU+5Zm6K4LtFJ+Kkmq
Zx2vTYnntK0EPtt+F9fBUxIDcd3jCbZxRHKRl3FeyN7MfiFc/10A/UBmNkVp3T2jZVQPPcqNGyO7
b2SEzibP59K6MHJYjQ/v45k5JmavIWT80J9KldLsDWFfN9i+xDtP0HT9ud4SRt7VvkPulN9T8H5e
ZO+NgVrjpS1NXJTmDQudPKbe8vcMKgaSyxSW/6FerH6UcOIuONWwm+VV+mXENOKyc8MBwA7et80O
XxYjDRRIuJSb6Tju+Jl2hnJ9V9KUYTespSmC4D3VeIdriVK4irMkmY5XJZdvJhnE4AiYXQZhtE4B
WgxuwQQcDn31ZeZW0hbvbAphWdgKEr+rbhwCnaPUw5oQ7KESk9PpY0pxIZ+uNd5C5FXx6iDCXJRG
eUsb1XTWxdw2RQqsk4ILd3sQr1VBqtfPYi+B4XsKg7bSlEC7H0dyPHpL69njkuMNck1EiDiFBP5Q
YBlPkB8+eGRLwhIt8SV+hnyp48gFiTTgPoK3Oq/3aw6nF6At20sdXN/TR7lsUzp6o/DOdMDjGopa
jygkP8Zb0QpriQguY9f6/jSaW+KALjid8sz27HrYnGm24pU/C7qUz7whBxCZbdD44XbclGspSdi+
5WzxZ8u9AgjR5SFXu33wFyqveEWMAnRHWCvPaIV3zhs3v3Q1NJvZcNOSD5sHXAbAP/I4LJfn8njo
cRErJLt2SsSeLVkvTjgkH7Jrt8nVaL0gNCSGvAphOf9gam026wLjdPZUm6ZugHGnitkUZrUDSnMk
HLK4hzgIiGC7o2gsrw0u7MxnoxDVAbyp22jOmuLUQmRPhrqSIMw+GQ99Alz8iZx7/St7sO44M8Xs
mvwmFcedPJMN6bDaRXk34z4KvhLilYuSS4UQZPxSQVYFnXu16cnsTvCvKSPIhc3ghq5LG9+CQeBI
/aD5i7YD1qJd8fpt0xSGwRpm6L0BSR02AmmARIis5mLo/KNu+eB48mVe6yEj0TCsQWgduMKfxy7v
6NyNwKiOgxKBdikm+GI95H/im7pirAVrbltPRqWeFFFGEaxAt09KnpgJ4cfdfuPvEEp1If+bK8vt
T9yCz+Oe80lea6ch9ye2hc7y1MiAcqxzY09e4n6zerjIB0xw7C0sKvvBfyMRRSxiIDMzPpNN7zfR
koFm+afKoIQ3v2zGy5poz1QHtCiFLLvcygosa38i2WcaBd1BtMvxQfB7b+zfgX9rEE2+52PBGaxW
Fu/I8Vepo882kXoCkb/ij3ZnYgfy3QMyY4gSAdwH5/rWydsYvdiTYuvVnnc6UAyNHo+YnqK64Y9Z
g+OWPrdZggp7Y/sYa9yuoYTbhigusaFlZ2j2pk+kR5/xA9P6DCC9A1RR9xhL8s258pgkADUmKDA1
7NwR0TD9hNEiH4JBlV/rdIdHhIdAYDAonzIzVw+uFteHrWGWVU+EP7gn9RNsnVCfrg31RLik509p
3ywd/F0JMsk/NZJkF5ihwzU+hlgzwoOX93wXDCb6yl5PSGHTacUynzBdjZy4WYPtQcpVJu4u8myG
G4xwjFROT+L+297RdgUHJdTlStdYhSi47sNFLglT5vS4WBuCJ1y6QxZQrj8lmdVVFTUg9/QwMIHE
ks3h84vH9hvU8k5qYUipYUGN/rzWVKgyse5GEVxp+t2ARmqyrM7aZBmuj79+t4/w1fP+xaOwGCKL
9B0vP2ACy8qmNYsX3Ofr2cIcnAA46EkgtBxVQtfBsHoOmJFJT6mOAWlBFpnZsMrJkoznLunYVWmv
S8Z+/BRuGwxYBfRhFxgnvofzgSQ3omy1+Ju+1tabvTyu2CwNGL1fy2Zh+9ifJfsbLTEU8vZWNWpq
KV72tsoQUZtVEe0ovAQZ8k0fBe54SQjZi3OKSRjPYhaSNT3jRb3R8iWMpZmMW1ZKQqXsfRx0OThp
WjFlx+3tG+CYTz371lqCB37imTBwfjk8z+s+50awEtORjW3DRmLhdvvGadlT4SA8hKU0vLZ0ROvy
PFiBnQydMZSrixmMg2VEdmJT6JeJe/2RjnrzLfOYQ/kjj2A4zwsaSEES1mhxMOrdelj8FzsFHs+I
yKA1jOJlDsfH96AVlLU50jfRg46Er4cmetx8tT5vPi0YJRSOP6doIMHr68h6LBKlZuU/MdHofI+8
vajlgkUY8WALVBTzUrV2/B8RiArN3Jdc+qbZt/nGa6X0AiU0qsKMdxFsWHNB3Gp9u0FgGa3uyXrV
ZrtDaxeijlIFoxA3+FDfUMnIJtZgQ228omOfR2TCr8tAdXimsfAIzx3Fezsksi4XLdiVIdd+w99k
NBtXf+CTwy8Z0VU0G4Xapd+I/JnP4opf40cwfY3DweGQHIWUU6lfvQTamzftQHxJNo7wMhH/Ydcp
ZDXwJ4k9CI8XpB1ZtNt5/OT7PRPsylsaV6OwZLHeWxaoHtbYUCKjAivWGEPlzPkKkxn1T92QALJo
JN7pWVHlxKUIs6e0iK1m5D5q4HM7nO/ZqACCoj5Gmi77mz5s+pEE/HhJ0N/TVl465JENYok+uM08
mSN5J49jDOcWIm67Z1wtLvkbJpAQ4sfShbWVDxOKLfXw0PNedkHkcmeonZTPCLtI1S00RjyozaxT
ygjmaHJijqXZL+GKTrfvwx/cJ79Bth70Q2viPBVSjE+YABQVtwnlGKQmYyHJEBBUxoSrufQyujEk
16brBYz4JYKNuWwpdfKU57w95WtzAx2MdTodGAK48lNV5d82B93Ta/jZQVirlZB572q1ezyIPpzG
Pik4dtYKgx/ECYUlfnow/sGydrRNo0j0ErshMHVehCTtWn45n6zfhbeZatdTInhjYfS+ho7umKsY
EHSkLtMMFgvbFGtL/i5pIU0eSIake556z0ZtyFqFAWq0NgpT64s/78sfQ89EOPY6p9xtXjS1Bb/8
R7zZmCFuXxST4N0G5nbVsBdLSvwFACXoNeGezQg4beDMU3Nlx1Ib6BVvfaYbaLeCeIXdqHeaowiT
IwMLmwRM+KcMfNd5gEMuqrQJPC6llh1olJkO0Ne3ENFVBAFs2/OaheQE4sWfulrLQgOK7QGfQBIC
LZbit7CKrBEf0FP2CWcs4jmxZr2ziDLduZWPBBtMOq7HUR6Uf3bThAKhXS0PRVmM67tmoFVz9AFQ
R+QHFa2C2fM4yiwphod8cPDQ+UE151svaIc0dvGOvJS2tJ07QYIVkYI53ZApA5/J88B+vbvRxIn5
sNQXyr8e8mjQRV/Su6LX2r0FeQwfbJ2CyXIsK2XkXYcmNKryYL4BLuaZUFBK7RO8Ub275YOmEBCT
MaZp3lHdxljvDfYnPJDBMFVaJCjkBnRvcW9Zpxx1z6vN4KEuF8D+4i82a89s5L1O5muEcGGEDsxa
4AJSXHoayTJVhD6xRuut4N1Ts0NjzSGRfoEnaeNSTX6eyNou3/37n9zY9tsAN5/QgllAxzwLs8AE
9BYlkjasaET0ZqzRybimrk0ZgYddMCh9BbSKgVzmNirk/44FumNEu4597Qbq5ZbQqY0WepLm7me5
mnNgBx06AD7dxEmnesIvG6rOkKIzz1vGOzHsgyrS5XUks0Lo3FabIE0J9EX2d0dt60RQZqZCc95S
X1nVuK7ZZODtFu9/aD+nStDFgIFMOr17pbLG6C7UMrluvzuJsky0PVIon6J//BjzcJ61zn9X42YB
1wQyP3Ozbx+Vmp/Vcm1tsvp7stC4TNFoDenCvrXM8d2cksgp9M2PoDeBd9sBA+5QtBO9ITFhwc2J
2rcCg7W9qd9CF0XNyaAx+/z+elnE99FlhQEKivxc8pRObpUN0Q/PssdQGCI3N8FgtgXFqj9AYoRv
zTE6t6MNAmKG9hK+gnpzKZDC5rZO5wsCDdyaGsFdiPzVoSo0JrEgLPl4GhDoOXjPIibPXN5PBf5+
oBGPAKi5VFF0uJweC/7XbK7AJZx01pFSUSlCQeB8Dwun6jhD3xpX356W6fqi073yiop36p+qPU4Z
ZMjtw2cmh/+EWoqmXqwGqZuk6nYyHmJyPsvtExiYBbsNc4P8q/LbcHVCZDEHRzhP2cRFZrVhVseD
u4dacSTTTcBCKGPGfe5ELCMW/fPfk6T7rqgxujZDikiB+GDBLfSvtrDdomR/ZcdnxVmsWXHlxTF8
m63DooKubwdVPPjodLwIBj23ppfhSKQ3RngfqYw1+wt5acaU1t006solmhnLVVWUwBVNxSDsxMoE
mNeIG1IeWosl1SgkNWeiIZ/Ci7/5/1SPa1GBWk/GQTC05Ppjv0vVsk7j5E7DH0H8gFH8tK3BxF/j
AiTTaMfC4qOxXDCawE/diYivdaJ9ZhKvFMzDLNhhIONVrrCLxohCq4RjxyatsWN91O1wmSJob+Fq
ZwYC98A0XXtsCzdbGk22fbClHIgamXB8UwO1sZ0tby5pSobX1eGDZmROe6lNTUOQA8xzVoXGw+kM
/mCis65CCV8LeQTaqRrrJGUNRn1bONdlTxolhoIaQV9iJBsIqVtLaqjwU83UApVvp5sY0ouuGf5B
b9vFoyxa6zl18VqcFXOa9R1l721sRjYArL/1ryVscalcJmo9EqjUXzmW1gexQycghcp8h/r2pqBN
wHPATBNTbuKKPjRv8M9hPBpVthEi5EWZ9ACzc9Ck9BJdTG/i1NjQaTJLcaeGQWzqTXDmg5/PlYra
EvAQ/cEe385/MkztqTp1+c/X3c4wG+ublucJ3Gts3R9kC10qi1ppIPpcMQiCkeDXN9STNnijVvEr
RRWdClTdM0J6kpnndikruoznXZs6AY6cjwwYGFwOflnOx6W4ziTgema/YviqjUG2YMWbDDsyXs/Y
9KvLfg56q5TVIAyMeRIDSBKCs+jLBZmkhydMpACjN0pmp/0PWYooieqFAFvR3dl8qgfW2EG2Dvn1
33HRZG2u0z8MD+XupKzr+esVUEsm1qj2s3yMoOVxMeIOiT4XJKFWldU2EWS1hHaXTW7DpznyM1KH
t6uH65LTOGkG5FSK0bE9Nxo4IqUQcSWJJT4ioZx17aKcolKZfDKObHsRXpNiUXJN8qC8TRH2sxiO
9QK9Wmt1D7piF3IiJxoipn7Ij3oqR90lenUY3Y1wsDGEcRizcskK7kOJYClaqSMkSoTzYywo078j
Dc7+ZJlSThFu0kIUDZQMOn/dsqeDzVBZROgbON81IROEi2SqHrjoV5i4musHilwyFfIk1YFCYQD4
l0VmDrYHTZ49CzRK98rpSgoRADKTlqa1eMMM6DL5Jj6ndETjN2+Elxhwh2GROzmEmryGRldCZTtY
vzDhQyA1OkOXMr/TjhwexblXFpIpE98a65og30mRpnvz6U8jdbMu+FeoXsxy1tYliuITB6glwcCV
fddGTY3yVGopiiVdQttfSDjL4pkLzqhLDoB7KbFvb/n8Q0mC8i/Frp+cjV/QoG7oPdclwGUq4OGf
8G05TYJbwtoTkTCxbZ3p8vusddmL4rMo6YC0beo9ezYHwTypvCqPUBJOnJPpmaBR4nwhzt1m7U74
9ZWUq6r+91suTaArLlNxC30hIbKzS3BytI2DeyXH/Shpmelr50TgXHuf7GOAqsldMX5zuISPNwwv
Rg8b+5nc+Kj5dONdWpdBw/tMKbXLt4T/rLJA36sHyXhBDG7/2dqNuJSKfoakYW68AEM+T6QdSYBJ
WUqVd0Q63T2PR2lWE6VN6Uc2zP7jdcOivUfUO0Gnyo3udfhM5ZxiG//zz8XbJOzqul8LNkWhyqoS
aGkKGe1ZAc3tJl8Vxz8WVAssE2dSCuxypnLlm0LT1ynaDRAU00ppl0pRApLWLCt4lDO7l9xo2cd3
8epCCsWOacUS5oC2ARBqFuxlS05MpU9ofPV96+eScOnTYJar05TIX6e/o5aV/JQCXtVHLnosxHa1
7JDMDOV1JneMLD9NhGq+rd9cLtfCe4cY4tU2fSqZAIuPVGZELkRMgsjLtHY0YNyz7tMG222bfSqy
yoClfaK38A3kaxXEwOpbHauORkvg6x6lVRIj/ytvjjp3wlcJXiWHmX8XhbvnXzdDJaL/ZHjHzxCG
qNvpeLIVZskR14KHX/XMHZIAdh4m44bmrqSxh/wAFwWeelSIMAcMSCE+GeU7N3MJRYQ45cj41xhz
tN1ZLjTqGk5J1oaeCUC8n56bNu9mJMWV/ADCFpQxefQZ7SnBMLE3xzg9arQfvnv7inxYjMf8STWB
0jJzc2yyNvWR4tSmzo87Rhn5K9jrmj+ucYyTOAQqIcrx2hWXe+RIjQgty5YfBlT+NM1JbekobmfH
Q6ZP+BlOCwrGsI/iFoUUPa94T13oI7gyX92YeomLfDR96tAFeW3vKOsY7K0rZEUEm/TFQUM4oi/T
NdPsMNSZ1csTGLPVbTQ7/rxDRmPKYHI5MbRyefknCBTaM+uhce9YSk3gZerShRlq7WMAd/WV322B
UECNjPvTPVJoxvtz2LUm5TFz6kTZXiq2y7FmiKP+Hj+H2AW2ddePEgZ3DYwCNhIkqwmrqiC2mq/F
8IN5EKioxnb6XP0PCUKrqkR18erYGHxyDYnZeP0VIJ0FYp/J770uwR6VjBvxsodX1UfzqoI8QHA4
kts5wQiGMjpdBds7/l+ziXbPE4CFrJ2UB/z085XDJMcp9lYTkg9YRJcShsBurLTs578R6HR7Bg2Z
hdSG7mKPTObDiUozrPCBEpLMpPHt5VniGIVDhO3MNTcf+T9ZiSsIflOyT9Zc6BFYMCsV69gw0tZ7
VW7FSmhRtCVDti5D9fdcdh81enUbuOjaehiQEsubpP2d9WKymGtW0G763rPcS6WfDcjqFYtHJX2f
FMx1+XnVFgqDn9i6ro6ECguBWV81xU0a+1uDlr0hhvb6rgZLJoEKIYUZUKDl/zzlwm1Duy08eXMc
Mkd/qb1ZEsdQvlB2wzznaOFksaL/TiAQZOWgONa0W9PTBNdpDC/kCzihvNwPPsPRp149QDfJqo25
d81LgNHci3poRMSYP+9kRtbRNP7QcRpQZUpWf+K+mtfWXqLQtNVbt9YZZEMJLS1S+Lsjrm0wQVmA
uhUeUUgSex2bzhP+P+8vjiti7ZCUCmGk7LXC71x/A41aJFlZwUO5360Pasv2UTlbB50Gv/qMQyX9
/SS4jg21wokHQGW5xBLHovqKsKe0A/7c+hFkaVr/iVh7bgNSIeo7s+zsk9yoEbn9BVe78ZSFvTCB
/wtWTRB4IxvWIg423M2QV8t84xXF/LvkCc+/PCPU7XDwZ7Z17RTzGs2j3q1SjsHBl9i088CWhNDe
g38rYiEqBIzgAarKb5ilMESuUbj8rI00RkK7uh4jylTZ9F32uYRMiVdlzkV3bpeY+UW7kCP30R14
Wi6Wx9cX+AxJNpQTwinnnysA7Nwl1aeJNA2JbQMjA3IGIiOGUm2EhfYTdGts3lWc+Ax5f/8ogni1
VPKJ0JLifk3MtA3z82MH0R4/A4FVd8EYZb3zw8b9jJ5+kLbybXk1v2KScBCpcs2GllGWnH5a5p+G
SD1t4oUfYEuT2T4h6yNJeKssAuak0A6JUzxnPF7ejK9An9vYvXnCZ0KrBoq0YfhFVE9vFAtPKfqw
Y5dIoTAUWiIlyFPYNDSnAWyj3dQPClWfktcpebUHQSiPz0DVgFO9oF6i0ezjCAYk0u8ZIG22/Sqe
n4R3gISTEgYvnWPSoMo2DR9hENCWkaMyNg+zgi8zWYfK/GP13cBxae0UFucUQAd826UZXwQyRwB6
hlfCDr74y/yY0MUI6IgB2PhFxXJ65HMYXeBjqQ5FYa/31AUjf016GUdc3Nr21eITdftpKjok+6OC
0/r0/UJ8HQQAJdpNV2KlnNmtDAU/XF+rGSarw71nBEo2RK9ijfUxHCdlEppPLt0Xt3GxaEeedR6N
LXgt5DpgmdSJfLNM7BRN+0EM4nETWL1lNTWG8qiA+oJI4ndnvM0GPESSU4RHgNCaipH+5eh4gmQf
lV57nJMkZmY4qxJJiCdYeX7HW3arI2nc8QL6kwRy1Obj+wsWEjR5osd1sV4y9KXowh0VqlL3En5c
/OAE481X8divvTXfQnSoPL79lUcy8wFkMvPMM/T7QVL3jEm1cfcZiwVju+jsK8xM6mm3rOrKzmSw
fg3Q5Nr0Dh3Q4d/0x0Nj+q9pl6g+HK/2NJg4k0Gr9S+xu9/PAABrJicTUEcn2VqtG/Vgb4u/rIGk
8HQ3tg9twzO1VkZVa90JpHhsxfzGud39RnUhTEcuBEKHtFfPhcTbe10tDJeWv6euD5iUD7UeQsNq
nKk+Q0VW3kx3npHo/66ranJro+2bANY5djgxmqAL+mdx37gfhnlczQkv6jtp4sQMmVMkVOUbhDKb
sXKiKjhNN3hyv7NPTsZ2ktyYyMRp2zLtpvGbv2sae05ufZ3/Pg/T9tVl/OFQwZG8eZpBM+E+nMBY
+wnioFcLVHILtm18sm+vY9+uJ4pLZkntFj1F2LvgTbGAs2JZsPgCifNqDGaYIUw3liWNmVt8Fz73
7HYPGRdLQOuPB+Y2j3eIZU3RZyq5F42ZGQf1D7XawjG6Nn0SqxJTMbh8g5xMrb8SCI8tBViaA5qz
HNaSOXfSvtWp0BrEpf8H5ttdMLD8M32W4/aWiHsZqY9BiG3G58M09Aqr1TYA8BCs+he2bvI4bAqA
eLbe6Khz1bA8gdHpCz6NMLF1cM027dKh3MR5myTV2T1ARwf6dFGIdOsfqGBUf4lotXJO8jup87Fi
gaWVXEffJlYzOlfjQqX1AYCyQI7zr2Q0p9YMAGaeq07zdad1qJfQcWx+S5eL+aKFB+Fqu6UqIGS0
wcSDONDicyHA5BF6JtTPNhkBGj3v4ZtZB8b3M+W+YgoLCbU4kN+NkkUYtoDbZ0q831aWW+S02WKH
yoTDQLXYrc1P+yOwB/UMRvyYTKrFKitHesGoOXRVfGB1j3Cgu0suB1TnRK1ylj3PMbnKaH0viA9r
I7LhQsDIzLby7BFVibt76OmO3yeDV4O9iiLCW2r2RnGoa2948gEG2DyVBFtQaUya3P4F02zde2pD
+GNoA9NJnvQK914v7HfUL6lpzsPynDwHj3t9rGxwyvVoThUTSCrCq19+jn6BDx5WfS7I23BMDlvX
2M9gp2uh+JlBJq9vdhvcbiRC4rUNbuMOy7Utn9fImmoEWshFSDhNB8tubvB3QUuBl42OOtdroFkr
uASlIV7hn9s8R8Fx3S8DutMlB61Zt33P6cS28ajGLnSEPFPniak8UvCV8btwLs1cb5+6WJOzyJrc
cAT50qlMSYx4cZViLNAzuONzPxdDplcKx5/81CG090catSZROftAusyszP1FrG1YWr0ISnY2CQhU
SQR20qiKi69RKYUtOxCUqVes4fgXUZYOmzRqzAkIbOgWsL6+EjPldMGnE1wFYO2zQALHjpFXNLtG
Ko5G94bRix9RYsATSA59gAAosJKD8pln+z5xrg3S+apFB4pcegavTlu2SRKn0HJcPtKmf9r87pY7
T4S/GkRWtp+Lei/WwlcQgMhFQ+/vTl878wyg8FvBechkNHpvhINx62VIwzgoVJ5Ha/rosQOFwjgb
t/t2I56hKw+3RWGrWk37mFa3mWUvB2kIDYkx+L1ZMl4lpseVRnzPvj6tACgKaFwSguJ98imA0+uP
x6yhMOK18EyI8R+27SEYVSPuSbS376meSmuL5ByaO7/X1iAeIf9IxIHBbQeNwVQCs1m36A/y1GaU
/QLUkrzOi/7Oylo70Up50doVyI7TWtudNTltXVZKdHQ6oYlSgDNLDPOE16HCETEg1R3H/bK3uh3a
ULnUobLJQUfw8uRXPwS9yLAkejNrWQdsIWlLpcI0qBHdXU15qZn+eE40SeijC/TvnxfHV2wmWUKv
qg1PQoCdb47yPZ3C0sDb79bEhFFefH+lK/z2MAnzvyojlYV64vhn8O5KBKQzOvI7UFPtnC5MVUnq
keq3gJA+451CQ7QubVhMcx7AQB4N1gqNyxGuotlUdPB3InAV/14kfn4gE+QaFqULgm5jeVUwPk6g
zPiQaUJaiW+olw/c1+ABjo2GiR3F5jLONelXQfM2sBkDON9jJuXaflaT/Ct9Q9mpl11my4Lh1Tcj
U+ikUtKEGIY0ZAiN2GZ3kQtOeesN56vKUIvbplD5Ik5mdjhxqF3b5U7W+NnH0o/n2FankegYETis
CN7O+EgiSOaNqijI8OGsd7mg8SHYV/ym7LFojNK8VvkUwVwugqhuo2PkhslTkaI5y8E65iCjP8Yj
Hwe4tevxzeHNu6pAQjuleW7uBQ8IMHlBIB0r8aRCqva6xeGKkmsS/8nG8t3vEU6sAWueExAeP/N4
Sp3YoGwlfLkX1oLYsckku3nCEDenCpACl3CFmmamCm+bYpWXS1hWKl0/97hIphv8CH36Eo9J2dy+
N2CTmqWu7vYgH42mH1c37XORvwnpbA8wHPq8Sl6buOoBbpToV9oY/LA0ydhCkQeyfy0i9NErNS4a
NN+O55KRGtm/cVa8dAO6gYjmyeoEP0NluNuKox54unWXtIeneJw7uAMV5o8xgUIp/1vHn/WBGdLk
LNqNxQQytYTVree6TrKop1R4Vj7S0L6STnx7bDjm2+l0giKNj50kfTkJ0ZWEbda83yYQrQeatDOY
ghS/sVRzOL2Se465NQTOA/e7/oNygKbDOLnPv05J5P+LjnZ8Bp0afCibei0bQVv0idbfryqpHcAq
nIg5G8eokc/EpP86jzGEHSxyG0GBPEaJcUERSnXLEcyHauH1pDq5HginQGd6Q/KLKErMmaqw34A3
eIdr7i+L7bGW4x1Du/JWX+Z4EyiPQwSyXYKF0jgIYQBFJsS5TultTS0zQT7oaIt39uZ7AHRUVKMZ
jJeiEVbwKPvOb/ZUB1aW3ZUMHp1Hv4XlDI/33cNtedDJPPtH7KpaCY9RXWxSedlSyO7ehbsXif68
2Ja6oGqEKRncPLMxJafCo8W/+funITVBl1QJnhE294YYtT+SzrEmH33+PnGv260u3h5ZqMtG6hFx
ewgBmQd0AjEH+C2lzD2XV1yL+0S7qJAAt9DlhHiKESJjJcPzG3fcqKUC08FzRLH9hWm5LoJfz1S4
hygaeCugGN4NOeH4dLvJW1f81uOAcVBqQrdfjiP+Vx9Wyr2Dv6GhWUEATzkg6LRqzn9IeAzTQz8F
kCrBcI6x9yEXK6u1t9eewkQrXNtVv9mofhy/Cc422ywJk7dw/AV47PfjoFR6f/qrD8bPE5w0WkRo
5uUw+/BVL3N3TxWB0uwZVSpd4EnUJ3F77otlV5+7k3peP5FDdysUkWnqDKFncCVjgFslBCYf8e34
7pr9nw8iME3nUgpTawDW0+klC1I2QiB8dGmruNt7X9I5zN7CsOV9pWbUDZVYYsPsDMeTa7vD2LWe
SktiS71xTlVx68sOrLXapLM0GN4QkPYGrp56H0NPCXZ639mO68R5fFiJ8gzLwdY9kyJfJVbI4Plz
PyBt2wM5yZ5wkQ2BNberLZXWgYopNtuNIuYZAerGl1tM3qLIL63BPwl61KBGu1O2KXYJUZCsW9F6
SvWosrfRkmPvOR8TuDgIdbNJ4SUB3oEH0cewD7df1hHw6ylv42jvn2hDNtmaZ2hjxLDEhbQ7U8TH
QtDQOX5qTDyrd8Ws5uyDdM2UdhpUjQigsMhGMMC0ZKixu6zDJK4vAk+aw0hpVTTdo1hqJf1JsG1e
ksQG9CXOgBnj3LbNX8e7RWBWh0fpbfwGysNjzGK9+oSjSfXfzSfYCc2u58PzESyQyotK89bEo3Tz
+ratz0HDWkG+hWMxB2qf2KCm9hXfeUVKTeKyxufC4tBA0Cwh+vkgSj8pqcG1hITOinGAs3NvvMlE
DdrJwnJ6HvedRO1XsRrTmC1n8e880BejKIrL8IebZFoYqw6g3JOYQ4irnm8WSbVQfcl4AoWTK/uP
uH862qZ9HvShz3hbjxs4vPisUiHnKNGkHyIrB/vZK/l8PCxvdsqjTBxGkFgykFDhAJmsL+dWm/Kj
yn3bWhmW5L9N7nET57WukEPw+aI/1IgvjRLruaezjNp/nkOu+9rtsPJ8NpFkJ/u6bkPADvbL9KyD
s3nZgh4eE0tt/YfMPl9wz4IgRj384YXtGE0f4PDh+05tt19C7TuNCMa8aRSGaskOtkih0yeoadpQ
ySLSeFmENAix0CV2ms9N+1+ZaTnSnU6lF/SXv4Fk/ohnmmX1zfY5ZCXFDJ1cdZBpDaNNjvaXINI2
/9knbTRE1RepW25ESPdSHcNK5Zd4sILjjGyVBYMVYzfwc9cKUtAeKqj5zeuaHI6PN05wqGhdb62p
C8XYBOurgtKIV5eKY0Kmra/YI8QhKcLP6UtS+QhwbM/AvVK/JgmKzzD9GUYxZiJrKAXUDn2TlKP9
ubcgFx5BF1FjV/4VoEtZU0q1197m6QdkssE8fHaMpOqsVcE/do4mYf2Tlsz85YgDizprDW05vfhz
SZ/4b1FZy1Ykxaq1FbNBG6g7YdZMWfzj9Jz3DDW2dWxSlKSxycBQiItybPp15Taz8Zo/a6qnzc2V
jMA4cKNR60Psv+VJUd3MCasVo+gNhtOfokI12yUXNYpJiIOog5ikO2OyS7xBOjJjh+xBB+bFJhgM
gk/WauMrNJhXWD/0S8v/owo6jPX5pNdYmosrvzOpVTM6G1iVgHrMgJgkJC44e49Rnt4uERw3fsGL
K5gZe/Ud5UTChXhYXVDyzFGp0hIqbZ69pSTGOpAUxK7JSjZNObP1xklCQ1Ru468oAiExAu6dca5h
PjlDBkkkWum9rHtLLv9VJRiGcI6H4VOijTMdFYlKjEstbapGPhJ9B6l65iiuwb1s/VWf1BHwNUDN
JuSt83vU7rYDZA6nq8jgTn6i9Kcte5PVLyZoV0JDeWE64GOYujdmetKJK4sOHlosnjEKK97ORt9S
B8kD6wInzuxcgpvXuJ76avuQbqSK+G4ZupCkFBOqoyRcPgfoJKNpjBcK+knXDX4sldv/9X/5Ol/f
LtMqdyhGYp1/Z0SucWiKwX6Zm0NYv23skKvR/IpRJGSMDFZL0c8tGyVrKxgz/ukvUJgO2lQb9G14
eqgk5Dlx9C/PNrAo+4maHTA2TuoQtLsLWT71E+XR1DpoWNXfWg0fMkavJSE5rfhWK/P2gyhZtUDL
Nj1zEsYZgPfKOwfT1IJaygamnu2mSF+AkUGmvf1vvrjUNJ105rDzEHcuOEcL0tejvvG9lkOlaSM3
g+pQigN7XAw7zFf+qsFLY8Sc/bAq84deKhtozRsvs9WO2FpAzwevLxdI50+enfes9ZBS1VPKqRVX
tmeiBXDfPHAA0MQ8F/Fdcsy4H4pjFEATmZGlWUfgsvI/zwT9odqi2s17k0lpPnrj+ScVkOo3dpNm
4tG91AcofY9NpEBWB2UJsYKZF6LT3OGOQ7ZzNqFMQMDEDK8gEmj/zU1yKQ0bKXktXQa7E2BxfrCP
Tu/xWtzAMpe8H/iIj4s0Nnpd7FsJNe3aU31Jii2FtxOGcyK37Dc72KNmweEdlwFiXVYhqwD80bug
bJwLFHXwDoBzrycqrQIJFOYvWTs8VcAr8sy8RzCS1MM49D5XAJkumbQihGAGT7lUjd99Hc71+8rs
ps9Dh8TIzIleaR1wmZzlXrLCWq/v+42CANpjihStSebAla1R0KDX57blptvUabJAxXCCVe2/X7nC
xkWlyNpLcqX7I08lhTufT9tJ1G2WQj1SBakWwV3FpYed5eBLIYwOQhMv55dHsBjbBYhpX33sGb3k
3adi5k+mnQDooPjNcxg13E4zA3DgMjmzJsYT+CAJvWs/NpjK8XzSqYVQeOF15Gm17AA+6Yl1HkC6
h2HxoVhy7i70rJdpXjpQeXShjJ4CFHmq3ARCB7yH29jVzKWsHOAi0AkDAokggL3/i9jgs8x4s/Kr
0HS4f7HHlnEKSVA+am342QsVIC8b2NIUPdqWgQ+cK1+l38fasX1X4mNAKBkLwIHAyyNFt+G2Vbd2
z38VuTjIR9zcVColL6+GP5PKiVz/SYomSpsqOwDDhs0xakGjVD7uTvgO2tfO9SNpDg8D/ZMLRXNc
yYL0dDnT0Pr9vF864RWTTkBZj7WA/vSRMWTiY8v2xDfcBpArFalf7A+Y5WA5x8AkHG0DBStm80VP
s8M5kxYW3A80IK3j2C+ew3jZDQWh/aHHWQE7stpgtNUMdbBarlJ+ZNyQ4ReqCBcPkwkVX6892g4A
WmkqReK60BwxjQ2irkQtiNSVp3FIXl2zYSDHwwWKoRlVvtrVKUsiOqy3WTgGUkKSUlt4HC8efJ35
ZCSqxKpJkeTMHAn0tiDI16so7ZEvrsHVlP9Z9eO6/85MgydUDkWy3PS7nHSwX3SSMD4g4C6hpiih
UddUFvg4Bq85UIw5Q9GaW12geH1wpK1bga1DagLX39HcrMUkCe2PBgtHFzCmBX9FMQZvUVmGeA7l
iIfOul+4QhU292M8hUyWM3OBlU2szbhrQL50ALr9sVY6Vh3OrTJRXud+bBTA8teBjnWx1UUlDncF
b3Q3zJEChu0GBiWeygD4AFTYATQFwn8YtutYV9eD9KDSK7mD6YTDp8QZQTrUv8K4aHLeFbw6SIz8
7rEWLq9AaP+IBNRTP/u07mLeink5UjLGi1t0S0dh7HnfOzQEjBx4CYCVL2FLQNfo04O0/yMSq+Ln
DAX+tcXFKALdTBifvb0C6gM+5vtYD/kBezgHxp+OWOswSU+9b1+t56OrKg8UsFSXgI9Frcq3BUbL
S+YTDgQRERy77/zexUSQZktK6GuuHNtNZnDl9fThnQxxw1ZnrysKRpMaf6bczJBvkNktakVE+KD/
iq7fm7/OUP2SL3VBeTMclomoAK6DPnMXGNAbPIGO0s0/ibDfn1cIW7u86d0jLHLUlUWDEmz+YjuH
Q8fVNRoTl8MnxM272q4g+J/r0kpFMM9lSqqWoiRfvPFD/kSy5hNre/V1QdVxsnCZaRdevO01zQIj
bu96yOWARUECCri974O+5PYkuhRvpz4Yu7QmZ2xI+TmKFC2joSkfKcernrlLpp+Z8lPlCtXJXp/L
0tyHfRdMXBMXPoj68gSjHH/nay7t3LC2RjJjaP9mEnQxC7UwN6sBe5hyXWJOQTcqmUBScDjmiZx9
Gqu1F7Fj6VTmpX+amY+G6c3dfNlFsVEjXn/fNp3HoPOX7XCf0ThNKmMjJyxqxVg3mA/0H5rMFOi7
JCSh2+hAK613MKiP7NslsuKHEh5pY9L+BekclRZIn0PzuTH71aRhgyGwgqkh21VEPS5mLfcVjlZa
3Krwpj/tB5XCU/RbBy3T5imVhiQj1j/BVzTk6atnqwDT9//JMuNChDfZFKHXnWCh17n1jNi+zTU4
mcC/e/RBS1VA2l/lswGD/ljl4ulLxPucP1L5+MXOh3AiPxFJ3VWBuXf+gOs+5TEJnlbMIhyDXNM1
MPsqoMPILsWUvVK+SBTRYastGVqSpBmQrH+ce8VF6iKrnPOktoVad9NvDtmmBLVF7AQ/bugL3Yx2
eGJXcMuPCQznKCgdIlyZLfAZbTkcSV4zhA8AG+XDIFLwmxmuEcm4joydi7sNb9XDRMhTR5nFsRxT
izOj47eWyzX8qJnXa7Wk4C4oSBvKjzoq/P6qUrAdZeOLr4UITsEytoCh0lo6MTfrFBF5YYPtdMrF
REQ4rAjUR1nnIsCySRUXRyG8h/TwuIt43HfRL+tf8VsB1GOP9RpBydX2zjk/9R1ktN5ty8dGM8yK
J87GdqBN8DAQkXsegnbaPxuXOPj2VtOIXZQxhtqrADoE81hzxyIQKPd2PTj1yXz69NI7sc/arBBV
iuRUNNOedlyDWKxpHRR2O3PNQXEvrwb4nocNxYPNEEe35I378Y5pW5dVmF5TU/qi+Sn1LDhWjQkY
6RMdwDP45G53ElHGH7L0DyGb7yyiPgdeTQmekRU1BfZLGgBGPX+hQqv3pjn4FzafdYisn5K86ZSJ
/TztOBM++7SGNIdcUwjB8acQ12D+n+iyxENgI4RoiPKkM49BzZVUL2cjQTpURYQvn+owEtloahXS
+t472SniXFr515KGDcGv1T006E3JVQcBkj7KwOjHBhOOfq/tOYk+rmrSteUcb7Cca1n5Yq2iLSp8
WAmTIHtghHws6Dw5V8Elq2RQgb87zJLOuHxzjzVDwU9NtR2QzjYcbGwrUMrhKeFi/FZHOJkh7ihf
rcjtBvJqZSORy2S56V/h/9lENcazHQCeFGVsJXGBi+ob0PP7Ta4tSZMiKAa2LWlo9u+62C8bm6jC
e4Fvc0R65FJfEumavOv62E2zRA9FQ4oUpZlBb4PqmtsR8TjDsGMtyMw5fzTVxFCWDQdWlhAGvd6T
a8A2FveZ8/qfVrlmlx0+BT//7sjWxXbZ5lt8OJNe72UwxkclxN70DxP7Hcj7TCBlCc6dq7uJM+U9
lcGjpe6a1t6YGtv58cKQR96JD0g9kn+xlHVS3L3h034/KMyes2yOcMYgJ/AEOosCYkWF1gdMzwIK
qiSM5l9OAmwfUzfo/3flPvJsK+ZASBvt8DzkFShEUwvWqp53CvyzSXKzh6rO+5VxCkDWSf9Yt6Mm
SVajfnCQdUtjSbbVf5Sa3iB8ZuQNjnTKtwXsZT0iqm0ClukbhEnVwOpp2tdDLOeExJcneEdVZxXn
gXaPhLmE7yt3+2ZgDyGFNo1CN9iSF+2dynDy/878HsFM+REwFpobSuTMaqgzGnKfci+QoMQFNXsg
PHjZIFXKDQAtpDCYTKEBWorgv4pNzK72hkJAFo60McFsMuZwNLoApIGnDzHJW4R5Zh19SguSFCEx
Cd4jrKwVXVDizrL2W7zMxpXqKTfehBT9GFZvfDBgWj00+hPAQFfCi2vw72EbvQ3OLyg9Xd72R+vI
V5Q3rzmx2ei413f68y6hr0aBV/bEjHD3ccWkHC50nEXSPfvA2bUtz5zGTZX/ZPXeiw7bgG138OdZ
eIKJix9aOyTrvTz7eIS9j03UfKlOruZQBzbn95gN2Q1/c+z3xaKBEhcm07sKNOgNRWnh5oWQ7EwZ
AlR0WFQnKxDo3WFSZZVV7WUDBclO96mfL06zqhmQTYv/p4EZ3+ke7QRgn41Pl+mO7cd2Y3pUrdIM
5gVwQko/5VKdzrLs8Bn7wa49FS2su7bIx2B+LasvbclxaC5D1GCzL/XsK3rvJyGqE8CrNOS38ifu
Hxdh/X0lwNVY2DgMhOGnrlSWduefBSVS4Q/FdSIN0SG79GvjtK23yZNsItmB+pyRhynlFonlLT7O
eEOiStuvJMjH0tHPPKN+8G/032QtHcoSYcfp/U+HlnpRyIG1CYG6I80kilSihaDIxOgER28wz7O9
SLDawv5msIAxn8QxxUterL6PVCSBVVj6JM+tCqzKMjb6QwLigQFyrMNzGgD5sxMiE4kKZoeY89nl
cm/cLN2igrI/Eukav3K492BF4D/w4GH3qX+3deS4IO8XUBkMk7ULUcc1fZ0H+Kcw/d7RseBV+Ff8
rlMC6qH4d8doLuKOztpRrjqhEH0nGISXA31NqMBj59TSQpIoRODvsh1I1huwPAzEZXRBFZNn++zk
pBHdetx+wmus6W1T6g+7QKYesrz+9H8XNmMJ3vaI5iDx/8sSEhkvWudH8edu5d1dGrovLCYAuS81
riv0x5wsuBNSVKepQf+38V8s9wgAdAgHP6igu3am/kl7ZroO3aRXYvToByAhid5XuPgPokih3uKC
R2+VacPgP0lBBuaKlAOBRnKiqh4IAoQXJ+PpTWminRK/+eEkve4/NUV1M/YqyW/PuTiCJFFjpc1g
aIhcp2cboY0fZl75CTX+ZdYgvmfA7+9yG+P5xyMRVC3WI3mmCTWBP7tpRrTAEG1l98I9KSfGAVv1
D6hwpcLFTKeH5VrYwVLSkfhvizPsd96ATOvGy3QR391Dg1jKDEo2OLqh+4MDjtvETxkRsH1MWwUi
vRc/umKlaCus7QHylDVpjOX4veBmawxTMgcWUDRHZ4mgkKbQp3bwmQdS/QJzibzlqbkGAcw0gZkO
qrRvaMsiKu0iqaqS0YvJ+oSDVPnYKDt/H9L1A7clfa4fJh7pF58fXlnoOWS/Q8gEolr+PDabsqOS
0mDF6b0l0+Q/wUSpKPJrk1s0x9+bVTpo61dLyh5AEDJRWJrVi48MpHeEvgdz4oBDPlQnOH95ok7h
d2smS5+w00kdFs5BT7DCfjCQMvnhvtHCDTw36SpV2UQ8z1w6+YHdgsYCXmT6ko2CtqZPYn9+R9Py
pPvqG98i5TOpzhhnJE//XtL+rSeRstl7QbeIgC1lV9Pu1KBO5DhVdoccJbS8rt7dyV3NPMYYhYjl
gW+cnicwrm6NiKrqNNoMKuxhLc75sdR/lxBXm3HOW5CcOd45BriTwlffnTHPU7PWJWIxHHzw/POc
r/AtxkBOTIe78oRbhf9JnpEtUDEirp8VwBPRR0nwohCli2gFkFzjIiolWFH73hHzmk/AYv7/xVEr
TmnLkeKic4HK72S5eSsNmv8EPf2k4oGDkao07f8g6v4n9cb/QKxWILHt9za4Jx16pkbS1XeDMzNE
nWiv2+h3C9k0q2uDWuVZc2kwGIh+rtTN0GY5swS9JgPHt/eHfm04WoZisr4+JmGzqWsMAsCPvcX4
PC3lXcM4twT3noOYlqk7/Y/qG041aJeEHqDbhYLhrWNAPazrIErJX2RoQl1ahpnk/8bfs93JhMWp
5vTKmWaOwUdwLYQurA2VCbtAxmshOcFyeTJyfruHfJWNOTLWDqF6/L9thSw+uTl0toUAnu4jtSv7
fCqK8ykgNR89toN/sOVNX5875XPJcLCISvZANOO5vxlXEvAPQQegatrPRO/9IKFpE1ukMk5IrFuy
UDxLJYDubTytLzFz7P+OciaXoJdfWFxrR7EKmjhqx02mthOZJkVQaPPupq/bp06nwx0x4v7Hvibq
hL6cp0y2HNYFujr1sOlyaxQqKIFe/d+4XUj8r28+RAt4amLVHMFBhLIm3zn3P1Yn7kculy/Vd7Dh
+Dy7Zu0YlGxUgGIeMWi3ywM26rEqYgv6ziQsHRoHy3xibEilzesZ/0Fp5hj5auJ5qBpw4Ows2qSR
74PYeb/3TyAlYFcmEOzpO2CfAVpQjj+odMDfqNM8qn++YvSbqThKws/aYGTk/O5rSm0eTWAhipav
zDBQTXr3eCbTrpE46AAZ0DD2bswb9vmwlmAqNlBM+5yjqF8atN/Lk/36MeCWFXn7fyXN636vnuB+
2oIuqck5cjeeomQlMvlEkH3TZeIRIa4K4rLTDpRCwLPOGDzjYOivwYefYa4Q75MRegyA4iRcqu+3
O+kjeb84n4Avcxfsvd3+VU698uOrYT+ZLg4w7cg9eu9KP02tDC44RQ1BZq7cOtn7qGlchYuE7s7g
CYlFQN9UqoKgYn2YF2w2GgWX17n4aVmkjXM3HA6ZnpeBclI93Ni6Posy4OlqQz9Z7AJTFzRrtcYA
a1riZld2JCekOTpZTqqmOPCXUFIpdlJ5Ytf70ZVXy8G+BVlnmdZzMXOyRrBGWX7xxmZJHVORXaoo
ucn6XZXakFXnj9t7vTXiV31Y+T6I/mk8V51lhdUmId7CqXZEqVurXNkpcxbK6IW0/56JzAlqLDrV
EqHqVDnZZnvCJg9anxGl+BSWvxiWYGhGJZXNIjI5pA/PgVyapu3mZ53eCvAELbG78vMk7OHm4CSC
UiQ4hJVuaFEGFTjdN3lxKW3heXYO9pq3/SYqwrydM3h2ax84T5TVlHeAcl+lYw0WxyTTjAny4Ubx
eYjPbuq1lDNoi8xUXezp2/VJwMLi13HwhZgr+GVJ9XN1suhp3pyhYN74W7PRhykJzxJ7i9wNWrO5
3vdeXc6AToKvSr5Cz/2RvPv3aF+fu0LQisOhsCpE8KP85XNXDQS9Kb2uee4ZJQM1dfxkPBCyfnHC
NMxPZ5c4YVP+AMma5gjK6t4ifRtOUHvECZaApaqfvm5UxWkLZWZEPmhs8URoPOXJy3DyZqTHOmwm
ichwQqsC6oWd0tjoBpMSfnk09i67nCKfVXhWW3sYEqrutyPv/rhOpSvemADmud0VeBBKhdK3jYwN
p+FvnMrdf1Cz/S65NZa/X5pES1DoEJj9q0C7W9KMa2j3k/YiY8eEdGmuv7BWccnc5NoQwpmaLkKZ
KgM/8UUqXtKNXit0AyxoRabHIoV/YUrxpXj0K3DS+bMbK4o8WejODm58QVmOUKun6epkXj0xx/6S
b7VhnmObgatxJ8lGS1vmVLeC96cyV3wcr++tKjAKOwduomcEZwUF7ON0IU96XdfraQOpoW8FNFlj
/FGVFff1Qv9Fdd0m3I6XZXpUep6/nXNFgJXYluGZsQn8Vn1pc9I1HDySkkNyGRiUWONne9zm+kyq
5hqI5vU9KNTbHwO5GyckaYHubaUQt+5rNgKXNVkjdxuInZ9pDlzkpvA24Nh9DL3UQiAMIFnSdUQ9
lzmz9OZh01Vdu0XxlDIioSCaC/t4U7Y8iuC5eCsJukFexoB0/liI8Gw4tFKz6ER+YOToNh19Ouit
a3w99uU7vF0kbWNxab1nyRHlWGkDdaNYiZ9DixU15F5ia5EkCvhf7fUuJTWEJ6MvzLj+mpUd7O36
9yWHuUNnvpRGE5Ul0rCbuA9mr0HWTjzlpAbSzLpTt/58vV3sQDpZ+qkKz1ZYg3MUQzHj/tiUToi4
C9woI5ZEazYZngeK1M1UjziPCzEWEU0csQ3+2IsLRWmRtST7qbVhn+3nL08bRGrE5eF2tp31vfbF
Q/eSl1Wi0gmV7X2WDUTD9H6n4ksHa2TE9f+0b0PJwQ6UuuyPWuc6gM1tj7IrGOgwa4kzYc/761zH
Z4waJeA8DGReCAQwnScC2O1yDy8pkNev2aLJuPUpHFl6ydPL1m9RgOxTYPqzJyL9EfZhIqN03X2y
TIgfLagWhCixP6wFAizuCC9EgazUL2dFdtNy/jrmAW3NOZHBD1fWKtwCIV3W9q1gAH+gXEEMUa3V
KPOog+X57qchg0pFIp1Plzye5qmuc2dv/1biVJrrjpDobD9a1rHT1rfDXUMmnAJo7LAxknt8uHy1
7d3hLSIrYI2wPS+PZ1j3cSAAtjiB31zwO/dQm1AvBbtALvDlKztDzoW2xPGcnalnLko+LIJchD14
LNB2z6XBy8cGqJYbBYOfBwSASx/JK+ZWx0ELglRu6+UmpEOF2jXfIe8CMha4XVp22uT0UTwljnnO
3U3tXuzkLqntY5Y6ZV0NyltTKctBcIJK804v4NU1Mi77ckA+CZcAWmYAx2leoLBaJA48ACqS2rxM
LS1zBfRqhfUkxiRwf+3nI1lZoN3rrS2KllKJ2c6Lrii25aMRGdOF4jTYLfkM/LZ/TUbebx2T16ZU
YhGNKoXwrDKioQZ1wK2Z7AsYGGgr5ROgfhX5WplrQk0kr7WZSe5hzVEhrdaiaycqx59bJo+Ojuas
l/aTeCZ75Mq6uDkKHmRs6XjY8ZBFpOriOVC0EVbvD8RyOR008AHan8J07ensno6aF6+zaZtjuNHU
XsGwnYb35R63FIPH9lRfLxd87W2nEQaACPDFRch0kFS2T2/BHmhiCodYt9B77QdMhXOZIXaF/oH8
fPXtAbLp5x92bXg493+RDNeIMPDplWBQBzVMkVbkXzO6OnMISFfpAj92RPjG38jyOwj24z/A7l6b
rsIgM/fAfDdRLkD9APTV0TkSxTGdCC8Fw55lTxz5cxOalQ1Km0SqS/GpU03UOlrhYxXUk02QQd0Z
MtxheklEjmDbjqYWv22yPcq1R6j02HRPpbjBSUT+e3Xtu1ad56MhpBNIoeA9aROaosLqaDnkHjeO
CC43Pzm8pEoX13Tn4MfUtzR4Zt3/pymC6kWTCzUwtxTPA7aNSIc0/Jidm1YVF3mwcwGnkFS7IEUT
m7vL5IZgu0nPIHTQssl1gngNAfwE4aEJnwJlzPVorF/enQqt9G8ihbyQgaMO7pwiAPu3fUNO1zNv
c1VMYumJwjCrEyoJ7JTvf7rtk0f15ev+pptHZOEmBBCecntF04Wsaw1d6uUr7xBHfGpLUtGkDldo
np04Xa1nf1QIRZLlODUG8IWEEnyKjanhdH1lTD1HhuVQ4X6L5UAwPFlyM9RflGU1fwJ00ZpcyamF
rA+qo/eYvSLhXS0qHAFhAiGS8i9C2yesBt7sj/0brs/rEY1Ko9Y/lje6y2dRbZPuoQCatUrSJMv1
lB73KT3uasSi4NAGAN0s/u6/K45MAQhL3Q+EtIanY2vEVjYjMNWt3X5EB5wDztfqGDX3ZiOq/uCC
JWJJMNPZyan4zIyEemlTlnKjCeXr2ssa/s6RwAtfMJl4LTMmswyCZrn9uMJPQHfh+6A0ApZ24I5y
pMjqqlYceuhVcWp7SlVYWkuUXCj/tAiy6waXW/YdooK3fH3TXqSZmYL7VwnFOgIOu7NGrnC4UcGP
98itTDftB6yRC/rgF8P2HYOxXGNP/Kb2xMZ8RcxnxC5e7CC68DLJ3vzhD67YSEOTkK6BQmi3KuBo
DYhgf/RlVhaS/HVAmLLB9hu5h1fUMGK35vI/KZvzW78ShNDV8ytcQZMtAZveVjFFEHXsvrXq3iRS
9JtaiNcQkpaxPa/8OfAkNrHC/CxK9nJGUITf1JlO1q1phGbAQVE1Lnw8yfbG2X4ppbBA80j47lMm
I9pSSwdxodwOAFmA4UXN4pSzfhNyloYC3itgjYWIDLUPsnP71+/HDfn06NGkeRGZNUpMxg7bpAKa
94JJXQcks03vKunL4EYlrMCiIcrbIwfNm6IpjmyYZWscyCum3Ei2obbKsABT02/4wFbgFmXM3wiu
JSh1q6rOs5spz4GfxRHwqHPfu8J0RbuUkNYA+uEN2v6Qidm4L1DmKszGnBnX/ZwiIQY2B4WpqLVq
zik39VHNwT/+BNKEle66FI12UyczqD8pF52enqKryY9wPAJYzrH0IgSBukEN2F968HPg+JKBKl7P
t8+bRNdeE/0dkupO9LQzCaJrtc8hAEkQ5pgModrQu84KaGgawqprvCokW8S52rdH4bgj13oaPeG8
phhpXT1FYAHT8cQkMU/cpumTIzJzybCZ2B15hYq9bG79jtN+jElDXcinrLw+skN6VuafrCeRYO6k
X3v4lXrjbsFrAR1sOd4CDJsa3gs8Ae0Rh56K2CxLWqhTpMc/iBNtPvLizZiBrqCRwpHmB8ysxa8B
4XA/fYFwJkgSJpMb4plda7hUlqqOJDeUWT2Rz49TuNLlhiHE2K8KWvX5VTeNoLME1PtPAvyPu7x8
K/mfAq2MC0TCudaOdIBLbUQ5U2EnPNCNxO6mJc2IGMyOfVz8lvyTazwEr1YM2Mik7Z7R7wPyUymN
AGkw5m2ulc/Wgaj3AXj4VQLAZ7TrGqazMrK/fUBdf0/tC1zY4mt38r7wxvGF9QZtOayLP96IIA3S
eak2v5n6OcGRkyRfhujg0WNGpg4oTSibSOoCZxgK7Wti9SQMJz8PVx2XIDWj5eWcy0PzVRn/Jzk9
ak5RXooQGjsl8MwRboXLoBJybHZeCsYUfLxaq7H6bMRnA/Gi0ty+/CWtON5heWH8ptICbas6x3uV
hWKHEdVNJUuLaUHmbdbOGMyR3z2t10/24AjIJe9kcGr0vH2Y/NC3mg5EE4avE8wmeKpC4Cp8DhIl
adhQmPVvhJJ0PQWEbFtAe7AdrCGZ1slB54ouB3KU54DuaY8GbUGBMh8m3Cfh94OgAN+uLZbKd5q1
vrG67jwQRCQ9+KR6Lm9TglsquH+t8bfAQWu+i02Az2bW5NNWUyP2Uqqu/w+Ttzxwxysk6SnNZ6KP
YD3DNnuYSDIaX1fqrRPv0LFk+Z4ckAuor73w38YIL5dcUVJhWG0FYKTDftx30XIkrbujfixcO6/X
85wMVD7gWm/YA00RRMbdJpRtSGjS+twTRQ8hgzoXKqn3sZz+8lwQaC+0/zUne44NGVZi6UFSccJv
9IYvCqvZCQ4Li2R/JwIjgLsFP/5iqtdX0L4zOhZJMZ/2tRqAFBBVhr2cj03GRcF4tBWQEn3zhrNN
lzYD6uth15mejItWehjyG9TYJ649i4GuXYNp7MUhQV8xR4crG5sAS7IgOA+qHtunpUFi9W5zRNRB
Qh5Kq/mhF3GTCqWBCFtqUEZJ6IkkeHHjpqsecHWB1iP1BtYfx4pzKzFkVPlkw09oE0XTdZ8BeX9y
kA0krGNnlwGrrKW9IfIy2xABjiIb+3yRuXDRazP2LB0vFqW/Qgm9etgFGw8nqy/eg0b+xVLpSGul
wlvwxTpg2ofQm/ivab6vC9xExSj//xcY5KltDkVjDbNZP+cJMjGQ24s0CRr8AeixDoKUm6r45PdT
k4o2CqRxBP4lOn9hUrL/6TcHIGGB2mURhGzYNIf3XidSvzw1mJ/B/yt0BiFKSsUmXAEbBYjE4jYd
5/hqZ9cQz8SMiQ4olvdKvV0+hcsjtyIUdV2N+Y0kcsh0KUGFsUSLChsf699X48CeMsLQ5Jt3AZCE
UCuZkCBq8LgxROUrx2pBB+iERMUx8LpvDaW3XlBsZw+THv3SZW3zQoEnXIGoRAMRYieNW+iKCxQh
tqYkkfujo5Jk9ZYn8igRw2eDM07qW8nsi+67eHvQ5Y3dJCrmv9GxSO3xBf3LbuVsY2FWAU8jtrY3
4L2JyBTYxImnUbDPfYmh2ZfLomFlxntgyL5odxoBsKhKFAYgPe7iqoKa+7CAStwAUbCNSkXiV9/h
oWcTms4rHSKdIFy8533GIp59xxprKGOOyK3chymVdxTXXWXVRnGYx6NqjwQXRznPPjfpBTS7Ni8N
Wg5JVz+iYQXyRAylFHjzA46TlnJmIVfZxg6VMszY2a2BFFz5iFGphXmPQ9JLtrTH9TVfx690MB9l
l7ZZhiuXlfy5W+L5gdu/LgKXEDxs7i5htQeHptm8hh1Ol1As5jJD7wkh/hANv2uPcWrBnvUBTcWB
MmjkBT1mMHvJ5ulHlTTqb7V+x04FHgCNLtd0jNX/H0QuLBOvzNxbRoJcMU7QrgGzJFabkaE+Eqte
AM80ZZX+7A/XH4L3jbvwrHdt7n7e9Lv+9JTq85v0G6lZo5IlPKYO+GoQkBClzTGa++RxKQszZ+Of
ibp2W1wioBP8wgq3Ro66g79nDXEb3tV3/uLoKgfBhmQFyFxy08IJXE0b3Xa17v9ZbpgUyAX8Nx0Z
bvp6AX5xvheM/rycfV7G2v5/FdPObZWcvgESKKIBbGBHokPBcNFd78OtTG2bqIVhMMGZx57lcFA3
dQtRUONvagV4VLYDIERMU48/9kE5ZyYf2FsoRrO64RSq+pBvaGs521wjYj02Fhzkr3ovw3L32Tat
rRWk3EZfydaqYYFaqdR/NlUC+GPH39RyTMLv/t4ec1+AIpw7HTLPMIT+5+pMSjcN6gkwzp7H+OSx
sBSLjdR5Mh2fb8sgtnVw9KnMomJzNs97KIcYOwdXilqS3qOV6goCpoBQ5VnljmU0n5TdJMXUI2cb
shvQZ4st1g1ZGauhmW5dvxUxGqA5F9RIO25gMrz2srVN09y2lR39nh5i1e1nuAj1JoxA7HVr7p4c
qLCPKbXu/TQekMscx1drNzv1i5QUp0OkQedBNFQ0MvT2StyPKHel6GMqxODuCOKq1YaRkqMuaPzs
4Qt2rdUUchIhTAsnRWU21VE2zN5YBFJJCSbk9NedNwsuQAycszRmNfyImzEp81qGHvCxRUWD3RF7
8b4jQgGzeTCAVV/7Tcltkpu+Q7ztlh9obW92mrNkBD0GpeZskgT4+3QM9emb03qAIPvSRHYqfRCM
oegjgIPj/WMOjjRunLaC5wr8Og4jRNzRITjH7t6JVWv4cJXoeFytJOfTRrZUhYLizio7R2JZfEaf
mP/xH/S3CT+Q5rQrPUYKj/ZEmujky+tiY4LBJM7L/SgnXJl5gdWbEjADRbHznGheqAyGP2bYWefi
CC7EbbXblONORw+Y8gA2wimamliZtHk7KKeuMUIRdA0+N4Fns9OMaGlAg1boKs/UwrlzwyaJ/xd4
jdzJI3F1KmsBAnp6slsC7Cckf7fE9658800UebMhmP6Utw+WBQtGpaTKj5tGwCoenm7zB56zfRtf
YP7WmC55wKiC7FGL5Y20mIQ3ynxxyqLFVvghdIlqfEBPy7uk/6aefWLXFSHL6jdp1XACrVMLcajM
SeQYK39980GnwOxD8dtXn39is87ncdRkPrMSlGDaHSQN+yHLykH4p7d1EryepmlPDvJ3YMtIKQlQ
8YklUDBjM9mDLkdYdMfhH8p0h7KGG+kED3LNlti1xq4zxnNaywc7QHejgDdXPmu2vRLOx6B06spJ
c6cGPWG9TlFCTYKT/GpBoJjJ5Mkuo/ETP3P6ZOeeUKiT9ya9FzYYNzaRkDI3xv/EPvLjs4Jff5D+
PrTaG4yU5jcEnurCgdA/GiR97XE8lMXKjDZfdvHQdAn6yLEXaXvmEJMq2gl1OvHhUZvbi/IPuHw2
rwmaZ0TvqSHVHKFPm3RCsLQGgqMXWvVVQ9xn58l9QVgxrP/a24VJTgJBG+09n8wY6+eEuJ/2w9Zm
YnLz1CkRfs21CH/O5lKiPEk9sFAOu3vu6xyuptUTxS03u0LpDPi8qRSVyVYlG7iKprAAbW0WJET5
iqKU3fxB0tcBeP6ycEo8uD7cUqopeqJMOzKwUgxo4gS/goGrlHuy4ow0+31am/rVUBobQd5jBFwn
kCPNhhciFyD3fGx73MA4VNBK0JAFR9BWA43kPXHNQr1Jd+XwH2c8B0B7td1ugrs/GuQjDQTuFySD
HkRdWh6j+XFBC4+DzKFJ5kP18crutuZbTRtugEtifhsTw/fufW153k3CEysEBJsRCAWRpqLyviOV
/AsDQUh6VNzZVY2U1dqUHejOfntWZOJ8AkI7VcRlYBHD/mWpM/I7JWuEKudLU9uJxoTZvfQqp4xG
XC+v+KUmjkaAaxpoFag14NC+acJQUcAnSqyJPuU0HNWNeoYRyjtXloktdYXhQ+z8E6JeLkc8n4Xm
DOoIwhVstt9NpWDfGBdNdvRlmey1CcP64/UYR2gcgetcQqHXkwiljyu28aJ2kGhioPyv9v7ex3H3
vR/NTRq5/FsNYueP3UX0LT10H9Tby0RnDGhUHHNifcaMVJUqzbchmFFCPOquelz6lW6Ch6DUPy13
QUvxrufGWpPj6jliK9ICn+lcO+FhiX7s/OaorKiKopT5xKflOPfX92pjhpnQ4l1DAMre5h4i++2Z
/OpskooK8DZkvxH7sEDmJ5DBCPHlAeXiTwfT7RvVoGxY4dcDZYDkKyDUtKO3h8Cz6SdnlTFIWEXY
NxT3q/TMBhpnBF+B1T6zWkuC4qfLR7XhS+Z5Y0uG8dOSCNRT0SpLmwUtpVX9VVPDu7J0oT9+Xs9P
8oG+GqU1pBaGb+JOUB6x/spbFOWU0KIDsrpNDrB7ki23dzJm+I8pBBe9StUVePdufIsY9kMlzRB5
MzcD/HyjIvqdID/U/ZeGBnMyOiMb+3dhIr1QhwlBOxRqGAIcxENCpIxVP6J/rtnxn4Ub3FZxcmOW
BaOXUjAYAxJsqYXQvwuY0BXaTdqMRW8h+TcDs5iTQVgLud1POcbkgprC9NrC3MMEGCUY2bbi17Lq
LtQXVOklN46L7Y5FIniWudK/1NLM4mMP9O8AmYp5LhLnc3VvBlv8Pni8pFP9ioEcC7jrXHzJOpdB
tk7oUUyW7awgHAanAxsGgA9eIMKleBOegi1fzUNnPv84A1rTDkaS67+N7Sd6NdWm5wce/AhsIeqE
6PGMpPwDLexuPvfR4Q+djuialZ5SGvoei3lmb6nK3NNrNSngit81ChlOV7nR7+XJZdvv5jqgeTiO
rODVtfKLsT76rekoVtInUfrMpjB0r1NGg8fp///fSNfO8AXkrz+w1A+ZZQa9zL7XV7jaBd8MRISI
mCQeh8m+yfx+t/DvYFPmhBtyeMuSgiEnXHDL5aSGyq+kQ2C9gWix2jal+22oBDs8ffu1ikd5zz8/
3t4f4Bgnpk3VOsVQlvAf0e/RJUqUdTFZ6Cyi7pvg6Ja9fIhbv4x0WNLScfFNQswdMyOWl2x1VcbJ
ZIBIjSzC0O2kW7nc2LoLI4a+a2DL/79uErL48KioQX80EjhPxqNhPAAL2QCOQiiKuioVHjnDgAFX
GVIa1o1EGqnnNh1UmTMMh0/tLFW2+hkPldgckQVJM7rbFHuRojRYVekQABdKLqUn59t22FGbestf
1Bv2TO4H8dIy+megvBZWfSUdjBVHHwDwS385e/IDdq/EABhL13XK0X5lR712OWLj0OO4BZvZmi9k
gfi0mQvoD1XJrHr9qEaX90I9rISmrj3PESMvJK6u27CmKGoDyzTgpNGUdnBtrARH/z/geQhlATwj
qxhi+BBTB8lrjGT/O9/zMQ3Ymqq27MyqRpPDI1twGSbI5Gt39jPFP2ajUO9w6QKd33bDjmw7ZR4M
tPNjpTnLhI1MiGVolTkpV6DJNnpRhCJK0Lkcx0BvLIgKutwXQdBUo6XXeCO1t/XmCgypRWRo3bJL
q16cu0D5CpiY1k+nRr5ea/Ah7J3MBK4DzhQzesUoowi1MgPPoILHN/pX8GGKkF33T2pUa7ZCy/uB
cBwLDWlM9osidb3EZ7XYY5hJDQdU9UQ/Ps+gN8OolcooXwAM56a5VOcHfZri+z2Zt0X/jXZOst4h
4Ei90BEsr8/lZpnJ2Eo23QSLsUqHP+/qE2GeQ/ansmTaMlbBPVic/neP8fAiIsr+a0jArLfgoAw2
gA3j2hEkcj30/wEv24DRlGH3yYjgrQ9xC1ZfUdaHdN+w4jW/HxcfJjCkvyU/CtaLPgJ+hdozXdFu
070xReq6LNyMwMDCU7i5AHLb1Z0C1wHvzIsZ/yb7mvWp0KlDczUhN3aGLcpk48dm8UgdnXleKNd7
UEFbY33xu12W3AM2lXKCsywnHsEVIHCgRLSgjYjj7ay1c+Wcbm3MU6ILhNVSDSAmKrqR0ezHndQr
vn2WM9Ze7KHUPhCoorlEkKxqkfFJ26X+TM1pjC8BUcwkHv3D7StFRxQNOhFbs4HWXQ8h8r/NiXDA
3OYqXdrM3O7KLORmpr3e+WvFkuTkoFmFXQvqpabOP9aUtb0WixNyoZkjWpiI3MFn8I7X0Usm9rAT
wDa7fxQXR/JfYCjUBqnv5kKpdheNa6llPc54ap6AwQNbHeg9Argqv+nMsCSrWsob2O95h4xZIsw/
5lHDKDeqNAYIiqlBK1eatFXtPDJr+EazbKdz+yeWpZp3+ILFQw948mvBipvmL16Jv7gVx+Uoj18M
86X9J6xKpMP1s9SHPRKnTFM5w1jKfEv8eMLYLo1Nf+1Q7a3AoqwkmmqiOcqfAb8SThtbL5Z8x6rw
qe5zPo8VfYxGGqp/3/0PItU/VhGp0C/c6QugCGq5Nt3aSuAr4L7RnX5ROSxhq2IrNoCmIFu9CtVw
0WRmy70Nf6VsP9L8jFcbkGDC1rGzCXHwQLS8kCZgebvdgIrW5NYC2x5wyHbNmdrLQKyYyllusJA8
YYZzS1k+/Owc4/z/os/2aDzbXFWO2T+pdUPDAQEI4JSXyJx3rgXQaRst0VtBsxErztIGQA2aX1Qq
LXVDU2pfra46dh1t71HGKjCTjaa4sISw1NF7FnycEuLjKVJtd5lxVqFgXz0w2L57/Itz22IOOPra
b67dBIK0EK9T91Q4+CsMHCfVXTfazjDeF6N3J85Als3tTppGKCvSiic+lS8bh6w+L5R5IhjMD7XP
3IE2KTAuL4QKuxCqJ/TbIbKCY0zg367a3jRGw4Xbwdpb82dYjSvX6Bq4/btz1kseMBmauCMlu8SA
xUHzLmRkorMGtGh+b8IP+aQb9dnQiHZkWzWl5UryjfFxRGdcuAI4oTvrWRf0PjJYT+UGFpCaxv43
IVmx6qv1IUHr4FVaDw8yKcBD04PzGKJo31NMWBhhegMvvWdtg2/ntXMaVlcJRzGuiGbsEASasRCH
A/Aige2oHm64OI2PuPMO27oyrTKjBDeMAZHhnoLTHaXKu2sDDZMkQek7YI2fAn8PuXwW9ybvWklZ
tVuIQnELz4H5wmZSiViGQycn0gF9VaBC3PrtcJEbvnSC4g9vZP4P0liOViPLbkAue+zjW8WyRXf6
uJNPvE4AIUd0tritptjXgbo2X8K0fsPueHLdpULYwn9ve9yp6fY54oSCglQOCMYHWmb2GFDZRs/J
5yeK2EICUsf3lPOV2EF4jfTo4CrcBJqNb26+3aLTEQD+FT/lM6RV7Y+o5UEICOB8DvXu7d7PjvHS
IuBRGxYNTFM4vvJNFdZiPMW2A4kN6m28oyboqGZNqd56bSsvL9eZHCvMpgP9wOZ0svn6L8DULoo+
r00NHVTkwhNMD/wGnAuKySncVFBXc6I4Tpfvu8vTKwC9/C1JVjloT1UuxJIm01t9QQ3nU8HqNHIE
B85KkG1Sg4UWHz3TWUFYX11Yxo/iQ94IbKE+DSCzE7ApTr8VylrD3P1Q+YxaQuv09x2m1eJ3z9zk
V7aLLqZ1V2+dT7NvPT1Pl4JjUblMqfumTD+V6uiWsbpA8iNhafrwgQo06TipyEGMNhu9a20f5Mu6
lswl/JlNLX9AAnCpMEjht7cGQB7pSou7z8oyadbnDeMK6e8o9irfKwqiFZ8xairlUHJ1yoGwTYff
FlBO8lGyxufkpuXM04lFMglRtP1yhXOaMJ7moHDpFt+3YkbYKRaUkuPmGvlVMZ87CjAcLvStzsBV
RNneNY2Xg9+WMRt5K/1v8BD0MgDslTVnRlj39sPdEjN6vFjC8gheUCNXakIgIoEEL5wIxQN5bLvF
81qkuQJYlz5G/UA9PBYZq50jV8rYCQ4Ws7iFwlh7KxFgQNmcbNH5xrT2cNZIUnOVMs8SnqPhQZm/
zRDRoFEd5VDPcG4FhdjcHh2fMcTzI5U/+ee4HaF6Bc3XmmfdrLps8YR8RIoBjiv86/+WQlAxf+Jk
/e2iQ3a5qMk4XMtVe8508Rv2uF0pthb3WrEmu/y8aFJbTfaMMTZdpDU3T90h0O/eB5ClXCi+FRLI
DJWTRXHO6kjpJ4MXqcNjykoq+mQvC0tU9yi0jwr7Kz3S1fnj04jPxRkE34/2Cuje7VBH46l3otbJ
0imNVwhigtO1DV+9w+cwCTz9b+tiHUCdgg9JrjI3MNVZwtNCoTlUcRuPGNgq+Rag0SqNZN/s2H+h
4RTDxqdlpFQiK6kLAgn1GQW4+apQp6Ej7dXS7toQhsBZEqlt3qlQz8uASYrsAyGsDqQMVJtrgJXa
vAvOC0t8KhHPpVl+IV1v4FUwxRCjoZAckNLsmzx6vD4R0u1qNbXhfcjhs0jq/72aUKCr8QHSurWN
y5iooU6nC8ia8yJgHY7B1dk2dW7UHYPzx/pOsnuhPbz5aE5PKckiEfzaRt5LOasBMRQYv3EqGPqa
vj6HnZs7uIbL+wVt//Gm47qiKlhomjkx7DfvXFG/Zagkyp3SoFEdAd8vsghKRh8waF1l7G3p9zZ2
+csj0o7g3oPcfqmcJxdnXuiOGXaFn7U10ldRJ+8kun31omgW7PwvzqPk5Qi2wX9o9fXgOed0jqdJ
N31W/X/uBy2qfmXbL0sfO93OZT9MknUCTWTnRS2fSUjdscyGWNJHmRVQrzHlvxz5BLHiQ2BOptO0
DC2snQTEHgTOybghw97+8m0KcHIHNCNE0+vQoDd9AiWAQSSX012+eD828Hc17fkDzV+zfnGE3UDr
UKFMYTAYecDFhSfkPt0iJrJSPivjgQHbumtLzhkN0unRprVpawJ0vEkZ37on8TPEfxlCptZlWnLn
kOb2dzEsvV0Ma3xaMWXHlscJKcO1DXkV8Mhmpy6AKVM7OeC4AWcdkNSE3HzkhFLBGauh9tqU8T3l
CubomnjfRCrMBXVtmJJ7SbXO167Dz9DnG+2roDr/gJbzL4gIywe1i3tenL7CxzIlEd0F3zVtzXNd
Re1w+1QEsGfZQU6fIOnIPI3tZF4S6VhlQcr3X5K9+Uq79soVZLGh9xmtJTWESX6kxskrgKRDtAQN
lZv5ntjTtsEuvl5gPacoRdP5soWBwW8T/uSYAU4If3WgQ/RieYzbYCqi1rTVW4Xme92jBiIs9RA0
VRWmlHtHziQGX8YzOBAUeIQiHThhvbLNudz0akzvdJjaJhHgIc5aE2+aMxXJVnMAg3p0jZKWHnso
Ts+y6KNjcCo78fHXvf71bzV8nV3yuyEWDDIyaP9lU+koELAFnvFq02/rfEWvDgfP6dKk7hJXv1Es
tWkFeDZBXokepSufbxOAG70I12nVOoznYuh0uWPaA/p5kxSbzvxuqA+lh9tqbjFpc0AgQd9S4lp3
7+MhGgpUbU1TNjou28WFAnKqmDDtXuZfaMeZDOEVc2S3eWdcGALpHHWktdd2Ubvs7yknVnlWwKoN
e8XKCM9eBAbLC4HsTfymX1O9VRCLUiD448azE5RnRaTiRzn/fc0dGTJEAs2Mc79PI8bjrglCIiBB
A9vY1+3vuHPLIAa+7XtTZwERuXylDhBXDoJIcytjdthsmerHfTxoF2zj+v2vPoxc9TjJ3X90NCaw
33yZ4QYaaEeil9EbjRglGrwoblhno5kDxOMMdv93HrYsf1BMP4P9itwTgwq8nEH8ecmDbc5mzGYR
rX8gv2n4fBr/hi/oppJOIUJgy/XI/BzDhc3xbfef3+fimooWfMKCObbjwLY2LhVh7wMYPRLP7Lud
fSsZVsuqGpcyD2XGvIzbVuKPE5kh/BOwb7gRdyLXWa2s1gdRF0gY24H+Xzm/+YKwkxmuRqa7Mu7C
g0QvI4s+XjZtPfKW5cKGogeEM/eYjvGufayH2RK4C6ZWIZdlFAbjNk+fZvZqFnM/5Gd2XJuIa7oS
6oioePG95OcFvtD23Hoq86eDAu6f4uWuRBHDRLYRSyxtQ5h+U9qq6/4wt66OTiLyREqrOgMXzWpx
eD0/myJW3c457Sp71KQbd0MKyz1aDkRPTtalZWA+3v3/Z72LAuqcZ7fiRQzr5i/bJs7moQiJUfTU
F7PdNbBB85uQn0LP2QWakCOvb2rV+m8mDwCaikXMiUyeydpiFMavt0zDPGARizdO4sgTbuTpyEzA
EvHusrfJcT3vnulCbWai+vEIq7lvf3DGWTFI5aeF7jQd9FPVD8xPoZKFkOxPBOHIi5a2CJ1zXVgi
NH6RffUnjRE/7mR0BZLYnxUAYu6PqP+V8JMngc3pnZuTKDwgQ8Zg7wpMa4P0wJNiDVSSwwxM2lm3
KXJx1hTiCY0PdnkFuDvfUj5VK8tSx3neemqpMYh7W8T9Z2wj297lI7N8+CpixMxccMcyb1d8fBXF
3iGkSVGjrdbkOEL7iS5TsWTb8RRIpUSTFGUsyNFK848Yb2hWR7m4PqW5DIaVv5tnS8pVrTH2u6HI
NInYLXscDBGaJWofp9MOSS6atCEExX+nN7R1tW1HtEBGbuCNnBX3vXbElEgu4xCokt+sbI/09aF8
6fxP2AXaPXNJupwtELvDbgDvD4VIEiw25IbCbMAezFWhY0B5Fzd2oMLhp4d01wMa3m7pdAGOL4S6
jU2nlIAQlxbZs5LRa+oFN/apOj6Kk2tWCAnT8cz5YXSMuH7F+LmOLr97sSVGV/rahk2+epqkcH6I
I3AdYuU8aFix2FaOrUOTV6uB2XoYtN+1cy8k10QHBSB6WlFVfs+mpZlBdcLcKIawir7pqTCzJz3Q
IlzoIu+LbTeUgtOK1/346qCMLDrBpXeWifCaEsUfYEGve6HsXjy8h1aI1vi+yeGTZFCqpIeTp9e5
1lv/vKEUCW3dc+tm3X9MkvrCZXE6Qi9mUKEfl0L3bB732SjZ6Givuec+aB8rImVdIZCE/2DZt31D
Z3dWV/L6yIyB07nRLZ4kzmhEnb8RaMxP61RrJoGcOaatelm62ryqcJ6yxDVlwU39Flrj3Zs582Rt
MMsBFVYnpQWYldyNBNAU9ARlxVq55OxsulotkNt1VrfwCIWpfEIdePy8e96f+k74/7Tgff9a0FsD
E62A+25t22BXkFEZ/WcbXPI3TKyaiv0bMjcAtjV2Rk2qvrcZN6k5/guXi8B2zZSr0i9JcKFG+YB0
lZYES2z6J6YW/bW6SKodh0FAm08yXj6IP6b/bdodn+yPgcIbmoIHXrCnzBFUCyE8XNbRCmtBteFb
yBbVI6QTkmsKs54zuMPMK2n2BMLtEyUV4ds5YYIPHdDANmY70k/aW0mn9tXBHhQyz6HfSG7UmwPS
jsXZEaq8Eim5xBNcht0Y4QaHTkPqn8aZGN+SkVdjGUGBSVsEzGso2sA3x5jHjmEI2dxgOxy6xsmg
DOCjXqC/S/4tI0H+Pigz05Z6YJ0ZppOQHiPO1PrQYN+sLX6S56sSNvZP/GnBjpn1++LYRY5HFULh
TwXV17lzCq3/ezn91rRtaYqryvGdBv2JB8nauvjga1Yhx6cQAbqVsAvUi3or6HGP943Kq8bhzgKZ
C7DYoffn48SOAdimJxf3KmHA2lJY1d9gbOnSvLH/3DDQ1p4kmr75Fk996xRAVSxdrOg4Nhs8opi+
3qBoHdmRL30J/7um0qUD8XKtZceBsYKBSUC1z3iamtlC8bzGxFCLUgSCJeeKCAVWAfKgXZpZL99R
jRD+L8EMlwLXdEGxYfKqJ+ZrFlgW1rQQEKe7CV3Vxu53QUv6239ONACZ7BaGKOKLNOdEQ52sPQxY
/LNm8DV/cIk6szV7lEouq48jTwEYUbgag0nDE+5E+NU+fQPv+aeiwP1fMAmGXLRgq88DHyoGTI9E
B16kzv8zkTVjP1lNOUEf+oOUTizFtKveidABqtdFpnLE4W9U6yGdaaCuF9AYATmPpiJAHsbNFaRV
ynJXVbzuLLRmyqukdWD4bCfsAX9SrgXbuieCpePd1Y89h0mkeYDueJam+8xeTEpYYcgkmw9DF5wm
pYgA0GZP+EYENXLbxEiBjjRsjvpom/ffjoeysu88YWVt4zF3FHvGrmiP1Rq52CmB0GyiYyo1sdIK
pP/AFRaxagYwPgvMoj6uYuSDuV2vU6eMJNo0ZSBJgfHGu7U27RqGZpBTHG5sKZXfXaHMaoL+6abN
ed8DxUQNXtOK2nn0rqMRs2OpT5mzPj+ewiG4tFbobyTwGnqP0//xdY7iUpl7d0U57t/UMIxrruJ5
w0of/WNX8mFQ6GuIFvFNgcjxHNmmbB0KGJeg6lnmere7OzR6/mSNVeVVW24OtKfAzwd83AuEi8W/
a4cFHjdQ/wxN+OTzZTgP+6z1W069flhrH38mExe6wpg3UfcIv+kz052jQip6MeXR+rkYgiA1zUy8
tgz/16RLIatonJOfp7OHTiyOK3ZNsiB+ZgZu/TOA8rMddzvngCjaNjo38xN7YPkgHPseJgVDmF4T
tblOh+aGdCiDZQzuJA+vca2mf2bFPNica6RB9c7fDIIX/bA2Rq/j7BGVukjpbUeem5CR9RZTrUtw
fTV+58QPEscrXyf1la0jpeW/KB1O7yal6CV50XgaWcPJCgWWhAV3MjZb7lanJHgAMOJ/AWv73M7z
WzGT+BIN4IIjcDB+1gG4oTihNUAgdxiNDayU4JUyGGNtj+ly0Ba0sHFxFsMGmgq2CqOs1jPv2bvz
QCKjgQoJYkvjXyN1UKRT1IXL6ta32VCXcQV7ja4eY51FcZztEwXO8Tx2OhgNMzagyGtJIp8V5FMy
9c5VaH0Pzz6Ia4/HkVg/5uRPke9bjkKN4SKXhiRwnHxyBSS6QCOCpvzDwDLHGZupA725/rI8UGVn
6rcAN++1jDWTGIyuo/AH3MEPkwoCWiJMqfaO4culDJ4zsoh2TD87So9qMT6gXS/VMsNyPiIHGJ2m
YjPoRzQGXj/JuGGFu3gEBmiV4tYqjazaPZcMPI+JkRN3lnT+13rqd3c4fEG69D8PnZaJlhzhVOPS
EHL00BZM7imFaW5FSunotLK3lSZFr8P51USzK5nkHPqZEBf5IaZ56n/FmNGwmmbYPIDljis14JII
uS6L5ahm2RiDM7h9AINHLGJOinGmpSWvp6U9aJ1HWHOS+S47Gq6kEUsNVjVVnDNQUfU5wE0YZAWx
SFcLB1oneGBaOOYUmOP+9tr8nXMbqH8lbMfNMZX8fMNA3xcPCbLDbn+gyIAjs7Dca6K1e1Pyggp5
20y3pHCz0i6mgMkfLm4l8EwJs9ZGgww9XmGpIrveeVhNUCGHP12YqNd42H/ummvQDnTtCyfN5I7r
sEpwNfh912UHQ3KD0/SXCEB3V9xq5TFOlEQVhiykoBLRxT30ArrCnt4sbUfNIPsicBYOXLcTeyYW
eq4hX9V144F4YdDqEtPDuTnKL5JDDjbNzdcOBLl0lk06We8/9LuUI2nGfieTkY0F30u3bPPDt89h
HgKe9XEhZq7uvwfA1Xk2IXnNpDmdjwYsO2mOPH77dtUfDf3LhTxiO0JXZu2XT87ktu0MHP+1n49U
kpMp7QyliJbGBXh5Ak/KubkIZDqSQpdaY4kEXfGlWpt/BjFofQGeGtY2M7yRFFdMDtHmNVznEGff
Pad/kUcyGcETJ/CFt7f718lP5R7K65iiiuhcsNepUJnQAi1c5MarN5/rWYaXcq+E5pJNS9lqNdKg
3LQGonfBLp2VaPebWrqrGNmv/gbcXzY2ki5vvoHcnY/6n71DNOYJwBvKplDhJ6qFMFEqHKKpdPI6
zSFql4Clm2hO+HVW7rfj5zTFs4nOvR7X4l51ePN0zoiV7jX66aKEKCMG42yht58ORkf/jV+4jaXt
qSENBm6D0oyCJYMv09yjJZrttSHqpGQ8zw3H2CVDZ2QohOeXKlaeugqMKvXWPS463dj2tz6c4Edv
UfKtROP+kKDwq0LNEHE4X+HCiA94D4m4MIQAxXGlvR8Dm86jWCuJQxY7Ijjp2GfBWQ8b5eQDByFI
W0p9D04wT8dTuCff7vE27nsi6TkNjr1Zl6zZ0wdG9pM6V058RS/FE2dZVnX3/xJ7KwjTf0VtdkhY
rWwShYxFTqdtP0D9qBLhRv/cx8tOe69DSCSdvQsDctuDWXihlYECFc9+85NoTn2osCM5kswogHVM
nlfQFC6L1PS92YSQzthAdEeeFcMFqbqhRfNYpC0IFs4TKf0/OinwqQ3yCjaAFKWA34roEZbJ1bPO
hXOUdYQigv+CyoTv8Wg0EzAi0JxBVKgaMvI0k1eEFjN2smIY/YUgFBHNgSSvcKFVc14ORgZxNNDi
TB0CihgyPynNecSeGmZZwB15HCmj2BDe2t2cQ1e+6KzdEXfIMQNmQAZ7GULAzIAXBE7E5c/0x0S6
Thpz7N9TFCWu+DZBt7rsPhAfaGF7/xHXe8BPpXlZIMm7373OYbZ12OKkB2DGZ/OCleoB8Ek00Z94
TguR6dhoZfmxMLe5bP3iadSRFXiTvzIAEUhnxg5kv3Y6nGVDoNkvJsg7qAEp11Uh469ArKoFccEE
lc3YIxhGw4KydbxxXpCn0ZgcAz8UUZGBvmv3+rVPIJv/7o8Er+KgVms2siXlwDsDJASunzHMRhEa
d2ckRs1js2QGRob0F4EJUyBs6f4n7QZkPCGCwNPWq/qNPkzOmCApfVCsjRmEQpaH2x2+M/J+e0eS
jyCYke6aouY9ErWk0T1fJEVVyhSNT5Kt8s3GoAM7gSH7xp2U7ut0NEaBcmh/lFs9dFktQ1FkmJys
cTVY2O/LMOuz5MqGKJHp+ob8qE3r0fwWbdX84l6WmYbCU6YTHUCxR7JG2R511khn+g1RL7/qAb2Y
WEZEJdfNxiWH+TcPMg43xV52wSsMRp5GqsX4Ol2g7PB0J9FsqTNS5sA+HwAxN0T7ookElLLdXZq3
Q94jKZjt6BL22Ja7PI3Xsb1ScG4C1EiRmcS2/utkxMLFh0uC0sXK+KFQGFJ8kbK9mUiDnI6q7qzM
S63oAUbLYoGrPSyB79DFFkLuYw9P9tlhtsqMRwswNLnqVX/Ceq5O+zwrVYd/+dUW+rQkNsBUr7W3
xZOCv77l0jGNdmHBcNGyF/s9TNnVfe0TVU6fxXe9nD8olR6KJR6X7u7nP3GutjBBGV/uZQ5l1KyM
7u4GGqkyFB4nEZlGVgZSB1OllUesZVy+8846azSUJd7fVA5TtaZC7AFG9PXqeDyNORsjRddqvh+h
Irgg+jiob7yeqouIBFPMx0ef99cyfKRgpf5d3klbWJ+3pI8NKQT/pVy66PAhbRzADuCpTED0pnQ2
l6IwSmNyivfEa7Bj3mI9gb3gxCqdguj+rCZPfhEgTrLo3wTVAFszL5Rb/AkV4SUfZiNcR24UIjdU
Fcns1/ylJJqmPgc0Xu5w4LvoK++wugJ3S3BYrAryxsNKNTd3w/k5EtGOC0e4tyKxrxpDH/vn2OM7
V4NntsQQvcmPT8z/Zn1kEx/IKu4QUpX2+tNbCvnz8UNSXoWXDLvcOt9oNkNaiHbBY72BN4TTbte6
8ULjF6m9BEl9jFedqUFg33+mGAMSfTKEgQRx2QlPRDb3DHxO3IpKy7tpS9t7sIE9aXmSltlT/NvY
NTVLDAU2lZQmbAfYEw3Hj1YIV0RgqhoJkeU0D428nlA31zt7C42/2Sh0LG1PYNHJISGUMNR8g+vt
6wrpuS0H8dY/lo6sar8PYYuSnAkQ+Zff1YzQcHJnmlN6oOrhbk2qiQIGWYN3BwGf5qT1DOf37gzl
6qIlhlCipHiRnYta3kLBZ+7zy20HRFY+pCZ8LZIYAlcJ/3b1QEWcEzpW0geohrecIauCltQtn6i0
fuP9LJzaDxHqYEAKiV3rPH80+qNLehnl6B5UZa+n9ndcRJtZeYnzUy2PDUSQQL7Cg0CtZgeqgUly
k1z+v+ff7BToAZIoD36xpRQV7orvrx0ekP/1IKMl8QBzzuP23wLxkPzf+Ms2CbGNG7VNaU4rZmcm
He5sQ0tRVTxpJJ+2QfaOW2b7Da7VB5gx7cdpR0qVP0zoBzcykHuwJmSiCfoNhRnxIDhz66obbJ32
HfEJZnNTdgfb2mZkXoBz0kodIZ8wi7hiqQpHMpdw2509vbcajBnXtfCuTriBhxwqyBcvO4O3rObH
Otbm5T9DZ+SHJdFmt0jtZkCke6hX1vsICZ1HFNeaKADol8qQBxQSG70NxGLzvrgepr8A232f+4VA
lEm1AQIVVdRwgP/G6CJsrAWj5lmQuYhAWM5L5GZJF4gGQP6OiRzwuAuJ17QMBv1QBawWVz4/BEL8
1cfNeHEMnvj4DZUdwBy7bU7X3OAKTTCBm8v0TxFtX0ULeg6rlQ+QivI+/o49S6JBy+zvuKlgT899
wvklkQnsUQYzR//EdNf4Kh2jPchTYPZgLFVLOtejgIN4YTidafROkikTDugxXn8qhmHoxszKeU9V
70VdnSO550SFOclt3yqi9KdNWiGiONRyNm6u3kY61uOVLFa+6AXtt/fcS/c/f6Itw+dAvI44s1Bh
8ui99P5oPnQJcppkRiAu33u/magaK0tp517Qn5CL3sQ7v8WxyPJZSXo0itIpFyB8QTssJjig5aiM
XEIdQcqqh2YnGEZyONZ4YpIkpZEKedMHtiSGfTZRkwhI6a1o1ag9znUVMz7FBAG7KwSar7RypTsw
ZytzC5GHzKiNysIVSfQqcmfqt3YkWiczR4WQKBCKNs4zXN/XeHKmQbtP4mqdI1dgl/fH9JifPruR
XEzA+dQY5+1QOv0p0V17hiwguhPJoyCCZl8VwUQjzjWLG9oYv3fnyEBEnFOCh4A/l8HXIrz7khEn
7J1g1E+axeEUwI6dc77zS/3tot+avb0OcPKQ3WWSZYeFPrxK6wywh2R3qTfhtnSDbpWaHNnaQ7tO
tjJklxs/MvDXK65Jt14zlq/c90KLnGcu8JFi/VpEqlLdx7sW6Rgy61UpqMdW4hg/2E5rZJL/uPad
MI2OodaViC4fq8BYMbJiHIEm76cjFPaXWIN4drDtRMT4/TC+eUcaZnLzE3ANEobgTM2Dwg5Qx64M
Q88KHzdmmrRVYbm0a82dNANAbxKknakAr/e7MEjujkOpCUHNQk4xy66F0mNPeosT/kgyu3rx9PRA
QJZkymD9PEakVW+tFEUbqKyMx9jrkclqYMhV+g5kKVWY/Fh6zxdvI6Q+0vzBPGMBT8n1VB9FBgel
DyxScfPUD+H2Ef3klRsjFSbUmbgpI9CdOjENIZyflwdBNpmUNPVgMmCwUar4CIrvK4xzI7gnapCx
dRXGmHFNlzTzvzyfZsay3xpOc5W5d3MsREp2FmBxiEMVBRG7qDotI7oFsBTXLQ58wfMmf11Ti9MW
1zHK+sCaXhwZ2My+Hyha4+fU4EeSVci/5V1ay19SPmcZiJPsbO/mdK1BArft/Ms7/lFt6pHP05G9
nmVKJHyhQMPSSHXOPNFLwcDQFD1yL3vhqtB9qAqgfM/5p/6vFtxHipbrPfw545XwKM4caXYopbgE
xq3jJxRMyFZpiv7hynUZ5eU60r5xdqIVlkgoKg7y/MMu9CE3Scq7jvABqv09gw2HRo7mNQf3+LJw
VS1Nbam+4i/JowokaeKCTUvEq9IID9Kkrq4aDIw84rXM48Wow5/o2caAruQROioO9ftE+AOUTl3I
j6TbhhsWDaJ6xs5gLxJL4Nb6unihkqqZKPj8KAnR3zlMHQR37h4smCOTEntYDcjJQrK+Jg4U8+OR
JdLWgWSftNTY3jZGGPLZ7Lt8RwWvrSJnSxGm8KXm37baZnN0nBjSLKuFGqWLG7xzXLftd7EG9Ht8
AzBUduBm1R1ftcbLzxzNss/vBC00usqdWRtH1O1/TG1LGIC9Pk58aVBtpYnwYZUqGzETaBdSXa6U
Vu+lv4GQPPsj3QfEkdgiR7jOfWp2OHcTWa4RCNcXQGkIN9aV2uVZBROJSfpKDk6V+NZhyV/xaZI5
prAaRT4bmjG6CY1WIf1XKshWIcDGOcQlOP43QV67xKN8vzrfuTtbkg1ib0TfDVqTRWryu9FZ3UkQ
kAbtN7JWxPoXBh3Eghw6mz6T5cHuA1tREnp49EZ/HLPBO8ycsORBiIaGwmHU4raQUxVPxs2ERVk/
0C/CQi3cTPhaPtNUSYtyQg7nU+D/1emNibeoPWGmHmb8oUMDMGhtrxCXZfiFuzyJ45joEjX+8oCT
3L9q6AnAnuhrOWb72Is8fF75TwXh2NuKFFrrPNvHTxptJD4Ddf5I8Z9RWST4w6cS0mHcQAf1wm1g
1b+usUdNJKTIgTD4biY0sahl18cc7tMY6HnwqYbTXnPQdkh8mIOWQd+cxfAxL1YJ2zHzCqkCW5nK
zm9oG56HfTJ6cYL8xrmLV2mr0ZM6WRGCC6hRk+Esdcblm4rj4yRxuBqeSXNpEFimv9YgHi6QS+6i
/+FDvLun6la7u/owA/qVZklUkaZBV60jOYqfB0kK5JEOd6u67fP3IX2zwONnS4BdjV6aHbOvb4k9
98AygBAVcj1z/rX32fNzlfnp1HENKjRrQJRhtY1tJ0XIKiZ3UOhukiPKFsxqbQ2yiY10R7/tS44x
Yp9RSVEzQAZHyjhddyEWysv+npVLLFvLD7ZZZwqDOqb5+11NEX00w/8fYkibN3go3eL7Bzkxrf7c
/p7jj1GMTFoJ9g0pbIZHZcg4dsX6zMzgBRD99eJSSaTAHGBqcOEGWj8Lv/lECwuP8e6Q1mMsMs8r
rDRPfpiNY3ib2EwOWR5dqZbp/O7b74/jLUanT2k8TqtKYpQw7Ee7JVUTm9QneRzQy+roFkxDAotX
j86LPOKZ1qJd12O4a1wiwRneH0xTbxnoo0AHnuzjJXh469NprcUojeqmg+enIO/NYjs1gCVPYVlw
ZeMDbqPZjxv/itEpS9/496wKwQDP57qTXEm0j7FgGikXqq9iZxJsiatjlNfiqm4tevQg+fvG7mCn
9sRkp3TSY+QC6r2t0C099FHg/jxyOznZ8pkxMA36ow5YeKnWryDYUMvz1mUXbGYfY4X2PFDM2nnK
n0H9Dek9lcUxMXEUCLrSpSEDQZ8iVOcN6tjjrv+TXqKr2P4iU6Iviq5a983V8+MjDlWlbkXnWgYv
UsSYs0VF1HUf8UhVgRdX/XuDLU0bmqIgzQJCR98qeEQG36H+cYIkpZczyGV5otn7K9NTKWg/rRbc
+u6Mx5meF7MtsOxBMihW/Ng8ZlMb76SIysk7mWj5LDJ3gQYZgZ0ICgQn9zmwq2uSOka3ie5o9uBv
s8RyhjO3W8RzKyxVeEQ4oJU/zFsD5wjS/dLRvF7rfonQoV0E10VzENiUaz0/ncgAAyGCRbUx4Tob
eDc2umJDV/GMzcKDO4AhmfuEYOgdi6R9/wJBShfYHfaxKS7QkMU0N3rAiMAElqiqtOB1gpv0WrT0
htVevKSsV6JbupYxp1wcNEsts5EtWZ/uIH/ALaKKen82enQgIOXpRjiqD8bbwOJyugL15GP2M24F
vEHJ5ihUurdHL+nDk55MKJ6Z4P9gTxUepv/4hN+sH/fvwTKGgphj0sMiaCppSGKk0ISIi34vLqU9
+MSeruYt6pCwxv+TLJqjnWJHjxtvMqQMF4milSuH/e+Pjz+XW7Yyip/O1EDTLApoiP6wkIwHHBgy
2MkKyHAdMvKoZKgTc1kqEhtPnRiz0p/5WRMRINe/1+zVfnHNOrRnCmBZUOm0flo2Ga/74Tq7LBKM
UUvS0r07bvpYok2tYaDnfwM5BpFKIshcxJSdKUip/ZOXookRu7S4pzS/XyHp7XklK00ZDW9OZiLj
rUKuwg7+SH+puDVAaMFzVYdDkIvmAK5dDulJPvT4jZZyPzN9XYODgJx6cOmvcMUimgQT11sQ9Dew
SBq17eRPVPw7m+5WlQ1QF4G91L/ac0mAA5EcRTLlLJkzV2tHaoqoV0MS1x0NwznXWfqKqqOk/oH0
c96y6+wIoWXrRhpko7058fkqgmoKRYwIdTKIg7OSX1HR8h682tDdNS22f/fiSXVQggJqUhUQaXYn
QnMU9ZqI/6WdTt1cr1Y9z7qU/46xSnKPsQYwJ4ZwRvA0AGerM0eSIfCSMwpla18EevE3JKqFVH7o
1GRGRowBclz6fqxjtuzH5DUW1DYxmYYOlaHbmtKxNnHjXxU5oxIv3Jn5Ub2Gu3t7wio1Bf9q17KZ
smB6Yh3GZGXjxxindTZtbray8pIEeaOOu+L8AxSSFT6MVaN9Yp4rM2XVeIDkMoNDwbIoEs2QwN+5
R4ItPFeGrZE2ToUe0e6zUcYKbS6KrZ/kxsFXjv91k+n8mI40efe4BeFu8c0Mr+yb967z0SmkbF9x
jHVgY6899VGrXo4JWYeD9tmtVDoVRCG4ZJk+ft1/g0g+uMfzaI/jWck9Scv7OL/4e+KuoIhByGIZ
WacgDt3SGuR4YnzYEujW9/N8HDIHVpFIZyhytqo0x0W/+Ca6ckjzBa86gOj9lK4q0Z5AD1iNln6g
4cxRtTejS9A9G7tVxlV7rCFoYP01jLqMSam0HCSW8AutaLJj20AYiwDLXrwhKV+FL49fsaffJu2O
kHuVaJKgjI5aZOpg6phjNJ5ZvwRUNxBpO5SRFqhnPQtbmt8qgVSubm5q0ouUnWonFVnsO/Sz1oXM
lCm29JC9ZY2LWVRnRU9qaFxJi1SLhLx/BI3hHqkCePC5G5etuMhkVsOt+ImVbO05zI3nlcuQY/MF
lB1qwbvlN2oM8fKe704AgAYBxC23mBf3sOsOkvJ6wb36QerovejxDRYprq5V4IKXK+33X+vqfTUi
voGn6Rx67JAFNpxrUTkjoTM/TTgmYqgd6BNKIt/H6KpQsPm9nHUAusqCz1FNOU7lFiO9w/+GIm4H
7lssAmH03SLbt9rLPgIP13g18AeiPWUryF2/po0NfdV0eZJCx08J5DghdE+ONHuTSPYIocV+nkk4
IEBwHivTYfIEtsR4bMemtbHwACpNrR2UHWelW+ckbM5tP0fTkcHv72D/TwnMiBN82h+wWTy8blqE
W+iS/N08aqpf/oeuT6izaEKbpS94aVGEMz34uw+Gg4IVs7NI9MeLaJmJsLvmzvztAb34mVKHz4QX
MvP0pH9ygxR7/OBh33FFkMuzzPj8bl+gRDPi6M/w5QcutUgxJJnfiLo1tLqfuG3BLIHLaOl0CkDE
pTT+LLwFisELB7qH+8KdO/U6uZ7VXyCtj9avVkEO96/ZNXb15S3lgxEdXd6Y3/r0NIOJjif6lgML
2WPqjKDRzvs6NEesewMPQT0MlzZX4Nq1hG6bPh7oXT+d6Y+LkB+NN08eRKefCO00mjjPMzittC/A
R5wWXVTdGA7fd6JNjx6vGjzI2eedeacr1fjyKwqyx5rbQj/L+BkToWxGS4a3ZMYDXs++Tf4w7mg7
1iIdRqRF+whjYLh1OiBRKrt/8CvFAIHYLq+d8ljgkP5G5bM/5vFaCinaHshilHhlxPuPVItE7di0
pUfpyOdA/sjPCT11Dox2/CO1u4qA8w5BXJn0fHFdIKQEmVofm83gCoMk8WxCrtSEtMxvLTHh/d9H
qMXdDgnDPjR1NNa7X37GzIkC3BogDDVPgSWhu6do8YQotae6+QRsom+BZNJbBXudpSbb8uDDdkLj
CEeIQOUsctDwJi+qJ6ckKuZjyvH+AgRQ9skZaIh4p2mRf1Hg9UTiFZvq8meTZtLbo+nrccUHLQhN
ojGhaZRjaTRj5yLesyXmms0mDy7gAtAkfVKQUQl7KyPFaiNU+xncMna3jhEWcaybb03rbbBf9lcB
QvyVw4xnTInUpvdfd0Ui2P3qH2GpLrUC17YT0ZwtHK77qiYG5aTKDtLzX9A5Dxl74gpV/4kEKyXQ
rValhdlXMrTBiQVFjjMKoyVJjLK3cI++Aw38bAfLwL4TpG+RUB6coTRM0ZAZUq1n6XDITOS89990
19Vn6ujZrmV/5mMim0tVW8flluFKJ6fY4yfubE8w1IweBbQpPFMuG1D+Vl6+ypszJTh6+21cn3w3
QB2UX5qWm61yzA/ViYdsfW4GROjr9dxp/yPkQgE3gSz5+4Zffu8lTnuNWajOXeR9IVAH6LCgBhGd
NNYmMxF/32wp+CAxzoSv73ZVTuh1W6lvuS/OdbiKUuU9WTNowvH1hbdBJpgkIUzC1z7HTcXE6Tfv
VFq6UoLKtFGZosWEac49plBBDrjIhXqhE026i9gTyjNptudrzqfV+o0xhmJLP+bS/7aBvelASiuB
Gjc7mDzkD9SF9RoH+GiCWUCs3vRufeXtraI7N4SDhSq1m71S8ztDp7oKqOw/qZbmvZGFT8TS4w1V
VJZldt3UFT1KT0AXyXwWpd+Z/Mh8a9Q5whuLd2XQIvBHYQ7b5O7FCs9lnZL8l2/ezQV45HzRNWhN
OSNJ9VrxGVp/zbSD6BJDTNHyrT/9jnz+3zgXuU1p853MZzdWvjSITUMeTpomEM8ZrlXKE5fSa1Qo
IhhQ6Y7d+kbKLabqSf78Sq6zWWU0wf2OPjbWVL+IWEMTOrCTxTTD3c6uZ/PN0/n7FsDzKuZaHqoL
/g9w3LWLNdtSv+3Q43C9raN9vQG0fSh8y5C9YAB4Ip6EGUnbaQ0h674GTiVu+c0fMMdUAIpc39hw
px/QzLR+GMDeCPiG94kssily38MIRZ78/Oi9vSDYsKPWR22Mn6vzuEUgJfkDuhbkaK+p+iLXA90X
JKBq/cb7nimmUZAGoJWDB5kRhbCflx8vndPSbrsIYOfWFtKzj7LUJpie//yCEB0P+Tc/YcXEZniM
ldLJyQTA7ltnerN/y4/LLB0Jh+RjGIv0JV62XEVsmoESw91SnKhuFLldhW4x/RErTZTh2J0z5WiN
uD0m5LBjc6S5cZfUeYyb8uiR+9VCxM+xEOt9l9TYTG5j2o4oxOyKvoSkgixX4ZJrXukc0L5P/X7q
/o18vbM2I3m3NZ2vtzt+Qj/gkIuY4qBWeELWB0iY7FLMkIKJLSLvouYXYBZL3Q92wPKqI+0vZKZ/
HSLqmnNO4FzvL82bJBdGrV4iKE5oPwPemfJ5zdu9E/2+p2OzhIdjO1lqxNFik+UT9x4eRIgJLbsI
34QsHWJ/LSOuppMWb8HD6So/IUC63eaNeo0xFPt6WyDX9xT2GtXiBrkEHggp++rpzlQRs1mml5bh
B5bMsxV0536bKX/yGVsn7ZKPIpBn4qV4neOEI5uJ0EDyIf0/mPPALAodV92mCvyskEL7q4d+uWRU
zH6SuOEGz42wF4HL3Pq9IxyEb9kvG2Rirv0B1+GEu2Iy4OXVSz7go9uEkjXtXpKtjsX8d8EBKVXU
PE0aRxTjXBvqEbx4nMJX8xc+HMCtsZ5pWE8wmD9OwArYOu8bnI+wwaKINMssq5KHe5x7TgpQsW7f
cXOjY3F8+z8D7zDueso+AwwdodVkZUrM+Vevm4+nVdvBd4jKe2vxS3GGdCycU8qH9DPW0WGeWdZb
qncguSdwTCURQ5pcOTfXMFvcOQtHKo9pR5GE7gsvw4jfVQyE3+1q+IxPXbDIYcqWsRDRmoRvvRrY
NVahxXgMcRpPkCyq0YTr6CdqKqE7exPDzFB85G3rQz4/rXMNETdYYXuCRRH7dGwJUQi9iCE1e2HN
DX2XkuUJ2Nlw08LowhBcitjUVlgKu9cEjn98lKALPPj7Pdm1nwl1v+5QCGyZDHgSU16Hc7szC4GV
eOH3NKbCWYeeSPxHjQ7bPHmPKrvenO9boZEZnvur/Aw9+3FJjuMYKxcLVxJItnfb2D3eiFEohTrz
2AzCTIZLKes2I4MEpSiLsTikVWvia+ixykMtokl2c1KbzX03q5CEMpv7A3I4RvcaKJC3TeUpVEFF
HuW8Ko8gkw4uIFmFa7vEqlJ2btartJKz352WuxACPx0htkTxjXYK8GPH47E4VIGVBZl3RxGWIXsw
m1/hcJqZi7CuOB+ncJTsslZdRpsq5xwKqi3JS7cNG4vwdg5bpd3ZRTSF+Y1qhEa5vOiaXHwG0Z6y
OKSnVMBVYDJm+dofIvedTGDTa31IrZJtlzE0pe0NgiHmfa70tGCvvmKyqIfbZ8VjPwfEmUd6hsSZ
qSKElWKbaX11hof5fHsMEKgGMNYLRyY+mmQQD6KyvMBN+g0bWawWsVdfBWmoSbMWxA1f8vPPDqdH
KcpnewnUCqOZNTd1wBJ8nl8+hq5a2+Cp7EkRG+hfXPG9z4jvZsqMQLvb4+b87ezenKN1V7GILUMN
SUc71ERMBvARZIfi22v1fP3o/5kEOFyOTTtrf8GlsavwAadxDVL0ckpQEIONdhBloL6/KvzeBlP/
MUnQdPBe5ZiA38D7UX8yqSN8tGEKxenHJuYIrqitqqyjb2FO/18KcEX7wm8EeUxqH1yd6yyEjruW
/0fRilPTdWMaoxfWxBATjsqjGr8T
`protect end_protected
