��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���;$v�V���KC2h�7�����	t���r:~�6t����<��o��//�͊>gY�.�_�1�.����P�ȵ�,��ᴹ�X�<�F%���3����[8����;��P�
I /��W�E�	�X�W�Yz�4NjM�e��p:����������^$8]�9�20�Cϛ�v�Y�<�ۗ�Sk#�S���	��OdV� �O��xp��l���3�@���y����L@�}q��q7�}Y�C��Ԟ��q�P�q�G�r#�PMi�߯�LJ�zu�c霝�Z���QM����S:`��LriWlI���3�cI��.�<������d0�o�Z����47Yx���bB[�ͱrO�M�n���ڠ���8F�4�U����3��`_��;�� ���o`h��Y���f�E����
����8�Y`�H\(�����$��>��#�x{��	���Z��6�>���V��ahup�H5�I�Cw(w��q���f>6�`����1ï 7���*�A��3Y�Fo�xP��;�,95z�*�I���ܮ�p�/������L�P�{f���� �����E~?K7KY�X{�ξ�cx?G���`m���C�b����4�����LQf	�RI��\� u��SU�N_�hO��\��)�W*���@�&������U��S{m\<�A�9U_�L�rꎀ�L��%�<��H�����ٵb��O`�G������C���G�����B�}�掚��8�gx�W�>�hƦma��δܭnd`�����6y��-�Pꗶ�7@��6�ZOWqh�ʙxI��B��P^��3�r��CjZ_��v̟�}�e:)w�*
�)��V�
ew��j��� c��q(��e��6�D�Q�菙�4�+��s�T�Cy�:�@�0���#i#�6J�8!��F��3^�'�Y�>�!�Й�H�Ռ]�����~|��Ym�Or��k%d5��������U�ҭ�	��'���ӷu.�$�;0i�o4#J+iv	�����/�qi�q<�����1��<D{�b�Pq��!/����:[�ɣ��J�-){,��m-B�	��&����_�k��pdN���a�dc�7Qb����(}����M�> A�@�9&�'� ����QMX��zH:��d�w) $��1#7�&a/̖W(�<	X~�\�-�>��:s||[/#�o�5�Ǌ�������>}�]�%,�n��J����xO(e�'i�i��ҺP���D�"T��
�F��-�	q�4B?w�
#b*��l�
�����@(�)���^�Z{8f#�P4��^�q�,�ȉ����I8^��3�?@U��\��_q�n� ���"�b�5�K�ӧS�1����d�����͇Ru�����S)d�{�=��"���*LDJ�AJ �mf�k�K���7pزb��E�34��?�Ǯр�<b{�.=+�$m�"Bd�rDd��6;��5g)u�zp��l�~�F��y�#Z�HCŭ(���$*#j}	's=�u�qӈ��#
��v}�ejI�X�%ʍ�>3�ڑV�^�w�p["wS�Lg<��',��'���@�k���z��Y:4������PF9iI!�/U{!6�`���J��}݆N/nS�&��}2���cgIˍ����G� mI�!��'b0Hz����H�E3[�qPZ�&4L�����Kت�E��0�ၠ�'����#�gY;6ղ]s�����d�`�J��������Y_u_m'nD0�@����9�B����{�CVy	*�,�#+����]��
TX��yo�"=�C�HU�}�v�5 J4�^e_,��Djv�Ͽ�>q#�M#[Ձ��`�l��	Y���q巩����y�a��p�D�ȆڭaōqN	\�B����r7aLM�ZW���/��מ�=��⩓u,���6�`9ߪ)���sM�W��0,g�u�����5�\9�t{r��w.�a�o��l��P��4��6j��)B��d�'RY��8�٦M;Պ��_����t�7��<AN�[
���1Vt�U6|9K:�mң���1Cm!@��C`ښ_	��LgZ�d�X�q�Df�?'��H������L�AŲ2Nʪ�$�t��}�'I��v�?
w�ɲ�=���Y�9��ϩ��(|�@��x��Z�,y�a��qu�>�g��D��R�#.���B��9����7I�=*1
���2}M� ��Q'^�x��][H��Ew�	��O� u��P��ǭL;���hJ_�5�'K�=�1��;�-��&�p�B}��&98�gߌ�·;jbN�]2��w�v��Ǣ=�����X�;&�9|����M�C�Xj�^j���B�r $?k��m��ǻy�ZV��nŎ&�R����]nD��5�ƪRO{q��H�k��!�w_HΌ�l}D�8��I'1�n�? ��m�
�r�rKaW���{��T�e��B��B+8�M'D�_���~D���#��W}��bQ�aUŬ�賛�O=�]�>�n������
�Y����i�