��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h��[Z#�ڒ��4m�ə�p�7���?������o�;�{��36��aI�.��ڞ�S/�"[�D=Y��G��1�ZG��kv*�����/0�k=mO\�_�-򉻡����֜��(�
�h+\P�V�J��a��4�;�p�bD{W�{����j�QA#�R�^U	F,���L��^�LBt���� ���a�;�/��*��IWy�ϝ�"�%�'���N��\R�.=����c�D�ϒ��7�l�ܴ�?������� �		$�b�X{� ��d��u�TD+"@.� [B�F�If1�(*k=����/�q�`�u�W�)C�a�� ���p}���H��0�y��B㡾T�A�h�Ҟ5|%=o����4i��/t�N�Ɂ�KC_�t���z;�s������6��:3Q�.�$��+�b��٭���#ް���'�r:���\_��tNs؋�ѧdF�x4s?H�x��q��eb�������z�F��^D+6�e�r�ts��� ؠ~3VB�s�zX�Մck}��)��X����?�)�_�+��·w6�vhMS������:C�g<~)��͔�Vh�.]?Ԭۛ��?�y~Y��'�|�>e�w��R#X�`_�^����?!���Z��*I
�L��`���{�*�Vc�(��)�FR6�6�������i��\�+f(1C�70�`z[�
�Q��?in�⹞D���jT]��*��N\�i�oٙ[>�Dا���G��Mg�|������m�8:�J���6�b�X	r�k`�t�׷�����R��A7yS�{��p��K�G��W��;�g��X���'c��x�q�F�_�./�RՅ��dw9Mƈ��>��d2�w@����i������n^Y�pm\�d�#��V�	c��Ks���"��=��@��#$n�r�*�fh�nB���r!z��W/*C���Y�y�Q*�	&�m���G��4x^��*�A�ld�*�OW"���])�PiW�'��	�;��Lnj��(J�����o�j�ԺcY�ƊȎCz�	\8�קU�9���}C��������_(e��W]���5�+f�d�5KLJٸ�͵��;����|�F�:��萤����9Mاx=��+��������)�V���pO�kY� 4����#��0D��址�O�U6%���u�������ާ�:����˖�����w��:��)�z����j�G�DL>���uGf��J��o��_�����E��fJP�_4?0,��Y>#��������UF�z�5V?��9~�ŋ{�B�:�# �a�[�:�q�Nb���"�fT�g��#Ϙ���aڀKoz���t�-+T��2:�S!*�nV�����bئ�|^��X�"G�B��p�(]
?�|�z��!�Do&	V�"���RT9i��Fj�ARȭG�2�A|���&�x��	�Ӡɮ��"�a����vx��1����I�DhBߠ_�+�E!�%~X��F�!��U�����fs�6/��?6���M�@�e��pI���f������j?���	$�Q"����MQ��w��l��X�Q�H�k�%x�2[�eU	�#?�%ό�����}@��l��Q�!��P�NMVڸ��j�+X�AY��N?ѷK��y,�����{dw�@G�k.�^R��a"pĮ����x�@��1+�YQ��"Mc��[�}��HP)c�h�:��$+�*�������_�߈ �U������oBtk�����|VWdɷ<�"����+:�>�^����^���F��<V�^���b��)8e�ē�\S3m� �rϤ��t��k�����������8��\:)��^��;��w�T7��
c��`8Y:���^/Fn�.-a�e����LJ_�c�4�f�l�;Ukfj��PF.�R�0�j�ȽT�q����)����14F��/k�޺�y%´�-���?^�%���xJ}TOo��χOn��
��Qh��ǣ�/��`s������S5?ѯ=�|�H��j��8rc��)��["(Yw�u��"eh;�=��=	�	̴���@�˟��Q�冝�	Uo���2Z
�����B�$OǌoiEt9��3{�4�&u�"A�j����M�.2�A��c��hY����j�g˺e����y*j�%�Ӝ>u���Q����{maR���f=�E(���d�h1�#�4_��NiT4|�iӘ#
�E_K:'a�9{X��YX1U�C�F��^�x�G���P��0?�?�1���愿�9��� #�L#J��'²���	�uI���"46���<5�-��`�r��RT~�j�C'����V6�љ�l)^���j��+�t��6'Վ��ش�1|��>�~�̒ &sV��0�AG���v��$	�`_G�lv�������D��+�
���F�-y�	H>�C1�4i�Tр5� �0 ǟg��� h&���x!�ٳ-�E�������X�u��	���s� ��k�r���.w&�Cc�e�ȕ�ɨ������]��6U�=�4�OT�J 91��`e�?q�i�����������@!���=��͘�Y씗�㽜,v�Ԯ��,�N�7i�K�vJ��Ht�,$�`y4v}v9FL ����z�!�����qho��8�
�K�'�:��=�6O7�.�
�<�'}D�A��g�
���P.�y5wc�.x��Q�0Oǝ=�z�P�g��j�����ò��w���Hǡim63i�I�^P�2]��NMֿ9f^��,�����3�+VJc�O��0����I#3K;�Χ^\�PdsƄ��1�i�!����[O��� F�zW�ۙi�Ѭ�1�c�<l �PL4��0��\q��	��p�Top	بȫy���K��#*{ߛt}�L�F}�+��vNz9?��hHv���z v�ǶQ��q��"�'���(�*i�X��{kH���j siE�!�am�b��ڈ,��<ԢV���E�f�,;� N0�`1�7_�yri��*���Z�lF����ڎ �`���f����<����h3@����F4�N�8��Ka"�$ƃ��f�����ǧ�_�ىo�ư�������Ɣ敖v,�A��?���ߣZ#Z}�aS��=����x���;l�� �T�L:���C��.����l�Z�[EeWX@}V�b~���I�^UF#-u'�������?"!m�@Ġ���g�b9�����q�Bm���.��׬_:��
#k}����A&x�?5YME�^k�Pj �V g��{$m�	�h�����#�x�@9�Z�>\���$��(�1w�zhP��?G�H��T�):�;�&����؊��3U����X�C?�X@|��C1�e��)���湿���Ŭһ�����9��6�]凯����]�n#J{Lo�˦�9����j� 4�����Tv� ���M6̓��1�j�#١3�b�	9��J�{�=4�?1BEh��	ץ�aM�<��R�J{��>�꽕W��m��K�q��x0� ����,Bp�:d���#��������(����ْϟ_�%���%��Һq�fo�zQ�<E�sS��K�ٵ����M�(/6��JzQ̻d��g��2�o��hv�"b�I�ny��,{�+D����%��^d+�`�C\_9rʻ�$(gU�q��?�@�5�{u�!bכ�$(��٢�[��s�i���_]!m����GP�v�MĖ9&�QAH�OR��Ӽ����s����D_JI�R��k-+З0AE؉�7��aS~÷)����z�A�l��zWd:����Q�}*�&-.�|��9w�@3b�(��zė[�2��ݼ��ߎ@��3�=�y�oK�0����N���Q���)��R���M��݂,gK�J���}��ygbSZ���,��ǭ��o�V�2j89�7���*�}5"����="�KB@$��E�f
�������M!�eNa�NM�r9�%�e�
�����y�p|7�T*��J69�iE���|��T"M�@����06Hq�/�=�N����*{�R�}KbNZVmA�Y��L�JR���NX5~s�e:u;x��]���LjS���A �����5xC�y4v$�'q3FD�r���1]cOǋ��e�&ģUH�4B�1[����%4$�Lz� �TM�'�ĩ	����d���3p��l�kI�N�E+Ŝ�S�u�jUS�J|<�9�"�����bs���;�Z�*R̗^����"��&I�$�|44r+��_��mk=����mv�}:�~��{�v��KZ�P�4}��j8e3 �4�~;�#I	N��G�v�\`*�>]��7a�o�A�k$Q�	*��Ɍ�Y$��:خ�����r���tZ���V�X`�'ƹ���]n��_̨J�(�k��{7��q��aQ���>d�&��Y�E�z�w;����b�y����_�oX&�C��!J��;⹏����D�REs+#��K�(��m�����?(������x��ϓ2�i��i�QQ�G׮b�[���)\�E��l߂�bx*�L�6�$a5�<�R@�i��)[�vۤ��}k�'�
Cr�����x.WF�|�,������>:��|~�Hb3��|�5�h�~�6�]F'���r+�����W��a.�Pk�;�N�E��,S��\mk����}�j�tGW%ᄴ���	 ���&h�|���M��E�7x:��w"߼y+�g�l�{|k}��׷�I�{�L^�y��ܹǇ��q��+8����6)�(<
t�9�m��_̤.]*�p�*P��+#?#�ӗ����Lf8�W���\�~��J���>��3�%��ʪd�wq��)�@�+~��_�V�ʵ$6�"o����_�$w�z2Ȟ^ at��e�!�͘Y��ZV�p�a�t�i�V��y·_��t�H9�Q�0�$����%k�ʥ8�pg_l�����h����a?a�Ӌ�+������Y��g��0���{�b,�?P��|�j2\9��hR5H	��a�21d�q�ˬ^6?mY�^�g��iH�s���L�].ib�M�*�˙3��ms~��Q~>�ɟ��r���r݇�"�] q��ޜ�C9�f�.8?��*�o�BC��=U�9U�� {��D��L�5i���e�?