��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�?u+οG'�K���Y�$/��[��1��[��ea�b����̞Y%~r���&Z����(����u�"�l/��N�I�V�>���@
��s6���,��G�����U;�Y#W����sA͍�D�>�'�<�����+?�5��'��_��"ɡ�m��� ��8�S?I��^��1�5ʉT��<����ǲ���0׊7(�&d˙E�9iI���d�8�0����Q����S�=Õ%���Y�)
��Ӊ����#{��p��|Fuq���1��פw*QS��O7�4����$���6ݜz����2�IU`V@)$����J3'P����vO�B�/�rڇ$t�����5G��c�nNS�BE+0����i�jg\ڇ��\3����N\�p.%�p=�~�)&�0�&%��Іl��8���|�p�չ�;���9�0�FW�ވ@���� ��p�}qW��3�|
�Ae�be�!X��Q}��G���g��/RNZ�|`�r�#��D���:�rf�J�/�8�N��SI�
D�h�U9z�|��YD��� V��e3Fs��7�(2��	�� M\�4�^)�+���9*
�B}�5����Wª�2:��8�"ru@
��c����4ik�?�`�M��e>��W�IJ?喝���fhd�b&��#<ڸ���f� �"HiJ�Ѐ��,�	�˾�f�{�g8H#T;�OB�55��.K�RL9�ݏ��c�� �SV����!H�:/��<0y!Im� �z_����d2����1SM��/CR�>5� �{�/˔�`�%��~a��k8>+ďtY3���*L�5\9n˃�Ȍ�j#}W�~���T�V9��xKr']Y�"l
nE��H8�a7`�t*���<1O����_q$a������SQXb#d�l� �j��{w��J�s�.K�w�%0d�7܄��H��|MQ�eC�����Z�*̌���+�.)O#�lE��	�=���p	$�(�`D�OiFO͍l�Ks�U���P���c�ګN tϩ������D!bu ua����pa�ݺ�M	״	:��ē=�:�+E�#J�򽘰�X�l��������}�� ��Cڢl|�
�K�rn�[�~�<C,�E)��W�K4y����Y�
���2p���n���2qb�8�L�#��r�Z�c�l�e'���N_~��rj���ǡW����Ey�#:�D��8uH�}���T�>���7� ���qz�d�'=��{�|gD����>�X	�^��^K�ǃ#�G���G�f/���<A�!�Nc���������*9��#����]1�,tp� ����+��A���nX�v�\���_c�W1Z��F^Z2J$]igjs�����趁��v̿M iq�X�&���]�ά�	���t����g�$jߘ���z����_i�.��p�ic菇��S���ȉ�=���C�V�h�ż�KsA��<��\_r�L3��ڋ}�d� �":���A�毧/X�C�"�gf�Df|��3�}����]��l�#�k� � oU�{t��개����6*u�.�X�s�h0��t�&����?{�09'�t+��+�K5�I)m,���C��c�U(���q�iW�ڛ��k�5t��L�Լg�z#������,�0���ɘU%>�[��vO���OO?��Z
8�=;�PE�r�^8�L��c��{��2�d06e~jI���E��O�E�)#����!&����-���b_�l"��lN��*INB�Y�c.9U]�ᩒ��(wZ2�ǝH\���l�"hX���x���3<	�qcY�KjXi�6��ܲ�H$<*נ�h<\^�ʝ��|2�?��i���z�I	�o�B���풔�lM�r���)��]s�'"����fՆ�,˧6�eÊX�"ulե2���,q��+d��09��锋?
>�S%���!: k�1\�A��1�I��Ņ�J��󁷭ah瑨yC2_0]S�\�Ԓ����易�ҙӖ�	���(�s��c+��a)�v��ږ@1#9�!y�].G�wۥ}�����/��n�W��'������)W�C���a�n�
լ�ؚr�kY!E,�����w�Z������0۬��G����dt���}b9��nH�����J��eR=��vc���fk]�>�&�:�?�:�_��y	���ˠQ+ ��y�`���4��;�&:}�"��}ݭ�ח�7�N�*��Z���5?��\�M�A�/;�Ϥ�i�<�M�dhKZ���p�`���2OIn;�6�	�p_	s�}i���?*,^�?�l��/U&������u�� X�
�z��o	!����(���,�P�z�`�wy�P��5y����'q@��u\:��
Х�P]VA���qX0RA�����hf������`����b����~�v�5�5	o@���:l��֛�3�Ts01m0�RYɝ�.��K���B�V]-q�Bsfۻם��CV��58�~����{�v��V@���gN��3��j�I�@�1�	�)�J��b`ON݉��rG�gq�����=͹X��/^%�w�奙	�b�������=Gx� s��3TJ�x�3�n�u'�c~z�*-��arg��F��b"�/CbGM ��)��A�ӏ?�L�tB\�8��Y�+nc�ц8 w�|��,I���n���x@��a��S��LS���A����ì�H՘CL�\}	KO���<�!��Ehˇ��1��|�u�H?�O�1���$���v>о��H�fAgW����7��U�U!�0�9m�Ş�R���<����lA�����%�a=�t!kQ<]ETasJ2,����y��^ A��u[Q��|ϑ��'�H��%���7��_����v���q%d!��?��r�y��(�ڤMJٷ�S$4蟕.>=%g�,Y���@-���SCW�����7��$bR���Rs.J4Ӕ�ؓ��De��rBح�)�L*��3���4bA�n݂f�-�0%
�X��h�(�w�A�l�BfPJ������,�^`�(��Ӄ�
��1R����?�E��V�p�-��`
N_�H�CS8=����.�qt�L�Wc��
~���)=�L�6(: ZU'������D��ȯ�M���J4����z���ɫ>����u`��2X�ߓq�U��^gN�l���;g��Y�9D�"����8�e�����	L��T��ELf��-�|����!�^o����F����.��<YS��NP�V�����U&J��/X��W�$,�{-2��@J��Lo='�l�ҶN#"۰�7�Q�>Y���h+R�� V���6��ONM�D*����gS�&!�t�w^ �E�2§�A��i��y)�"�����
�D*�Ñ����3�x�^*r�ι� ���u]>��׻�G�	��ǫ6��| ���^�}��#���V|7��=eu�~%J���5/6(H�wA��%��Ò�е3{{/���|�b���;2�󎴶!�������ɓ6�0l���j�ϳ5ٽ��d܂D�q���Մ�Z4����N��ϳ�z���G���=z�қ����`�n0`��%0��j�&��M&�hI���%`΍b����OU�~}�3�s���E�!�e8���z�n��$I���m�A_�S�}&��P� n����RT7���Q2��N�!��`}�͍�r	����=i0���[�ʄ�:d?�0����̵��f�D��/�eP㻛�0Ǔb9�	<���}���yۉ"�RvXzN$�پK.+�P]z�@����}{�1:�E ���S�ۃz���ڽ�W��;G���{��e�q���)0I���X�#�a�L��S�{Rl[M�4`Ճ�їG��M�B��<+��X�Zg=x�����y��ގӿ`i�������7��������Se�U����pJB�*��z��v���a>2
֎}~����t�`�7q`���&��2��t��nyj4�" ٩��r�'k�um剓N�Ƴ�rhv+�=���zS�p�+����=D�׃��U�P�ߐ�ʂ���Иryb�]ȉ�%1�Sm��XQY'l~�"��Fsg1��Zs���l��~ȏ��9���|� +���Z�{=0�O>f
�����O�)gne��VD����%�
ά��ntt>]N�=�	aG��pi��>�䝇�l;���Rf1�η'H��㰓A�2Wa��	LP0h�[��*#��uG�N�X���$��_������q 8��!���+(5��skZJ�9�g�,A�le��3Al\w������ݱ�C9����&�qq�� �!���8<����ʰ�O�c��W�q����/�/�,�7���EE �Bd%��(���p���7cs����ĩ��X൰I���'L� �ȿ2�۰	�j.JR%w�/R+�J��鯖?b2�)���ҙ$$�%�z�:��e%V��mи]�]!JC�>�{F��< �ʉ�~�ﴖ���1:�(�E��:x�=����APo�r��zЙl�c%�L	hqd�<�ת𨡄t��y�:�[R@��RPcs$9ݹQ��?��Y�O�(9vM�K��p	v�f ej"m��F�p"����o!��o�Ԫcc(J����Y���	ie��9�ݙ�b9�8k��0g�Fw�פC����0��jTz8Z����F��9�*�A3ʡ�LC��u��R)]1\��vT@_�Į���tԢnh��i;Ѥji�m�����
P�K_Jtw:�OU��,�	�`ޕL&�X�B��u�h���jc�XB��02qaH�Nzs)y��������a$|�l��^��	���FVT�?��}ݒO=P�x���0|�
��������p�􃞄C~$�)�{�6}�6��P@1/3A--�YiĕW��b�_��;�zy�e��I�s6�S�,W�C��a���YO�5*�C�bd�ȥޢb���7R��l�n&�t�[L�ܜL��Ͳm|��'��n̝Q%��E�E�Y���j��+Xu��*�A%������&�Ŷ��%V�p�7�α�S�X|lM�M��N��cL�>�n�3������Z�wL+>M#;y娤�sؔcy�׎9k!���8�ȥ��Ԉ�z�i����ʗj���:���4J��9������$�\^f�(�Y/v���|Q����;��b��ZH�:�|��F`��vP���Eo��)$e+�mCJ(H��R�F��>�Hݹ}���v��5QC~V�$�b�O�Έu/�7�m���Y��1c,�ĵ@�`5O+ч�D�P�:���9S�M�⍇i��p�,�S���_�H]a_P
/��a6�E��M��Lf�6��L��*}N�,F��?�q�q
��D�v����9�]��Z�U��Uf���f�R��@v+�!����|\�Րm���w��w���R	���CS:=�l����6�Z��	3)h�4i3���b�J߈Xl�����zo�%%8�P���f̶)}ZVO��P5�<��s��f��pP�4�� �!�ƈ�`��'{����{[\s+�>�,D��o�O�q�(fMQϟz�����Sk^��z�A��c�I�bx���(T����A*B_�d����jeD�54i����$nm��*�.�P����z��0��e��� �r:�e��dxlo��ن^Y�ZBҼ7\�\Қ���@��a�����L�5�����¤���Ʌ�AK ���:���*C���J�ܶ�ީ���d:�!N�<�Tnm̀�72:��6!qඁ����d���ͮr_�</����%���37��U����k�	��Bu*�K2u�,K���)���Z�HŢ��L�c�T"B�] ���Jk�lL�T7�����.��=^9��0��o�[]��_���|k��h��R`�)�+n�2��о��%+
��R�8�*��Ω��xEWuI�T�r3��������)+I���=S�{�5:��ӫ������s3��$�I�`��tI�uw%��/5Jw�s�y�b�^��~�)Y}9�Ot�9m̑z3U����ض�[����wF�w��`�E xS�T�����g��B=fF�TdF��[��l�+�����3|^A���9�����A���D4�21%��|7EK {$y�:R�5��*���f ��d5wko�vh�	?�H%ȑ���b�,W��"+�<t�K�1���3_��\�q������UA���ф����$�^s�YUj�����נ!�t�[��m� ���7�Y`͕Jmbvu���6������^���ft&�wq�0�d4
���m dh�b11?MkM����ؠ*	0��M3��3ɮ�I�?i�`Ԭ\��7�2�
{,��؊�Nnt���"\:S�,r�g ��˖ے�U�_�p��N��Z�z�?�y��|u�0�`��P��6;�$�Kt���I��(�g�1k$�3_}D|�z:Oy�P#{��e��>�.�xhU;V�dt�����~J(���ae����8���"q��g9Ɉ�QN��d��|��~	�c�����
�|)�t�B�Z&Ct�Y�A�aǃ�	���k���(�z$��j^f	�3mc��a�|:Pw<t���ՎX=�[_�>�E\���������+�.�]�ڝL�.r��H�^����`��F��*�����^�\��X�7@n�g\lH��O!�>N�lk2��j�lOѿ3�(c+T߂�_��y"����[�,G��ƹ):٭�j���(+�Y��>.\ߛ�|�ʧ*W�FG䛀)�,���mg�XK�}����=����=_�*���n �̳&��혃 ITF�Q��!Lu�����ɤ&�BΔ�;��*��&i�6��p�G	��UL��֜���Nb���Ȱ�0�j�ȼo	2��
5�=����HA�i5�����yiB{kQnbn=v�A>G�
�2�[�w{��87_6�^0$j����?n��p֛+fV+�eR���aŁA��$.x��"ђNT��S�$�H���[��N�ܓS	^��J��� �1�!|;/?�TyM� N�b|�Y8QQ��Ty�����ރ?8��'�q�Z8G�4�g����W��F����Q�D7����©��6US�I��yR��_a3�5��/AO�&ܦd��Și����~�^���[0��\f�š%É{�3���q���Ke�G2b���p�y���,}w�s��W!�e `��P��'��fZ
�m�ʎÄϾ�8	��}<�A�%~uzj��Ō ������D;u+	#�j�V\{ZݐY�<��rb[f[_n�����Y��	"����9�"���w��6�9�@�#�JIn	��P��)��0��(3D��1B��o�,�2����:��f�C@'7"����/+XƁ�x7ȦEM׻���7!z���Wz<=���K�;	��������o����l(K��tO����XJ�>����KbT���\d�B�+Q��%!]���TN^�s�4��NT�aG�y�=�#����b��~��2[=��G���v�)��Z�]X#�ߕߔ& m��	��|{�$��x:���k:nB,G��ږo��;���{�� ;��Fvr���ǳ����7���ڟ��Y��t�r��?��{If�����t�O��᧣����B��-��DJt�7�b˕�����n�v��Z/�r�Z\����6�}8�Q��8�����-Mz6G�)-eiz�zr��x�X#���_ͥ����G����Q�YsaI�w��2eg���ē��$P��֗9�_�zQO��e���n�����^`�5g�1�����8 ���-�L��u�#<��s&��@]z�	i!���#-��ݩ�J���`M7��u�� ����[��m0������Q��	�=1x�E�`'揨 ��?�4��/�r�5#��(~�����ׄ��
����A�y���m� �᧙C�LM~:6��	T������X�֑UvE�0��r���N軟���G����$��Ǌ�d�M����1r�l��
�Ō�7���|�4�������g���r�∫�����#�ҝ�.&"rQ��|�f����#��A��b7��!����9��W����f�s<�r1��&��ѯS b`��,��%���5���S��������� ]%]�4����W/,Q]�'�eX$u�2y�̧�ւi�ꘪmh̊�2�%:R�h��t��o< #w�����Fq���һ�}ܠ^oD�P�����';���Nֽ-v�GO..��"��V8h[3�eel��X�y����v�u�S���UϚ)�:�UX`%5�V'V������"�li�	�lj�-�.��K �	�B�Hi�f��ʷ:�M��NsL%
4��}}^�_�Ҁ`�cps�&��v�?:y�A<BX�M���5?l�Rͯ�D��TdڬE7��]�pRJ��T �a	����KJ����"f뫔qn8��"���?:��QKVLyI������"���J�A_)�q�G��o��kZ�Q�����*C��Dz>>�dt�?���cb_�r>�d{3���l�=gf�9�����!�\�GO��HW�
%w*�~�Sf�y|�+FҚ:^�?�vt���I��-��l�n �b{L#;��.y�o����q�=�7��j�"Ebҵ�ߠW��)��Ƞ�!x�/*צ���"Ҹ��?����πd�gƖOͤ:HRp&�J��п�/�7�am��m�j�DN,����m0��x@)���ˮ�������s�䅠���o4��}Tt�8��ˏ�d�:�z��@���l%#4��=-���� �_��`� 7�&��j[ ෦�=��K���9���%9M���9��{��4��AWTV���"b��(��-���⫌���!�;-�)ٳt��O~$/�!`A]���ި��r�4K�{�4�{h(�y���%	�~�i�`;r������l�N"=������Lx"����T�̼4���B�gkC؛��dh�"�	���+��%3��{w���z&e�5���p�E]Kݤ$�<��LdC@������������f�B��f�1�.���Tt���X�`k�-��'��)]����Ohy*�2��0��@�.� u[�Tu���d�}d��m�<�=1y�\t�(���P�LT/�^�CD�<]��ޓ�����x�߇�Ds��~�Ƴդ������Q 4�%\= ?��`���?B��r�5ԄCm�K��ܠ��iu�٨��=���f~�����&{,�˨s�ۏ,���������`�����򱊲�R3;!JR����g1�ƿ�C
��:�?(���\�;����҄�WS�`o=)FWa�h�p�8$o�U}4ᜂ,N�s�r<Sp��r�����r͈)<}���E�h
@!\����x��'+G���
C�����$�./�L�f�0 G��bu4�tㄅ0�B{��� t�+� ��g�
���m��C�X�-5�]k(:b�I�ey-��Ht�>r�ړ�O�bu�6Ղg�n!��&*����&��z]�Y���P:n���2� �抉C��[�Dшe��?��t���9�N���hŐy_�`X�3j���cΡ�^���պw�]������̟�F���9�|���|������r�$��˩��d�+
��DZ�G21�\n67t^��Ǵ��k�fn5�s�~i����$��	��ʲ��vN���#�!bb+�?O��t���Ԟ��(���+*ŭ F�WP��r�/e�Z�ڬ/�=oL�� ���"��;���fC�#���"h���G�P���ǜU���p{������j�yr�\�=�2@	_��NW�ם���Z��5�O�O�W� X,�[]w��1=E�����]�s@	h�t$�a�Z�YHǠ��?��p?���nq#��-��=Ȓ�q�։�цC�����.K����,��tnN�G��O�A�z�O�BG�p�{��ޔ��\w�/�Y�����oc��P8v�������h���δ�2��o,/�,�<Ɔ�rm
u��W� �*f��;�_⅃�CqP�5zN��׽&�Up׉��������8UU6��yF��(3��R���Mt�#s��J0m�,�[�\]��-�YXa���T[R�l�Pf�6�iT6�qݐ�?�H��j�Ӝq��r����x���G�;�S���F�8c�[�i )�%��}qekH��7�*��@w�i�ƙW:�T����O�,+)\x||u��~�Z�qH�!��^Ȩ���à���-��;�ja%'�6��E^�3���l"T<a�((�`R�dO�����"���N�U�+�S.�sU/��C�p�4���,1�zE���a3���iaC�^j����ő�d��ox٢m���R@8�42lW�ɹm��
�����&��?[	��� �WP�dC�QS[��_4��|h�K��b�R�&�N�8_q��lRs�K���貂�XA;�&��ϻ��E���z�y�?��L�2��
@�8���ݾ6�vzՕ��i�mI�3e͐�Dl9h����i�����ġ��������ؤm�_K���3�����uL����@?�����91�4Dxg@�ZMw���
G��*_�����K{�4��(R�{����"�)���
������"o��Α��r��Oav���hMv_�Uv,����t�,Sg���*�v2]�3��)$�#���ׁ �"��]{I�>��*��)m<Ś�80�R��umm�/��\��In���Mـ
�%l#qW�ӹ�����5c��W�HA1fM��*�(&U>��Y%���U}d�"��-��0���+�EB���(>����i�ەߔ,�F'֘