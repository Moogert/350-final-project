��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���a��
�����]�1uΩ��!ܻ�tB�H�!s�O�\
.��V�W�}� g������*���Li�ĉ�3���R�\��0}��N��i�b�QO3s��N��㐝p�W ��Kl]���BI숹�(�a$����=ZA��Z��<e�TrRd���t�o#��K7�QX3��O���� eT�2j�Ŝ�5�| ҭ��\���I$��Ng��^�i�cۣ
,�P\��B:�CN� z���� ��hc��GB	:b�[�5Rf���il��.Q��</4X <�Z*�Zv[Sr�w�P�����˘��C��\&�η��zR��bA�AE�Y�w��\�7¿ȣ���p�A
 I�!�C�^�@��r�>�����.H�"���t��}�k��e��n��(m0�)?JYk���:��&�N{f�wLo5���X�&�H/D&��e��'�g�e�x0Ҋu ^1G�p��U�y�z��8U�L�q�&k��7[Y��K�{ޤ�.0������K=�m@�m�s6?�\l�$ӡL����;���z���,-�	r��]70�ߡ8@n�_���
e�`u�]��w@ﾒ�RE0Jz�Jgu��_�/���Bj�>#���p)v<��]�j
p�C}�����n7����gH�Rِ|\3�z����eP��	�X��o������:,��B����G�<�K��~����ɰB���W���NB�֠MfX^���!�?��{^�Dx��!=k`Ӂ08.��O?ٚ�{$vx�HH���OA[��(iX/�|j��u�p���J��۩�?&��ZM@&�&��H�&2��uy�
�k68
A.�b�G)ꅫBh1���:ab|��؋R+E]�iސ��h;ݟKBZ��[X6�jy��M-+s�t�@�������AY��ё���F���e��y���Zm�AfAB���Z ��Pl$�E��\y�׆圄C�N�t��pu��H��l`	��0�v���4��x�-���a,��UMxBL�F|�e�M�)�2���-n[8��"Ljz�(��X"�2�i��;�$)d�m7��=Ԅ�ك澨����3[��7�n�@uo�*����Q0�Q$�`�
u�%:!r5����D��ǫ�SW�l�����[�3�����8:�M(>6�Ra��o�^z���(�k�6��~8ȩ����ɳ#v�_���ys�銃��l-~�K䥈�G�8�(��p<�ȜT�Y��ĸp���r���_t�B���xu`,Y`�3��]]���>ӥ�G������F�B���
F���D�N��2���!��Q��{x�78�.c�*��f�ȋ�ي�騕�K{��3�L�.$Q]T#Ơ�`p`̣�5z�G�ŧ�#�js!I	!l��izZ�g����i������Z!��V��N	JE���Lk뤟L�"V^h9��dJ�2`�?'�FK�ʴ�wD���]Q.�����f�䄒;4G?��ɣ%飴09N"��B>�ɑ ��؅WjAhy�H0��̙~q�gW
>z�ٓa�8�Z��K^�I|q���?�_G����#��D��%8���jМaOrT��N�ۣ6|��E̩�e�^�u�ijom�u:5V*�9f�֊��8���^�o����r��hl4��[W�oz8\�ȅ�5~��+�ϕ�>
�d$�m&I*V)����e�5�u�c�-�@!���~ʦ��.�y
���7�/�7�nvM�������0�.$sD�"7�z�a��Q5��R�L��pg�'c�� 4y���d�C"��,yfIY]�
�����ͫ������l
���ۊ�}aAp��r+�&/۟U���%�\���ƫ��BJ��7�6�A8��� \ʷ1)ۭ��-&o	�qț�L0cEI�Dݭsl��(`����'i�<�\$Rh���4t>?���	����ǘM�hY�h�o=:�K�-M�y��Ƭ��֫�0i�� [���
�IE�c���!�{#�#u���n�C�O��c�k)J�����袟�k�ir�=�'��K���L+�=ۀvN`�������Jr���������^G�V���(����+�a�*o�zq%(�	Թ��s���2jPx�0�9��-5}ǆT�:��܅D^�M��u�t�mM�*�Y���kmMH�U.F�6��r�E�5Y�Q5R�#g��.��@�\Il��#�m�U�H��������%��*�FӭCF5��t�EB�`f�Xd��q	��ad�$�o�����iRa-���i#%7��P��E��j��T%��vq��'de���?6�wm̇��O�Xd�4��q=�	�
B�`V,#�݅HxT�{Y��5V��|�un����B���{��̪����������e�GI�u�T!�Lf���@�&�2��L���
��uk���Xel]Sc���n�!�v�lGef~~{��|�{aco����oZ����f�Lu%N���X������o��8��d�Sƭ�QT��w�l8���Կ���{[�$iq,�<?\f�����^d�མ�ږ]9-�B�ܮ���RlH�#�0�?�#hXEF6ꪴg1IL�5���I�R��m:���e&����	I7��V�����(�OE �C0�ߴ���zy�����p�W��IJ��e'^ߨT?���#$BV�5�PF$���d&g)�Y�q�U
��'�%X�?����9�uw8=�}�c[>g���E�,缢��Q�8u^��]�v�5�7���@:���e�o������i�H2��>���x�Е����,��[P����D���Vlt16�p��|c��K�Si'�ӹgG�-�C��Ԝ�0[*`4�<8�
�����F>��p�,Q��!���{'ޛm�4EU��:��"U=����>�h�='��ց4"zUe�0���S���%GCG�06�z�%r���x�*Y�8D����s�·����n~���<'v0�r�:����ʪQ�+]W�Yt�*�[w�K����/��7��0iP��UM��Tm�w�E��m�@!���yΏ���;tȀ�|��*=Z�K�`��!¨o3�Ǌ\�?#Ve�ȑ�� Q7�k/�{1��%{G�Z����tb>�ٯj������+
�60[P�`ƜJ_��cy�m��JQ(�b�憍�V���r8�/��M	�@$}E��؜�lI(���.i�[�>q}�E��O�i�OZ>��KQσy9��d��cZ���7©�٘Q�E~XK1r��l��9��0�_��m-���R�p(��]�w�^#i�˵AY�{�]��KGL0�77��eO��3a����o�Г�/�ޛ�>f�����R|xo��>n�8�_Aru� <2@�ŗX��Nl�#1�t��u��C5��X��0����M�i��&��<-�b�|� Ì���_���[מ�V�&�0�	�]�u���ɟk���f�.r{�].���������+_G�ǃ���*	�/���o��r`4�R�b�79�|�X���q;�	����r�!��Y�Y�sF���Tnf�2lV�����HZb,���g���㶠Sn�j"lѮ�i�C��I��o�yn�x,��~����n�����d��I`另q��{�7���5��:A��T+ql�uy �V�%%�uy����3�&��l�(V�9�����t�1�Pn��IE�r֚���$/Y���q��� B���/�R���,�sG��h#�:�`|H)���]��Z��c��ݖ� �n�ҕf���p�����O0���(����iw����K�6/1�,�@SU����X���0s��8]e�X���*ؚ�2��O�tL$A;?�PÅv�r]&�DT��8*�erݰ��d�v�)��]��S����Wȏ�t��l	�� ���셚n���@)Ҕ�5�?�G���ۥ�s�B�{�GE4}�r��E>7��Hw��1r��|X�>�/y�R�g���t#^�(D�;Zͼq:�w!/ر�k��<����R�]@!�P�P�Ɩ6܂ܨ��p.9�9�8�T����R4��#��x��y��A���w�XH���,k�g�{9gXUT���E�5B��Ac�{���z���E�]��H��_��yai��PD$���۝;=�zw9;s�6�<��?�Ը�%�ct&����φ�ꁕ�]~x]�ȅ�ْ��#��>�[O���H�� �2̤�x�}����ǅ�0� ��t�yh�ǗK�JJY���%'OV�;9k�8b�L�p�lNj��@i�&(�~�7?��Ʋ��d�a8H�y���ι��B��<�'! hl$b�{	�_�,tpD����m��!�B�~�4�_wQp�&~Q�3��Hd�,pͤ#I���Յ��쬙xIt��ܷ,?�	}h�uR���Em��c� 8Ў�������,����Dj�v�aQ�d�p�b	����ջ.7�=�vqX�����u���H�Z��bC��� �Ȏ4����fn�ϳ`�F���)z��!����7e�����'PgT�0������a78,��MA�ۚ(&i�� �肩uTPv��Ny�R��b���1v�fU&Ds%ZdӔ(J��FMG cg���=_
�;��D"m���c03�%�{[U�3%�%�4��G�q��L���<����"���(�=���Z�����uW%��<���?b�{��̺i����V4�*���Eg|�������1�/�Խ������}O[zO;zܽ��O���j�Wi	��Si�͒�M"�l���-jW��hS^���CY�*�x�^
�l� M�|�j$��!Y2O��Yx>LnK�� �
�g�a�>�pz���1�'D�^���s�^�Q 4an�fQ� �l=�I����&��.���c[������/�x$�/qL,��po�V�uB<���?4/�!�H7'�׻e9���ܐ��M#�X{h��1= �-lGJj���Z2��+���.v�jP�\f�'�����Vn�/>�'��B��b�bV��%���b�����YI#�͗���f��r6���Q�n�5��;�,]�����
 4�Vݡ�8������Ic�{�:�]v���m��񸙞��=.�O�����'�?�;����ڽ6��Msx΃�r�4jQ�'X$����r��7�����z�C2(�����'�����]T $��L���ٙ�Y�.x,:q 8�f�1o�����Ig;�W�㼿����wl D(x0���ö�������!������Qn �Ly'��ˮ"=�G�ԯ*���ݑCw��S���|���1��_���%�\C0�E_�5�
��JV*��^r�%f��p3�W��bB[&>��aK@��!�uL1���e��rg]$�Vș~�VGG�uN���x��DvJb���we��RO4�d�_	�_�:��B�렲��ej�%�8�V*�$�!qKPX#cb��BZ./��m�e��{L�T��t����l7��-੣P,JrBe��YikU�m�x3������1�-��0�=j���}���w���_(mh�ҁ��,+[��db��N�q�)2Ǫ�=�jW�9��м�cY݌�uD�lN����~�YfO���-m��Ca3d���\d6S_;m}�����L۸4�����KG`P�:(k��XifwTJ\+�b�Z}H��V�ޮ�Ƀ�y<i��XT��PcX����]�n�pa6NUM&�n����W���.%��O�`s�+�Tv�σ~�h"�r�ڊy~20S��9�*��v%��l^9��r�H�@Ny�_ �Y���,zZ't�����L9�2����6ȇ�����b�)��H4~4���ysN���ɽ^j}o���B�.&X;&����<{$YAR5�[s6=2UZ��/(�[�Vv����	6_��SB��Ϯ��Mu��S��~�9�"b|`���`W��Q�(��MrFN�k6�٭�G�;����} Ŧ�x>m\?��]�g���_s�+F_!�,/
�8�[K�<�������rD��'Iܩ�ވ�3{/��{i�I�V�T�4ʂ��n��HK�(�6׈�U����g>H�'�!�^3uG,�Jtc(7�Ǡm��%��� =��)��}����e�A���u��=��:Uf�����CbBo㷹�����=;r~����a鐖o��������0|$��1\/��C]հ��4&Şy��IZ�_v�
j_p�[9zp="�Z�䋑9�!&��Ѫ�a����:t��s��i�y#�%��00�]%�NoV��f�H���GN����M�J4�\�R�L�,7N�P�sTљ�KT4�g��f�i]xy�t�NcX��� ��Zv3�G��'p;����q�<�j������Y0�DK�b�bѽƻJ���$-��>	l�w��H[P�@K�Wi0�L�Y!�)s�ϯ:|��{��%���<h��v����ՙꆠ�l~�����K��\+u�;��"�q�0�,�I�ܛ���a��y�ߢ��v�K�R��,�3���g�tkK�ٽ�n���Ҙ�����f=o���7��er��ߞ�M��cp��*�U����W��n��׶Ufۮ����My���Y�K�Bً:P�4Zy�M@��"���e����&��q��5[����A�@�L�P{m�
���r��!�;������ǁ q~�ĽR����,��U��<.��ɨ��?�+/����X�T���!+�y���N>�౏��,#��6U�����t�S'�9����$���E%�Ks�P|���i�h��X���b�3����f����P"Q؅�J:��S�k�˙��V
��!��p�T4�K6k�`P���z�����~�ɱ]g�}�"1WL�c�|��@��cc�YWɃ���!t�Rj�� Ŧ�Vk�U�z����;�����;c����ȉ7]]��d{�-uCz���b����6�<q��$a;��_|5F�hh�L����׉��O���+�Q��R3v�u�X�w1�/���WÀ���oP���7U�qG�Gou���D2�ӕJO�M�|�E'��Y(��6E��T��}0ņ��Tq�P5]��C�o �t�<`�h$W���k�����[ab�)D[dS��|��&'L��uȚ�~O_�T���$+T�3�o�1��A�Չ� ��a�&|2/ꢊh[%3{Û��&e��� 9�/��╜sܦ� ���!��N=P����Ds�vl�+���(zA�Qe7(`�Ң��G_5���-7��$@,D&�#%\}�]�86��}����EM}Ah>R����a"�����_�������.�҇�o��S.M�1��'�d�@]�[)�������ho�Ҝ���+�͔���������ZV{��a�s��t�n����4�L`D�M���Y*a��k�����d�jw�zQ�[*�)�d�����kN�ՕB �$T����>"�O���/�?{t*o��@��)_�45Kre(��J�
��ƛX�K�*����	�`:}z�w�o�Y$  "EW̰>K?���JA��:~\���k�.G>}��[����|@�17�h��l�z�y0͹`�ǥtO1L�������C�����ꑓ���1?�~FN����σs�$�Ô�Z\k������������D��!h�����:� ����L#�ʪ n,m��E���	�>���&5t�F���]�Xo��X��#kH��M�}�D��;.����k��4���<�͓g�>J��eRcCy�E���6J�G�C�Aȍ�d�☻\I�3i�ӺB������~3��{7����:*�	�_K�4�F.��"�MoŶh�(�Fv,T�F� mT rA���ؕLx
V�b�l���6h�-.�je�}5�E�i��}x��#o���4��5�"N��gR�á\��� =��@�ɸb�2	hLg��2篂��l̟�c�I���/� �?	�IZW�XZ�ޯ�N1vx\����mY 2G˜�,[γ�ϙ�[�iZI(iS�'ꏳ������&�i�\N>FN�v��f�梅0�¯~i���~S���F)��d���� �qd(PD�V-�/�E��Li����N�y��4�W��ܠXC}L�-Ƚ�辍��$����Z\A���b�m?�}�Ä���b{�I°*��$n����p3�$%^���i�0+�k�V8�p�'}nM꧷���2�:�n�7��Uz��U�Y0$)���0�@'&��$��ZWY)��ۤ��"�.�K@E�q�{~���/��p��@y�CK0�4�B�b���Z����&rKk=4�����#������鐱��̫)��2-,h�ߡ��}|Be7����i<`6��B�B@��6@���1е�}@#,K�ě8�l�jPD���v��&�f��|��,]����|O�����-^j�r�B�� ?ς2k�<��Ny3�U�3��^�a�v�6�!ռ2��)� �"��	��X����L�F�o*+bN
媹����P4*}����:�'�|&���{r�D��O��%��߃����:~����_��}�8}�;�.6eV���8��rB��ŁJ���Pl�}�SBW\����ڙ������v�M����u8��|:L�?P�z�	g�t�c��İ���Q�ϐ6�2d�R������%��>e�Ku�S�r���;G���u#��0d�ԙ(Z���Z~�k�8	��+��O,��jŁ����W�F5����"I�xy����0�1cu/g�@z3�-	a��T���W���]�\DN���`�ŵ�I�=~���_Y�Ŝo�"߲��~n�/���|w]O��m