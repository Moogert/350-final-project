-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UIw1u+ORQN5V3HNwIl+3UP3KCO4TFbBVQUyveKYT2qO3HNYon2/802FL7tQRAe8FETRsoklkSXsp
mnQA9ikKMySEeCenaIUKi7E7INTagfMwjuFmT7PRSypa0dvS0wMS/FMydsG4Kf5Zofhbek+eXdvy
qx0l9WChA+honYPa23CmwC1QK33nuUQOdiC9+CZdJAytjusLqEyMyJsRdMyC8Yu3QupBfeP+61KI
v4jyR2Lub2Z1LvcTwfw9NfaITzMFfiosWPjC6sVjS0Y3oDqIP+jg/4bjTljgLvkngymEscd/bk4F
E2sczxOXdfmbi+cOGhXNRzj7Swp5q9NgS8Sj8w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3376)
`protect data_block
+aJVQNhYu8NE2pWmNnAEBUZr6A14vC6azX5VH/f3TTylMvbg1jAIINBqDxXvrKvPMmLenf82Hfho
IKaYYC5kP9/viKEGSARyssGp+JoJCCapJEoutA/pzWsEWFzcuKMeyrzOWZsqrdaVsPq8GrhF4pAB
lE30ftKm16J6z2ZlosIX38Tw3TTZP7ckc2n99nEUFO9XFoak3rXYWQwgcyfGIpRI1Wti+8QrAQ0N
pMSR6fiN/nvPpAGmxTPQ0QbS+yrkc4i/AY3nJ/UVtgswkLHoXKNPWrvoDFbAAeRYSAuAso24pWGP
6l3tIiRqsurx8paimLr7W8gRdrhc2qC/9lKrBDI6BG2ba++TD136TMGcaVzFLMrnrXJ9zdPngdMN
iMRYi/ROknDXQ8wR6v7JntOuMiATMB4lucG/SQq1IOuPBMgwr86H9Fteqz4DaFdPnmL5dnr6GlyQ
fGZjKdpVs/6mzkiRM4pyBQiexUDgZsV8lON/uD8QX2KDvSB2dJeKLS7BgmEZFlOcI3s/F/Nx43Sy
OROtc10DQh7sWK6voSVQSbwJ6i8PQ68QOmrrT2V/9QpqRlGPvi4bbK6Neycl3/EFsDGfmxGnhs3g
oOvbB1/4UBJoD8m67V9MpohbN+wALkAY8R+SzEfy9Y4sOqEZrXlak+z7YraxQoOwXxZPtJDXFgbm
Rnpli1ozAHgNipnwREyppmKELemq6TNxRkCoEHUEfkIlDZ/fvbLUuVVmGq17cwNg2xQUKgeTHme8
Jp9fSlDk2nP7SkN1tLOoy9h52wt1MXu2rAbNmK0daRDtsc0haY35sfKmqzvE5AFgyr9zaDF82LmT
Poc1paPS8nYH+o4YtqhcPrbzVjRf0hatoHe5N3IDflINoZ0TGltPdIpEgWCyivdqK1r9EDRkOe85
5/oTiJd+0GHFXvC0isNSt8VCx5mbRLM+lu/tgcVOGj8LqgJvPl6DsTntSqN73Y6J0boA+1pAKBPy
heGLPeNMtEd+1ZR6X7Y1AZUXuiBi6fYNa2CFBaIVpbg/LIIjV37WchczGdD/dbK3Q5O1mrl8ayLJ
K7e1d12PyDH+phcYpy3YOhaBUNuFc/mbs0s3TVx/6f6GHAtUwkKK0hOjylxF6f3oqH40xKBFKPHw
jdihnDjWKLv8OiV6fhPuGfqsis/BUiMVK4FwRKM2yrLvwTj0uucRHdckeKRyHthSBGi2w5JYH7WF
ZK/8TedaoNX9VfLeNLcwDUbEYxVyzwXruVe4xpIdC7X5uz1czA2bQXIazbFOqfkkwQOHmjzbph3H
c6LcZ0s83yJ/7WFPhDM5dF5j3z7GY3Rt9Q6TM8vt39BMKvXqLmvOD4uWS7NJvI8VhRHVFnyPYliV
Vh0aKzYCvYVUiUMbTdQXRyUpoUKUq7O9bW7v+TWop6o9HpRddX5Ps1xcpSoZN7KtZiEOO21GzKMI
hrOuROPJnotK0s/zKcY0i2U5Zqfn72McleII9Mo8oHUCLcLgjTTCkaw7thbDgnA7Tzeg5iSSZGf8
zzGckrwxhxHUvP5FygT6t8+wuadGa8F+hBQVdRD62aoenz4S+z7+tDpr3TRVqjzm4LklRcw4Uc10
GAxSmF4766u6zi3yMaaIdqBKNYvv2qTzNCCJkYPqnwMZahlr6A+3NBM1eXtfy1MwYsAC5PjhU4mz
NBd0WPCXNzW+kMg2No4+WX077N2chQoRcdlPEDk0quYWqKCL8hiAPSiptDOVKjgxZpeN23v68Xc5
MPmW4lTv14Xe27iOu6DZqyHyA7YER0bdIdEmZ+Csxu5TZ8sIZ+errPgQE+YNT0PZhr28p06hgCgk
GPdCkD+dJNJdswVpomNxgk50xuAaZZ3SdwOQHYRpzmof9OMenoLANEynUrX4Yx6lCJWIB61uf8Cq
zyFzb2nbfcaxttymqgCaDYxPNhF7evySEaqezHGmv43uHL/9kRc9nNxc/Sd2cTgtpGud3gpqaTqu
APPsbVYpD7Edr9IUatXqfW9tLAUcQ2CThKVCt91aiS87mBoIRWtJQQQmtNDmsHc0Kn7Ms7R90D4s
KoSPFBUmtJpqC8ZmqUyWVyckgVEGe7Fq4hHGXlZjQ1GVeh2l6Y7cSLjNiUIriARc8u8RShbKGX71
SAFDOmT6jsQOefIYgOaGQoU56dFJthvUpMa9ZOR1fi2zqPp/z9hkl52fMlVzaHd/C8op30mONG6P
mA8bI4adoGoNQiKHNc1ai+sV4tMPjX/sCyyZqcD7MQUvhN7/Zbqxw/QXS9+vdlfFa6eeeNrsRK+s
dqEhoXIfuDhnZWRoWjlAQKR5TsT/DAjbxzRmPUE7lKFCog2xmRhjEJ1dj9u9xZYCYtW3eHnFtGsL
3dlHvb2Dys9aAkwx+ECtqOZ+hJe/aDvbCcj8SS1wxLMWJNVQlphWgVMjMjm885hWljptfbTHhZW3
BRfgfLhu9f1mL5whMmo33KzsMZw8F1Q23dqftVyAkOO+AjDjXuvRMSZjKksoCONDi1qtT6Q9T05v
z4ZzpVQs6r0nD9odipYbKegCDyQalmrB/A4OeZjkxnbtX/iN4mutfgG4iKX1lS7pcdJ/k0XYZsex
A4C1s4IZYlIXiAaQFWuTfbcPWNYqvVUDbD70dqcQEEg4nraz+LPPA5lU5QvpBT5GqgdbhmATGPs0
9Uj2oZ22X9UGYAhqRrHaNoP8pmNkgjclzq029gjFOYIfcSfqhbr6BP7frfMh3fB8Z93bD76t2oI/
JvELsgm5Uvsj6IoDbDvvrNSg9kBX1dYE1JSQ+CdEvzqHpFH3C6VayEjbq2aaKxmsjPBHuULA+CtI
M81tWCoqMbrVq5Ccv7/QwO0xbLjjwtsp/XWINTtHrCp2NlQsy37Naggv2st/ekg0CvTyWt0BhBzY
nr4jKRF1XiUaUYjsD4301PdgJ2cgq9SllQc1k/Wk1cyDPFTsRgP6A4n4loj8DuvuOgSbNSlcD850
qBvABWmpbTvnA4Rz1wTWFUzb9yWvfcqJu8t5VZQUscBjr1t7jWozLX9k+xvlyh7ixr03vrI6MNv7
1k652hZW96smUuj4xmabQvDN5WNuUnrtAhspCEMru3ZeUFkz7hAriSe9FLtx99KGVRzuPc5Vs6+V
qPWeMUsPiUiWa3F0CV7g170Oh4fehmSQfW0G6T0bsSt+F9k79XzekD63yDGVFVBHGK9zrupjRO7X
rBYpahmOo/Yf3rOaAmkcZR2U4EPV2cHnwnoB8rvTprlUcRmMHDm8qvXKVgSO+vdSb6nVEqup6WBk
afA0DW7dKS8/n5uMuvw1iucQQ3bzg2vkReea0YuKBDNNv7k6VsGWdUfu/mOiVRPUox/vOj2Xdg6m
OGDsc7CyWIdJnsE0BwZ0NNNhLx4V8Ps4sIyg8e+uIwaD+T/Cde9crupP9mNEr7xEtK6qcQoplmu5
8tJHU7U/Jjl5yYBui07djRMkQrrj3rke6K1zdnfv1Enc8pucK3zekUqM5CDcwJGPmWdyGZ7nW5w1
VF26TwuZ8jsZLLC0LEMyL2kuOM9aCqZvm+9mpz8AxBu7kqrN5mk03KTlODk5sYEn0TlrXljdISiE
TmDA1dKRUXtE51LQgUGnQiDEoCoHa5xUNd6MoYK7CbpS4m6TmIpDtfgOr1rSO2ZMeyO4rLVuT1Cl
wmTAvtvMB6w8Egx3ECm7cHu+Gd/gm8LTJ2W1bZdy+uvZEn2JAcRAIjx7XEPkoKAXje0aSsHbR8wC
4CTVuv3ry+wKslqVZU8wsjeGrH1yQsDbBGLg6ooQqk15e7ZfZmEUHUdxS+/6MD63f6Dbg0nJy8uZ
Qx0eSfhb/HKGRvhFWoVBqXjwQy5TG6mW60eYSgqGT57fHqhcbeMBoDGOMXBRmpjrgSBI1dgwlrBx
Yl4T7E2LwZgULHXNb4Vbnur5apGA9/Z+uPRwAlB4k5bOgzMkWti+6dVElcuRWrYHKzZGw9UBBdD5
yCFkceomdKguxqZGjxyL4TzzllGTn5zANacgwzKHlRSi3n+zZz7d7lZR2ZtodeymzYth52d/JhxE
b4rBFS8BHLN29AM0Ai2v1Hzb/GkfNsZbfsJA9Pp2niM4rt7oFnl0GmXjY02ldruTs0d20b3qv+3D
zHWszNq54yrDWfqx1aiT7br2Mj0zEWeh3Ulrsi3P6rgMqDZhlcIwQUC918jpS722xIGSIsvM9Ef6
pN0JOURrb7Y3giB6YPof0njws+yccUR+o/qq8E3tTNv4agA//mHG329i++eBKp3z0wcRJpkp9fRi
aG1eTXp3b3/WVqGPjwTqc8CdmJuzXInMLCj/wijG/LqgUAB9UblZP5aeNLaWq8CNaPrwVl8O1xXF
0BFzq999ESygOPCeGmdfG7mymHSI5jqnAFcbsw8aXVXvLBX21RJnxdYCyBOqRjF8eaaA88xUkQje
3crqdl25MxIQZHcwKetkChJr7xnTozZ8WQbYxlzu9qNh8dbUeqO+BB5aMqEOgkyFqYGFkY2cctms
7GrbDfRCz6U5/rUTkQ==
`protect end_protected
