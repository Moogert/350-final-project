-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XlBmSj+CEB+FFm3vox6rZBiu0M+pldZB5fK2NYr/S9sAvgtOL5gFkJH0i6E1i9a15cC9p5kUVu49
MHYnTnEs8veZzU4Pw6sK2Oe2DHU/qK5+oXJQ1b87CkCq+W4303hSoDqK8v1AI7M+KNzG9N2ZElKq
+lnGRxtg54CEfTSJ9/xl3gc+MtaVseZVL8GLHqw6obIWwiwcBGWTZdd1k+P/coODdvF4S4TI099t
XacsiKuWnDryWP2NegmEgxLv38SMWG4cAqGAglSahjUh9W8UJT19rDp3FrBXymz6+/RFuos9qtdE
5Yvg6X04Wq2c42Ow/X+yZYieV85dn/e1r9FoXg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
h/Dz+6sGIxd+iuK3kAK2DNuF9h7JHdFTIRwNgwN8oyhZvLiXue4s68t3PoDIwFZLs/OATwk10ZXJ
To3Ps0dBfPsa5hbeS0EntO8LSVygraZyAiWSeKo58BXjYryzFVBj7EgTiMmx9vb9xtDQUdTp0JXo
6HQVonvsXMy/3VIccP1WDjP8v28j9NfaQ3ESUIdTylBIgTIfAK7vYZ4rlPf8aBqYxWMmsll+0emW
buOSwHMnWwPImSXnKCPNGgLAXGwbDX9rFnop/ydrVlFwudvhSq9rOpVg1rSJqiKERh/s6rp6CBfG
DhIDCtqyqjfrin8x0k8r0NX4W0gn/YFxLxYwlLx208ymKHSl+kbjUWsIVW4lPtCo42u6Rpbt1EiA
lwjnTXP+hgzA+XH/2tJcTAiSNTI65P9w99970wm4VMG8c8LzpFDZMHYv5pnXGgyt6PBwUF4RYnst
KWGHxWdLJy7eyLjvzL3xAhPdh6Ieyjuq62lqJ4Ex41Fh0t534XUcZ1m5IH184PiR1UAAb4hB56QI
Mji7RwAG1Cuc4rMkd7jZQ2/5JDjdvE8nvfgX+KtZ0WSqVmHliiNbhokStBVs0hQ/bwJtCGmrZstQ
CeMnUAbh82Kfu+8SexB8B4YXlV9Y9L3QFfq5+HaDf+R9HI527ZYy5dT0FIDRcbSuHNnrzt4bBtbw
MdfGvbe7CuO52qS2ppOmt7PrakJkgxYvKwciIIp9KBnDy503xyfBMSRa8pCF5k/fOUvmOCkXxYsz
QgrTJl8ZRcQJ/f0uyo7cdGg63MuSfjB/msbrZkOD9jqxwndQPd+HvKJbFx/wzVqVGU8mjRc2VImO
J0Bk4aHC1UeMPbfhy9VPHJOa/DSQRB1/S4cLqAGwXXupo6L/BOL4EQZgalwMA4/ZaTNdebClg7VJ
qGKzxVXHO0OgZ0zbet+ZDsKo3j4doe2cjlRC3ZMepgTpD0veAuBsgDjj0UfxN/pvFYlr45tfKbXL
FRiV+Vbd9oGpME4paOPBdnBGvi2UhwDKfCauTiMf/3xH7dryRUvbtO+s57O7qFdN1x3pRViO/5yf
50YHHhIaqA3WaC0pu7U5E4IUD9Mhyc+onGhOifFdNWnyi/GXJ0z1hSm5/0Zuv1x4u7vyGQ2yl3gg
7YFY44rhU067iIoQ9nljIbWkpf1gCVqWMoeEe8CBpWYW0Q/LwiJQdMBQnMBQgQFlQZYHp3PcN7xa
nA89fnKB4GFJbbWQ1K1JAbLtkdljqv9touifQexN5a2yKy5O5ptldVKDmAmqNhZUGzgzbWqlVhAo
g4hSHT5X/oMwS7NdFJcvuV0e0JdiDDURav4kS2v0irdxmE6W/9zK6ljy+KQ53sYLM4TGg1Ekf/9U
012N6M7ZL6c61+Ie4jMqMSbVCWEdt280ptIDhgyGKp1NCUCFBwtJwLxN+neyAnO1ODhqgjJFuDoX
6pqrUrUNVs8lfGd+KTqh2Yy555vRARQqwORjvDFoQxscSaWC9hKAK9X0BFGISWLUCUaYkVYR9HUT
Chuu1eHoj1OHTP41Am3gUhJxJkdwZIxcsmNtNPy/L5/ND7/YsycVjAvZ7RmHTqQOfc2zo5SH/hsW
a9AEp+i6WKvkV00EU83KK8ZflW9lRnFfAC7FwkoF8EfI82SASW53nrjRLBSLvkiJHz6nyaidXg05
AvUoH/AAFYB6tQt30bMRoeuuhyH0AQNa7QYsYxK7VIJ90DXiHX88ojUojMnm3498dSvWQZOWLsBz
UkBvYBgLmyq0Mvz2ToW9lFCnW9HUMEXS/UJ3qdU5rpnIY81VrIFm9FucfrQMAsZR18UhYA4qflb7
l8PpWjL23r25gtmp+/coq7Zk7ueA8YESRtprPjfzSO4o1lvMMLg5svLDJ1XtmG0qjw8SBjAZMp/c
QkAEoroi8ieS8ayzhojs8YHOVLCbVsThjfnZDbaVMWjNYuLx7Urk4CGli2kh7JBaRVtayb9a1eKH
58iJRe0aidk6SI8zQalWv5YODHJWiAvVttoONQut2ywcPGAlGJHnB4NLTcCPe+FDXHDJJaOOXvij
mL04YWZyq/ORK7zFoUyht04r0YVEe6fmFkKmtkWh9AvLlW5D/TDV7/lbkPPE2wXULZBtbHfzRs5s
CUG2o0mdGAbLRC8/+qCq9hbmJTSUgbukQ2ftfRfPd/RbW3tBuvPs3BFl18auwR6J7lbUAOUp8qDH
W1XnUvSXHX2ifTShXExrd40XNrDUXr6l0n/Z8LtFdPWA4k4+TTbHnFqpKMun8CH7HIdr7z1wgd+s
cR0I8wpox4fEHul+NJu7SRT6W5qq2lm52oJBemTLjghyBEfa9WA9zEi875e/mIMIRB9q6PJtnVoL
irUKUaj/dgqwSvQ5ZQ4B/jbg04F0+EzrhtK1Z6TZLgiRRswWA80y+y9egZ7skvvzE+DbEI47Gr2C
fanDLcAc7tz2QIkgkqmNlPOyrWcruwDK6imHWgU2MfPRe3ejTrwfywrTsCKScsMbkOYWRuAAnmwS
CWTw8OVcW+xCK/LTKWo2se7OhzjUdI4ap7eWbgSQ1wGWrWgiYidJkxuDJcaiL2zM7z8UtNvxjy9R
3Oz8ENXMePVFw9h4sWPrMwgYLUM/R6q2pNtu9ODoEG1grK4BEypQU/rAIL6sCVYqb1SROIDQ5vz8
5fxrI1otg54HYXnb6iiNpDICTzihzpiWhuuzMbjbwpZj0/IiPLRKGDHe3tgP0D8HMl5O9dOsM3UQ
UQK7it/bAD0yaAmTJaamaPnrK1CBv/fIecjP4L4dynR5cvNQMLZvKgEytA+l58SRCZDTYR5SyMWO
84gWcSOLA3DhFxY7XV+uqEizwZ7Sbd1vE0tqxuNVgg91a/J8sEdXhSoM1BqDFzH6PLniXOMO9VoJ
5bT85QA/iB1QaFj2s1gv+LLwotGIQA/zY4206lg50j8dE/siQT6Ki7oOgz1b6FvMGAp0hBuRa58/
/TdOMM57raCQSkvEIT7RZLhNLQV01kFR2SFdOWVRMEfxfluUbQEepbBms4RSwn7CNykJzlbmq4ex
usdtVzM9C1YiKiLNmcWRlkwOxUxTqcOteohs3s6GCyyExyJs8CQHghAsooBc5fx2DZyzlZp2OsIO
kOmECx9ftSTcRI76kyJAtdsozkbZ5uJt2GQYD3fxvqGxgWEgQZsSYyFgcUQFN1nWsItms76O8Pec
8/vKX93xTfEjpOtbbcac/BiJkkk8fgh9c3DlycyJWP7/SidzCW8cRBVoCmxY+TIog9Mvxvx8yr+A
6xMiGTDM9fvUxK59PjINZD6q+I5U2oaUcVixJntXmEWOLHKNFHDBJXo2amWB+zchDo7IC6+CPA7t
E6+n5ssUSohy02C/3FL5VBZa4imF6GO2HpQYH1E040x883Rb8x8iZ6lzIP/skcq62XPP4mRa+izn
BOG7jRKsBQPEMWF4ihLnq1nvsZDKG8A7JzY1C8iLjjpH9jvgNINCkFB7f8P1zOJRSUvQ1wN7O5h2
9H/hkzHCoOx09nnm/AdWGqZ+QqlbwmLa0CmELP5B2z5a2VyAKMio4A6xegbsWYwl9N6J9+YeG893
4FexnVNqpFG9wQkZPY1BgVknxr1MQVfW3MHhHn0cgpOlgO8tXVcCNMUBUwMzfOJe7foajoMrZI7n
C7LKFodqCHLKYOomIAtfZeIR34l2NQZP+lnlt4iprRj/OOnAqyQiAI8Chbhgz+eeRj/gLEmMlVfu
nLBFV4qgmllIyY2On5Dnv8C5Qrb+DxiaBM3Py9TChT3VT1M1TFw1EHhF8uY0ng4afXvCNDqGNf2K
cqi56O4RWhI4JnfLwhsgGLC99EB42xWcXxnZTDBV7l/nSA2MKpkW4CQxzeQWnXa3pAeKujwM8rvP
Ue62la/y9dt02iIytZ9b0J8eYjkj22cmPovU6w1LLRymhW5e0R3wWVbsetiNce/bp8ON8rahOp3e
9/n/HRoH7BOwhRBxjdVAz4nZz98/wK7ksBNou8aM76E9wSlKRCYw7mW/6cG/ULVeb/bBlC6245Yc
fkedU8VlvjY6dYBqpjkOiZmMIWK24/SwJpm9+ETosvnb3/vrkP7GA+dox9Frlp9CvmMtOziyVhMD
T/VGDwXR+HIbHJyYSVbQJTsO97ejDNhWOxo8iYrzfdRbNaHiDCro8/Nu0HOlsuSX48t3PDqHhSxA
2fUJRyappIo+E72YlVUVQ8Np+1ChiivGa21bN08JsZcBavChVTi0uJT90Q4vuiz3a4y2kBAmLzXl
fnuExbEdtbQNGEepn2LWHsEkd86xMxSBRuj0AfIV6YMNUlpOXVX2+21Ps0AsG354rLuySrb3AJ2e
cJa3Mtun5nIj8W4YRMc9QVH6xy8I/XmQiAmfBts87+okDJBqqe2hDvAUS0zSu++fmj+BSlIo8R8X
j3t3wxTro3b1CGdJFcr99vO74k0PnjPSBAq4hrgrmTOR5ySaaomrKohox5a1HiG4rCw56dbYLWlI
GZh1UgnOYIHFWAVRARzIN/0vYvcMboQCapeIy4QgsCISL1JBcno/5aLrKSgyZWagmqn03F7Ox9ge
ZAo0w4H7ua6I7TpKmRJoFFIDPXUHPT+ZBuFXEUqqeKXIA8U1OHNhVL7f8YZTcvaWFTcLfCtOGSzz
7fdtxiyoSUFy65mOWIxnTbouDFBfwYV5v8gGu4P0Y8nocZis0o9T5jZCNXRMCEkwGCQ+H1A0i9Ab
YwdeH6A6kijPGhdMRgHYr/bhTj1wC7dGtGeGheFtEEaMJdrayiEkrUuAxiYjNNaeTBsgZshTzT5S
mf2ue8QU9nZZBVTA1ulAuLz9JhSK8x2xPBzU5AnNsM7s1S2ivpO5+80PEmVoTgOspVoF7VT4zNNe
ip1Rtw6DfFpKXUFSf712ZnObIXsbbB/bjvejTshuQPxeMoG/QZHD66hgz8f71380id5Lg8C6JLyM
V0YRSsgjdtNGpCGutYSlWwe3r1ouGK+0JXWq76Tpt0J7aLjL6gIR0kLcKwio3jKOqI/PNawhUUHB
+2FvIJPyib+LdunOLCEseyY71OsPsXUZNlrNOQKZM0JX8HNnW7SwdoY/Yo5AGIO1dnS0FBWUlcQd
ehKor2X2emDxWLpc9iFW74N5F4U/2oqiXQNBZuSK2NfyvDJ116MHyxbcdReVNxcOLqxpXI8Tr5BU
uNHd8bEwH7Oi0wrdkbYS4hIvLOAPXQDqcdKTT4ldLS8hEjwmJNlVLz2uJK4KKLTFJ/AyMlO3oxDA
eX8A3xob3ZTP5qOWqk5ezSDg3k1/xMwr+VH2ulkrYF3vzbg7QNKRc4DMUWttFEnNuZ/zAjiBytCS
kai/aD+HMztJq7p2kmxc1M5MtOpI4HtTwmTbS2LXzp9Ah8aa9u3nxc4koolBrrenC4fUOwo4qQyg
Tga0MxWL3vS+ToJTxaKKpXsFbk/YFpBy7BU4iXSwbSMoRFdwcJ3VKASl8Y6tc/ARnSr5lgj3XDQy
5WoBx2injnkoqJQrlPsasn7d8oenQ2m7/5dm0Q7WLCAxoNv8FKMgtJaHobnc6Z5LcxSuNDDD/AAi
URsKI6T4qoYyne4xTlmeVvW0klsWbIy7rFOkNKtc1K1pq55ReZ4TRHGsk3ABqePPPJ+XIfZPPMrF
Dk5BjM0iTPxM+oaBVagpINjZPLUlJr+1GNfeThppWDVb46qRC6lz80qRd/D9wB8dc0UpOmrlD33O
9PW00BAsF7IgVcUpR7CJqLo5KGgFz2xUgJQoZJFsQ9AsBXUp4KdM1Y5wykseR4NSYldHi+9A940K
FtasTnbV5ORfP53lwVPmPOhpg2l1gkOeGgo59ONxEQrhNlsUWSSDVTrhGCzJ3aZaYpiq9agJSzAS
PpXlXiod1jC3V2nI4fBXQd/pX69Lji9ZD/06s18dhCIsISXHlgNT8XT7aiC6vvmaHzvnRn2lk7IR
Zw9F5FM8vo94+Rnc+BIY8bhF+a7S1E48aYF0jDfku00iaHy2N5dD1Jp2STb+2C1ItJwfX5IxatFj
kqGwyNRqQEuMTr1Uo0teI1FX5bmcDU1/uAOCHltiUtrZIelCPBxSYJY01xDC2sJp2EywjIS2v/rj
DzRKXX5YYHG1h8j4jjtmJHUhoZ/QSSdcq9+Q/wWuhqs9bnLdcyZT1UwNGvLINea3aI/VJm9elI2V
7CNALDBKStqDAJ2GikZ9gpvH+xoL2+zWeQdEGzQdq+SmQ57A4fUtkRm1TjYGbiR3RiHxBblBhhVY
b9XV+agZYNsDV0SK67BP+0S74eNjd24MguKB2B32UFygtZb0B9PqXwBtnXU253JSCyP0n3SBNI/P
A3tpSXgHjaaloFA4aw6hs8eU4C+wrmK6a9lHiKIClj6N8+ZhEhL9lWI9vS4yuIvuDDHA/P+RiNbh
alp9lek0aagsN9/V0cPtsYVBS4zZtZ4Gzoy+fmNJ0Onrw1a2RLwZd+Z7GdhLS40SE7A04HobKaOz
MlfPSnFV9NhNeDVnVMiNB1uj7CbvUkgR69DjQMfF0/CuJfSB7cZo9Lc9tvaHsWF+YbQV2aL1Tojd
B4hK6wK/xZM2Kma/oggVl3zyQJOJf6IlFSU0FTqPlN0pFPdgCNz3gjLV1VztBJAIP0suhSCUUd05
36uEauBEI4274Lkcc71FUBCe2eygz8e2Q42MPu8JukRwYqnYhFFzDHGKPkXo80VyX0MwfjtjQcBR
vKbEG7bx+dRcAa/CNwVnc02xtvaNcHicUmJPsqrUA/1eM/2hEelE82O57jKhUXdxGaQSC6KpTnVl
c6MVYo/ckfIY9xDTF3bGrv/93F7IH+5eB72h17kt3jvQDTZpDu0UmkOreIQ4rVcmUCthsFbHZIXW
pxA22689PDvMate7H2oWqTCfCy1FsXmrLrAeKpvOTdL2gkieBjh5bzClYdgeToF2oMLFB0X7m0I6
EtB/53RuLBe44gAaX1TXqKNNxzLdk0h9xd9Ft+uFTtyvqb5eCwuJerE2lIxKaoT0ifM1qqtKzHCy
REHwXh36SQ30mqnKLurZV3BePT9rF8JjCShYc7QqHmUpSVkWRZQxeRlbfk7dPSq84hH3/3QvtxNo
jRmTKQh0h/OPuMYW1JA+C49ky8oBVNfwFTPlmjwrs9Rahr7RiehRblTQRmUzsdb+zJDn3XITgRZQ
33CXoDhIY/yl6fVWUEIiXyJjUZ/ksctnNGwmxAK6OwHt/ECkKkNMkNCnUcEbmyrawheTd6GREfJN
88Hr7MsVSrWzm1qbWS7J4wiCXnkpMThwKqCjkd/GlN8nvl3otW3gcdv07lHVWPrrmrPDvrC/v+AE
lA9zzpEKXES011wl80v2tZgSchp/tjEHFdZCbidpHirWWhVECS30LUj98PV72e0Lte+ue3EU7upU
oPGkGF1YtY4HuusvE2GDvo5m3H6IfSmW0Mfk7VrYDSNJFFka+fPgMhJe2l5oU+YcaMYF+oKWE7QM
Wm2dWrkzb6bNjGee+twynG3I5gKo7kAB1UwJo+GhUqBXhXEDWSCeehh4F4JroPCczUreZuGBMNkk
MA4Z3p8pM62cSOssY2d4ve1W6aPu8f7e6KlqObD4qGfbAOQgYl956VDivBNO18TQJZZx55vbvkGl
G03E2l3OxdteHEedNK8MUZ9qu4lsDEFt+VMc4m4Bh9aIEIzZV1hqBvd7IGs148LoctM8FEZscz4x
eLPRiVU2NhLHhlkjkMyFIZXTOERs6maR2qak5TdgdsnJXohF3/zx2YBVnOEyZhrnGeqm3nWAbXZ6
6XAxUyIUx1cVGC8V/Ah7DzcpjBmE6B88E0BGaDpr0XQ0NU+Sz3djBhaZlkrQgQXFR+c9o9QG5UpL
egAQ2voSIaTv89zH+5vql/r2e5EUoDWHjOl7ygjbAdKjYK96P6xcdqkBIOM5GnVgGFe+j0odtYxX
qXl6FU2xzcnN64ffHD30tbqdzu1/tkJQrfPQbzOWGPGmAYy8eMc81ZWj87phW69Mpvr8tJeWEd2N
KQwU7SB9aRn51uq2vGNxSl2lbB40Xsqw11Vj+Ev6WljBqi9m+i5EnppunDL7ThOc8yrMyTHOsCKH
0NKl0zCxCRUp77QCXyTF4bjyLtsnQNFeDej9rTZZ/vJiwLJdO74aULVMy2pAhC/ymQ7O876SZpI+
+dZnf7M3Flu74/KB64nYgGSVvTOiPWmixsSmJTCJ5Sc+UkMtupJGtXgColRekfJCysvaGVHaveEK
Xs1SSnP5dGL/JSuKFrrnJzxNc2uiIKVqVBgvvgdDoryOUogEPOE3k/k2PTeZZqsbEntVT2nyu9za
HkO/1+8Ngcs5AQNkGqbMTSYUCbR2nmBwZJMiSxbVZhsPriuAb60d6UY6lhoUrKXCACWtnSsNiGCe
MNvvzp7/RewTfr0vE/EyFPo1kt0gnrnzW2d4WGQfGRxVkFzEfCXMeSLLLKAMwJ714oFYuuw0JeXr
AVv0o/LsnsrUJiPIJcF1/CO32Gz8thmfCnhLC5hPSt/YArXpQO5Og8BGAa7MggsaqcIQSd9XvOhq
B0cfhz+MmTHg3+J5k+rtf8vm7I+X7BHVZWCAyxT8FiybQysIg6QqBP/Ghn4w82htkWAkmoMLaF5e
8rvQ9PTmwW3WsFbgFnhXUZTqUcvCprGvKiAMAWxZiVe9C3YIEBymJa5odAQRkr2q1NJOIxkqBO5S
FYwVGrQ7+nxugpvOHDTvHUi4O9fIQtXTHymKUHM4q3x4DWKR3A7KqBE8KSRDJQ+MF9sEfCiaQdYK
OxlLsWHasTRAo1RJG2iOsFwY5q7Nahn1E/O9hbk92id9H2/X9u9+jDr6vtXEXr4hNy2CfjECiB3X
UwUmpCMyyLngoypZkuYXzNqvsAfq+N8JIYT6WRaOKYBMZqJ9rHG/KK8r4IqxnVKQXPb73zWGBFgQ
T8tSkXEF4DyjNGfkILeQT2HYRguJ3Bdfd3iX7AH0ulUsibXVSIl0m9eKfcdeV7G3e3KT+u8bQbXh
6UxY99HxpyZ6XuHm1WZNOstMthl2dbJnb4BhkSE5+mxCTPkXlfwcICBKZ7qPQG7/YEs4g5PYJLCq
WvXhvjij60Udrz1ILxGMnwKob1mARJYGdqKdSq8ukozqqtyIDrTWwEPeICmgsTDyVlyVV9n47zCF
mVpDGa62rE1M7pNbEH3Cy6X/nengA1d8IJUuSIKZ0FB8cx7OT4sl2VK0SIbi65PSD5N++YKWZ5eQ
RcEuBUd6wj7Hx3whCCATvjSyWCqxwiiC5fzQxSQp7tzwvPLFTWJwUxJ8/6Y8aAvxlbpditYsX6FT
pe7vsDyuY9qN3R7sIKlMpUsEWzwkUR3qknYTC7oo54VVQ3EUUd3e8oIOVN4Uo0r4z83Pc5HTr91A
Jd8E2eZtbpAU28RJdJGUkieZmOBJ070Xhgs5rmAujLzBWoKfhjIV/raiob8QlJKcNV54lU2zzgRj
DG8WLKaY3zkbQY5VKepXlDbdt86d+xAcgIjTgH7BrMZyBR1wBFI5zOFAd1zK+mpLIpYoQjwHUqq+
0sJm5CG4BcSX5hfvFNAWr//gNv1Hmcl4ig/lhZTV+RmM1cYFzDcoruM8BC9DLETYgdHJoiI4U2+e
B9jimmVjy3d2jlUBfslasR5YEbpdG5spB1SGbdLRw+4rtTM0luQAjJNXcU8Fg+d+DmbSy8RJxVPw
0gNSGNh2sCCm0b3Yg+Y5UT+qnOATyqRtBWTVmRktPp+bHPjJZ+e5/e7aizrlp+b0cV175VuJ5ltD
Wf+bt4IX01RFC61nIDoFGkEmi5cDgoSmXDPWog9/npt6StCLIYgtNZHQnAnkI3JmhuYLJH6Wli0S
gejzHLrLvNBxcuJq0Z4c7r9PAlaGwnT3XN3w4OMukSZqEmQtnoWKp3FZ7mCwu6lnUzVlWUSlPYhy
O5EmjWx8uZFqtLGAdjOT2MakGIenpkNlu4OKwmlfKNIWc3/2exi4cf3pGQy+ZBmleYGCw6D3W8xQ
LAmrozPVfexHpiRGzVLn0DVfDxZcMTVJLbWTREEsLwxZoTDKsWPakdOoDHxrqDZebFDeS79WKPLm
mqRC6OMlFQNxfs2LGma6cBQVvPgRQp+eMdaQsDTXJmys5HMpY12/ekuxOajbeYTkURkWR7ohleYN
5fapsB+zY3lIzV/obTga7RjZU0lW904GvDXO5uxDe8lYNv/GGBwewNxJ/MM1mqahjoY6eXdYcZ/n
dRKYOKXufIwCTorLhBfYrzKUahB8o/QMNLTLZSV5BE0WsBi9P5V0sByUlH/GjcqcuW6i/FL5kF3J
xFQQ958+1zv3vnOGsS8/NPW8eCa3jhmjCBPYt5u4jNo6UP09Q4o9AD+g1/YV5pCVV8AL0bsi+R1f
1+FddHsnUZja2XhSI9qf05ll67GvH5KwIZOq2ugosI+40JY78/umR3czIOBUzka//gKn2zOGANAF
hPH5UoOyBHW0u6uKvxSFCidIp/42VpYrXfYElKoSHPqlpGeR0FFqsVHmm4Z885Kkw6DQi7calyMj
jdTypk4iXEWNVKl7/TNuLTBbxd+AWZR7ORoDD/IFGdE5VY1NCCFE8b+qHbc0sWxLnWAuYaMu7At6
k9GpDCqZt4npTSosibdT6OvG+P4YR6XOMirHXv5Tqgb09mJ9bLR52P4iL/hMWP7J0XnJ2QthjGHW
nID6EBOTIH+2BRkJlZDuMzIPN68Aoo6x7Fmt3f6KTYC3Ut6Yuzf1pAxK+v9klXL3rzK59kSgbhQw
GAU0EBnUv4gu2Sz1LD5rdGoFMXkLULb7YCLpQgPHoVMATxHBxpNYNhTcmyd9zRQ5q0Pi1cUnwrhE
CqgTZQyOxJnD5t7bJcEcV82U1p00IZkWGPR0Ln1OIlEJciBNU+oQWNuG+pT0dz3PBUJ4gtDAIzBo
xI9R0hl8FSbF7nzHCpS5+w3DvcFeELRMMtCnszBH0fF0CAFDPOCU4JfOBswUnM75k1rbkflJBB10
2yRHI5DNAXp1W1a+QXGQ1WSzURn/MNeYhHotqA3GeFrQLfyiD2lUcfj5ItQaId50Sx8Iv8n4sr/R
t4o9JDys6yX+gyoljd0IinxvudWY3optpvkq3/wqYXg5MxN1mOZyi1NfxTgYNBOq7FUj9LL+2lsg
9znRyG3v7tPjPFseZD7Zjd0wuKcEppzp9QghKgx7gTfoYtyjLddPopOTc3XKk1+szROsxgPgzSRt
XvO20B/NyuRGz7p6MnPeCbxNdJhkd6I90owkpBMuxVyM/4pSqB5mKxXr4ViVXJMe3zjggsWo+UGz
66PqOVPOhofb6ohc0303UFYIRfSqSK4+qQnKrYSBk5DDpwScd0P0j88tvQ4f7xr5wxQT7QIgXBkb
WrJt+41/XNxRMOx/HOaxoc5u3pZ/qoSV6t0RKr4d/KA3NsUMTfO8KNtqh0GmOMalGw6jsefsGMPx
q3Heuyb9i6e0AP1f42+F+o9nEUHPpuGjyt+CSsaJSb0ESZdT4bR8EyetROJuNF52w9Kf6Wbv74af
RbwgS3gI9/lo28kV3P/fF0E8Yb38jqeB+G1YA/OI8nBoxB68FCpaKWNgj21jn9MpDe9wa4YYodUB
T9xm7hNv6aFQurzkUoUMzVRjHZVmpCaEPLOf52d7sj6wFpV6hTB/qhits7tNc7N3Rx6a6zy7q9oH
fxtAE9kWSLieN5Yr/3Gb+T15VAw7Yxg9b8CGzyfWd17toGb8zUOXaCitWTsXI6G83+5KtvvCnTAP
diZe7CJ+Bzg/uJEeBJgHZ0xKlZ9N1yHYYYa+2ffbWb6Wh8kj9xridiLIrYpwYTcvm5PSnUAWHI13
hQvkxkx3gnukIQTTb6Pkf6kaUpdxc+D1C1SbUZtUsrucTi++JiQSTnVUME35nDDcHROGhJEpd7Vf
Sf4SaKNtBo16DaAv/TiCPcaHC/s+26KmBp3Mx3Ci+UUDc3H58L2QKJG+uUDhVGAiQCfJT2enWenO
+6WQAhqrLAzq5bPjYxcA7LGGX7O92V8TA3y3/sk9146muve5nAQGe9kFZLzqz/64KYQZV/Sn50b8
CkHHhaITukJZtkKFFpYbX28AWxHAGe/BpUprvAICgbSJTAFr08OATmbRrw5b1R2+d3smgZ+WvfTo
lQX3wvog97ZcBz2yltiEwVBBSJf/wXvyjvno9zBLWQAjoa0V0LUlEAILfsi+XQn5w/SWEFjgDqW4
si64Lhjsk2LmTQTFGbSWqpMTeTrAz0k/y6fSJOsaNjPW09WRS8DRTYTYBn7xWPCD+9mh11dL7fg0
9dVMggrLvKdsXRrjl4SiD8jhQMfMuhj54g+yP40wWS5RUhyaezePmF+JWVhNzXSvsYozYibAOm+H
RpRvMUiJYYGpKrO3R6CtriTnJPftmEbc9jbbqMmMNH7UBmms9i1IJU+lzeAahBOYdD/zeBlUE/fd
DEvngIq2oM3UjsW+76SeNoPLkr5hN8R5nHjUV+G3aVgy22qgwxWhihBv/8ay7FuBXO+T+vCNvgzo
Cj3MwiziOZxZH6d80ODcUERkv/NHTwL3Ti5vMggPqapUIHB1cIaAd2GyCncWSOn40OwGm84JE77D
EG0N+gmKCQBNUseAtl0lfF0JEPsg7DiuBg/70zuzg3B4HD3ypl4ByWJJ92O/rfYuiP6dm4F0V2i+
U7VcX7F6NPeNbpqW2WfvAgIPM+ax8s1/SPfN0Qcj8TLsqaHSnnlUcAQQvrj2hm5cNhRudpPE3Ygj
H4bmqqe/YVX3C21ZWmD4NhPp05PZEtfBqzP0MEpjM49432LdFLhhyOcL0UZ32kfoHkszK1mGRylu
vS6Si/4JwcNVkdpYx3lNE6Z/8USl2bpUkrHI/Vuju5S5Cc+GOSuGs/z62ms1tRryKxR3kJsy3c1m
WSGEc6vpBRTKPxPjxYb9ebUeehrA4RRehCy41BD+Y1i6xfgnAnhyv01kYugxsgI0BIUWYWgDCQ1L
kGJ0GfI44A2l8JvapUgWy2iD8XgRMIqnSL77F6QAGclROQhSzofmmhC7Cz9g5QDh/Sef/fxiOUXo
tBmerEf17iTyOe1ZxVqmrZW8M3OrPq5dU0A/iS6QUGig0EPvIlGq5fBq654vo8sUSMkw7prdEvkF
uNGLHACKFeQ/V0ObazdrImouHZXTdGfFWUK0/sWC2eHFV1C7vEunHkeUV3loAs6Dx+hUR+gJQMvg
qaGV7jdmpInTyNig7Cb1HjEl/mw+/uZ4JYob3VN9NbiUpuIGLJ5d+2UBBLS874yhOuFuzMzyVC0e
Q4iGwQrWmBfU6ICAc2lFPAZOC+awVV8jA9wkAKHt7kdfu36K84xFDQ+xSboFu/7x1DUJerKNVJ5p
+fDWqXuUTiJvGBHai7KbPKU+QZHP9V4OheJ3/RbffMRjEiD8gzMMujA3+nkM2lTVT2lWuuw41Qdc
FQMgnzPOJY8HfSmkBPjcirgT3ew8ECR81Q7QiaUNjJoBQaPgdAMKBctvu49CqL84OqzYH5OgjHRe
bGbD5KOFrrL9UYUeDb6x0PUKmfNcLoTdBgRD3L6RmMaD00sY0swz3007cuMkxyZETYsjY7qYwH3s
PUtf9+Mhbs93QdRXTRkYLo19wNBPq1Vr2vwBf3a2fuVb9ygDKUnQ7gixnazj9xdSzy/u/s5RPC8m
gKc9Pm7bKMAcaLNOLdphKTfU78BqICF9TL3jjqjA3MnQYtV28V9gDN7AqI7HbTrqDRQXZVEDxy5U
ggE86DTXM4y1EyO2KIeDQKzFBKPc65AH9n9bam3Ipp9CfPnxgXu/M23vvViyTEjkhJEZzgWfSsBN
Rij9JiQgHJXScyb4krfX4SYLGQ9HMtdIFznQOoWP9mUIHLaBz9ALXedg+XwecFd4QF122HwyUl+v
Z19RhxUtqDIg4S1Mk+mBJZIy9m9iy/UXFs0Ws9KVEXBBjRr0cPVWrs7vOD5pXnI4WArsLp6ykHir
RNvThq9WFtjpZGrz0NcVgQjb09HM+me/7dKA2TcnMg/gJkiL4sad518CMc0AsKcFFYD9HMDki2LD
hS1a5MTVELuOnuQdUc/mmBAVVCxaWE83dtWtBXnB8KxvNM0TnTQsH03fbgwGtzvbaRhWwO/hBoSp
9ae6qvi9xnlsmhwyNB8MbPQbKDyqD4BU6oV/kC9U6P4ebsJam3ETMtl3tbpN681Or5rAEWQMXLwp
BE8Mgs6OB96lJXSj/Ly9a5wbHFcPP+bRZI82oSHJBpYEPybFF5sB3k7VGLJ+aM1RuEc3vaDIHyrw
wSutpkMKN55gPylWH0IgRsxbfSc3qn4+RV2Lff7WQt1DPZdo7cyRJjYghTWDpaLDK7b+GnBatYb4
+Eb+mL32pCvBCE4KcG6rDHtbwUIYgZXikZ9sJ+OoDE8qWm21T0JI2RLMhluf2Qfpmi+Kl8WKdS1d
VuYTBNzz/A7NwO9DubYGVYGOaSN8GvFQCCeYYYlIkXJGp8QgyniR5ZmJ1b3TCgmjOklyNr0WMTZ2
/eao8w+xd1kMaHLs1nkVFJkuGVymx3TXdqWStwselh1XBBBD2HCOJ6CiHKewE3dhLWkC9q2Awcva
0TeFG3aWx3QVt/HOSRpqSNWH00acX++6ynDd/mPIAYfV9/ddJs2Ib8weURx9kgTHp79U7mGhFIAR
l2r9OCj0+bj9hUdKh/8p2/g3it404k8h9AJNyNxka21T8uDCy/iPtYeXTnOm2L2eOUAlyqLW7pTj
Dhm9PBqu5YuYTarTY8HL8d1uhAoWQDvALOE50GH7E3BesOxw9qWxYL6J7G+dxK/uDH9T1DhMrmTj
Hs0dRxbQqu7Nn0HWsCjwXDrXSnzfKRATGvFfdpLlOyA3mjyEyMP+jOBuyX7ciTRe9fJjZHQNFJjV
Jana1CHHKZ6GsV9SGNoW3jBhanYg8iba7Ai14+qvUXdP0dKRghh+nSYZibkkiFGAq0lxGBCZVX5s
hgXqH3+yhKokuZRted45NyPXN87OW/0dm+UmNo7WyUNOg/QuvcvGR8tfr275zSxM9v1HL2WWANZI
lZ6rAun5msJB0o7c4TJ1vp3XH9Em0+qUbwWUs3hIlpnIKnU3J79O3pW4q2NtIguwK1htRN31l6fA
8zY3GYgZuokWHdWZzaK4qPDq9BZwW81nfpm49Pkf8zA8/D7YtI8B7PeWaIlH3OUGeJ3+t7zFPHNl
a7eKOw2FFXg+e9SdtHlt1QwQI7ko3uh87x8LIgsVbbyJLEJuycxOs65X1Y4Xx9dVVr560ivlWuK5
zTa2QqDxSCw08v+1Wh/e1I6GV7JKnIz/TMXvTjl9M7XLzfmTAfJBJ3flBGRmrVDzGVC3j/JV7sMJ
InOpHTLIFa06RwkQoH+Qeu0OT++6xnDKkOULd+qtQqkMfyu3cJ2wqp2Y5MdMD8nPa4bTezl0krzP
qV56dAcEdXjlxeH/YTru6Nwp2/LVMiJM7GUlNSF1fPZY5MGpeBLcKMErL6e+WPGzBngU/tGb2XXf
c0GWwlSE3JOyAzeHis/yUojmjCfQBj69Q9U6nTBl6s1XN+KUumV4DvxG2xomgd9YWUmMB2quu7tX
fNOaky0T2iN3Nvyc3KwVJ9trXd/LKpUHfEXGJjM0o5AC2aImxj2+shx3ldaSpCQxkUSdq9ZRBQd5
7no+IK03wbltAgRKMxm7ojiefO6hNkX4CZBzvQZ5nnJ3fpKMuMcsGpTTB1+ykG66nlvVujiJ2mA3
ALZmOyrK+NMgIvhwXWwcv36PbHgBHSA1y95cAoZpqDFf1yeKzMx9bwCKoitB5t/0OMXQ9NA1ARa8
Zu/OCX/7B4fWk3A4S5fHUs4/YFLYebXzt+1q/iEQfYm+CubqESOaOmIMVKtZlaTgtgdUuohwyW/+
FnctmAJALK9fABtyyN+5HBsI4buB1yArZEQ9QTOZNEUry77s5USHaw6vcUMlwUZRJXd8inEURRM1
v8ddvkUdzIpWwWXUOkB2yv6JOZTjY5YGpywY3guexr4Fi3R+lLOrr1Y5j8e/MizSJ47AMWvwUtzm
tLHFrvR9gFx2V8wCsZpvFG9oR4Fv8hKT4QVO7iAe0aeOIvnlmsajhgA5QRTDZZfDHt1MBDHjxUGC
cOR8A4pusFOwXX2aRK6ZwphNR1173HgR/3OeQMHdNbdPTKlv7P0BIFXS3HePlhOCmp/9H2LAc9Fv
ewp/fG1/nflijUPT++4ko5R/b3wAzgb+sT3lrWUM8vcHezRbykNh//MYTyG/y6qmwVNUg6Jy5P3K
dlSDMhSar3RNO2AEOFz445Slq5DnNz+PmqiX0Ixwf1hvlk6jAbiXiMgBhFcLcxh13KBBlLNDkVZ/
fJXaXWkto8Qu4lF+IUMprFDdaDZEHhqMF1+7xzXnV8u/1MpIAn9RblWx8D/UulNxnCFmiPieMDul
S5+6f8Mvbcq6/tJBM/xswFMiCyIPZfe2nDIWqBbvTNiYtyq/swZrkKCgRJj+nO1576uvqc9opm90
0YvkJNYR23Iry8UQlhGr4cFV15f+AjjZxns1FFa1oUpbI+p9HeOMAHiipiXFLBVyaClho0qW1YRR
3CypSJr6fQSNpf1L0tan70a3VPVuLxi86RF9SvwQspV05hBvuxNLb5h8a179vG/dud+otQixUd07
8eE2m+7CpfbW/dBR+sRNLe5SBcPjL3CIPi/QeKuVMATdN/FcekiEG9mxeZiEBC+JpOczeicexfBR
kw3o0KVVVG7byi3Tb673TLUxz4hqfX0g0WkNmIXu4yHhEIxxozjKKPxQ6hlGmLrZnKGnk6HyTIYz
4JM9VdS/MYWmxGQTHekhxGNkmvwxwRlQriQLojy0DxF+E/vyyJdAK2Ud0RGFI94ehBvO4hio6yEO
e+jCzgGTWjG19jecxOSAtug+j6QRN4WgA+nC8yomi2OQv8+qqfC99DQih/Li/rt5lczSJhYfaOyZ
H56tTbFpowwh+mu3E5OY65Cc95EqtHInCR8WuJXD6uR66VCSUw5yi8OpCs6jPAzR1Az8uWMVNav2
7I+Tm1SOmS1lG0LDmf98TmlxvY5L9vjZ6l0/ISMSBmFw6sTN14L1u5WuZKR22b8yEOeYchUtpkR3
w/Bp2b2Woodfgix84FQEUaEX+BA7CZZ+8pUR7z6rb0yzUImvPdpRumPicD4qsKz4OhGNra43i8Jl
UtAVTkWPu3BOu1xw8WxfsEyOF0ruyS/8eWc+VhP+aTKOcuyv/ccudiMAWXLSZEo9NYPsubCYtV8f
pTLOLf95b2+4MGjzKZu+6tS0kOxQuOueyCkijuFi15GITrjLApIJMpc/d3N1hXAzzmLAQWm9IVw+
GHfkvWE67U3iTumm4p+KntUNMxB3E3Q/NFazpezq5eNuMS/kEjfYmiWvCyFGA1EiXL7qPIPV6IAt
XTmgzJOAHdWDlbVldnHKcVUJh8VhpVkhckvtv88njvxNqhI3rZ55mQzfPTvYQXPcdo2FgpTOYFj9
VF8L99OZaKwJBZ/ubLZCQN4RTfB3gr90jvuibyz1n6BNt9wXUK6cAiYBHr5B5dK99sH5dp045DjI
joVCNPTysG3yic72v/Q7nByn3XIITH6kCmXLCUwS0VtBYPB9uq2vI6scrM9A+dELZdYqW/KFaCyz
6/29pfVOVAci8H1PEyvoBVDuuqCDjbBOSo48H1Q0Ir1m+gj56+zl3MWfExD1tl+iDz0FjmuZhqVO
aVxnbQ2jfIoXxmhy0MBTL5IkEXPJilVj9gzOhfxJaWTpGPRAgpLlhwhWu+4fmSpCcmRqzmjHTsap
LE8zyDEZbH3HSXlS7Fv57nvZYVzh93q5bV96RzV5S7ldBrJSPNW29V3epfdR+LrQDecMBMgwZkXi
w83jNwY5PE6RFIgtg+E/mzvHLJtI5h+ZKlllsTz7cygDhN2O2Fy0q+kDOhM14osn0gIPHdGFc8L2
wuzP4oBcWEP6b0CQ6qD3u0sngZoCBu75GKvDyk+FmtDT5QnjvCPDZHutWIlIprDHDb7IGduLCUw1
wkn2kw80iRDAIkGszQWDZ0IDOv4hOSNQcaCHih5UJUcudEFYQBeSyEXpS+0a22U05l5Xe8fkFPnf
amRRJAIv8LEEJSYCSpXeezIHbV06uVdZQBwIShs/PB5QjawqIz9rDWMdNjeMFOREPhe27pRBcsFe
jVjjRMkcMpgkEoToiNJwM4CYyKVBNFBn8toFpE1L3fJP79p8w1j78lkWON11PdmMhF2fM9KPRkQW
OCMHy2uU5Vg+n++zY1N4z8g9NNntAV+JoC3jyfyNR9cl8cUtEjs1YJLDMf5INpJcECuORa6/mEEh
c8mQZHuW+Q15ESiJvvPdHMk5BQPI8RZlAat6AjD4noa8gLLVawvB+Wvp0K2fYersHAn58F2+RMmT
hknx6/1PLb6j72xgRvVZWS4B9nvsh9AY+vleDTrcaykZ0k/s63+Cp/bkz3F2qW08fVzE+r9Sxe3p
THh2S+0c2m0q2J6E0zo1rKg3XGiQ+SEYajOxmrXCspR4LmgTt64SKCJ7fCiR25hKncUPZ488qWB/
ZA5TUhBcO2speavHCUKNciBtHuOSzDGuivOn2QNw2lqxME90B0oKZeTdE+FNiHhRK+GBw50F1YtX
SsPQPGzUXaQHFOXY11fUo+p58oZFZG4FEK+BvkPeG8xovKRxXdC8+n0ehQalP9wsjQagB4kR4z3q
Mv4NPDDsvn1f56/oTBzmTHvubgSRft1We55axekOu9SEElxo/emUphpQWd9loqqjkh5wHT11yoKS
KvucY84p1ZZfIcqFvzpCNAwIR2aObHjDV1Y31sueoyC3582Jpdkj7gknCZorHdyByAhPqqrZINbm
M8UjkcOav3VkdIb2zxH7z8JP90PqAZzlr6MczRjYp+9eE/2vEHgjl/u2GlQcRHSoi/zhQpLgu2FT
gGRM4dGzvU/+FMfBUCJZX6iR9gg2olURUssCjyCFPfyHS8JNiDrpUks6aeUZVEq05u/7rSQKJWkL
mViDgobgrZo1eoERwB/R0WPDMNfntuagjPevCfJt1OqTE2fbUSdNx2PDtkNziYeEAGRFfmOQw9Sm
ynjSBu1tMkwEJw7ZBm0jYy1LTxjFiOvnTGoHgehYM5zRuC8CZw6bmMthIIQsFPgrlJgO1DTgucg/
TM9wdx1ml5UcbkbciBeFCnuASZ/Cm0wpWNCEEDP5EFJQiPc7DJcx90vXRi8GRxKn+n7WV9DhrRG4
gZTPuZAs98BNoSlJ7yERw+2XZQ/rOC7pXIiGTS1cyWr07focPdFVq2GGcoBfeNO638ZTDsxi5ZMz
S+FvOMSnurXf3m7i0qIhH1Xcz9SHBIIF4IXhpGi7N2c9U9wdeAH6VK3yGAmCOn1aIod7oJgo9GtI
Phn92tBDUdM8yDxW4vojUTQC0/mtN8Z6obU+aU/VgWWKyDm5YblBRD2D9J+33EkoMirksM/Sn/xb
d7m2ju/+/tqFrBSEBv6HPQvoVX601ytef0UfX+127FkBYwou4rFWBU7F3snY1aponSpVG7qnSxPe
yld/tAd6saW6b7nS4Cr1VntzE5nue65ldMEnza7GJURXDmOaQOd4ymC+CW0h/JLaxTyVHDYdBrBp
++QQGiWPgoCeO8TCrw40lXqMCF2c81g41U2m+2IVuYz9SNlwoZnaU/yqNpiSDv/OzRo0ZSPryUS9
674AzPJETExaE4cnDrQg1OaHYCOZ/20A+meHRfRludeh5+sBX4abMKi3dWqlWfNDQ5/ybTNn9tei
FDC96/VzSuoNke39bjd+HGPUerO3SB16WHFmnft7no6UxrPn9QyerNQ672quBvY6tR7BGky0bq6T
ahYrAOmZJlCvT7NvQhxVDCsevgMl38onrht81h/NM5mkSVNWpe86c71GpJJ+pDVu/5KEa/zSDKg5
yiZW6V9o3IWKAHxIrg6pRlyekzYAci+NBrO9ZuaAyLQVneCuKn4WbSbkBcaSjujbxEYCMOZNfqug
AX/zlDZJ8m2fc0v1L0G00gM4H8cs39Bqbden6TuZbstek15cxnwGHwcGMMt5bp7SQllwAGF7GYA1
hK+nfeDXYykxuegGfABm7c420lfWvkx42+CoUwfbaO/LOmho74cJk6DrYRcAx7sLW1eeKC909Y18
PAEx+CR2IDxHTenY4a3L/d4cTRXIcKv9ecaUAWBp6aWyJwY2c/cpNZK/vL+CySYkaj+4XZcXgw6K
KqBda+7Z+kF0rzVLVeAZz3/UURC4losNtutndYr+olZMjyZdrlxEZ5R5oglvRsdtoQdSHmNk+sYA
Nnki/Nz5Dxiyqfb7fj5+LptvLhlplL1hZ6TNV9tOz2OfzKBN5oFOTIXvOYbkxCj2iQGtvAx2cM4J
v6QlMGLWeQ+Ep0d4Pxj1Q/LoCmus1+z5JDdVfARfrnRJuWSnPnhFzd0l0TTuvF6Bv/rFC0gtjmqJ
p+5y/0oTMJFoDIJE2vdkHv+tlmbfFYEMGPtKXfHxWvvDsMpMWsvDvcY0Ea7IYpr/wC4alNnf1Fx4
INwNu70k1wm9tQK+fS/g+Zwqu2HNlpQhxdC78HIqi9WPvRBY3V1NVDfMxwQxkUQUQ7H023+2vAuu
5LvI8BRAWI+cNdDMLlVvhYSNtESGKZQDFFiQ8lxRHQzgoRjGeLp9Xr2U8vhnZ5cQi9/+Ia4Gzj1f
0XrKMxH+up5TQ9sgkmFMjdsi30e0k/NjiyWSzpMWjlNYROpooi49WAw+41/GoOiA02p1HjNlxRAB
8FPs6yfEyOn0s5DLA6scw/+ssgDpPYfTzLAY4zZV2YQN+HOy6CYBfH7NSjolmbzyKVKzc5utzR1W
0Qe/zvP8/yqlKrMFlqG6dTT6zCW0sz4/o/XSCSBH/MxoLNmefxSt7jGJk5G4fYwSzesYvC1adv5O
T2ijvKwKRNKfYAQcWX4ioqc2zx+f1m33OF8IqASh08RjUP/cHFAb7hcQJ/diOrnOAUbviVkHFglO
O102WvVVmU4P9RL0NE8GrnhklZmQW4s5plQHNPCfwikTz3HF8XSnv/Qmp+ltcxkt98hLJh76y8Yl
GwnDTJ8QdWnh8rQcLTGwTiK6iDMIjyk4GNtQeHFp7t0xaHXpALEYcFqGCGTkweHY54BV1csIn7FB
2Kj2c6cwtGFf06kFoNNZcdPcZGpBZvHiIbWjFrA9HtK4cQg7CHDeRaVXuef2ctAWRZjlITpGZjA+
fkpbZu6vZhTyL67G5QEv1E4l2B353rVBVP0+U2ptliXeoVCCFF+Zf7HOAxYFEVyphl4acDUnr96p
WCUDzmWEWsnmw6EPE30ieXYLB1OM1bSaaRFe1bDrJ84Co/WVEsMjN8Uliy7CReBFETII8eZRvn1O
sPpl/F6tUxKMARo+ihzMKXoGCdvjxApXyw7pWxkjpFCDhEdLD8VYTSq+FF6T1l3kTc7nLwyuYrjD
bh31jWaJtR1p6vL1g3XYVUdzhNI+a0BhO52B3kr7W/clgdV/9D8tdrtN1G7BiZ+19vf+Z29f6riY
bPluMITStyakmhPK9gbXGgqle625Tnpp9POIDP6LweMHY2VXF/lUHQmRiV32e8Je7aS9IXTBsf3L
P3tvn9zR6kOHYjxwjrV6e2wS5ehLV6zTM3oNi75KzCVWiJA3Zs3whz2CmbQ/3po3zeMF3/NdgsG/
Ucb76cpKhuHEndBtobU+UwJz7KziKf421WminP5g/PvRoN1QcICfHZ1u6M6tJ8YoA2H+jyASutVJ
lq9pEuQNloCDz59OSuDvsXnTiWLwX8t6NEQyJ/n+R1ClNOmMD00AYMcQLOOiMji1DI69N8zfl+ul
v5edRRFELPW2/9IWOjkp8n9B3bWG9hRPyjZG/LjxduZjhmC9wIZjWKD/zBNsUc0jj6zpaXTxnSua
KIpnOawjOxzuj5BfCNYiZC033kOeAIMSJUP4maU2S/0s20kEs2htPekF66X8F00MvB9kNeg8gaZe
/Ilay9dcdc3VlQk0B/V20Ldn/s4DmXjYEPdLvHRpE/DJ/tN+AtSNQPe8E/CS2Xw756PLU2XNMcNe
lIQEfXA8sAOrIAF+Qgt9+M0F719Zy+mZIJC8tdoWlg0Wq7jh33wcGaMupGZAEteg51kbQn6PQRLW
k067x4D/NFzKc3qv26fN7E6S815WmRDmVE4Iz3fT34VtUXPFl8nLWdDqhrTgiShjzS6LH3XjpUJW
1DdPCLdCX49XrT7d37Cid2hWbx1zVG+ra5i6gL/wsJ/gDs9qMxfLzgo8rAoJBZPquPUJN23rMBM9
Ii5MUXV+cVXUN0zgJueDnvZaR1h9kdmG6yrFYwmmrLQ3fvHU476r7yf2r5YaIVoa1f8JhQld0Grt
5RCbqoAvr1g/MRygpQIjMHu9GTd5ElKgksua+dESG0M/xR0q0XbeXT4QIk9rQbf6eSTnIJBrDIBJ
HXJevbrkvGy3fKKZfaGj0BFZ+43TjIxYCyM/ISfzOvUT/gFMvIc0oc5mJQYU3AJejdBwXNIRW19J
ikP6Xj9XP1Sz0mmD3oF8t8ZtyYI6Z9WrlEOSMoaxsoSz597xKy2iiz1McofkGJjJ1FRR2BXdzjgI
Jewt1xEOt7zi0duC4Z88A07k76yeTxrBY9PjPle/Q/CVqgsMgv7NwOzLIo9VYQ+tL4lqA7oRLtX0
nmrabOBNoQuLk4t3ZNUeuR6aQ14X2Jr5WoO5fR59Yfh9f/Tbh5f6dKgMlz6dJqz5VY5crLHDu1gq
QS7uajaghvRYSzrYM3Iu+39moNJekFdO2BbsuY9wJKM4bh+w/bOZNMIxbN4nqj7mB7HGJKtMYQBE
70+jXudKCCUNU/4u0Cog2IIryqiMwdbrhqp/6Gxlatt7i4GMvoV2bq1KopuHdXTQj5MTuA4Edq9N
ERI7xpNKHVjAY5MzPx66rGd5JAPLTAQSogWCD9wG5PWp2Q4b8Oq+OZ63RL4kW4g6gw1odUGMH8+n
sEMuH7idtjB2ROtVrrQb8h2/uEWadq2LBkB0JxC2IG72jXIbG0Zm1oWagfds3aq92SR/yC8h0smY
sD9ymMKFQPDE/o8GXQvNWFrJWMeLzpN0w4CkDPgerYuO7ImX1hP5zvSM4QRE2NoG3e8PHCVRyQj9
E3wO9luKMMsnGtyorM6u4GaF85TdnJ+K0X6asB4KA+NyHE2mQT+I6N63FWsbjf9+yFPWZ1z+eb3F
I8D0I4MP/W8glmSZbcZJIDju7FnXwxPshyDzNzm/KbePSjf/CS+5gTpVQ4Y7yS2PUKODuO9GA0Gz
2UrIdPTKxmvUjsav7w2I3J135jkO67tR6zLl6Wgym++6dBM5GILyVnb56uZOat45ikdAodTb/mrY
+NGjUbAbM5x+zoB+da0DylHAlqz6WoQR9R1wxj5KcKxh1qmOkJXq7NifqzKECQstiEr9GdT9nBmF
Mpv9F32yt2D8XKZiAEPlaTLCJ7W3pViDsQa+9QRFmIaJ55epoc3Hb7r8i0ZTtfQJG3OGNavTJKM3
587PlQHaLaVAAPYmGGThL21muuUsWTkhZhVtGxLreuCqqryTNa4Tj893WEgpa4BHt9LwFrXiMQnA
3oTeyjM2NWQm09U4o4axg5R63TSR7KRySLjLxR/k/bbsQrRIUUsWaX6E0c1zsdCPlYNo1BXMDyVn
gf2oMYXelcKz8F4UfFqV+6Q6IDZXii2kx/jt0iOf+bKdrwBf5NVwXbzyIGRigUxtK891QNLYHXLy
imIOQJbhKZxu5SN62fQmbzQKDzCtJaLQuDzBjKxOW46JbNWYOX4prJs//uQIvsDTKA9KLE5gOHOp
h1mrpGeSN2E2XfiwTJmy1tLPl2RCZlPXW0qtKtPyy5bmJjhUUF2LLXnQ15ADR2YGkPqu4Gm0QaRA
YA4ONqp4Lg1BdacId6uzpeJHJxnbhTxkKJ6UVzu7EFv9iK/6S8VlIXEwnZIgzjIgw9eZWhAqZkbE
6EAaK7z/Nvga9DKAMmLUYjB2P7V+6HcCUrYnPO0GnW6u1KdxmMi9JZcaJLpy2mCaX0zJIIwNbyto
+hvDLC4gVggxFjaFfo/oi4EzuylsHvwGXyj9Fft91YPzRRy4SjvvuexKvUm5aYLr9D8NMUB7P+BO
Uj9UKfu6zGU+35iXdWqxOcGUNsO1cDRQOhEN12r+blluuFPXNQXpwQeS3f0vSsmQR0MMUVz/Ji3I
NVxLH0T8kBvSByoCdaAxVd9ecOb8GcAEK9V2oEQn4mPput/h9bH2z51FvTo6+boLU/DCkvnJ6og/
pdij9p7gquOnuf6rb70IQ9+odKt2FHaEdsgeMeURaCYZBluJ+TD8M8J31sPYfvcnURcPcvSqIMI+
N+rz18+RDubbg9P5V3hZiV6oARLU1cJVdZrhgyEXUJ2ViXmlrrZE62j4g5mz/oRxXObgQ4t/4J6Z
ahUFJ0qmkJyRn+iLqmd+9fjEiE1Ql23rgHtQODOX6BF4m7uhqegEoYrxWnmhmhrmLg6ADiHHlkzW
JfQq2wc1MZ5VrikFzocnR1NKH+AAJ+JATQP75lxslgcGtRfe6SyuWvviva7izHnAyVNjUTX9M517
n7ZWUbor3gsZwDhHV0zUMXlKDVSre4rtZcJCMTwOW6RoQaa34Thh4QwWYfDQy8SRdyyDKhjc6/zF
Z2aIbapWXk5EUZfe0YPsiD/N8mL+74s5LqO2k1VRaKUFN5sE/jl2485y3T+3PpAvTIOg42XsnY4Z
E9ijTxQzB06V1An5kd9KlQZfTFioHhQrg067B3IXTv9OLHJYW0j/YGWmL2loyuIWKOaWGbCvPSfw
fnrmNuexHGxf6zgFnPBO9bCj+gxhK5QlzQVmz/gJaTH5yDtBQZBkHHgeEZtgDEiNZhLdieZBX5v1
FGlmkBC72Ji/Q674VABhvlGBwR/z8ydyZKgsH0exLIxHI9UM9P5NdkSVOls5Z+SG9GZGJE4sMcPK
+Jcv6sD/NdaWevXewXAStt+IQq5lBC4Bkb8xpankcDKf6rvmNgizyQWZ34uoAf6OoSOSsp6Qttyg
dUpS38182dHTEsyk3PxkHkb4axsI6I5VtfSkBRJpWq6JXez10A+HZIrmOvSBzqanSeEt9hX7Lqlx
wqX3kjbRIPXKCyGMpt6qlI/Ku6zncQRyqlEWuII1Bi01oGc6nWNPLbxQUmcUO+OcMdHLZVVOx4EC
AXVpqaJtkwpMZwRrnM8qDZH7PIE6uBaRuokbn/GN0LAPXW9O/LPfibXbyDpjJFAAuygqa8Ui9P1J
OKM0resplr7k2zIQsUHpp1GbtR7V4hdQdu1saGP66tQDeWWc0CpZHMAJd5nMsFs23jsMr3qpHHcC
rpV+IqcNljrVoQAvegIXUiWIaIwiB4/Fkhdn6QuOz1MGwKpH8WreG5Pupcxc03DrGgvOH8t1dNZR
N9ilCSk2AFdGPLaKh/yvrQro+OqV2LexMQ9z6SihD+IWBIRBj/po+w+aE48TWlH0+tC2xKrHCwA/
T4oMNTs+zjjJZtItmK+nWUHA0luWmHnb3YTtG/qtMah+RQKnRRLAa0jKlAaYOCnuuTwmQ5Ai/u1L
toZNKk/9F5A7OIDYvavUrvROMbHTxtulb+Jp+3Wh4CXPWXL82i/qKYOfuEtpW61xn2buNIFsryVu
u+wbgMS4/AnfVLsljbJDbBv92+iSmUwyizVdyg6ReRkjJl1IiwXGDx1jlfjdkrhvaJK29hAzuvg5
52yctRab8UEkqfQKzi1fPS/91Y1lJT7UXqWuUTbT96591XZfWIBiuHmErK7+EQ/ycQgC3g+UzbzK
nFd5XsM+eplzOhKev0Nuaa/mkSTBBX5n254EhfufmVq4yK/c25DvaRSpwBkml+Jf6vcIb7os8q2U
uKLPlUrcoAHI85dsTcatnENz6RRQXM8PAbZqrCoIMwnXLu0x7JsXiwC7Neeq32MWeKeid0aAJulU
NLx5r1UpYkxDXez4NtzqrxykRU28SHtWRWzijbOECTSWtx5jixp8ZVUK7TCV0Ea4UJQKmQQW3oGj
GjRU5dpICoW2Ax68iIwA+nIx3fNCQvoR7s/8ysldrmLOW+7zAV/x8E2lzwbT1175U5kX44WW1GjA
5t5Yge4rmrsDRqu/FvGkzNbdTxa6QSwfl4tm6xAmoGQ3WFIO8fw1C8yVqEaE5VL8X0zgXSg1XY54
2rcfd0KpnJR/7tzZAyYyHfVus2PYvkYxl6JIdHamSQC2Ez03VIf0F3wXrc0f20iVZ5FCC2zSIqsW
jNby2yacTL21P1ouTm+SAyFV0Asf3sIIG03M3R/l+Tm1gakCV5OWrXZ0j02HlcVOmCkJpkKnDOqC
H2ebvOVIV4SeWnXnRHGrzcImcQ5jGwih5pYKF7QhFdACfMYNihDEPItt8Sj8Dv3KWMyxSA1p/wKF
5tesLvv9QtBBaqugUI2NJHpgSLLnCXOF6+xl57fxZFHye+DJKhc5W+PH2F8gtLBf/6EWqAYzqIfz
uwv/qxw5X3IpWKnlpMy6tRdq5lsEBFCFYwtn1DloOY7XEdGhSpKnsfn63OEXQ952XLDfoD/Lrt0e
wt8C9Gam97b2Dofe8xclhsxFwdnDlOgBwegRE/lVdx76Z/rjlolBplt1ooZzQFbM4D6NyCQ4nYkR
3DaEfPQVOMXRUGnUggYN8hIsY37lxXdzBHxWuJiQE+LS7oDzalK0pRY6M1vdIN35izbgrMOPfoYY
3EVmhwDg0KMjvEew1unzUbZ0JBOX9IOAdbr6uG422VkwOTZfUkV0qDPx9AmxmuVcM3IZiloqSCMf
vAnD0u8aYTEWVfHuWefw7dJoi6k4dZf3A1jl9DA0SUyG4W0C0vq8FgE4WJkPsvpD66yVvvAX4zEh
R/09CTRgPe9ELWh7Ya/0lyUQvbVjGQM3oTY4/5rCBJQ5E3FEl3sNRLb25fkngVtQ0SNs66nW8fER
f+HFtxp6eyk+yEjv1UdgI1cNntTm3WK4SGVNpqE8zuvmUESjgaZdw6CxRzM7EXQRK+Fe+ibJ5oPI
tMil/DYmkWFwMCEtg/YCj5b+3ezkMXwKHroFrTAkzbsKv1GbSs0C1DZszwLDC7GHo3EI+ncbsvA3
NGflNVE5rnvyvnDyULTos3sdSI/l14LoUiHa74dYKF+cxLGrr1cxFPUHbPINLP1d6sQQP5j2w05O
ybgMAMgfQQQDOQk/sjAxM8EbHNfb+lzBgol5ePN/k9ZE4AZFBhVFNMbbzygKM7wUfEcjexJTugYK
X3geDUOSFlu2+S8Dt4jxBgQ2KN9RfeUfvS7mmFYqsNamZmGXet8Loq20YHxAb3aEjfF9AfXMKeTt
tqVvxBfhFF8/wgO6nMjaMEnvR/UV7sPrCZ7VKpq9f1wiHI//zv2Y0aTp2aw+Oin2wcl3rWEQcmx9
+rUOUldTxUpMQEAARl/Af6JrvyEWPv9fjn2isDK14dySmdEIprtLP7LGzZN5AqK+i2h9+08COqbU
XHa7xQOnAgQZaBkyp+ci8fJiTy2Rt6PTG8zdtaNwOeW28e2zX0conE0FOC02lxDHLuk9MItDvTjO
SLPAegoPcsNsFY67A7rQSaEqYI2TA2Fl6WOy0lxMU89vXnrPNNcT8mfgrjKMb1TV0TSGA/jLbTvL
Tfric2WGG5NfFIYX/6TPPmYY8UA4dd2LQKZzRIzMFOyl4UyIUNrVuQGSnwR2elJ1UuC3dmYIvq+T
Med+j8eB3CgnoMqW4iw93uarp02e+TY2Id4PIHI0a1DlLwc6Q7RqwZLyeFvAZQuvDt+zcp40Hd5O
M3zEe+A2NH7rVoaFCxwQGGXE9kp8LIh0FtKHqCmNRFIgHXZatg3BNplESyLfPbt6Awbuq66eQJUS
ocrhLeV9H1ThIgUAPqZf3iCo5kaPrPCUXVbIwFXXDPLmzbaannhvHEERyfdjiL0E0YFclu9AXN8p
YGN3RmvLFyEnt/ZUid4JnkAg1KVGg/co+1OZHM1i3qP1vNhpLDGIs7emMUvEv6gzKnocpyJTwP0U
Sut7VXsJPctXL2CABx+2Gn8pvSAjLsCXyM5BD/+R0raL+oS6FVel2kY38BPYFyka3Aan97mebYe0
lSkCkQdH7t6f8nD136gltiRcXXBV/QmRJRqqK7TLOH7J1gHAI45HVWRc1ea82MNcH6rNtFEgfZWL
TZ4OT2VLgRQecURXwUuTa9AUIumzXaPU+T0KTue7RB8Mw4SSvsSSK+4eSGmYTILUPw31ZZPRueTq
PtpPEAFecSbuVFBrg83ZjRPO3X6j/XyGqVqQQlSORIFt4+Rk3g0iyAr+F8ehAspbWxBRaTIpZXQi
P1ZalLByXKB0H3rcMti9VUZafOpCFL1/K0UN+SsAm+OgR4bsGQmkOdhSPNbdw3fDylplGou71oPQ
gBRSVvzhYPIBj8UgtOvNkKfsT3+N+OK+jEz910Mh9DvUbQEWymrpdZCI/NA1TZNddOZvuFo3WiMN
dR7gK8aaaIUkK6U5VAUqd1FOvKI2LnpT68Y5a+7g78vIK7jJn+gpDnOiXKnL3CbznM4OY4solnE+
jSGJ1KsqvdZGJSdbx8JwmV93JDMtN1WUSvpYvUCkOOpF1N/dRcMDtTW2TyYH0MOpFCulBTbhwEzv
rO77g7L/gzfqV3rd8Pu7WlyBcVyttdANNiyqOqSF5xqKXG0hssCOeHS0exWdtiZX/FBs8sNey0E+
5Md/WGF5KuLUqNQ7gTc0zkVVtH52s+dOKFmD2Fx0mEqbW6KJa9blcThrpnbo1OI45TDek14uxTIy
E2skSWA+1QEu+eqoaTunLj5cjkxEpUgw8quluJlZegnnanHKtoCMtMXOGcIoAAVJDUnLjjEz6RY6
DQZXkmBF9Du/dK0hTvI5Zg8s6mSlYoo5I/kU7dASLIwGkzVTN6Bz6r6CDMAGVUFU6HHtg5aw1ls6
w+Q57tdBVMa++W2idspRepUmLjkNtZ+ZqiklyGPBGn9yIgDusUGBF05ZBEkPlJUutFMbwdf0YuZe
7hEA+tvrj0u9s6LzUleBCj7bYJAQEHlJihPofPHn8W/s5O2lPNYreqMk5ZWob1wpH/oqPksVQl8V
XXFui2Gvjp1Pe7r3L97Ed16S0q0hJXMwGtfmpzJv8x00VtiU7soA+NURZlePxThHZI6/yuAz+10q
KzKV4aGIZ7K+8zttm5/JShLjYYadvceRDjDyw0mRyfO69SVaYCd4Cx6NWDXvY1qj7APOwzPhqGIy
KO595yOvIakYs04zEbzrZNm08vxlBX0ToRdh304OIB291vEJsNR6Ew26+Kda5d2u5BonpQa3Mn8d
kwbB1ZEIwVLNHdJsgtNNtZ+PLwoVj9bW7MpoJHBB33r8SY/RcgSI+o7YZgusSl2lFT9ejc9YQej7
mW7wTsqtUKMtP+5YWLpDRYx9WhAkpbCWG+2Lz0Pf22qJJlYjmZzS5OO+i7C55o2x+4Fl0JiwGPHa
vK4xjX23ZpU+oXI8wrCJzSpwx2Fq8c5CqiAmzvwKjhkqXlJTnNgiXHqRKeHXHVCh3GQHHyGYVIvs
x2Mv35cofOHxBmALFDZO4quvHAY08+NoABqLIjlpWTimWrjD8LSkXMBdRjG3sQiI5pnnz687f2cS
2Y5RiMbp1C51T0OFmKZfb7qtMj5jpTs1JLxwM0bXpvmkizwdayGuPcNXexRKeSAy1YTTd9M/s0Nt
fNf+tDiSe5hUdJnWpfZNCrr3IXTiXMT20Sd9GaicZ4YIj2Ql388oNIjBDw28UoNzEbTZGJmit5FP
I4CIjQTdd40EaXbt6pFQD0yhYcfufzY6BRog+vdv3XPILs8AZowQlLKwCka06t6z56lHRC7fo3G+
wyFqz7nuCvESAv3KgnGv5HTgP8iIjM11j51kaLEyorUPwkiw42+oMK9EEHbkz40gk1M1HHUU9TfK
3+jz1/wjOMV6mY/NLwQXC0gz1Md84DAYps17kuN7/rtMJHHu1CS4PP77S/OJdcjAGDyI0FE6MgYV
xggTtXYVMRpyONwI5fvcZKoQob9IvOoDoSzD4SWiyvswPSCfgwlWGZWuy7amscRuSxN4HO+8h8mx
bXmPBoGWIvSgqsmvduENxf7ibp4PbakUACi7igXqnggdow3OpD27zQQz6MVFI6foyWhKILLUtUeQ
S1XQBpNd9oFpWZkdbMX/2wrOKRSaUjmhaqLWbH2H6TgJDeVoy15FSI9XQYZbwA9YBsEaJVwYkjhK
uTV48J5GCSiogjfUqIMep29UJau6qHs7NPYEDn/HJAgB/14TonXQwqPtB7VopblDAd6geQnIzBZr
Wbo0t8QcXagitxUMLWqaHJeZJyIIzQScOMgU3NkNVYGsJgOvBc9awK7r4uqVCxb8pw47eNeSF5Wg
MvEpLDwC//nWWP+yhpsRHHxH8deu6jW2txzciyNfUAjaWMBFG5QAeYQuI7C9/ILr0ei4eyuOjX5v
W5MR4GWWs/SqGoq5q8R+8YrTJBXkgwUvRMExYivL39tNTuXmUsjRVUdq5Sgpxayn8o9G2PHgww4z
xGz3bnYPNfsBdYApidsyn6UIxeWjAqbXQg7+Hkzzzwmgr27Be1am1cOVgl3smeQOhQNvQtO+RgB8
/0Ly+sCCLYZqgA2ee6aq7TAJJ6BMcQ6TtDdJET/ik1Q/gAc+tHYDxgGgnQOGuKneOvablSOWAP2g
CajpJ9HgKwmUkcAbe4AWIsm2BDC6MZWeGz8A/ATvAYkykB0GTVNVBZaTs0Q5fX8NKea07eJR1POa
2aVnndrvGt6kFrOaSygxXoHbrDMZZ4OY3trjMISOPEp8HnTUbzilFK0sY/A4KEp+34veqWL63tNb
sivjOm5Fb9hPcDF0/gxG/7lCTcNZ9jMPTRYDSB3GQPu8q/R3FJ9aiUmcdPxmuE3pPoJkVRRozoLk
KwDwNve3Ec/oTm3noxq4qSvaOkSGCZub3IdRggvcd61Qt1sx9EDu30JPAX//xUdX+tpsxwSA/CEj
BC3N4VROnUk44LmqNKGRJo3tO0bfsm/kH1lEnaw4EuIn6VZo1OZtNLUIkEbTdpwxQGR7p+sMh8fd
F2x6mozKXJ9cGZz29T/f9FDuyaq1lbT3wq70CTb0Jbpd3fQgtLkwWuSTF+GoBgJSkJE3W/lKxQU2
hLzwfht1+nxjhY6qMzl3uWSz00H1lnl2pGbQ+kVrvkniGOhZTMqXWyWlGgTHp718L1hfsyCQDe+0
/iQUpavLlzX73N7S+zBnm5x+/vZCwQpCxwbWxtXMBJu/fNgrjqZu/3NEfSVxPvzVLRUxDuRH/HKq
PSpz+MfQroLFGhe/J5TFVsGJgW3SrLH3ygmYfCobBkhvBGSejPn9PDK1nogT1J3vbnAJrNK9+REt
6df6t1bBxgkyMNtpeRWX5Iuc3if8c2mt9xAc1GBoj6IXedHEWmOpdwDPCSQSDdrrGcA1rDGWpdJs
Xi+1amy8c4G4aBLxhLqc8wYIrCnw+BY+dRowMzefMBWVvdvDOwACSKk/MhV+9LNv7wD85ALxOyZz
DEg+URQ3Xiz3Mg/qZCl91CfRlIXynJq5tALKboZfuEp7YoBPVQxjQfKm/tgJdS8NAPFC+Z5S91gn
Cf92Itbhwbn2cvKYAcBkN6Hm1fEWmgBg16bza+7aQZPS6C7B0qRGcDehT+mD01aDSAfmCd5E2zx9
NOaphqezTC0zheUdImN+T16aUylMz46jM1/mI2u/RtjTEtx2MXWPbC2180eVfohE7QG800ztL0BE
9VUacb5jXR4tnwLnyEgckoOH8tgTqwR2/gcFoaoWAhzdw2iVzQMMTGTai7e2q6aF8VxgUucUDEhp
+GCRqIZgRnyV8nXigEKF1g2rVYAl6AlbqaLleRQ/2XzcdQ1+c2v5cF7Lb5niLiO1qIx3x4NlsA+L
NLy0pdI0Qp2uf8imWBrjuQGBA/J3A0R+/I1rOSJNM9xHywYHAOAj2pOPm4sQpdiF0ExUYkUWNKAk
mm9LtR8Unc9uGh4aUoHdsJRQm+At3jdbV0oDfb0nrFUw5zqEeNx8jp1SzOCdBgF65wh3ZN4qcac0
+/K/cr+KDUOcLikQ3uZ+vAkbd6k+MwJfX9k3c5wvmcwWs8zM7y/qrqpZkZ2cZjCsxzfVWy0jZsWS
ij5VxADjk1f0IIFJhc3aUTs7OnSegLpv6sh++r2S/PWx/oTvVR/iYg9mDAOQsu20jTAyzRQcUrzW
zsSrYX2lHF9Gcl8zi7oo3MSQtSR8MOyRoRj57OEzqXWkKEGGUiX5dzy5gbTK7SSMkbOeoMt8d5zt
iXhq8yawNd/FDQ1raMnMyGzLV2L5WCthdRZm/4U7lEfnm1ifc1i4yL2TpLDADt3f9ASFSSHQSwx8
o+qiAmmQjseGbn2KgbhQLtcgJouOi5gVjS9vCxyu9YALnYJ1HA0PhwVxquqVCyf1eZnKWoEZ3sQD
EevIbQwkfM6vHz0AJXv5iG39X+gqR5glfQ0y4DhjhTp02yvegxO2UYc+Fvuzh2aAxFO7x9ZtvnN5
74Xc5qgCYFkSAgqGL33QTot/TTpVn5wDstXuIN5zuidAn/FB/46oIjwwKv5zmAbGbO/JVObhe2ri
ojAaG6E3P/ndyQte+Z9VE6hWu69tf0oOcLJZR08IrAzyHM12TJ4aCoYUIVLb3r2itPv80K3nlz7H
sdcRtl+woPIYkDF4NL6hRnAW4oqpoal8fW3gQ0fthL277d59GFIt3+kozHI+RqTkQENkKXIVtC4Q
YETWSqmj4dl2nnuq0WHNQw89lkecMXnZUJZ9h4Gf5NzayVOK0WhM8N3HfTCcIHNGz3Z3YopGtJiY
ah05DBxLlXVpvKHdG2KJNCG9Me/X5pTuOqnAzku4MMDfN5VttnSdqIzJzO8wG3GDjwYWqY6I1opb
U8/SVG7RYLdQ0/J7aa2wzLevytLwF7xRNF3u7u56LJCgAqTrJc+GnFcjvy0G1dX5fpyzHga95mO0
pm5T1I8PP008owdyba4UzSdoepp56NJLNfJKyhYOSkuBIUx1f8cl1UUSddaD1sWnHmMMbNwZTgTo
GLVXr553FSFGtF3nV1bGpwLZJpKeU8afuJ7Vcut+0b4LPFLH1jIip8OTEZX3VKrbOGDsZEe3pdjJ
o0DZwXVa90upCGEbssZOrZbu/tDxqF0GdR6Yrljko+sbq2DFJPNp85KcePwVskDi2huo9L1I7ibe
xdb5/piWzpwGC0aqYEdzACG2TgLmJk5II2NlnOArWdXW8hAvPwLRSBbI3R4P84knJdR8v3gsyq9O
Y3AgLSkM8sPYzU5OffzeCrAOKJgEaLjZCmVuFrTMbA94uU7aLHqI8ySW/mc+9cOmhZj9M7FehHrk
eN/tfhDPR5TczWm4/qDNxRdMSfNMHR4TyF1h38D4os8IT5HSjmOth72GKaD9lVGXLkKF0DHUT5z0
9No12aPWlDRoKA2gg6oWUC5k8YjP7AsCTm7Nfq3zNTWk5GsmlIgiFu4YW+x1cvC795j0tT3m9c+N
Pan94g89zhqaHq4ZH3q5ojs4wKew88Ba2Rs9FoiYGegzuMrgZkutfcjsU0q8hrHbxbZBp/xIr7IL
LR97sWEDEu4X5ZJnjrek8adBn38kTElqH82ajU79MLLD2blINMaaHMHEFaG9Gh8N1Vnnc8J7wX3f
DZ0rvzDNc+T6o1iGiUwNB1y7qwcvP/UbcT1UZ8ziFGepmKCyRYdxuAV43sjWzJ4ujFMcgf3XohIn
+odsDgtYDiCNLuP6JwmAPDZ1HxCBC2bbzkUMwkIwFCQP4lxq8lOj57+Z0dAkneLkdKOFaMu8mv/N
Gtdau5wiGqCpkRg5GH9DrKqC77Pba5CiTF52ovLpOcUaoUQKrwjJaV0ckmsdfdax0/6vKoCX9w2j
d7iilOVi1D9VstWSn9CKhQ1erxj1LxPXz1zjIYlSmJZzKANeJZiNtZJF/dTl73fu7X96ndMgnNK2
4pRGOjmkPyAI4a4b306n+1G2GW6oMyhtWpgDxUwDbkw+BTcrV4teNVv8ehy5b9GNUegqenYwgTEq
1VnZONy42JEHID+K6j85CUIBmZxRaLfC2T6TNKbGIug8AVWaXbRfC29J33p00IxmZl6o7CikPisP
nyfRMV40dIp1aye0K3FD5GjfwTtzUMVebmOeP70cUNunYfmYzPcYdFa3LPEShrBZBaJ5hVm3H2Iw
ZoMlaW+P571W6aUNZbUaohhUInreMEfsVn8zV2m9qdA5mAedekJWdMriiBL5EsT8rPSewAfWnotG
QfiyJuuPWZ3DE0xmlJm4Oh4hLpcUCNTR7lFJS4izrwuz1TD+KM9UxoIHpFBwI7rhzXHmxaLSHKuh
+AHsPJI6UtTOP74Fvohqu9zm5xRrXk0rSMclYV58Losh+HbPJigVmXdGcN8PeL+Yypq0IaVCmCw+
hkzaWmQqEQ9LgDSshbw9xgDgEz0n+Jw80+FYXQyG+hi8qj7OcAz4uf+xw+ZS7XzrWsP6jcBCo76F
uxdC4hURH/0XGbqwkaDHx4e5IO5MhmRRdcs2jXbk9gNFJ68AqAZ1U3Ze9Vh0Jn1fWzb4hdGEgoVn
cSaI1X2Y6qkWqA2xNMPTYXUGYapUCofg5pRpdsQn9iwqPwLVsECFEMndow8oUsp9wSF58Wc/VrzA
/pz4kmS1iqjyNbuL2SaBqAWw2gDU68Af79NB9720teysEixwiVSu3j1fzr+VS4N+ixMPDV/nvuZN
pgprXkNyvHY/UpipnIAtTUUgzWSDnav6pJBwy1yDBWlHjCL8qyiF/FZ3f28nnnqJQZN2YsEC6I7S
3DK80gx+0MeJoC2KMrNCmWTJA510pApM2RK1STanYuZDswwGGAaMP8cOYRRuqednhhaYvv3OqDeM
76T9PLXUHIootNLdHa6UGfDT5N3FQxn5yiIFlx5uPxGiydbC1IBh7cM5DGKkJ/e29mSbiR6v6KnY
LT9EoZTfrQDSJJiEJUPuiXEJo4NRtFVoKaqL8dbUUgVP4PlxH+tuD0VRPkSt5dTynaeD44KMA8hw
Zry8EfzwCq8Zo8NjwD1KpF1nBpvYcEkLymsRqzVDZHq3Ry9C72FgfivQrMlh51HH0R0yjfG333CI
uRmPUz1PgXvK3uW/lkBW+L4QM6DRJiIKJQsf3eBzXHz02fChNW75hb0oJcK8t7N/vdPWzKqe00VK
xT0PgSAi9fAld3VmXoVGFFLtyc/toEico7oAVlOVG57L9kcADiDSNqB3Ngl5seCr5KjdRYfDES3g
qvFR0v9DviSiGa1mySpoR2y6UrDfqnGlt7EYePe5uMZEt9JhytVO/1im+dIFrPmnYpEGqLqQZLpt
7x8JJFHOKgebCZ3P1ym7V4Xc8oM7HrGX88qtmTjLUJWZLuln+RP3P0jhfQHXaSMEWNouMCRalDpv
0m6o1yEn2Vv9tr+rBLfbnxkvsfaUXvB4p2/MJIbq79nvaIcByVHyiXEy/T2hd565hMEO/d1QfR7a
qw3dQlxLAkZ3flIHQfRo2/fs7Km0e63ZcyjtlYZbYPBoQ6LNTsIDbrFHqW88XC8PtaT3y5x+yQv9
dJK9kZ3QBdY+V0N/XyIQX8geXtsbmfR1vm4nYlEG4jdwSus/88zCdU0LTzLukA65floLBqNp8VpH
oyB8talOmfR4JTMSqrOTuyERnt2rVdiZn4KEC6Wgswp0/LYbxxJRqpUWKiRZbQwtknm/qpncQpVT
n25K+LbaynE0dysQjD+8HzD3LXyXUUzdPBBeqBvn2K9zek3IekPSIQBKhvJkvhNuatsE/pSUo6ZJ
A4yDNn4mz1iqX27SKnwGX36dDV1lN0j2qyl6y+yeQmUksnUaIEmEF/ZyWu40ic9EnF+0deR6dPJf
cpkZxi3QZDLidQil8wzcK517izvzhXZXENLxW3ZirCepbfLIuPfY6vWtXNWch7Bzi5dpanPKSWCD
scsRby0oNnR6cD6jxqd1mFx9QA23OGZfM70TIvGK+HNLjJ4Bu7sfkcnk0tEX2G9LbWV+tmxFYYbO
tcCK7zh0EeqNw8FWo0ayMlhWSW+i08z/lS7QskMvuD2BE8WewXUebDwSmyIXoponJfbfkZ782o5J
pteq/JC0lUIDuMubyT+kZKSoenfo9a5530TJL7VmERrj/10q4zGyDtweI32GA6lUZVQtc+6Tsfb+
yj8rCLdnTbbkKtq8WamO2gu9XuI6U8r0FZwu6MXZLsJo3TX7lcHy6NS0jWlM23gw+DIWcnT+GPti
xeETupUhc6aHVae5HRCaJySGm/tJmIPIR63dghgrLWH7zzfN0krTjHwlp9HVW0uSwiI8hGVC9E2k
v9vT4DeKyQmZPAeeA1uu5QdcYroRwVV9ZUISaLym77J7Km6QZQOilnjZNeclwb9pNMDkDcHxNHfe
9/HDOGMGbailULX5vcuB2K7tLYPCh0hpw5ypyAIjT1zE47FrLj+NYOuJhcjEeEv74w+daPWUP8rF
wcuENZF9HnTxYuM9Azix4pIrFQy3YN82qb7KZENg1jHfwurLOQ1h0BXnRc+IIldintbeTaF2kjHH
hbEG/tlsBXQ+DSfpfaf1vJtBX9T4G61BL0w6kfrd/6cejchj10n09dA0xQVyreUqvFbwnL3H8QKG
AskuWqE1h3OTWouexHEejUH4BVvLiZyHXjkjr0ZbOYOL9bcmRACj6hPTseyBvpU6xcKMfu3bYYsm
LMS5HxOICMb4Xc9DSYdJVwH+/wa82TzTWNMW/UGylnnPX1uA2zRmX6CGcBc6Zgw8H0XMb1w9phkA
m5MWH0czGvzqiaVDmwyTFT2dKencTUddW0TjJzZ03UsUdTfU8QWKCKSfmDbwkd0QZBcO3xxArZmC
Y+5K9m6kTuFg+s/b7sVomVQCTWANp/QagigEArsgO3SZ4M9K0ZccJLx5eAExlCFkLEkP+Z8/Gko9
WSKimeXGDrQCjMQPk9z9BAEa2pkKm1O4ScUPytttqHNCW5cWI6Wlt9t6CU1UfsBP7WO6XrhS010P
Bw1ASSfd9t7+g0MGxdqOxP+Bt2bk++Bu4K2gb/TfSBqrq9dqcMI2fPYpz+756uPKOiKcooSyu6Wu
UzwnQTdDWlxPeQQBUjee6Db8++ZGo8eVT0IeReRt9j9YrYpLJYg5KbbErbBgktfF21F1HZp5PDc0
qPP0C4q4z5D73x+bAVjsh7+1jGYCi2tVlaKzFEyapu2gN1HnH1EbOZAd+wANRWYKHKQ/cNIwSmMq
L5GqFv7QltQ3kk/Lhp26P6tsW7ouOUWcHeMe0SMFCVAsLuGEMY3ON8Go6enmWYhghDfVa6LXy9FW
8UdrummCayNeYFvkMmW1MaQW6kuN1o5lqHFfVEsg04DEyjMLnWMbuJoRxn3SSq//y0NhReYmaths
6No6D0r1hgn2kqLnjmu6kg+6mZz826ajsAlEGcestwOBmQ0BfOqRVblCzsLGBpAroLnTbg8IGQAY
90JCfEmjYcQvLeWvvT6BXFmhYHa+pP0NVwH0hhJJ5OS75tEeHx9/u9CcBOluo8sP0iQaRnnik45a
IHDzYAwC8P8F3FZELm8tc/SoWZp4p3wwmuaNDIVQJFFbufF+vmB9019h/UgPqKg136ItNdpkI0sC
MyLwcjW6Gd8Va4yWT//mlKFBmBaNUYi1L0cVmW3chl+7kgq5LBA9gPdC5Y8budnDAbv1hhiQ/prj
soEpOIR8DxO0ABoG4fjdqa2NS9QMYGvaDFkDVFvWXRxaMCfgcPST62cEtujpfoL3VQitOj/syn+e
j9vxBov2ZrXPBRBrllIaQN38OdEuJISD6B7KMKzFYFDzjK8fsPT9Oh5np1L5423XIyhoCRVGwVXJ
66WsBh77Ks4uaPZhxvWYHHEEonSGJV/BC4tSlSgRs9YH/h1Vv7bXpuF6YzgBGyoIBUOd38wSBkLT
ToEYoTPMjjGvea6IPWBz6p7AszL8DhiG1rnqMEzXTQcaKrn8mG5RFnGrWe6BVKoMmlR9jg8si0Ls
RWWXMq0BpK1/kpEL4vWm6A5MvtPjgnX2AmOOY2yOEbs9AvuTDorNYRXoBgUKUOBIFIPbgekahnk2
39tkWrZT3BHxkp8aBc3ydg6P2kzj6GPFh8CFZ2T28fOgjSAqDqVjl4eg2ixPwKYmH7/xoa/Pg5Rn
ywSyXyZ1nZTZGFAU9PWoa6XC20T1EFNHIIr32tuRdNF5R2WHAL0+m6oBhEB4aHTZ8QxorjSAe+gQ
V4IrKyfU7e2+19vh4ljYUBKHsbaIoKzcjseLef2wGpRVzbPNuy8Wi4+8peMSRrVJ0B15BC1lMHQI
zMX19VPmPjMHETWVhpaR9Zay7ogctJ4S5QC5oqfcvBcBOy8O9l+p3aafOhjMO/hCnkbufXwjGiIK
nLQDWdX7j0ZDheVB76OSCJOVE17oqsWJ7SIMBMjBwGUg3AWRZRTkFeOZiaBNtSAAB6bGo7u4bc9c
U0kt0iqaNS96lNVA+58boSoCmSICWHG/OwE0/A3/PminzhWJTKANm8SdHqyXiGHw5zSnWpXjTuer
QoGwcmdxRSj+gcOd7YsBNoT6GI0xzcvhHaD65AGeew4LUGIyQAnRI9cdCZvcMhYQ3ri7lYRup+qZ
cj2I4AYCvtKX8TtWQsNs0/vWaVmgG40DaJOBJ9ecq3U51LGOCCVHFEIE4STVq2ZCUMDJ9naGLOl5
MglPRo/1D+eDnHnJuAEdXY6i8ZupDVQGhasOpZ6yBK60C0w18KzVkR7ImNW13TDC8oH/+Oz/zhj7
VJKgpDq+MHP5C8Mlpw2uQojeMhveLxTrUY0ct1EH9PXwYIFIg2D5f4TtP5Ge2ensDS3lKLdnC9V0
40WmVwuqrDPoYlbuOyrTKwn97FPAoTr101vb2g72qqIq0m3gHZYr3Gwm3MuGxxBShqn9GY8vska/
hvQ7qvoq5OdTVuCEcTJFDSmTaCRjs3ReKovICOqr2X52crNnL2fGUx/W6meifAcvj23JeiIyB8j0
eysbJBjSmjUvO7h+hla2yTkW1CXxz4azTc94KzonisyCh95LiX7KUXipWk6QfwJCDHwqua8PILF2
ixvBdiUYZB0lVMoC7RfL7NndeupYCf7mGwQeHXrXKoY3Tf0arjCpbiuO9ZOV1Yu2BH2SpM7IyEsb
92Kbmt7JCCtPYg6c2Shhc4wuLW+RUQ0iGeMWXm1Jt8AHR9zkLQdbuCfJFb+oHY/FaQIvBicqA71g
7WBJ98WaPczDJ6saheYo1uCJ0osKDekK6kLHL/uNPmsRP5b60puZOLs7JYr2ZMBc/aiSRGWJMTFY
T2X6IIhhWlHFDop1YelhLBY7fteL5+ht4M/E/G5LsNbYG4aVj0Ufxy1LLUclZHWnVSZsRcVIH6Nw
QKX9mBkxGZoDV1hCptdJ1IYIe+CXmT1u8nJPpkiXO3+XVhmotT+TMsPuTdPG7nj150WJMQmDx30s
USDBOwzGQTmt0+wE6ikMlM3iO8dljnVhyJ1D9brE5hDM1gXIS9fASv6+kA84Nj7duL4ln0XWBgSL
itgOigTd64YQUOoQbwcjIBpZta99TutKSVtUvN2jsLCAywbknGbUJCs7jU9aYEBV5BHXR7fyjqrH
BFtDaoaFMmRHewEsveEjDcKgW+u9jpckNj9ii36QwbIQdEq+d9beX+ycW+yf90pdkrSVRYl1DXxV
rOtA8GBG/55fmxQdKIE3Rzx0Rky6OGYwYGPfU+yY9vBw+TNFYtgYp6ziKua1cWx3cvA+NJOCIfx4
lwkLX9/3jNh3D/GNbjHOE2f+ahJOCmkZpcDDyNlfkSHEe6PiDq2RTKO7VNct3mKDm64EJvqab5Av
gXDr5sl6ayd6m9IptuVOjEaPIm8I62N65NR7jr+S1ZYz5KTYP9UMCZ6y35N2K1RzxIt8ZR3QgBNF
a4yoDBrRi7MuyUJyhiV0K3xf7L9pSvCvyK7e1b0R5AZ/iFKq7pgfObW7xOAHmYXpcGVVH+9m+Fdk
dRd8cevVHJyAMjNQAzq4fFzarbWa42ZyV1ShODrYVT8Nv8QtBx1wWqXtjxrs6UBfF/lD55ygbDxa
VwfJV54l5nNxq/chQM96cXvqPk/+YHIMZa7pEWImiVE3rI87LNLKNVJj4GuJ0AJ0/wKRiEs2lUXU
RsP2cbow6HumnrKtRcX0EBZLx3aAi5eHDLFxKCX5EZQQ7i7yRvcU7e6C6SVCGlaXkAjimq2Y5kma
E8OzuE/TCTmacCDUy4PQsSHNDa6G4Ib9xDrFYfuDs7rD7MOUBK/TJlZ7bmIzNp6hh5QazEPo0j/z
4DVVgIWu6jxY3vUlZxt+Lc7osa1XKDXwQwjy4+NQR+ak1rO42K4YGGW5z4qVyJhmiqyXRstRd33i
L70Kanr+lp+UbYN0fchb7aKznmJboZouPjUVxsP46GM1zP/h+JNaULnZi/Zn53lNl5gPj7i2kkPr
I2iZSD2RvNgjHJFo7rjANwpP0Rpr8dgMUeL46KnevgpFtE0C6NzbJzcXtvkYbAh4Q4870qLvjWBp
mhfn6vkCfS+Zo1kOhfQmL8weDnjkLBYBjIVl32LvTACH+s5SnC/9t2njDnHpkDNR3qiekucq7fQm
howUuHAFf82absocOAt3kr7mEBPYMloPEtcJ5Ks4/ovme9soQ/px0ucfRzKvbarI+WQn1GEWx5MI
g+dMB2O233+7mYVMDUBTvDwNURoOGqK4tJlH4oSsHEA9tSq9kf6PPiy+Eg1wDiA0wkT/zSjor18i
75Nkacaj+zqGll1MqDfALk0wjZGQ/UwmS4+xlRi83+Eplhat3HCJn1z1J4b0N8A+nmSZ1XB/2Iky
2wHLfZLWWJ+hu1+ZdcT4f8b0GI//YqBTCNFavsZOGEO8o9N+y/bFwWOo69woAfNnuY9BLBnd0xIw
XPE3B5ORcavyFL+cJHSrzKPd/qmv8UAjn6rMGdmJxDHai1Bw+6QBz5SmcxHTEr9VaUXbB149NfSh
BDC52YvbtqtNk8Tcx/NM9jC6UvwjvCmgUhPXR72nmuVlQy4dk+NnF0sSSnKeHvshxYyuW5Iz1Zpo
0qSLqSHVaIU7XTgEX/Y81F5Bt3a5k9YBhhmfXxan5NmoxdF4uBEcWk/JVw6WrzrqXAdD6hKwzpuv
Q7Oqj5eLyxEynbP5N5wimZO1e+ry9Nwl8aw4vu3Fbfo98snab9+OB2KP65gMm1NrXe2N0YblpYFD
HrpCOLA5SkfE1IVTlJ2fuc7fZOEwtUlgoT92BFbU12B6g3DPq+n/5RTsymhvKSIccjFgGSLYkqa1
6BGmvR43sQGYON3IhOFOk4UfLjyWWP6Ocmr3FoQgxS+dJwH6ghzAzVBesfzxTXt+NUOrM+IFEI8F
yQM209cByTU3Fu01NOYXKZXZa2y9zMecRa1pU98LqQAfrlImfOXX5waedCEN8pYFjPPPLJwGSNnP
rtoHit6bckZVZ8ac7U9klUGWZeIN/Oo9BEF8q2IZBhKjh6WGz+UhjrptlSSTFvQo4n44mPt+xKAj
uglw393+SVzQNF3granFdourTUwcZleagrn4NBk3N7OEhHe7/QJy26xcTYZf05Ta8bYpfUepj/e8
uFVsiUExLh6JaeCA5F7dgiioXQK3n4+N73L/Apd8i84ZGhUe87+tdXVAX+iS2yxoYJyp2GGtU+bp
yNpMphc8CU1xq4nZfXHaIRxaust/QgdfMY1DXE8T1KwDDrH7CN61g5LIkyayerPkapOml+Sc5i8z
WeQOHikL6J7Ixazg/M8wLtBhxfBJRwvDCMPnL7zYZiMTOCS0ikeaGRWmS54l/JXRVQR6vIKo5Z7O
x6wqT6IiFswH+9KCNJXUkGMwkBIz1Lk5y80/HnmOJSxLQRm8LXeQt1DUc+m3i2YK0f/JNO0IhZcK
uKAa+AqUPE4EYTnQK+5u5DR3mYjuZIK6KUCA70yGs43lIGIW4xK4ueR1IKn9q67+eOPpCu5JJgSq
O1l4i+mT+rypsh2dH244RB/yUQpbv6FYBeOsSNfZZ5INALXa8Jg9srv7MVa/Kay/rOqAXLXPmurd
zlMgO2vdtJDvCabqY1F93Q6j9S2SrwR8GHnLnyVQYa9XWrtx5wYi/R5Vhrtgpr9StFsLr1xBw9k4
bkVCeM+YlQ2OLJhc6vuOe1jyM2TxjteW+09gc7m+I4IJcN2dxjkS1SYIi3kAnYffYrvpFt0px3VH
5i+BUc2COHAyZ5l+B4AYD8QDrpEGyPhVMLiUFt+gCooB73bS0uUyGyipymL0FFx2L/OnK3cDnjpS
qrF34wg3SveVGHdd8zPaLyR2RkrfiPpR76BUg94Pe6PoOTRhqWCjWpooT7+EICTosKmooxzowVNZ
1Q1juhnvTJy/Qw+KLYClxZzV3vJt8wk9IhWy9hFpQLDjMiBwR/AmiEt+aebxESqcDmnnqC/FrquT
SA9Ny6Awf22fHO09/PBFkRf4zj9YTZpHuX6RLuNj25CFVT3/PHQDNDEXcu82GQDGmlIiHl+MXto8
b93uvyOVrqyvRQlN3QwXGUZhk5v/JvMhXfsKiG9Ysbdno50OBijjQELTHhfqxDUUntgKqz+b1Svl
N2GNbHPIsu7o1DXk6sUECtaBiJMng/YfmCwUue1rpYSDpYlEUgIzVYg5P5kDGj/Ua9D6k/wTMka5
dpdQjrdPea9Ck6xjCDMTnar5yZLNbSuP2yN0MjEHre0oVO8rxcpR4w7490WtkOuxQBPZzzBdmpeE
ls9g9uuapR3CRaw8P5TDY6KPFgloJK6scjVuLeerxV90THKaSYud/Y1PYipky9pnltEvVN9g15AW
cHHU1jnt8E92esNSrbkhIaXWSTggP/uMW3XN+K3s3OZtcLE84ln2KFqjxrOeI0GA2vBaddth+yIu
F70v8ywrhqyhirjBqdR4y9PDUQ8kjdWWsYa7RFnax0+/lsfdN/chBBOeM/mb/eCuQA185ypGJ60S
AdlV5wqA90N9Kyk6jqz7Erg6Z/LOCb+q5SfqlWOz3BObds+3qdU06CET33ZCvHXNWXoDNkaPK6we
wimk96aIdzIJzcTIQX6sqV1wH1kcd0Hbt/qiwCYPRV71j63tzELgxE0PcQaJnL9x8h3V8Zz/37S6
I4D2qY2vUYa9JHBF2ufA8cBAKFrsAs/v5dHn3NzxNlkzS4B2ltkFvZG/DmQTxxsKmrEnonypYnQm
YaCHJIEv2c3hoZK4mpl2whknBFb/m2QZIZjR9yseD3Ao561jsTVWVTovlml45T0/rznOeIeshWbW
CCDGZabzwRy2a90JJWqNkK9soVYeyZlosKeFQxiyP6E5+4lYt3UdyyQHnIgQgpE1MxZMJ6LXyREA
i0U5KI9zOlVfJq9WVEgzXU/7TypFfJCWX4uL996cv3wbfutNQmPyeR9qrJKPIKdZ84JycQIsr7sf
0kYo6sbas14SbZgjyCmWZc8iKeWhzePl3aL9K26w5ol36/5Erp2Kpw4kAttZQTl8NjTdTC+d/GHx
7x8Dmic3S31k86LUlZbbhsSzvtCfliIHflvdDa1oOrA4RfIhLn3hD2/9kU2zE0ixNNLCDv/A3Bcv
vHo/CxaQGPh58DPbE0hW+kYHJvmekP4C/cqs3jhJO36fWWiAetbvGikEuEgOTPrVp7kRbOxhH2hb
6xNj+/wPykA+qEUz47R3vkrNYzcJajrdLC4j7wL+zWGqGBVMAZnjHJ3hc/X2xeKHFI4bzQ3XUiwQ
kJpFQOPWqS1gw1rrH/PM9SWBVmahGt4iHIg3b2PxPIENP+FEkjglTHysuT0m7rCBptUfA39Crqr4
tMTpBsF6bcWnMKiAugemaDCziHCEDfP51Ssee8Rwv/SqheABPq9aeLdaM6WKmYnXkE2ydkdCzSfx
n924A0qqD1R+7U7fTVKht7mQ6HsmRBrzX3A6uf1Gn9VmfybI8g832oYEETAoHKnqx7KrMHLXIrwN
DU3AmL8TlW8qvFmVOpPRjnemBX+ynoPnUjmO2M19n6riJVVCDzL4n9jsktYTpG9NUAAFOg6/mIeJ
wJxVWPg9/RiFfWHLQiUoTNORiQ8HbuuhnUSRnsw8FLWu99d6lbV/LJDeEvl5am7YBANVzNLISvO0
WGtafPH+56kljivtvCo5c8BnPT7fzBCE0DoWbUkCjbsPJYkpJcHXBm1+8Zgho6dA4oIASomsYvfK
Jc1s7U6Z63dxIbZRey6px1c2lNS1hMs9lIPUMJxARLR9LEQyRHxcTTYVWVcPCmG4mHZ5bv42ce+K
qjAjFtQBb8g4ogPqZrv8xw4L4r5b0cO2g9Pk6+bKprfgGvw2dNsiZAGh2WWDx64A9KqHMNm7tR+a
Y3ImYjFslydUh/nFUWMP4GV8aenk2FN7yqjpdG/fk6gUubH7GGDwgbJc1k+7xH5WeUGifJD9KeUe
DZ68W3N9USvr7R4LHsFOH9Euh8LuWf4ruc/TnQiHlsbrMZKxgESekdAlrYcfXMRJeAUz68ydBf5G
5RrgHJwzHp91F8yxjZ3RtTRwEOgFDW3eKMBCK3/fTlXSwZ3xdV5HqIKPAEva27465rW6TnM7r0O1
NfG+rmbBnlHSXZ8+imEZhPyju3fsymtkKEr+ebFq/MQsIy8UGdJCHjalrhCwWS1QkG73je6njJb9
92g0m3u0ql0bgXLzJYAw4yzS3oQh3V5OGm2rTzgTnmqUD7zE9PVmzrKXBl2nELMw3R4bay/suUJN
1Z56QhCrHpAFCVTbBnE881EqD7rU+ge10SuA5pJjalEiK5ciP3u0Gvqtp1VDtLrcb0JCwq59wfFf
iEzAySMuM36JsoBFvyQYF84Bd/vDAU0GV0UsNsyJQxLWkT6hgcm0xfoDBpcXVVccdEhEz56NgT3d
7dJIfhsM0wD9Obin+fFeokBuFJOdfEjQ/g+uOb0e9lBKfpnFwDjgREhAZ3i0Xq+EezZyP2sBbqOt
+Us01/4C72sUPauvQBsjF8wFXIel+CJ6Se8Ox2bpmzHQ+Klpj8+ZmjeLpYfYmiyNaNPmWvUm3Edd
H1DvWORTo7odjK7wdnXR7bOrzrZzEeYSzf7pkvHMcs2OCTZIREqWAx24DWPAd6nS6q9UiXtfJM45
2LGrW3f3p4GeeaBdZJj7Vveaei7997aLxUllhDEOL+42lHhRN3U6SV38OBcElRvZ1gtQ0RTJNMO5
qUQdPBum48v7pDGHCU8ap+YWV6fcNa7YakzENCVv235oRiNpQ9c8Eal8fPpEvr5IiyL9CVvqeAVW
DvZxgepSD/JjSEdIarz0WK6VJz1GwbZndBHEHZEGzNIQ256zs3H2jERQGurLN4QwCGGIPf4GDUn0
Ogtfy5Iz96mdCiHz0953wlix6FK3exYpEfgcNSfOO/hs9ifwfCih7bWDTy6LFDXpk9SrsoGbd5Le
era/jboRzdwLUGKPPiYJimrPj6jE2610yBlztcE9B6ahczVg1qpmfYKz6Xr4OSDxv6/Cu5Q0hsYa
Acx0WSBMtWPzApw+C5EXOBfUYU/jjMiprhwQfhXwT+2JEpjZtp5Cn92YBWfDmRffoWG8aHID1u8F
hofbaa13s6VUBwKtkCxC5UxEGM7eZTuguqNCecs71bbTJ94cGzeji5flkMrNh0sEDKN2tir5hkSG
9LVumARS6ol2hIyfKPtqtD5yqj9CE4/2lAuff5lOsE5Jb9OuNzcgx/+pIpHco50GUiyMIpK9WGsR
G4LzMWXxm7pLgStWkYcNozdCRbGgiqkorVI//pcWt83X72ymY3GLfx2eg7A/Pp2iwqkak5UEba3L
7v0piP/+YTJmskru6R4+SsHa6nnFZftgUXnNdi54aOqjled2HBqpUiphzTzTxZe2wI19DjmsWdbf
aezp8SoKUx9EPkv8l+HM+HPB0NZhLltBRYkJBCovB9aomh8b8jW8wFCL2x9vumy58YchXMeAUNa4
fpCh1oVwDGCge4VUTVbjWnySvZQNPyvlR9Ro4HhrVIKdRQWYI5168XXLB9OxmPuHWTR7tkcqV0iI
TOrCH5MvmECODlA2Z7Tf8ZIDNWRUH379qsYRJArfNKWYYy0ktgMMQFz4NkvRvw3h+kQrzeaADrYv
Zlt0/aMXlNNejZnon2ebqkThhGmg4Mrle4AdoRdDL6bjJW+3PRhamSaeB6PI63djbNhIvpaP4jsK
gVE6ew5cMWtP/RSGbjpSQC3ZRkJlib5pmLyn21cqf2pk4xKVF1bxXCrcSndMfZuFKHG/PSzymGYe
GoEiaq7OxtIfI6cBb7Y67ZDN+VefIAei4egym8csoLDnhoZ32vW2XMOJ08WxKtxW6gEJsHe3iYIb
lqGxHIqb2EK87lYE+bwE5FtR1aTYJEQoa7n1VP84bSDfwkTHE6rJ+IhbeJ2PLnjdiSSPk8PGClSf
wU7jZYO3mBnCE7NEvpEDo4ek26Yyb/2sa8fxVU3QWsEr0PTnrkVyhOfjwb5UQwRv0tfnPLPeiAxn
sTFaEQb7+8RIPTGjtACM6x+OqS042uNTyf2cWkU7mQjBp2Tt2IMWjG0AdM6QJZI8kRAavw7p5xnS
wS46BXjbTi9wzE93svvGu2BYVBKRUw1/hwH365pELfLpejA+HzSavPljFKOdKpAvcHiHqbpQrsK3
xLs0iJvpZNDxTDpi0XCmD0kvgAcTAWQ62+Onal9pHN4q3PI2FDKH5w37Khu/uVAZ1pyByAod4GM9
QzHIKJLmhg51q2BarWthHRrbxoMWqTO2eA6Ee8jrvyNB/MIVNRvR3MmHf7p/Am4XhzeLzKdi9Jj8
gOHLZnT2jz+V/w7F/WitAPtCjp87JdS1Q1splpmPYk3AsewlyXPErhj/fifdTs17w2fkTaQy5Fam
L0jQYQ+sF+7rANm2EZFJpeRku52cJezduDTLWVZJ4AEWupzkjQrNCLw446ffl36q4h0FsyT+InBg
82CGXK891yfCEMiuszsGnLQsyqrmM43rUfzqzrKFCC+kQeaWXrPPI2psanYMSO6ycictAhLzRCp8
smaTB2n+P/Lzj/k182QqmsF2jLISpt4WVkhjiYxOlHTunZ8gI+bPU7ikeZWW1PHKfaGbbkNAG4T1
jb3nwPXqlQ9d9rM86oABX6cAb2uW2jeW+XRKyBTzrjTSC4UC3Cbq2sxLep+lJ+LsVlGUgeiUK8xU
/VBR3/bh4duFkLL6WOP40kJgegH2vDx8AiQJJ6DMYaKTvs8TU30rAuePIGZERs37u1KqoskdpnBm
MZSlbzSubGDJ7DBBHzuxw6OZsu2foZnAl1/YDYmJ3x6Uykp5wIUFQUPOkirXzZK8mDeIiGXX8HP6
8s6fPrbXy8Nc6fNguzzizxk+3939Y4l8Qd/tCILPdu4DGa7JB9R30HyHoY08oQIgPNLTMBWj8wf8
wZiAMzBOi2YsJ3oRcYBTwW88cEUCNLgjLpUDE01hIrvhzEgujP56icEuGFSccOnwRj9ZqMZIJOoq
/3waai6lbPnViZtm2cCl0aLV69tzmPTq+7vvsFUVadCUf07zsDI3u9sMDF0C/ZOk2FK5SREadIbg
NBHSCjv2M2fwdcyegK5tsdOeQZFLN3xJTHVEe4Ekjg3xNl8pq5s3f3GNbpA0CxE7iwBGolN0EWcf
SOR8x7QnKxSYlPozeNI71KK7mD9gjXIgmf6DN6nsGoX0iW+IaFDV8uzKcXmV80GQZIYAuK/HbUqm
GezAA+1JGCnqja6SGrMRTLJw+zLM3gdiX3lKRCCjAF+wrjN8NkVQxg3HvtMMZKrMUDZk//etsi3+
cKt2jUgNoXwwDScX5uTT7Q2eS8Yv6wTP8qYzkuyelAWJttEvY/+edgSSX1NUmdMg31pICd+m5as0
J80wlPbuBg8LxgW+y8DUG7+9DVvMjMEcJ3UFIbfgJtde8iUmIi69h9/TkHNmdCqH6PdB6lqCQl1x
fVTcikMD3K4q+P4zUAgO7lEkqDzaB0ClDXMXrtxoEWK5AknGxZTckmM1Wt8VEByrlegfCVqILyR3
dwPO8mXiAQNxzO/LmfTg8ZTHMxYGLoLvoXjUAuIQDzqQ7JqZqf6WOFYswBPN3hna8LZXLTSVjRKr
Z6NYBkEdBEYmI7o8cY4xnkyhK7noIiDxXnOVTuNt+QPKPvbdYzZvJvO2xHOmoQBgea1hQ6rOddy2
EXVvGNf1HXJvPptN/+I9yGoLQ7xCHgtCa9nBYxXAv7csR7Fwvchc/taZlph6npS/RbO3Umpq1bwr
2b9GbICADyRlDaxf3PxGxcNv2ougU1NHgITy95VpKAaI3/a1mMItsxAZg9mHM8SVvwt6Lfyerfbw
+VuUiRI8KfmE/0D9BaO0DcskeyC+Zm82e7wivfQhMsIu0z+4QiYUTej2hjmecP3jMgEBMGT4tvbx
jD7XModX3QLBkyJAYppu7kRFia6HmWL6Ca3s12WX6REbBTBt5xfqz3IA912hr/uYzrScDKUCuP2t
gTk/yhF9VylafP2DbmLMdaA4zBayGx2XhAw4HKdUjJVgDHRovYPHsNvq1ml2RqUW07oX9pPMwWDC
G0rbeBpQk9/w1+wcC9JmPLJbG+GBb8pMLBNFTYRUw84nSRMQM8EFKh8fwvcgzBfvslW1ux+sVqzY
hv0AzjXoVFgVzPS0j2W7z1CdHpWibJ6iIM0cOxI43xdPl+xnRCc9apRwSJMlywlTZAnYF1xD+pyN
yOs5/5IUDkVeKZOKaNdiIVR0jvmlYlN6SfG+t9a3z9WiVCM8tM/U+D2ule7ZlfIiuMCilqW5bDiB
jVC/kRtandB4g7gqj/5NLIRIwNZBgSh+wwaF+xzGcXq2Xecs0bqHWBPdHZTS0l0jAKTQ/wPu2tKv
XD+s9kAYty7JDnj3skhI5me0fhLhR7Ru4gbg1HeAbyPyZ57qrp4Yyv/DHmKbuOLW98hL4Fh0gVQI
sY5CKWpTjjm+twf8JQ3rHOTAGGq5c4qBKoDAmoPn0mSWUtHA6yk/S4Gt4F21VgSSkCtmNpx+fuRp
V2xRqStUxZ2BqGkC/ZRGgKcENMc5p8FwGh3kGpI0AlSzbO+932HaeNyrI1Vl6NQDHhl3mPgszzp2
xgocfiCrB+39k7UYxVLBF122GbH2cqg5wTstMCs2zix77a7ixUExSxYbjHtuI6rdzJN7BsvcwU+W
/pl56cQCHXkzTAxdNt9S1fVau0mNY4Lyew6+YR5DY8mHK5+7Wl8u362BXu+yLJ52aTsw7xpVLUiS
xf2idK9am1Kif57+nB2fueaq0O89U8XMFecA8EFJAgN7rrdBNKICWg3gPcepEsw4nUL9djnYcXpT
LAxf7SBQuLgFlRXoktY6FBtuofGoAuF4F0SMe0SQrQQ+CYjamWg7EXttQ4blfnvxNg/ilvwr4hZf
onfIPWgokelZm/9Epv5bzZVZk5FirDPFtRXq8+ObT3pjVBWEzEwmUp5Oj0pBUoWMH7C26U5FTleT
n/T71bP4aRQBkLmqCcSlXitrZrTu1PuHPCWewb1Qwfbbqky9lzOdlPq4tkiAhMrAt0gX3BOpL3sh
fSrs5QUc/mNGs1r0XeL58fr7ZWec6D5nI50bQuZI1tVlpMEn2agEp2WbbhcDDpsJ0On7+TJis6Ok
693FdMZzwJi17aTEOv9ZrZGz8Rg88vHTVz+R5mxH1HIuthDxUYdUl0uJOcCmBuqRe7Ef6YrqrRCC
guzPOBzRhiSK7da0hYvtnnOMsiHh31B3h+4DE/uoe4Tw/gIQUTdNUJLUmzQxrL2XFwrVSOAiS90D
gn33L+VkcPh40UM/PxIoyGpjkDxwkT/Bp3me4hyX6bL2y86y7XcCVUAzzYp1KfXSnpI2SQfePEEo
Wq6qD7DXLFoscA+nqQEOjEWb2hGke0NDM95J4+z+5c1tA6p/bzXW+zaIEL7SvDz2ojwjrWkAXrQv
jPPNv83i8IQm7F4syjmhXHAR2gUrOKDbPjQwjkOx2muUezuG/YKjM+OHhaJzJaYxUINX7D/swaig
wgQDupT8YtZRfP/QjQA0k5D83hkNtD1nEM44IwvhL3sRWMDa/xLD0RXl3lRzyhnXKHWebOtfSDkP
AySa7fNAShWf25w5ALbGewjSbSvmOr54QYsGDX2zKoKVUa6VTgUu2La+/C0KNfMIsOKJ7ULqQt08
UnNynLbiCxL9lkYv3KGXjyP+lm1u/yfK8TNRkd1CebsUi8j7lBwR90IHtX6wnldFXZ0qeFCNyYYt
7AvinwLcSqCNI3g+q0sgdE6p/uTASgtDF8wNRb0clXJy8I6rc861ZYINyG9LBMjVJ/nfdCio3zjO
8FNBe6qxaYv510T8m4cCPdsG+6eItc3WELIYGeCnxyKqt0LmYGj4fkzkSLDgM4ES78VIAWrad207
PmjRITDvBgzoafzTk6SXyX20BHju8YtgtbZhlC952bc3c7dqnqyhimhBrLS6gYLXHBxFlv6Nqk4v
Ee49gEGFJ5nAzdMJ+pfwdvNRf19+OLsMHk9VAzLei55eBvZTlbQV16PMeQJ3ql5ZZb340CvshL5L
8ibuN2gH2SQtWVFwETpzfcW47VcZoemYNIEUgJqb5mOgTXwKqsRIxQrw3gLYw7JFXyT8ZA2McqpG
kH9fkz1LbWRGPhg9y8KnL9wTQckpB+Qj/zOQcG9lmNcWwMxKinQEK3DwXJI0A13Oa2mNxRCJmRSd
3uXCR2L5juR9U5eXgbPd7o1nPL9/BWxtSPv/orjdPsakfF2vvbX0bdJ91b8vpdG3pcXLro4ceyDn
w9nwpkN3V/3btVYHt24HNYV3mn8Wb6p6Fq3GNbhmF4Mgs1TP2iG0l3QhsNkcI3L7kO+jXLmDjPhw
Fap/G9C90noMjRk6WXo5swb4yvArM/PimKejlWldJEpc+u0wDlxOn36Xo40zh4AMOS33J+TTewFZ
VMv88nKZJBkdb1UW5dGYCkgOQ9OlHvPQgxczT+k2/+NzCIBTu8kaFJbPSgS+nU3vVFs0zwpBcgLU
a13RNl/wKdZ44fSD6WiGoI1ypIIjHL3QkdO+X/vURfs8VzS9DYY5nTXgcbRAat8RHi7SEO5wpJXt
wx/WKGyaMNBPUDGh9vKpV506oMcD10AFCf8/H4B8Unqom5HAs9r/40xlpm3iyarbjWqwG8tkuA9X
e1Hbhj2bF+lses/LZDs1+6g/0bilioyr4uzTtMgtDNunt8MMiFCalrSuLMk7BuQaJmRja85z9INz
JZNbKfqWwg4GA+6N002rVhyneHfD7rdtvIm6oMKGVQ8u/dMlIxOXqpNZItSSAdxq1ATGuzAabH2z
6q/Q13Ln7kh0f/Fc68Dq330Xi5QnVhN2e1hPIOUL10ikToX1P81eRKi0XWLBCC7yj+6XKhF0bX5C
K+m0d2CDJLmTwxptQtp4rWdc/tTxUoW3i4IeP0V37yDMwFjOO01S1S+o4stp41uOM+rB4g/1HTIQ
WAJ+WgBzVUH/OL2V0YzzApquGLZNKQa8tEgvG+6NekA5mxTQ7rKRAf9yCGZM9llwh470cXN5Rhl3
1C8atCvGsHmDCiFi3QIBIpfXh3NrDifIzd6dBkqnJoVnHn8yoGcE3v+5LMbTykH+MCFngKqeJdwm
hXN+PFQ/wFSx+Hk4AAp/LmWVBonNph7QNusjOcOw4qZEbc5wCTxoPGKG5u6uZPApvmnKujKOXFsy
klIhVa+UufA5cj4CTK6A9uYCckdkVozYW6Q5A1daf3SJwDz931rEXQaVfCCzI2qXaZhiJ0Z8upjt
mlTfhb5Tntjf4paAEMI96yBw6vH4XCTyotYBunly49KaD1EprcaGpDzRHJRW67t/fm9wUj8dU1/s
b3i7yXW+GW0aK9YuvOTBtaj1I+TqkMD64Pw2i1mR3064bkCdGUlIrpRtdjzE/yWZK3AZo4jAjacd
uSR15BiTz2Btm7ReWL/degFlhrj4g9fip+XViqd3BFzHXcBMixQ09u3l0/9/8H7Oi0/AdGfIZdJz
xqaNAT/dGah5rTq2t1CxdhcHtocZ4ALovleWbKaOan21CoelF8iPgxZy/0xgvOyxGlY7I7swc1cI
jY5Mlq5jsoLDlZQW9Roa9e3+IWYqP2QZLxeIYtzBK/kvBdbYCs8ujLWgzcgUsis0ClY3fPivVw8y
fbrvB6t1uPunflG/bZ9NSKCk928vVs0+UejXFHAXBcal3XkR06cYaQOvAXYrKfhPorP4mV+qfh2Q
pWWaY4cGKyIuijXEVhRvw5DR/ZuL9oGc3oE/geEkM+E+Go5HkOI6tMTRm3+X1VGBuM2FpTyczS8c
drwV1SqvgMg7N3I8Y6UhamZiBgakYLHv8wHW7nIQqHvQ8+bUNQZYTTy6/8ytwftC5MZM9FR9577P
Rfysh/Vi0V9N2iHTtl+6r47WU8ls1qZ7FivhEgpLN+PP/vDUjC94ROkCGNLkieYDRwm44WioO4RP
i7z46/VzMqgQUPo1xkRTVcZXAtdpANEqx7urRftDS2kePia/immkFjnBc9bdkkT7xHDcy6yGO0oh
UzpdQ8m5ssF0xh1PdoWMFbMwpMKHG7mW22FcfeMSd++KIwkxHJFe57CqDF1yqLicpZhm+f8ecih2
KLkb+EHvbDpwosM/070qiIYedDtdfpDdvo9rMeJKfQdPS4lk0dRJjgO7UT21388+nXdzhMFF6G1r
UN64+DAtv807WqZeLbRK1UpK187tPo+C5vdwkKD+NsWCSYR8lS2idA4YClV7kwotDzgP0bKrFhBi
o4HBDteHXsAstfLeZ07Al2I91iOMOF0kgZFZog96pEw2rCmxgaJLWI2t95PhzcIUkPvYvY+tk7nJ
rntOcwtRGKepZS1b1IPAu8vDuaySt/fMKJ8U4JYgBieF6fotK+YfVTlFzAsCDnD9RGGGSfUEiglH
r5wY26SbTWFbOztrDq+U4fC9vne0qYGlDRvN6pou/6qyIkEVTOP9seK5dRuPtknOJCyiLj5vojTV
eNecilcDhZ8wJstgcKmUdcLo1uyaVst0mMD0r6jRutRImTgQDEApt1dnMscjDsLO0LgVSIBc/WN4
XCj3PA31t0xo2zFT1Z90ei9xZu9zWuhDvhr51P1+gNGPjvQJ3Mf2kuBH088XxBoqIRH0wuqqxqpL
ytOo24PvN2i11aJSVaG1t0vB8/75o0/ssrqU0g2YMr6vi3JLF5NIT4agwAnp8/eP35NaF+NBLSo2
IKwTW+TC12mhaVitMzTN8cS6ICqXyAj5iQ/oSV2yaSR+iMRjsvCTA0mNG0vxcmOMYCb5bK7VG+hY
nIiL4y14+BeIIFJRsUpw7kvuXDBcdFWxRKAzinfcGyXAZbYPVQXSXUoYNI8msNffHa0DdkPJPz+A
xz/U2923DFJ9vo+gOKVhi+oT64f5X0+11/8ipaEx6Ajq0kVxNsvgZFK+xQdYhIChWEqM6NZOiful
YVGhaj7yFZRyo46uffzQqU3dY0YFeNVZypVZ8ecZjGHUb7v2Aw81QTXReKH4CCMlGyb1w/jODz1f
AlGgyW4YIaUUadlLAfF9DO1FxPIWfWVSukG0Drm+UbMnA2zC1zqi+yShoQqN4dksZhYWKlp6l/o2
BJy6tq0CEsYdEp+y//JKWteuK1hYqslY6ZEcC5WCskdje8bH5K2BMAH+ws6tPoR2kpkJ3dYHjnk1
qQuuCPpt+9/c+14wGJozFuHK9M2OBpDsiOI+0lsOis7YQ5fkp4CwV8VroyaEluqHoMe9/2DYPRjA
GdCTW7zPAoTeBXx4IWiKj/VIxk5/lWtMkTSUzJanEbW4uvTsnvxg90kAtx6e+/0g2hrUbEY/mMNM
6lhrhWOQrXaEnTHfkM0aJEzaKrakhVNgZtRDM9dw8uRB3FW+UCsI9Z/ixgmiEZJxpnTvewOS3ad/
hF+b32r5f64aWgk1q6vCwruLUcOfGprFTM/DJQgof1yZeYcvCeOtuGIU2mb62JwMoRh8MVspUTG3
82Cjqdlp5filLSLfYteW4WrvmTqBsYjpJzpBiiaPu9wFFFnZkn9cBk2B69/YNOsEjJTIi8ooygQ4
EVkX6X32XkqAQv1jCMS2BKvPsKCLQjxIXBhRdWz/1EynLyRRAtqN1c8xK2EvS8O5uuaJ4HkSz+vq
gwTB/flgGxCoCHunMdre8eaayKyArqw6BQNYvBv1wnhqHDaj1uXkqdkWqGgaHDPEM4N35pEpVwQs
wnhL+El14drW2ORUc06Vy6lv0NyEM5tB7wk7YBJL8BJqdprlrr0ySBe3XQ8W4hSKMBCJO1JgNB4j
xTrZCrHK4o6AmhWdZaQNWEpGxv0mjEQUSVk9bYgSBjy3ys7xqFV/gX9tFaLMue82kQm2gRzU3+ha
SFs7PuCGpAmfFaiQDwtNI4Uo19u7mSnzq4vf6LKFdpyoYFBMtrwi7OpFuV8uOOSoIq7pGxjohd52
SaNIvfAyx+aWMIMVloigv229Yqihx4v9D5JRDtTZ4q+BbnQkXmVVw1ynQTV2UG6lmBGWt11pZwDz
K2i9vqGR77LV7CVXIsgM9rXGSM8/nVtx+xmdsRPw5e5xTl7i2M9XYXZMhNSswcstr+oo2qj7HDIs
d6cCiE5PNxcp1YG8QA5w3D3XW39GUxUXtOqbKy1uu2NIlysS1YGnO8NAiXD1yLkWsHbcBG4Lhd9Z
TR7uRPJzEUrcZfvVjqZX9i0fRQcCvdB2LeUE7RQaApaYf9cGP4damH+OXGFvzJzcuqzGa0VWC+8Z
CgJLeuvuY8UN0DCSB/AiEHHIxuyC9XyUsZTd4B+CM+GAIspN35i1vrza0PD2/ukBxb9u+nw6927n
lz5foFFzD60iwytAHCIP7HDJw6tfmMCLqLgRRB8IdNu6+6nnNTv9CTD/NhW9z4zm35HndKbKQ/LX
s3zwttFe+LiUcJJUjAbcXE7tchxLSFVgNeFH8+xeY8RHQkQTqU7fvhJDBHqgLgflN/ufb29X70Uc
m2J9PQ5EC2R1DPlQOoTyRiCp0bpo1hdvW27AHDmJ+aNiJWfWI3XctIuXOdqOVGHGZWSUcq4WBysn
6sc9Y+qDVNp8mMCs/lDD5ZEMep6qserGKq+sRKLnypZ+DJV7gyBA7P/yPNJc/CJMTE99yKwtGonF
cwIzrm7xSb+E4xJjVQIkesjPoCHuMA3oAp44siKyu+2dmo+UoDrAhz7iObp3lziJETQudX5JTTMb
IPfWqEFg93ZTT3dlHwOqsBrUgPM6rlbalKS/gGbMoken1/wvKMjFE2AP2IpA7OZ24ULy+Xli1BML
KWtBNn5TOsLiNpTcJSCoCS2rTXgfxnnMhmofdTSbUWp3SORKwCxJzJeD9P38kjKCn5YU/hW+jz9R
wOLuFCU/tkMlb8OzWwFTdfeBeTIYFu4t3VC0D5Nj6rFKYL0S91WfInWZHcKHli1rvGr0flI7xEaB
2Ary3CWR7dWqwOYMbX7jknnCqLqfNx1s7d2PiLb1tHsO3NMiDv3+NM+YKM6roMTpviIvGZiETJxk
hB8+CdhH438zs2jSJScczpaTxjquRD6xzYI10svYuwcu+9KNwxQvlIvFJVNjuM9rRLqDywtiyeiN
V/jNh+iDFuRiYPockEz/SSi9DUsOF7m3nEn8V1J7rJuDmheZV3ep0C5Ont2Yfp662VjURsVJ+TfY
pAaKcc4tgXo6feH4qQXe5UGFsTG22Xb8xqrC8br8udh/edixjaoxsc6N0z6mck/Nqf/wqrbYKGhe
HDzQYxWeOwdHDcEBeOvWsaRFSubH3gl25vAKjdj7jxRIqHh3kthWEWr3dn+IY6Lbwm1jmn7jVD+A
mh7ExtVrG0A/hhlMhMEDiahSaRJYIb6kT2i6tUl6xPKqY175xRLB094IZwrqVi1uT9rp5WCwJHfP
8b8wbuEFjrMCG7Jss6RENOnt+cfQKvrD4EX5PzpYZZ5gYJeAHHex5LXmszC8ZqX9gllmRnkJUYEq
Z/n8twS0reHfhxeiDZsNDSqR45NN6noHrVLP8Lmc+/cgqiP/ibtFbev06C9S+p5kZmtt1O2UjMZL
Q/aRnzCGHdijGIfW+Uqb/Czm2lQKCqzZSSe3ippaekWVw2pD9DsBDkvlj2NfaeupPLKA0GEUfIyN
wlM428FXKfp9IFbzjqZZPLg7sExDzsFQ8u6PIgvP4ZkuvvvZNnl7lVr8oVX0iXp48nIo2P9YFgkA
O9Kc/I5IiOvk+1XaHe8hsQnUIo/XFwuE6wquNozBAFI5BQ9o75/qbYuM3cmXz7ggp2S3jolqO++N
bY3Av/PJRVJASnvOfe+3imlcKHVzfKRpgLCtiBmA0q8DNalKu7nm8DM6Xt2CCVctS45bVBSzofb6
Ys836ydJcaIb1OIyzOZCbypGZMMzLjN9UPxg+9G1dAb16LYT5QOnDPJqioEO8zvB18CiBfaRmOEL
qzVNsCpoR8jAm2FxbO/nEKYtOKEIiueerT8yncES8xZBopJH/d6PG/6GEUhJXwBrLgwgA03fw6Jh
NN82i3msDLQ1NaOMZ2DVVfUMF2KcBOLBlpDhkDMcMayVrmHZ9v3DUfQREt+4QqoeZ+uFXeMM5xbB
+oEpBTKDa2/18oqkwZ7pGre1+6dzMtGtI+Ppnjhzu4A/w2s0vIILvQr1XXgEWkVbCna3upPHvh6V
mvokUHc+PrI+g7h/qzzEq1VKsSW6DoLxD3P50ELXJ+OY3muaxla3TEHfwgPtNgCKOm5fx23h+78q
gbpQQxMoypgg0lp/Jn3hHmEuVFlwwhNVvA3j7uJLYuoYMVI4dnM/Wf64o305FYP4X01Jp7TtSskv
nZs0AAgUVtSLon5HWUksVayjPCUiAjARXwX6SAUuofRKG4AuN9VKPMLKvz6QI+T0kUsCWBHXjznU
ihKdTQfugANncUcDsRj6YEYhsQQ9zkTqvuc8A4qMWVJGxPFRwMjZW2PvkH6b8qlUzVXstZ/VA+sp
jB48p4MScLD3+riN38RJIwCAv2HaT1zw0s9rLKz327mHt/YocBMsKSvgi3xu6Tn6sWa38oBWG273
pOAOZetl7GEkmZPquVBvhgICVuj3AWqeFJccoN7EzMg9ileMm7+5jWeobaadl8eOfY99xMylfuxc
MPm7YrFBO1Rtd4t98dXHfDtyfN6b2zX/zYDAs3tUcRrGZXqCJUtX/nhXXUrL9wkeKiyYhq8jlttm
XbIyGvcb/lPIanImvOuUuyukAncwgczl6ZITIh3pixsCPyjqZwwSEdZJ/BbHq1OYIEIh6PN2MuZf
JwrlrLwfYczXkyy+qIfR62KtJDqpF20AvM4ts3rhsSDK5MqahDQ+dolBxtQD0T+Gd5zFnplrB9iI
u1wSSj0QkqqJKKXuNTxvl7KFfIfw2fkZQiV/o3Wgjw3C3UGbgoDmcwhz/zpqYkG8H1L+ri1PKcpg
3tAWGgD3jxtNjudQYPvI/eEXKRlM4FxpYAT839y5fdcJm2QGQCNGx6sWVfDaGy218eRhDAwS/y8C
YnGe301RvdVodInT2PrmoYCRPH+FLnasynWnb3YvGs+fcdQdngMQ5eohoPaEStCCN/YjUqZ8jy+D
h6Q9C5yMfN8tC1Ss5rKZe0VygYAJq9Ge4iNHVelF0MeUi6ATNzSpAe+i1vdU3J4WOREGtqTA471u
UUr9sJlF4ABcDGjk1zRu496vvWBFoVPbR23VxpJf7hJqx6YLPmA4weXduG4Bzr4pH6ynFk6xAIIF
zuACZdXX8jdWll60u0zdslqOoRga3sTdvP74gq+JCqg/vWuxWc8cBKmW2Qc/HQ4RroY0Ef5bmo8l
Tgz1/DCcwHruIiRV0p9ZPVUY6CuQCFu6/OgjkTVd3g88VgMJfohyjvPvzoMSjXowgu2LA8XoIcOK
4uz48VmTRB9UVbJQomNmxjo8xhGNSiqvzD+IPOG5oh+6zrE/D4zrdKYRvvPtudWaQr9aancNlX6N
CcGaIeg7B2w3ziHBqckX+Q3H8HwQt+G5lX4wAMRaELHDISKPvYXyqrnpueX4YSicYHN/kvPyy1lM
ozd1DoTeyT0Dv+NA7jm/xvVA685TCMX1aJoJc4++hpXAr/dQJ8Je8aSlP1iX0I1dPFCP3d/kiDCp
Za/3tg0M8ZGh6A3OO+1DPJ5RmDbroqDTv7w3crTMOvlI4RyzqoNZYLthxkRzJEc0HNlOgs10Y9eH
w5Gi5qCHRZ3pYAGwrbqqfqp9pkIvNB63fPieWDLUaBU27JR9VpjeT4xeY4KrbaK370/TE5Zi8Bc4
lXfosHNR7sHukrjjZI/wRubAqkShzpypZe+nDU9hQ9YqT4KCx1PYRn2nAOZo/TbfRS+dmllOtVFs
6ZvmQSDei9asbWHokPE5duKUyUiAU/xfWsx3Iwf6dAxHg102zIF/p+dpl0TGEIFGgbJdIMKrregt
jD8Pij0Of/G8YEXugJo7zoLlNahzfSBRSDhYFYkWVjb+BLnIMR3JGsje5zbUVQG1ForkgZZNYcis
lmST7CCXtOHKSrSsw4Xe+ku1TRg/DeY1bo8ZmQZG+AAwW4pVrdSWn/quBllcZ8WetvyDYNBs24ib
5Hngqmg9wBph+1ahPSgLCofyKq8U3V4IiSymiwo6x9U2DFzyX/fKwJIQUwiWipLhh2F+vdO5W+3O
8UbDxvQ/jqT9oVXHJSY/iBkbYQ9qq5GScYknAuNiNQdwk+PbwN0yKUvTpWzYZkGmtd6lC9dM5HJr
m7jFY0be2o9AH6/B5ljvlBPjEduoxJKjFnVI4dDYPMwcRFfNoRmAT5IS9XlCICQPW/yB/+rEkuuW
qZTs7qn4xMXFImqSg6IPNcboZ31NSl8VBMxp5zpL9XnI+Y2lN3NEgg9VEFKdqzVS/V68mLagCQyu
NDkafQlgUu+kSMfVxY//WDjAk92m0WG3eEo0jQ1t6sMKAYyM3ni7Z/7wWj3ppsn7HxYrtab+X5TH
oJX1cgcyTM6aLLY4eoraDC1Xkfh+PiFEvfxDtuuEM5EmJCrZQhj6Zc2M1eYK5TxUDVmnOZ2+cr8J
N9vtQmBreoTCQcfO2qIk5c3L1wsDgUGy10rg5DUGLsh2gpIoFyvO3xuY45zO+4XvnfxYNmcbg9XF
aPXNpn/qLxpXxicKFYfQ1i+GwejqsgFKUKLAbbymuP4WHUbLxnDtW134R0O69qOozn0yFy5HHZNV
WXZeVXV43Cl0L/4H8vKTYhrvdMQ+nZ9Oc6NDkE97VJ9nyjtAiR93d/sXwWfdy3ln1YZvCg5sw41S
f3ozn8B7vqBBz4CVfiNHme4aoGOd8bFkjT4tYLQaFozhgc4UD5e0HKISzpNjFNBe9hjkV+BsD2B0
Xkh19BSIFq1MPwMuMeeSUihckZJmJku/LWBN+RGv6HyCJpiViORy403JXOBMc2/1xu5NTvWyYE4p
sIsBybkyIbrcZITxR2UEhBGHIajzbdlViW+dgweylyOTnwA2Rv0KpgAVgJogERWUHwCeDZ6WL37q
W8cOtiLmWDVDHzAQBQZYpOinVG2Af7g/pGrvJhXSZF30/r8ZpqOFbU065pfeCnaKZfxs8mtspMuI
btq6savFGMXt/JMaOwEvflnyAY0OeVk070F0shnoA4XsP5DH7PhlfHmisJBmByYQgpoBPOcQYE1x
GiFxa7QYxqkN8AB9d9iYeU4U672dDsBQkfkD8sW6F5Ftl3v9Fv0X/U05fylqzo6RSWNW4SJcg8R/
4PLmg+Y2rsEaWqbP7UNxQxQw0oRqRB+LO39YSpkwbicshu3APC4LfD1FOP/odm+h2OAaOvWSAycs
f+yR6Y8xsbQUmxlZ160fHGHVEcRCMBK6GL5A+jDHfe+xFSbpfboVUYJaf7CcCJ/LfdzW5qJ6NoW+
RUqVaWPzbr90TUdKCWkUyyjQ0qYCsJUXViEktoZKbC3dmo4ydpQuw6EMYejk7ThMv4kuQDEc/Fw5
137X+uskP+SZMQH99Lz+NPhIViGppkorgY6kSSCqLt7J3WZBB5IrHl8CW7qshlvmHchmNp+Hn+k5
cjw5hwuZk+mxDck/kP5q8Y7dJKKNOifKDPNQOpITKX2PRISTc2cUF1lZ+WfPz7/xYal3ZRqyixkd
LdaY90mpKrRPdUHj2XBi0CTtXIxcMu8YPJn7jx4HdhkrQaNiaZQPNST8qiI4xUrWscxihApa5k6n
2L+2maRIwfyTW/5yDmgu23SnU/yaHkoqULfF9x62Cmf53w7BPVFYjwe0Tpd6bmpKahLKV909k0wq
BOxkcgzrNx1yOJpie0BYUIpTBBqJn78yuslD9MNhenSQFYadwHThRi7OTuExlyVh6lqULTCaVmQL
rW3mJ+pRJxlYwDYyJwN1SeOVy5EFpTWRiEJ9etenOVLI3hILCiZfi7wXNwuCeZtcrixKhmZef/kq
xNotyQtca2zSMC21alnm3+N79TTop3PyYnHNa/mRiItsVc4QpN5tEAAV7rzSpCLHCv9RkFh0zqCO
gGGqVlPklDfxXdj1ZORUu3LCfSLvXniEqR56VFhISCtecWLXvbxSE3Uhdq+qVPpP6wZuaEX9NR37
bx27LunSA/mTR78w/7PdEYMvpyKMsOZ9ZjlYOGVDnw0yI7kLPcykAN49XEgL3zst3iTmB+pmJ8lz
3HdVA8UFZmqaboBNhkLXKC8E09bahX7MXSD/UQ/W7lW/Er17QuN7O9PR07P+4U5VdA4AqYL9L6EC
+FuoXJP7FvUD0m8cZTx0k1U3nunvrs2M2Vxtd6dcd/V/rfmfOi9pUhZbR9qOcyUivMhlGG6UMyC4
oUEPR/KAGWpyotBT4nYbIoLd8oq+bjubj1HxCE3do9zY7tg73BOv1PKJ9OHqtPMO/BzF7eWt42sd
l9jfxH5yfjNZatTRPG/D0VXPLabthsjLzP9gskM10jMPfDFqcyNcaqNfsr/tTWyh6gdHCP0/a2y/
rXstiiBQqeojvY5XRfjfxjRqRd/1yJqcBqNi/+m+iPlHUu+6J6uvyPFitfTnCt70kFkQNlj1UMo3
yb7tzIh0TU2F6HyIqvT2yBLMFE47TeuczfUEhPsPBjZnbJzhvImlIWvQKCikijoqufhUJC3Wmryx
vgFDXPCaDuiZxaB56LBZoN0+XJamDOvc8AZG0gpHWAS+QINtCF4Tq/3EHEAn5hDsdbKn05Fm+g6o
MN2KTcEZmW2Zx324YcWKYAvR5s7gWh5itfraiE8b6hDJrJoaotQOLHCkEH1nbLBW/S8P7pJxyn86
UHL5OciTM7+Go3Jjim7PQKN6IyZ+s+Tfzt7Uxo72DSWeh2h6iE4cDXlHR3d9cDg9Z8roAKYIx2Tn
ngiEJTs6cdv4rgxwCqHjV3ZhvYQF2qH+aigCduCalOYpM8Jw/eudYPA3AujF8Xbxd4R1Hne20iIq
Sqq+qEuwLN86lO3is0c3CaF+DhfYDbi4z8Pd7c8KAOJzhyP9ldxQXZ6Ed/Q1826emmh30sAZWTsY
pZVk+D95IHFtXcy/VxSv02JRz+8RBU/5rAx1FeROfad9aNdLgNwtrzRhYvVmkeXSioUN78z6fEQK
w/eb6Q8yYDsLkwtaV4zz4ccG5ATJbwY/mW6pPoMRCZ0oi3Op60VklIGyCzYthvSymbylnQthhw5r
m0wB2G+fNgYPrx2AIHiTY1cigH1lBvh8T0nuNkbdl2y4mtejQKy1QWldA9DDIV/yqtwBz1Zq0aYq
1ZWbL1XSed9tIx+TfJE+72RegsH5tN+HfnTAsmFCvTEySmTbgD2ZKiCjXWXiCgpuIM2FADPJFQ6y
irdWHn5rJ5Zrj3IUmCPT3i0i6WpHN11hf+AQ5pRkqqgPc5BRDnZq8vcqQRmo+3EjTVlLQPEYgc4F
cXVXukpT62Cyq7Qf4AomZL8gsTpzOavBdVbjfIJtJ7jeh6fZkFw06fqi0sodapRLhL3flhqFTbH8
5X8axRzP/nTZ7zVHGii2AxFqJbduApPTGomcTvH0870yYWaEo4S0BZ5dCBpdjZ3gDoVRxdJpbgBi
jpz4Bvm/iBR4PuviHMJ5tYl86ZQ/9rGyJn2395ywU5eR208WxSW5teLo+JeosZbnHFoYjo6lM54u
r6P38rhKQtF3OJ/CT20760xm9Mfz7GCd34xECqCb6Tu1lvIE2v5Mzc58RM2XVXTX+ILhlSVOg6jh
HD4C5Hjj13mHHWwDch9uTBHtSPaK7L/wpwPWSbB1aziFjHlnry1d1MtFFokBQV9FoNm1O7AirdLq
uG4jLrKS0OF6YkKcU5YZTmLmkd12EK2Xx1f0yB9yIu3UFc6XCClmb4ED040Rc5zyNPZHq5hxq6yL
UJzhVjsuZI6Lw3oyrDP8LhPuPLJxjyM2SRi9oBMr2HH4C7/KvgnZZnKFptD8YJXfnumSE2C2oBz0
d+7yZ4OVK3MODIuFoFq5GKWPMlkfIfDiOb/JquHq9B9V6BEAk4TISZWcIz0Vvu1JvpME+CqQ49ga
YyO/5gIdtyiscDo00EI3keZDehHoZUvUZgm9CngL58GkFfps744+6qg/sm3q8nXe8rUTkFt+5ha+
SRMFN5wPaaUziByRYNgIxj6+AXFdsg/nR24Lic5YWIBdZUGXYtLmFq4F28hnkSOEuw3bQ/dwWLVE
TsKlFBTw64JEAqq8XW86P+7gYVMU9Dn1t/SoO+f1zkNwcQxYfR50gvROfXQYvSZ0LnW9oq4ePXqm
EGaA0gO5mbMCH3vQVTJwwBA7fseByJn0ZXnLnsYfqgjudztF0L/JfhOPXrlceNzborXybkATCS4E
VSyBV1/JI5kRYhLT7os00rt4QqvTZnTpZRVmu2PcD5vHFoAJ/Mwp/9aRiJuuO22XXg+bPSnztyJv
qDZXQvjcoUl/k3dGIq+NzWq4G24Rb9I+XPNI9xVnc4uGSpEgaq29BUZNsf1ChIXGnJqopNmDFp6z
7YyGB+isRIXBe6VocBPWI3BBjBm9JT/7Qbg1QWy7npbVkvvlhHjDhD2xfn/HAc5IDYPIHogp1MQW
hLygzluxes+33b8d8oqKaB7LMAufNTLXo59IG5MsGdJdA5Zn0zMEcWnVXzIeKYSzHTVQppDH4UUb
JNk6TqH4YPkxclcU9ZL0RY2JeUeSPFys8rXH6iJPKnRZVwnCBZ5l2LGNSjbnV6ZONW2ksnds0TV7
CDoyYEu5ede+YQuG1jbIdrQwAnNu2Itiz2YQpexXYeIx4PqZWReMMnYGrGpLNUg5Y5DSB21YoF8b
RR3tsoKZ3aElZ41qs8Kvq5mk60wugquK/VWPnoPEG7xnGe7h11rWq+GK/ce0MSDi+29gOjvNtm7I
l5Z0eUh+yGj6VcZ5jZkNouTv6zj7VJ3qGkOd0t/AcGNgUxFvguvKtaBKFxpdLEEdlr+WO6M+t5/E
rAuEOJAwuQlDWAsYnF9aaBOlsDuLB0qw+3Nyb4NL0cvGR6HWzo/aooGg9LoAfjKjZQlvEnsWrqBC
nkrsEW7K4kmH8ENpz3YbBTsCsGntfViMrZvPdi03UB0wDrO/q88wpoqstTSxU7UeN4pNIupaz0wg
j83JSUzZC7w1HPFKOd1jDBTElQaQCf70dQ6WIEzbZuD6U9NrtHyTo2J3RR8kU/arQ/3ppgEla5RF
kseIiPuocNfUBPFfXSWXRjRAFe466vgY18Fq9byd9ChvIJ82gtZvxh/5haQr2bn1T1agQV2EJfBJ
ZCVr12xBXR06OwoApUfu3Rr6iGejbuDTr6jZAX+ToUsEsTequKwTms6XIlikRr8ESWKwUnyFoiTT
aEadC6orA0djjTh0ewJe8H1AsjaFS6QtYoUlG+X0NoAkM/8zqPyzSq7YVYntiIn3jk/pYG93OTuC
AU2aiMKtoLZUYXvVXDbEAb76SSmaBCiL3QurulA7Yuaxo2aTtkBT3Gsc7eFUtfPN4w3YH/xR4F4f
2N+F0ih+YSJU8I7n9qvpc7aNZds79krr+qAegyjJ9OTx4YL023ff9nz4mfEPzw/AafFDbIIXljf2
klRJ1fCEw5fV/iemMNqSxwarFvGGj5J34ccCzd1Wbp2S5ZI9dOWzYz8hTG21vIaV881ApXFyDMaf
+JusatDV+kcOrosHE0oXVYJavEX1A+Tn8NXhOmKz7i0fom0ARYNJ7vnyY/emyYrNCqhWuuIEwQtJ
Aa3NPBIq8fCjReLkcXAogIoHOjUjOvYp1gRzVk26RwkUtotZLB2WvjNeEa8LxKPV74TxdinbE0Sm
rg2DtangSTLNDRuajK5s4a3zKV0TKfGtXbDboGxu8MfFDsmtI+cZbzIPKuWxd5ZCm1kPV2fFgp+z
bHcfwp+2spCd7BEWGpQric/RZkhqFZ4U2AB1UTtmrKxu0rWjhs1UVU7aPlZwlfQyduvpfYfR/2zY
fARe/er7p4xRp5OQX2ro8dxMAZTnzeh9R2k/mSAPc0akZvrgxEDg5898r6yuABfV/YhvyByOw9pb
w5vWfJbPTJNTHwwJ9uT01vWzmcI/Hc64+bleLar7sFJqk6PrUZatuyq8Z/TJDiS5HOlF7ICJlYQv
fu2a2K4bsQag6MNodpfXJj/jadjT3uRmS56Efj3oM92HeUSoNykINefJIpx9sO+38WpQQOCVejGo
mGeQCrX/EHBUDlSXX1QFPHuBHGfiHWcsG0CeZej12kBpuJgel6dFUdM0pTtmz84j2Kv9CJ7ms958
1mmdKovW0i9Y3w8i6CK9vz+DU4N78SmuG31D2WKoVbPiZC5o+8OYGIv2O7BA+6akxPqID+TEGKs+
z9M9cbludkdfgl5pl+sEhmgz0cUqQFpW1Xma+9/iMZAjW/b9X/tHPJ9S0LAMH514IFNA3OQS3gU8
oNJuzmChOZy/+cohsgO5azZk+1Obz79fFPYXV+FQAM5zZdxf3anURgZsLWOf6GRmVfPzqwPiDHrL
2S+bE7vVL8CQBb+lxREsswqc7qO5XT2IukPyKj4oIKyCXal7h+2+YT+VgVdNocMPdPyQwvDPjCbR
vKNrtnzjfzaACqlNUaliAK0/X3XxEXN2NNNou8TbAt4q8VDe+biciNVa3idxYG5I1iE4cZLc33VQ
z0sLrcYPx7QKBaYXSnLiuruiTniaJcmK+Oz9Hf2/fKxeH69F2qOfbd2zZ842XW4oLZZ0vssGZH3e
Id03/BeroEPzEYf55KRPpHaxYY55p4htYQDBOpzO4tBpWyZC3oB5sYovhTpSWx7W9vwzhxdXVVJ5
9ELu+kji0/nHIUQFIWT5ZV6ZnqfqVqIQlnlyCEpm9saj5DmY+KtlLyIsQEWVFDo1fTtnkTjTtCaz
5qXQYAs859uZ+alx5SF8yM0oETA6+2nox6FZToMefxyLBy8w3ddX9B3OyJJg3RA8nDHMLT/EQVNo
iNx5Oq5l/epmc3E03vHU3whf5svjShIQphO/GrmuhvDdptovgu0fS8jf+WP7fsl+oyt7MLIozH9c
OvKuII/Or8OK/CCFJsQ4wXW+eDKskVjDeIZMDzLQuz0NukEzy5R0dCztnoXHbSzCpWnZ02X4eCFG
sLGdpfvxHf1MPcvt34YVyj7TYGc/ONHjNxWPo25PH6xpSkiVFbg5/wDaPWdUOxwRRc7FsghNwqTQ
Rg4ngRUeKgJZN8jCTPmSC/+bW4vx4jr14HRcpdf1Be6yQEQGI9djDA9D4SQ+v01IWr8RGVnJThke
4P4ucXeEWntzcs18tyWVg+V6Uh9M2aE3p7eTrMNo3hya+w4AguhnfkVfDFPgTXmiDBwXGqFMLwWY
Mb0WCGWLEgZ8X4zVy7R9FspdoHZqoMCSOnK4I3MaeebW4q5WLLb4ymRssaCVVe8IxPgeR6cDuw1o
/tRW3MUpQx7h+v19KCKEhswtsevxrMlBRmj2O7ntPHQ3tSkxwmvA7v+gBh9q+xefmWrDAkHUUy2q
ayUGSDFRlS5S0RobQiqVplVGufKMX6G5EOeW03wI6v0SL3fWV2VBYekLNlVFz2cPT4tbNqlf9Z6x
FaKvMTJxY3qZ64Y+wem68QQljJjqDowNYQ6B5FYe+IcVSQUbYtFFq1r2tmhdcBCJZCo7Wc6UQ41m
8wxUu7rdl+jB10A/G5v8Bjda9VkJCeuqnKe6joiWCcs5FPFIj4BSl2IBI8bCLotbmqB982LTszz5
1//p1oCOpDOE80uK+yEfWnegISAl8HgURCrV61MdsA1xjwrfAkcylGSPkcTHSjZUgLEXFgYmMQbJ
cep18oP+3qexdlg7B0S2nX8wdxHskT0vN6dNBRZU8N1wqzN6W88Chsu76p2TFTeoWGKtjuXNruiH
zzbyIUWkKe8H/1x7BU1R4w7X8LlrFeb2OlJoYBwDDEWItiF6X/2ihxPXimhdwVYL23gefJZQJlK1
sWOQ1KKiwBTmd8yH/Ufr0VY3BA+9cd3oXz0rS/S3h+yJqUwBvRh8CdIcqvK2RAzYuc5ZiUBGIUY2
8XnyGbwFs4hSnpFW8kCnH4Z8H8Z5cOcwT54LEVbVPMq9fPHcR7z9xZcT9hKRV3jJaFcyT7MkxD+K
fRcI6hPgpY/ubDh6hmfZ2xFUEwn12tnJ39FRX8yGgI4Uziqv5uXeu5oJm//DmETKoScbiP/HhLv7
+UKgiuAoas8hzc5aYXm4oiGzO5iaK5kRjdqZn81kfSffGYhdN11BpT7GjMxgQ7iD3M13dfRQwa9i
I7lbCGrm2I+V7m2v32oy3Q4/2vng8QW0w/GTHvskeSmI75uMTHo8zvDsYwqkrM5PCiP/uk5Bdq36
Dow/dzjdnct+Dfs3m5QpXfRT3LALCDuwpUgHZsKEh+fvETc8N3K6dARpQnJoUKMxg0VvE3nT5r5A
FSd6DvOYsZVQFQqAaXf6ybrKduB3YOUeLQ7AFQWm2grILNxS3vU8AguipOdzjZEeiOwroO5dtH3T
QH8jBlxLcnN1sxxMLWN/C7xRhrSr8cgBo4ZD2gOyv5tr7xCGy7i+ewKqTYd56o0E17g2RdeqFNeE
5ecZi7G+Y8DSBGNZ9qDt2yZt/0wN/RnuPdptTJT/wkzQC09bR9eOxT4fCKL30/E0TX0PCUJamhrO
vwZWbGR0sbfJg1pdmmTWDIZbo+KorlmtY+8iBj48ifZz+wt6pP+mMUXekvSTUKneF4n+H/mU+BiR
3B9dxFBrDzlf1yE2K8Xv78wzr24ACbz70TE7HZF0zBNDIeCdF2G5X8QJKUrmFeY+9UWTVQc4CIr5
OzEEUzosmS1stC73wrJHwy+DTbxFSL0tjT5Nm6rvIV6nmafAkvcsyqklxVPa0Qffh9tlPl+U+LoP
I7nq4PssM8o5fKsVyROwd+HTj5lHaJHzJ1mw20XdCXiMUj08YxehNyux1CIGC6rMrw3N/tZXGzvD
54WB+WIpqgkbbURlnK5oPWpF50V4wO6LYTlZw6pKWta4t6sp3WDRBWYOCBwHa8S8ODnGT3TaeAHR
Pq0IA86iEcVJJLXJZ1NFsdjRFvQeXbSnJ0HIvTQOlFivnt+v/BCkcvLqffs9ISCRMKSEUsDcGhME
s7y5IZkGYyJVKSg8pWF26fIxRJdYAk44TuyrA9+YWzpoVfuqgf1XGebtiKFRNK00bP9AIGGPyhJg
2jnf1Rk3nna/aL9yMOAaMDI+yh9LJETQOppDVAfUrGgnc5OD5vnuESGIG9hG+0jkKzpVQCtwLgoh
V1smhxpxlyQgrdeB6zBOW8cBd4LalFNjAT4arzoq8ddfA+zwIKAdYaTQDUIEXNtPMU6SXLfz8iKa
Bw9KCu3e65Ae7t5bF+/lRVeKVe18g2dKv0aLyQX8DvdbzBG9kw6XJVP7dboqexGTwBfBZ8fptekj
P0THQGa8N9tXQzldeZZZ2c2bEfDHPngTB4wzMA5kZgmTPXX/jM895fnP8GViMhZcTRyPCb1QVRe6
wj/gs+LHRZS4SU2DExGeuyXtsNZDAjQBQ+wjBNb1LGOXJm3gxAivEQMg3xJQaEXI91CMfrfsuouX
ZcHe1xtz4TKPO0xvRxi/OmYNHM2UKXY6Yz19ULlMQMAy9wnxA+olp0srW54RSO/o8b41BbrlBr1T
M6X1hpZ9k0geHBUAfH8k/8BlzhHh8VRlg3gt55Z4SU4t1AeFNaARcgRPQIYFqIC/H7hx4dOuPLIH
cdz2cYcluS7HlsbPJnBNTKieWXZjKl9zYFQv7l4QcZ6O7fFsa7pix/fNNOkJHZYcs4SW57wwIPuJ
/34CBcJVclrJ/VJcFE1AyjZBI7qqaegNr9wMbzLyaD69VR17FfJNBP6tftb+Vo6+haiNJRjsP7uQ
O5CUlApTMfmsyOzTh5oYJYycIp8QktZPBF8ufZUD3fvTvu87MnVpQRXjPLPM/W1sxQwm20C2jpaW
wb5Y/KReFAGr2blyZ6L/YscV1NgxnpPrF/dlzXicBy4M/YFDIxUXjoSHsLGGmzs4nmcbz/nol534
XOnxBDmprghDqWe1y/BXHLUrSxKFDmoee5UBvW8joUE1FKDDqxustJkg6lt0rZVBwGvWjqdNDghl
u47+lPonYtRZqYf2yzbsYV2LgVMlacBcFbLJ0b8Zio05SDS0ne3dzDYpOuLXk2txCGCrTEnWe5xt
4cneanr0chTzJ/Hbr1LRjlrA8BUnDzg8mBHeH0oIUrrr9AA3CBbAgsvWxwML4Pg2iGndMAB/n28N
key1OrE2+5LNWK2qR9ZiFUNGTQV1D0NgxxB0PK3q0UEwqfDz51XUHd7iJgqDTkEewMIRYVp16IoB
wsU7xz3h9mRR7nD0g9TbDHv+mV0+Pi3f3M+6Q7wnt0h9XM3+cuYxJ4/km0ykluTf+yC1KyhoG7YX
sEFtYEg8OStQQjpOl1rwKxGIrSaGZrr1SzEfjLxGRy4a5uySNWmQ1+4orNuTTU9LGTDKPgmefuZf
FNZitK4ZX9cKHrmy4WGkMFdXlS2PhUKCEOqHogoTqcCHVdEZt9dAzeUbrzpHT1m4BUgmmxbv/O08
yhPCq4UmoEWnFVku5w8Uff5YKpafV9Bgft8/xaeQ+rRuFWle0lUROJWMA9g6mF2C2/s5he1DbjqL
3c36QxuihN3DCGBAK19OuQxewkU3NgTJ67a/fCDtr8I9pEnc1iraTnUKokvm1vdzbi3tsA6iGQvT
4KblAgxW1slmItlMldUuXxScc3w4a+KLVhWlBOS7dl1GcZwkvAbxjApQzHGSUZD+g7JckeUfV9q/
6E43tVjCjFKfRb8imfbsdI6KSrv4YAenOgfmY2gGFSfoYAX0J7LUVpTGZiH8ADPOq1t93yZo/qv0
LC1ZiDSmHWcF1MCGu5RK0ux5nOVF3if9CdySbgUO2QTw2lkc5qyOtUDEpKiAf9ScH82FeRTUCxy8
jX/5Z3WaAD/8hyUG5I5VpY+GtF2pIcDj+ec6QGZpKic3HZoO1yOFMrST8ux7ZB71EF2t4vtkCFSZ
PAbhxarfzTa/TZhovZ5MG3+nj18IA4hViHlbpt5ipxwNTxDYBNLybvaEPg2Gz4bvFdAgJT0ffvkz
I2AhUfd8r3NIxAEgs0aHIzfBG/ZqoMYGWZwK/x3HXTxxnmmn58xReRjdZ+mKbQtzyV7wka30fbPz
1/yQ5tGUzLGBuJNh4gBECcV0prszcJZ59mXY9O9zrTd3Dh7yyfrbKKwseiGHBu+0D+1EoA9sBBkp
yl2I0IdUSDV4CivJWz/3S74cvvdYrJ2jgA2wzd4nfb4xA38v2LRgeNFt6Khbq3ZYCfjEHjlv9bgB
fAhZGyHZz2EDnl2HIGvq2bJ3Bn99lSo8m8XS1gRL2TL82UkUbjFwOG8FA50qDAIWsVWsUpSdHJyn
F7RIGWUftN+Vzbxi2Tknaeu0v3uEHanyPM6cuydAcCxyAz6//3JkmPK0yNJLOf8/bExy/vEh1LCK
rqq5XsvwaWZiM7Yzia0X/xQUJjTsM0A6BIeLwA+a8xOu5lRjgPWQ1KRr1S09W8zuEf+vppywJvVl
19n9ACDu/STZuIf1TLg1gMPNCKDqSLstB8lFuWWIDMOh/WPeulYf9irc9eeCpsFf+kJ5PFAzWn4i
EuK9THEeKiz7Pe+VIuA/B/76nR3Mf2Pu/MpVhm79X/JgZvPa5agspA46Lr/uahhwwev6tM86vn0h
PXEz4J+xtvoEzivZHBlZEo+9fb7zcGTDI1dRwdsviQu1K/0q/x2RRvUeOeTKcfTPtbHWEBP7L/9e
YGZFCF1yUfYMdcX35WpJ343m/Ef5C0d/7spnW/IxWc5jBFkpe/BbvpmaRMG6XfynID8tZqxEYiB8
/O2g1IEph9KLDxZKg575lBleq/N5Tl8V+botKszP8LYNv5P0QPhAInU/iL/clDEb2TYPYSMTYHtH
LNNCHZTNQCtBATUQHaYCFJaU8kIM9VtmqWdbJZtoe4ZnU2ynwa9pUo4PMNb8vBWjOrmwxo9CrPpY
GZjhI1McxlxqPYab/YeWrzmoDdtmFpvA+8BYWin80xJRkXg+yG8SP1+C6oaOPzeCfchMvii1hwmo
VtVfqeVhL++ZoNWwjw6pRI0uSppjbAB/kLXWwGjr/7FfRBvaTHyQZrAXlTWmkM4boXMKv91+T25d
uUx4CXGn8p21AhsGEFcR7Wy0LvR0rXtGCNt0Qcotz7zfOJ8ZNzZIz+9tADnl78c1t8yVyoZm2+wO
Qu6MWtUubJuqk3LFvIapp/9VlGTXmlptdO46m3nu9rh7jqtBZgCLhbajSNQl1sDSrC3w8QL2Sdxu
2J7f5OE4aVX5Qh/x9cHJibzKe0JgiNVjtVLwMcbuldmC9YjvSJHdEMFcwV78stpEi4y7ZbiPYs4h
89Ge79aXJZHCrGwckwLOjdLc2u/S8ydQ7qfJXjqMviecgRnPmYvo8KxZXpe/rZC5dH/zvTxackIW
3eVYsmyszyPdCC83IW6WdYQbz6Z8s1Bk7YxvjmuGfvzqjoE9EH/ptAal9f19hrDy6aRC+1FGdkBC
jBH21GE2CoOsnZx4hPSt3blOt/ykeqj/91Lg7pT28n9nsAak8OowCvzLamJJnE0AJOonRImhmDDe
lkZTXUOnshgmYYwMeDvH5VYma4r3n3bQs1lqL3rgP+vjDeouRg/mpRJGk6WukT4ojykjO02zzfL7
r/T4tIArgnAP2Y0P17cN0ZcLMYUXdzYiIX5b9VPSqCFtTF+YT9MsFjRrsHxw1ORdh62DQEjG6Enf
5JDUyijjD4Z8yHSWip3vEDw3G09HWGyCBRjX/kqtr25LehRIa72C9zfyw5y9cEp+Bhzm41W7vD/o
VUtLehp3s31Nmvxch/hvDwD8Way7ieMdlcJvNb1ij6eTuzRB23rY2ax+Xlqg/2H1yYAGU8pwmV0E
23RpkXFgHLUjbm6W+pHSx0LAKUUB2wbCVFahyXMwvnQV2gs3+e/xdn22cUY8NxKr+ixVm+xADJkA
+nCjdZsyjuYsnw0CaTxQ5pOx0pUQNgCzTUrUZRNy41jay3XD4VfBxsNm4oVOFsFwlz7dVLy+PuP5
YIgaKvadBo3WQTe370BGZ67VsamcGkvQ9+MEJSfEMzpuLtS9U67YSPc1k46I1j5eN10aZqh8JSYz
VgP6zzllAjBUMiudtNvmPyEuYme0tmmbYEZHQzm1VOqI89ILZqcWy99YlosHCWxWRA0YFkzTh9ZX
v8SsjD4Ja0WU3CvFw6on3BQCNjuBvggzzy2kVqtnuYcrR2HuQg4bbBJqgi5/g6+m9JoL3p7Tv+Gf
nPKf+aq1wwyjBRffoQeSqm5+1L4aQQFUXJDR47YvZFuO8+cciEb7aUCUufQP/v1E1v0SPCezRpFb
Ryjiv58w2Gt+v4yEbgbyRlJv/hI3guLcqYx8Ic10OIC7pgas0oB3gKyr0qFfywLpSDB+oD2udGis
5kX6sLkwmjTg85GYp3MH0CjhNK6J4PDgIVIXA/sU2UhZ3flQkWdKSS7Aeg7LPIW4i1rnM6d09WIL
JK9xpfEZp0F+Lu9pWTsCtRXN+je95dG1hFEe7ZO+3RNi3hC7VlffSUGqB46R6rpdHu/U5zTSywOi
DfUuHbXtmYVKduf4bH/EOSAh0xqtUCVi5cqml4ATGsMRYKXQVZY1bXSfpO1yLu7iT4M7hdeIQ//8
RFzQz/ZAJ1DK633xEUv1BNoq1q2ut81ZK2ucBl7b72/jyrMH/Ssym8NhRxuocVB9QVNWU4UBvDZX
PPeuvb8nMx3h95WLxse2wHzOIqRgjnkIqc08ewh1yU0+FPdBm/C42ehd5CsDFx3+KWmtsfAuV83L
QNqSF8jeULFHNxKqZfJnaakRVcTbs9SBofsFJURNlDDKurbuRD/s7Cl3D/MtxlJpgPIE6svIZk8r
3evg3FBh48R3/2RVXQpKn6+uL4jwz+SJGy74Vqy+i5EIS+pyoKNVkX7kATnyRI5PyKkig8GgjwoF
9A3gLLnPgPr2hZdcWfNEoI61pkE8nemGQE545wGXDBot6v03kuests/UToAXY+rxWi3V3Rs1Tocl
y/LxcMSsEf3m454IL/7oTXXw3Wm6UBZRKgJ639kn+AnlzLugXxnh51gZfh2UTIkHv8JpfIpk5CnB
2AOSsSdVNtfqlnIGXx0ZNzhK9VwYhWq00HD04DjC1/DFpHswzbeKnCCDXIQpT/TIPL4FSrGSIG+V
liJH5WBHdq3UdebQY4KY+cJXVZYrhqfDCLxKYUBM11zi96ZfPOBDT8i5H768uhrFiQ75i40sAh7u
aichGESI1mXVqR1c9dG11UZfPRsSkmGc2OKNL7Qc4COnEgVBnzVAyOv4AmKK5Y5Ibv6sRQT90/tT
0774FK4TrGoHDPKi3bQ4wsBRbUDvfcg2NBlasvMoLpQsmLrkoVhdX4AsTzYJXMLsKg+V/iHBO05d
K7mW29YeRhh9YeWqKr8HFl7UFq6Lw4w+TAk961s1DZWQ6hbahmP64MAgTdnZY8lyspbmDzYsfaIU
Td1nRWfK/m7HATzCiJeKHBK98MYMfXp/sGO/4p871lbD1+9YWTr4wlctkmfIygguuYglg+wrDOe0
xTZT6QGe2IqAWfWFxHcc0aBrCC7lDVYT95i1AUD7M0ew9xUO39JTCRqiNYtvZ1KRdtIqAqVfexyL
5zeHiq9WAZl3uIINF8KF3+89RspEv4xlZP1LwkqunD6Q4+YbG2mGr9o+/XU8AzsshymMLh7Ha06J
cAEhcsUvOwVqok9mAyawt6B38QE9eh2dqamRkAol5G64QTcNVXYiVESOpS8BvCIlWGq5kP7eY+PB
FrcUINYpxOZOhO/nKb5RJ/qbwFFRbhl9l8vhFV3Sns3IV8ivG/UQoQ+02MKIXcEgYcVi6ppUbC7G
7NihbqdgwqxQrKWyhcE/IAl5cOaeik+85/XEUAWUvZUTokbmZLh78E1Q3miZEASFjKMi2bI5rUyW
3hDiXRZHlfJYJEJYuxea/r2j1tzvvGQXFNMD6ziTvH7dhEJ6tBurfNxRj+QkrrmTxGmw1bUyWlOI
efPGCkuSqQwYtnGl1xotPNbMnjgsPnuLXVeH7JbJbD74vrHucIqYnsxEXCHZ+qWMsGFyT6e+sM++
B4Ot8S1jeTUIg7xFA4zv8TFeLGwP6XKamcWlQuqjQBWm/ttHnhof6y+FGXnq6nb+LWzWcgD5QC6l
CRVBj+l5cMAuueJcWm3TIx+PygqoJ8CY6Bydlz2KpQm1yOPqggdpCb1ep2RnF6uZ4yAnoIaJvhZ3
VmguZBuiQXP46eSoNZCDPlnByjzJXFewp8H1rVfieba3tGYv8I+sEGUEkmNj9RGqJaolRL9M55ei
CRs79vYGceCPPrgSHObmPDmic45IA5yYV+PZbVEMMt93nPGkW9MSE4cgMdppgh/+oxPzNCKAleal
ZPrNiiycyIVoeiBwidAhJVWmQPKwGPQud83J0AGvazHJSCYCLDP+ntXr4omDl8Y3+4pbZI3eo6Ha
lHZ4aYLq4CzwH72+9nhcHhZtelRi0Q1yYvYWtDSABr7NIdrEyX6GFZgkarDs++5Wg0o1rw0108pD
dVggkMjs/CaGXl2mRHv8yK2KBUm5pbPBj5jDkLf61f0sQDTHUQbq3xadMamzAW6Bho9VlkqlQufg
M4iE+c20BZMX8UmakpFMkIeBcN5EPOlzJyeg1G6azx/Miak22dKOe7MUtZ3Ad7TdCck1QzklW7Sk
OCnmtOoslb/hwxCqDCuQq4aflju3kS2fT1VEgLiuppPt7/6M4Uar4WJ3p1z20uRFFU3wilr2krvl
j5ibXYyhmlHWqflvLYaYT1LxbJzxizNS59FTej2NKE3A4wFXzCvXc7ZyNYZIhj+ZKsy9BAPcLTQD
sHGT3fk45zDmrJqXLvufS5YqU8dMW06UeozgDgae/kk1OTG7kkaWSNxK8sHfrHMpKtHMKWsTUdXh
wDWos/zUnUvIdyYNTkXA34N6XPXqxv7FEWdt5P7JSUyKFjxW6FdnK5Edz59PUBLRL8hVRVcy+tqC
bOFjFov0/XYYbGoOoUeprR6dsa+9BzXKjfB9/P3fhWkxnUoLupoKijNQAmV9EvN23+B1N8lo4f7j
lnV18DcCEdIuD4rpojAlDLICpCVC0dn1giqMS4IYM9nJBoRyqEwpz78FCJBCf225snRp7LiVXWzO
zJl2jUJB/7f0QPsIofkXyf8S01TU7RPi85dhTbw/7dRIF27uUr1cmHpmMws/tRCsfw4o7QhmX1b4
96CaDnSB0Vl7EVJeVG5AZvGUsxonrl+u5t9w00MG3Uo2pfpzHTHWLYoabzAcF/27S0e0ODeKsFQ7
VMbJoBSVj4nvuSVu2Ifjy1ZfIpUeIHddKrGoH0QJGaZPCZtm9h6Q1DaMcqplbG20a8vEPcbMBAFq
1MomXii2/j4yBIa/xJiHCc/lMv0oGZb/LFj4ppkUuVhFEsJincszFbSRlrb3PSHuI6XMOoWc9pnv
I4qYtDN2xlCXiolLUv49VKciiM8/nlY+J4VpQtPGINtmKBZY3JkMHDUpMP1Ds+bFhIR/lfni48pm
sTUmvIIuNBNCQW4duP8iXvw1lgJkOCb0nDxrGzRSIkFtWSxLhRjXVlsxDZZHZDpWg5Zuw47ByfH/
XomXnh+ukbKCf1nO8DLgtlWhgA5dEwEtveUkuHakpFRHB4pQzbTMTyEv/qA78MAObW2YqhB5hipT
OXdK0ppiwX2lOKdnkLU4+rnUhSSyXy4hnTple0kgxvXtpTw6YApfnZDy6EYtU0ETYpSKbXd3fuWp
EVmZWXE8HUkhXRDNMZU0eudNtUW4cgC4SXpkCt/NDRL6Unzd5US1oOnLtRpFRlyPgI3g2IHoHKlO
gmWApaIEHCQ7r1E7DlyUa0Mn9Xwy0fONsSCPZ76586+93x3CM7H810opMs9xtMTzY90FZfo0OUOB
t2kJ5nt0y4z6Hk/uTHaGBmTCbQtq4BnR8hcH4fKShL1VjdTaz1EStEJU2YODA4GqH6tgQXbGv1PK
2zV/0IxikwDLT1x1/HqXElY6wX6fgZtFb7WlzMoXkuUaZkPme916RO0RPseTv1dqUnB4xcgdGV+X
FBl1K8t/nWr1d0DozlEycoSuguY8P2ONW/9QE2vdhGQxeLSJB1glHcFPwASg1cEE3CbXvr/RgwQ2
lKN4/GVNjX3D2HfUqFKgoiZrJPzG6qRQ50Q+MIP7aPkxrTrgMkte1L3gur8IBLB6HMQHQmClvngc
AaTIbiffsSQjtA9cMQhDoT35tz9HXuDtc1HwlAWgVfg/nCQPY21Ms0MjTsa+4wHPO2JOpjumEZ8G
aE7bEx350hGt6rmVh/pHM9+Wyp8IwGgkL/9Mq4hTf1YbUpI3NzYfPs8mGPh6koHRPgC5VX3bo3q7
9kjjQeV/tKowuG8SnWQy0ltPi7KgJuvfZhYw99SH5N/GrPtiSkR2BacJWOehR4cuYwvk+IJeT0u5
vu4rL8q1rHJ/GHU8Bjy0HfJ6uwuXTgS7xRjWoXNKVXEoKtloigQV8LN5ZxSMS+I1ViWJkI94doQN
hyMxhHq41HDtNd2UCMnyICxXsSSZloe0EPLE2XE299sDt7mxC4pDqLPY4F6ugU8FUMcWH6hvh5a7
nN/nWDfg0ldRV1OEncVra8iCfkjiBKj7Uec5/OLgLHPeRuHRz22UAAIjdbCoh43yCM7ODlN1K6tG
gxnmzrownNci8CsCcR4QPrnltX5v36tSQvklTOx2Aylsi/W4nT4qjGTcki6wBqzut9ZVG/oEW6TQ
9YyuTb4BUvtzuaKzc8hlcqVRs9XpNiL1QckgLRz+ijM9diSCs+F6aVQvStrE6AyGvtUNxWAHHqb2
PC4705uMiYr5j2+nTUxRBBkpnueY0Q3WnD9k2cIfuLX9BhD2FDDHrgI/4eLz7OEtEpuboKjkYzka
PjUIdXbUSP9aKpKIVZ5sJlJ/pQ0kmm88CXcW9enHZTZRaXlz5VXrM6jgCz84xPvXX6+AhoZOL1OC
OL9jl2nj0Jpyq+9+reSs/FkvfAh4EdW4bnAy6VOaZQtoh74lfM6HERffSv9N06jbs3sJyT04miKe
FpMyWaAnAhylL+RZY+liUBH/0kEji8kn2IB19LFKU837RHns9h1imiNFXO1jqWAtVkLA5jHejhKb
6MTI4abxurWtfOT7zvafahOV3+pwhdlqq5/JwtTRqpW52fBvabOpo97dLoPAzDq7j888Dld8qMTo
f2fcVvulD94XEOVFsB6rhEGYbuofX8Y8On2N+GLocr1G0vuk8nIUDivRe57KN0ROGZP1TELEq91Y
fVjp9fOCM3Ts3gW9BGGnMUaMDxdspXnAS6yOeZSsGV5mgHQHwi4BorZ2fY1Z+4NngcLFru2VvDUe
gFRXM741DqYyBUCUiMXD8oW26dIPyXHyuKoUoBXIlY4zX896Mumt0RfMa9yOGv/8ucdlRdZZ9Mq6
BKgBIuFwihfhy1xFz8BYv3JAcCge05VEPFKiX02yde9ecgMo00E4rMQMcj3z875+6WdCi+KN6q49
8YN/vAVt9PpQE/lKRjPuqgcByxTP3S6RLYwb9lVhMDyjEl5vUSvyXbefKp+wvf2uElY3vy3tm5Lz
57BAotF9Fe447nTYUPdgTiAyMety8/ExP9m6dmuG1as87lcHUHdolk9TUjDVrq2z/kEf2caXAPV5
iV6ebTmIxO7kaGGy0qihTYgOYiIe6mqnrQbgydMiHoMsGonzvyCaGzKck2U47se20BeW0xpM33xb
eOBALVTcDDyMA9s3NGy00W3D5VYRDCA2MFCtcYeNc2EPY4yByOOIjZBDnfxvkCiP4D+kSLZQfTRP
gkpGp0+ObIb8rIeXUsjia18ytNuvwpei1Jigxa+LaJYTxRlc6rOSd6suhEt1oUHy8k+GwAgJiwKP
q7A4Hra1S5yBZ9et75Qv9tYdPixw46opnLUfAu4/ULbIsFNWx47nbPzsOIUiC2sH3TBxROwSGhkK
tLhqSs2yDBtpeQX/XWb5x+S/Hux6/UWLIb6Vvl+x0+at/p79NavLMnK++iJ/vN7RgN46JOSycYsQ
UoEy9tj1HElJXp/T/HYFjvd8Ni9ib1rV4E/ZbTpv/t+a7JpLGnmHYxjPmGE2muRa0Ick+jc1wJ6A
xbEZazle0whWWl6umeSAQrTbd3phurtkaJOEFevCqosmqvdfVAI0eBX/PeIVm0k2Iotej8PcqNqh
bpTrmJmAlpjmMV9Iww62DWeBcIJq2chE4vPmgvNZL0SCVeEw/2LUiN9p9yUOC8fTjcD8TZlVSWS0
212Lx+HMhesmifDO6yreHyqlgQUNLxpH+2/l4duqLUg1aatdKW9vYRdFmW5FJZ2dkX0bmv1Wimvd
FK8CyNbsFMMZqB/YmlQU42LsXdzAmXfGf126f9OE1mqswqXPoI7ja9V8DkInvHo5xR/86znxpKc7
u8zntZkJysp5P+Hk2pVXBSGC+wN0r5DNj0S2P4XyLuxatAsWjoSuIDIbyD7juttnPaFGq0Oum+J9
En4zqoUjyx9GjO2ecBl/ABzMb3Ac4eJAyIjLmwnKOofXt8zb4BNSnCKpQ/e1gjgip32qBKe2xvJq
wWHugmw2GbsVMvOemFSzZVk46hxfkoKjqRpPztCeblYcbbFa9QLQGb3G7wEr+MEN/FMZ7Fqo9/f5
ieV8zXoeSsL6w/vTHB3MP8EUcKUZZ+3Bhziia4Nw/JXlNczcVhNFKL1NNbRgtPiWrFxmvP4d5Phb
aMMXxQO4w7UHgHojkETyeOvWxvOxUB9fbg4DET6cJOzjLVfBQ1hsacWVLGiXSlfZ67X/YnpTn33C
0gO8ylxgm5zB2L1plKt7ENcC/1xAmEaz090J4pUtHElPHPjC8gvxlQgZyk2cUtAoUrYywkcBJSXS
NTLMCaShPzfXDH3/nh4z+/JONIqHd8P13S3O3GIraRV7CsZswZzg8bmW0rEPdJPsbsBTVP45KpqB
wRNPpxvE0TeshAC7nTghLVMFzIHurVcQ+fwg2lsxQOhtgDUZTt8kDLk937G3FFsAcbtidEFAT6hF
ChfYJxiozZZvwP0n8uRUm3JPmUZQrfFl9Rrv4GiHgq1hOXZEbfH10Tag7213M99te1nIILcUBMYZ
DXHBXXaHCroBlvL1ASNoNdvqfdnUnw88QZOF6CJOUYe/KOFC1V4k7eQrdDVAV4qaT1NczOcrxB5I
Ax3KmgqmYzlK0uHHty8LZwaBIhc62zSdDA3dKhCv9v1AilAvxHvl1FPRqexzTdUTd7c5DOcG0IKq
BRXMB4eh5n3oAt9s76FWG5BKn/za5o4/Nu7q5ulzFwLrkX8xP0UyD29KeeC0AEzgPsH2yom4n8dj
LXeUwHysL5w1lQIGycSJywJ5FFdY1yimDwUhVIUPAACG8JEGcNaw+ixtlOtevEa64jX0yl5l4s8q
OHJAo/iVSrXPg5taGCdX87Jw5RLfqXjGxKV+Fpmt0rBHIRrmpQvIoAvMSKWB6FnGbXwXQtIjkER6
nVuBAuckYBb5GHO3I/EJSHer3/H9u4End1Kilukfp7xyDQ049Rj4qqE3VAPWK/y++sfOcp2qsO4i
doZCOaIvHdVZpfULYhnGwxrpwcApGL7OMzTY3PURJRE7AKqjbR42Rz841VHJWfXDBfj2nWVzhOUL
970xXL/6AtAnH77DQqZVcYeLqvcJ0TENeMGIpR1Q+ON1TjKho45SUxSPTmrYNp8SYEzBxiSDP8mu
9kxCCiOUd9ziYcxzYASYcYzC/vUBWsx2d17mT27e92NJP7NFSYcmTR3D0DUMMqnNiELSsPSbKwgX
keJp8RYG7tZrm+2ux8lva0uWsWLkOBIbFcxwHrVo6RBp4BZGCqsUswPIgL29O4HqGiL/CkReDj7A
IqdmjHSGtpXYeKDvqK4/QtYDHSL3O/cBm3boJ9PaUcAxd1t6CtlSvPG2EK+4b0GSiKu/zdi71w6V
kSHoq1GvbiVMqsCJECnifpIPXD0kXFkP+H0KO8LeIbFAUiVcLMQKl3hbY7m9e+WGlbMCJeC+8FXU
lLFrY0NdyLEqdVaIEddZovQlUqV4eCPevrb2cT81O0Pmo/YUDnsaHIoAJragRrQCP6lYvCk/nm87
fNS/l90EuiO2b4DJ6Rk9Oi38BbxA3axpyPjVn/gO1b7IKsar/OAzwrtSg1vMji6aOjygFvDlTIHP
49SIoSoINu/FQIvkCXc1WxXJbkf71cJ3SjhjnxYgDpksQ3eDBQg4CY09byHq6CE+0X/BvqF2FmIE
lz9KbYU3lcw0OXU6+TonEJSkZ99caTgMh/r/x3Yk9zY7I7G/29+uhh6OS5dSHkLUoDYj13KtcG/r
Q9UYSGxQpKLhq8qGdG0CIsj0KdnAnkBQh4JZElv7k1TK0bdSPFDeWxh5a1QzlMn2FyHmUkrZNlYk
mMhLxmvPm0LX1FiQbgji/KmTyMkquhGg4dGtvLVWIl6fK+OZByKFIeTcNaUZXRJ+d+HwKOovYQEk
LyHTmGHAjZzloHR/lR/4ybOm4LAeMJPMHQSEj9rUUKuDTKI5tMjhwipBB7h9T+QPHoaInwQ+ktp0
jxwmYOabsBgOIZlBCf7dWNLRu/6Q65cuN9hJS4pC9fRTt/8zS+zivXSyrHQq07Gt9GdJUn8vVgUw
VApIoZLIMhGena4WCt8R/nC0AU5tSOs0a+tWm+aUi1XEvxdzZba3MudGhwb4BduqcVcV+WWr4lN+
/YPg1ppBY0WC0x266ABgd02/uBAHnL98CRIybpOPuWCOqUH7wjm2J2/i6BOiUrlQZprJcQFdWPNA
OKRMa1r80SIaLva3Z4tmjA/IQG7Au8DQXZL/Rgm8XEKwPP43Wjtyq5ieQnTOjEXb4pC7pUVN2mq4
sCaJxb4Aerpa9buVnTCfUoDyDEDIOCfw1QIhc2qQH7/Xz1rubBKjBcW3UKpWULo544AxfHMftsGB
GAc9y1ZiM3DqHQg3l5zgH2MlvHtXsPFtEBbFmDvM9f8m8iDshqA3dyOZv+BOSKLhTy0APq71RI87
Uv4PJHzklE+6PExK+04V+oXvidmjEviISVKCYJWB4evEQ7K9CPJzdvvR1Jb5hh8ETn6VrOzgi4dT
0AYdfvu3R2RTSwMi+uq8b/jc4HAjKw0w8pHV/nb9ZfZ1xi3wRNRzNbQcq5ibFXA62qkuBBWiV906
FMUFknoIChxiSF4Ew42h4ZVQGIK02hkunC8Sc2zNqW2fVr2BQa7qcOuiC7J70lqMU59mwi6NxVoh
M2y57zDW9i7ZAOUm+sW5SGHzhno2jlc8ySTqB35u/Gol88b/WWjJPdYS9FRZsADJOGRTZwSOjWs4
77jrf/IJrxToluXQv7G/ef83N2WyCgW+h4IJ3/ZHSrVWUyYz6+TPhJjeNxWRbpuag0G4MfFIgCHj
zpt8O/CHcCZ8TYlJ3HJzOqTYFa95Xd6AYK2AABqbxsDhuu09kaJcRD5Sk66QbV+lDc2kDBqRUEzr
2Jj0nnVSbErndpIGShBKItPkPNwpjBQ0iU/HEMJa/j+p1T8eGzgXzmJ2m+NPYz7W40ZCeYS+FdeO
ssFpZ7oj4eK/DB2oihEagi4SKU9DJklsp6R+g4R4TNxWiyYzKoCzCCasBAS4fZ6ctEI8HgEXgMug
kz/lMXbnPaiVf0IkwxLsoaORvhFP2eYf0wPNVHVRYOfjo52G0n3Vl3KSCGob1hMX2Tsah0WxCjY0
shkQx37KfYCSXDx/ybZepy+RfjZdfI+VENw1PE/qUHd7yA0G0B0/UmCxs0bl4dtdcb8QNbAf4qWC
U0KkfNKQXbdBQJVHYUlaqCkXDOOBqjg0mYsNruP2SRH/b1JpWFy4uhGdLir5JPknRLdly4fCchvm
1M5ovRNuu7um4SslzY84LyTz2QxZK0QfeeFyVpvhEWWBOK2481v6qjWupWwS8u3+3LoU8Fq7hY53
cR6XJwX1jkqPaWkhqO2KA26+Clp15k80vNqwK89bdMjqAEG2YH/gK2Az+kXgo5hBi7ROrYELwWsS
ecxuxOk0jC/HghEGxQ9IZcsCIlpcsgP0pavlzh2dFpGjfb+ID634TdMDm6Uo7VWCf/F9eGkmEe2+
jGQV7ugGKW6RxJOCxL8rgM0vcteNIoC5gotjinBr56DoSw5JwzScSOggS6x2F8ny/VswOITVZ73u
JigCm8NtaQDqAC/bHoM+r7aRzSSZzLJCp8O0OxqsFMMZ/oaLTlSTBEgCw7QUY2yrjR8xue9dAiEz
2YMA5rKYImpeNr6cq4IcpWJUPhCBV/msqFxplIwKfa+Cv/7JQyk5KL6xMIiCnaSPXcenIAtxcGDk
mOHqtc9pEQy0+RPRyAM0/VrAoBB7vXH5wI+w+FrDnzULWQPq2F3eCmidayYlvj6+0+bKxwymqANC
hRzpA1Epyghrz7xSTcpyrbkjtnLSfbofMiFyS0P08EjUiyJEL3ZasRoDrCuanGyRF61lDrasHz96
7/OT7LHNHIZdP5/6eG4zjHQzw7mHuQtAaiXdzfnLVUXJyOj3N9MRMLAUyYLUJJnV7+Q1XtNpSOXB
1oQb0SGHEeP8+kiZwra0YA8d2ua3cz15x4GQydjYvhdSUV0NpPqWF9cATBHsqSAasiccLGuN9Xe6
NLIsSdDcsCHgfXRPVzRB72lvC63jPcJdxmKxpIyOElDLG5ysa5uSaNleeuoIJfFF3boMygiUT4BT
IcfU5xPdzemJPqu8DPormUty07FMfnYIyWaVrcl5/N4wJOsYtfAR2nhGtXZH9ZazIdBBuz98SJ+z
ZqC9k7DzXgQ8EdAJmNgjii4rut27Z/8/nnvQ00IEpHEv6UwR76MEcELp9ivZb9oZVJFvMm9atcRr
TNJstDjVuCs2Z4Qn3BRHqyk3TiMIDwqlC0i4oHHWRJhcrckMQaYWxnDvYIcQx4Bk+L3iFaKSWAZ3
OOBcG0kuBf9Q7IUyDaYonBm1RulNUtvKzFs1g7boIQ0bJTXbQvHUQoIdxjUqaUYMxdUBC2KeJua7
eAZRmPUaI/+o1BUtoFmgTkSYqe3YYOkXlHe3kXC3eGjSDobt6vAv2NR2aISIC8NrY8ktgh2f1lzK
59AZ1YdqBrSoHzIGo6LhfFzVhzjFsUUAemCsZH9aoxTuoqvC+04NgmpcjxCdUNL93ZHvyiJCDGTL
FrGkyytQahcu5J5Rgq7HPfsUYwHZ5RwG9qpqom7mRZSqkPwWZFQd46/Ei7DtzBqKZ+TtzodLW/cM
NJb80B1zvurC8kjT31uef7wMXUG4q/5IzPSiuWYL7NRz75A/dQ+7AO1LbRw83D0iZwYP/926gypw
INajVddDUnANB5d2DtwszLptS5UOWuwUx186g/RFcQCB++26KEXaHunNWxYGEX/XYLevT/TWTGuG
22FK2abnUkNGrqipHZoM9VF3/rCVmh59t+09q52tBEBw1aZGCdRd6+baeSCWMP6sYBiN/7/mlVgj
OcZ/LuWeiZjpMiZchWwtriSMN9V6pN4xrCMzxSbfoizfFWaV7X3p0SholwzFn/WcTCuPrpIvs4uX
IV7FdELtAGDnK6GhUvcYiQ4ePG4GsqnP5BZAY7zVkxi2YOmr3OPuWpybKAZWzl0tCKaMhpPpxttg
/S/bArVNaNRkAUl3bY29+OuzidbAMX+bqWSua8wxqIDrp4Gjca4nPCASw3JRXrzxNBUezQk4fZ5v
rHEjN0QXEFKe2u/X+Vm+YWpgJMS0+Yz0mrnAXrbZa/aKEr68oWdnOjf85Jum5wYDdXxpeHl8HZnY
0NtCduHSsRbFjFD+NRmTWpjhOcQgdyVIXvPLTmY6Nx32j92tiqJ1A5BkjWd31lkhTfynsslgWjdU
10gRA48BUGy4wCqr1bcktqUJ+xng7GMPvI0o96wK7eFD8y6xcb8KJNM3y9/+sq84edxxwe0e2lP5
460JbFZ0h0qXtvva+U1IsqtcNIPC3CHxXnQBCoS5qio4q7R314HZrNoiRJlhMGUjdwNNL9TlRu8n
L+1agPigk/R2O8sYGjmmCS9qTB9V8IDc6HVrazxsqnb4GufF7hVVbfipgLD8lDRvyfvuOibVrPsD
PphQgunfFbtYXa0CtYUE2iYH87BhyKXTNdC5pPemXIBqZT1yNps4fj8kQeuQ36rgX747y7SHQpMj
HpMFofLAVHfNdGRxy0rKigSmcTPKOELobwQrMUhZfUHi7C/vE9fEVgfa01ZP+as0S6wEZskNqonw
iiEFJs/OQMDTWn/SD41hQWX8MTAI+9WdTQHuZlUZXAP8SXviCgR5n7vyMA69qQKTyr59vM85RigU
5xw3UR/A7wF4H9ARyEddWvfDh/Z0X86EgnSHiaQ3qlk0dPK3KaI8wdn2nyzfaCy5QEWf+MWl4rHY
bIe0vXTRthJ5TwhNu7xU3baaOZP5MdkTmT23ZvlFlTZJsNDyVDIwrzJUgBUleMGUSZte1M2qIAwk
ttcrHT+1jm1h/npyI7WQqrPZWUi28mxgNRhhRcHjEmRA1uE/GvRDwvzXdDINmzfi31/hULRhC1pV
1GxGLgULjXHxw9oVkfC0dabfbTDAyQt+UvmNzBFW/6+4TvpNi+YrIG4Cd0R+EDxco3oqwywUAZ0s
zKaHCaOFIHzhyA665HEjaJ9Cmo0Y2iw+jymuhqK6FZMlkLrLYxP8viqQHD0zqrE2CxBqh4Ym7uFL
bmUg5LdWz/iSmyrFlpccsYD/DuIbnuc6yl69D9K6g9tzf9Q467ihZgQUXJrLMssuph1UR195mTiN
dGAEA1FH2jCZ0OQilc/lxUSq1tNMMBvR9DhVhKJK9ealIV8LqnrjY4Iny+rVacjMsqp+cScwYAvI
lNcEiLDrgEoqeNcMDoDthCpgiqwUatspeFtyd/WWRvfxdkG9HyjkoHAZexWZ9Qkc9DBRFwMjLbnD
rVsdepji6ocXB4f6a48/EQ8ehCEb6Skiqo5Qg3e+D70vqsh7N61Ri33W2NBNOn7gR179xOpagjFj
Sa21jtC86eWFlGulLk5tfVIYSOa1AU/f+OapdWFaz6o8QLJScc0voGKyzCfsLz2186qBFvBAmp95
bJjm3HZlr4y27jR8t+vvCzftAqT8+o2GFzYdIFTqOaS6/hoOhDIhtDKjlof1BjWXVOaU+l5waHko
3UpkkE6XrDKPJpSNCeWKTo7Nz1eIRB/7y4AyuTRer56vTdUuSQC5iDjMSlKLI+dkR9BKoBPBePXl
eqWQ4VUAWxBNblFIk9gLbqULjNjwaqTSuvWI5C5b/+eq70qhHDDLYP9yNlkAQrOrVWlo5hAW6xVG
aS7nw+/RiU4KNU4JHBkf6FV9BEciy3675itVCkMOukCcQuzZPH+KMfHLIEfgyv6fBjfcn13H/0GV
/eIWKnlZpvqrvmmhrn2lXedTt+AeGapt0FaQavWvwuUeMHwLN36/85g194l9bzi7BT2EcNNHeaj8
bz1lcAgLZNL0im0jWl3XqvO32/16G2VVrqFCs1u66zWe/OrlaLmh6nLyBbUmqjlOfmRmujpnaijL
nNG1ao+W8IrUREnNJzzCI6/VeMBqMCqG4DUQq0WBUlJ+afmPH27oquGmbgIfgKnbGoqiguhOhTQu
TUHxtb+BEZHFlaMwDSuVoF0MUG3V3i+TkWa8ke4omXPNB8jwkP2yg441ZGxJbjSZaYfmx1dAssgA
ZOojU24SEZLR/8FW1R5sS6nOdQkF4UPBgjbd7knDYC/8LLufigXMKGaIEIVs/FXf+e4/0FhpuF6p
+DeNqKM56Ghjn4ZrPBaKr6JEs3Cbz41yqDpd8OM6cnj0d8Oqor/jCSIdLvMNtZwFa4aU8GX5hMzl
lk3mLAuGHAITXHufVFzkqe86S5N4d2ZDodTDPnCRjxs+Lr5rcBBpx8iiYcvUqt7xPWH/yjMqoGk5
XSxyAXNGn7P0sfVppKyDm5Q9638nEwQNqZ2q9M7nOzZ4BkvhA2ZKjNeXWooSvV56Pg9eq14yKYnz
6dJiMXv1clcsHf/Rj8LdgjaUHlC5llBNqouvWNIcimCX2XdHD2Cc2h5i5k48FlW+7vYdu96CZu9z
He+V/viF9fCJQhy6ux+zgRd1lA9cKxmbH0M3TP8FFqMHiZ2pu7iBiaf9jZCuVaYdbIKYX5ZDWg5R
9cIxw/YqtFwFL8rrTriM+7FrcAZLWhz+H30cwva+dooGHnHf6ddLBFXVsrhL5rzrcbxnasd+rW1a
TyRckNHoixZ4YY9S3GtWiQDqQCzqjqkhgpL9yVlxofeYIMxXBljVlTYyEYRsAV50C0Wh1Oy+fPMw
jr4mrc3wzKYZK+7ZEsuW+q8WvrJeZRnr+ovGUxBFl0gWUNNioNyXHcgRbHEbQTN2dGcGDuyBn2/k
2BGZUUNZzK6CgukWDpNvYHTr5oPeARJg1+bauw9/r0iVhet+ENmJFVE2/jS3D6jlsQZD+BodonI/
2g6r72Y3N8mHIJLXzz64ZiFmMoVOioLsSSWpIgEgeXtPiHi6tKPKj97kUzXY45VLg2a/vD03zH7H
ym0NarPe6sagW3eXpMuPuWVdtREqor1Ot/TTsVreQOJkA7yD/he7Y1NlznbzziMGCX0Rj0ZhL0fw
WVKljYglgaYEn08KYUMPRYPeZEtgqrsoRsZns7zXyPnCRtBAzvCfefQJdxN9XUZDWner75bdHcFq
w+3+7pQ0OMRdx74XI0p8nNTf5AEto+yHI7t9PHtQDyCKtnWhjRpEX5cyYyZXLl1Zn0HF9S1qz4nL
nMGtuuxJDXcsFu5vD2OkVg/ncCKxGaVwugfiElG0lC4Odg24F1UYB8Lc8DYM+9S9Ox1YiyUytjkd
5n944yovKbWWuJBj9Wic91pypU84YaCAz5KuXH5S3BzR2ClFcmkpT3nekBOgkVsdG77mCF8/jNXR
gRTOTiuINaBddApwhk7OOf+DjNiORtzWtpupDVapKsgLdtRmdsHMF2ETTOKKWHp73lLGLjP6im16
684l2YwK2bbGz9oUK+3zzPl5vTPdfBuZJBozEsNi/hPZtKGToG9K4n/rdgyllx38dMu54RPjuKDK
wUxL2QJdZQyCxFBUVr5Ou5vn9YrVzg9hlsZ/k81Z0iHumtJCRzehT2WjPH09q8Rw3oeygKMbUpE4
A/3cfIm3m7abjxEJmdcpQuKcbdTuPVf2B9CeH8GrU+Hry99gqWpw0m/dqsflPNyLEjrmfj2ioLJB
dCRttJ/kLyFLi60Yup6yVLn4K1DIMpzRXQO3jn3v3gzWG0qrYCykrKw4RnPDuuAGefPnsyK0clgo
NJgNnUQTjvSVhgL0Owv4j7E2XUQHAhk4zjAXmfzzORHPrTj/fhl8Le73E2HQu+fsqIuRPLm0N8yf
rz/3vQE3t8Z7NFaZUVuJfM/EA9VW6n31zHwc9WmCGKAa1fxqoMzb8wTsb7rzNUELyGeHsukfYrGw
5WcjSriN6H9zmb8IGUZ5J38RFd/TLpyqMkonyMrMYKhBblqnepc60maGMCrpIleNHiR0c6v7hH5+
9fnnsmQGVhPY6DqwGczbrWCAHjrlNpdY+MrArXlxuPywyRsqq7+Gm2Ez3fRFrKEvSM7fujJ76LV1
XVqgb5LriN4IF3V4xIJROkLWbdc+N1l8wO9yTaTvyXIP3dUqQVng3X937vdZaUM8K6aRH3IaPutQ
NHk4eZPiB3Ol9/dIfCl4mR3XknmVYQlcvi9YOmTqsnG5MWGye/sSSD+MbA3KmZI5a2990j6RiJOc
hrhtzlF9O7cNpznyt4yS7lIorpblGOoTJgN4TFL7R57T3EWlW3HTV/YwWUbQ2gXwqtxfDsZkMCIX
hzxoPZuVBmrfrYjWo31qpLYKjauVndHZqzIdQm5DpqC7mI3//Yqp+4a52SETzi3jWhjL72MC2B3k
WvfpIl8BJlirq0bZiG1rOQyStDgeENi3dAstcxFWtuAnlS6JEviHdxmiaHWvVGNPMuS9e6cCHUzG
zsC6theWFlCV5A2S0V4xAxsa4LLYL5m0nSJ3xb9ueAb/ECQnCO9JhDAAnbylL269xrVw7LnrUUOa
EFLrkTmhSVaPMcqAsf6Z44MT3XWTtRi4ZYOsDPd80VCExZpv4uxGpoPrE0kvPu7Xfz8G+0+CRgQD
9+/ZsrwVMXC9FNSkuqcx5UShIX61ifYICVVmveMVu4fr92LdHGmaYF7jGAekr9/IhEZcrgP7jFUa
A/7pHo1X5WWBgV3kgHXAnY1Uo5vzd5PCYAKOs/kyue0Eqd7UZFiFWLqqa4Ux1XNRYnSJ8qxfwu8E
3NenBvaUhbtRQRgKE4wc6PBcWR8Kws2EKjdykPAHjOxtztdiygc1v2c67KO4p3AYqclPASeaOaqJ
tx9UBtqehPEd+u/SUizAk0VaobymhVhW9G4lH3N0XQleeydZzu5eOhVL4ryoZkxo1b2vRi8BiVVk
KCnefcabKX6CGMbasNUtpRnKMEpjrgTAG3H090NluXdXxCX5gGwpHNQFHTSnKg7l/xTSi1Bur52W
Ni1DUqPodXJaVrKtIcVyVJm1Bnc1UYVnEmMklGyDfeFcZ2TqBLUan69ulKZaWnQJa8UIAV2w8ZsH
p3i7tSIdPJTDp+JN7Jh6EQE7+/NUT1bCQcMYjHkxMLxBf1cUx7gJdQDTNJimqXFmcGuItxBGW4+x
cUxJ98E8bI1EkyBehLCpozO/0EsA2L4ROEB4IRaKxEXq3+lqE/ttRJeFAONM9WDK1V6c4+5mycRt
eQaMoBlRtQjZ1IJAhz9m9sy6kvr9MPYMW7qbFT5NXnHzDRFxPy0FPNFM2tXVKd56iIlERFgVtsD3
zsQoJPvwcrQUG340gVUXySCzWm14hGssOEjfgkgnCyP7Uo+Su0T8CvrJ9/CBKYDIsrMp++MJKhYE
m45j82PWj8mbJ/rXL/9Wwzfze69yQ1q83RfvuxmHjx3Ex8U42vrSv7iDbxWhtBBnGAiGq8Qlq4wy
uMonF5v0C5/a13Nit+9njZ3JBKLbOPO98qd36cCfyVF3W6TdVlMawCyVKa79zyb0m5UaCckEDMbJ
hY/dB0LqmWZdCeCbCz2cyEtKFs7QTtvGWJE7ESlTxATnMKzCv3Ii1rnKpcoYzOVcbtknp/VkjRTG
F1nHz8nbzc2QCDgzDs9oBRgVmhFDGwLn/y88B1OAJuBDglOMMUH1PUDTs6ehmHX+2XvFvDgNFF1D
x0AiyYnAZJbyQ9uGi9WaA8tHVlrGYzhTYEa4Xk9GCISiiWulRj91ZsiEeGCfZw4WMDY0Sk4vqGod
DMq8c7xqSPN/NB319E/ys3rgcifhxzCzSkGDRRw9k9Ich6LmSIuG7UBWnjFZPBP32QqXpA1Zoevp
x/qITE2QfskXlGZg6GSyG3gbKhMescpGC9NShk3/gwq9jsvlizWgslkmtwHU5zLGMf4TIJA9OYjw
9hQn87J2vY67wMwmOaImcN7hRVyqXdBtfEVdUWtdrcu2iEqNPN6gTdoUQF2dqnfuJPFH5WvIgc9L
l9FjlVMr9onYqFX+6QMkrfiUBNY/hXh97UbN87rwVM9PC34ht8epOcH5NxQXH9g03ArGTTtYlJ7S
ORwbSdoOz2jIFtIMAWa1suzI6az0JexygkIrDhH0g3LkavLLmt/ma03PWkbSsBg3IqotIKUP8bbT
awD7RR6XSlm79J581ykgFvbx2ZMg37Oxf779n6GE3ySd7Otw/MSB67aS6sZGk8krUkFzAp+2wwzS
CsGTzZHmYofbs7RCYUXN7/ehKwDnOCY4fQv3K34n89sG10L7DTEQifE9/daJggrn/KDqcxOAic4A
lTfuQFsQIJ7d5pH1NGqWl6Hp5O90U+ABm8PpMpj8vjpFYeaiQaKbLm5GSRjlMftjOgEHfKQByJma
CTxsPR4lKB/O1eERIudz4+XzFwW6Coyun1j1FZGeO+IoI4qhh600nutn0O9nuTtOROKBrjHz2h7o
JEFmYuU8wAFpK0EDvSxa+mwaisXxgBJbP7IOco/arDv/Fk1nQugSG1c0dPsgzmN17pVG3EQY5dq4
sGfuFcjesWNVD7SBF3dZho9KT5ri26Iig65R+B6qNVFasfE3ZEwXD+uhl9nuH1yfND7+FV3pASDh
+gDE9IhwWUtFP6/Nt8K+rw4+E42U3fHIb9DzrpOe6jbTUKkNawrVASO+DOu4tzlm9F64hqXvqvbV
uB4+sR96190ifR585eaJZ/6TragRRd7/HdlGyFBSyonoscFpOk01SyDMjkbKpzaGwDKMoFyuCQV0
iuCIivC8Z1+gr4gmw1bGjMX3PzP1ZPYNAVBhxSjfXgUh9H3Rz36MrxHTIWLAkO0P3H8lKvcHQOSp
J8dHlJX/GPzVwVn/3HI1pWy84K/nToG+9Q0TecmKUuOZslN6YCGLfO3l57YX7hSKHrKAd1tdeoxt
PwdbAaZApnPtra8wd6DV34YEk9bK8visvlWcdbMchSXks28damSPxTHQGyu/uRxEYWb1hYevLhem
9rKcdsYeQyLPmaefMEnye4LQxajIPxwxp/3SU3vzPOuHLmiNbxC4U4UKiShKPU4JBRnzj74yt0zG
ZCLezJnw+b2w+Wap9iGcSN8EUgY1K9qIUT/RFvl0Tgt065rQsXDv+g1Z5jPNMG+DNuky9J3MFals
Hjj5yXAzVrjBhZW7Wr6btc7Ntp43cZRPk/J5rHxpBKbvxdsZNk1AAgh+hsP1Ohn2HyeXUMTfHsZm
mV/ntHI6x4rrzfEXfMQ0mJiP7bJh4fGNqqjMhZD/vPDMIB0nnLp+hHQ7cpse/gm2G7pmRi6WU/5b
srcvpuSTpo+/oibZPBg/iy3mtlaUy5BT5uA5phD4XluNX+aamaSHT1BipHU57t09sii/jJcidE85
pTzszovACm/kACX2hHJPk7NiJpFl0g2noWT14zT0HX61OCjv0/y8p+C2rPY6VU7Kh2epiKeOThVV
kAkYeycFBfGtPF0aVNl+oZBZItFk8aSqL6buUE+3rfoBqFEfoo5KKjl+UqsZH8/YaiVcAHDIvF6W
/Rl6YhGt75KpepZFBSPTw6IVForpEeKa2wA6t90EN1+o9Ol7IohL+q0KBNQJkFouLv5rcJZcPgp5
fJCNE/7Qig9r3injAem7vsUGuImYTJWeXfoQ1LshOCuoniQB7w5IqxJHSj2VBEvINrrtBSs/zhqm
NXKlqEWnB01bOsGQo/+OPxvJPsOevDMw1DYtAA1FXpnZa6qO3wKzcUp+YcVRn/SOfHhr0qZqmMtD
VgrZmzeDssotF1XJ7dq2yJdSKRrcbVNjZMzS9uQAfqrEb/Swp3U9wgU1HosbTOL1bRTROQwnE5Ch
etz3c3B08CTf2ASj+6p+VXtG9YnE0/4RxUa4xQV11JIEiTdO4Ipp7dPNkbUpGzlqZvBn+5zWN69e
8QTxKXZiVEVASakbkJio3JTqsc13ek/fQ1HnCl0VSOdK/NyDNGpZdr+LdGUyCC3o8OAZLILiCSib
ZAKx7u7D9SvWKU9xBuoVR+CnFuU77EuMLGryPcmiGNvng/1eKrJj+62zr3r5EVuLwpyPm8E5z0ZL
7QPcJB1X0jkv5K7NQJpWnvkdtCMP1Sn8S46IJlXVxPHATzzXqZ/AY1RERVFwNTbx/6M6s1oWpgz6
Ywr1uRLDytW3AdoCqXlxEkxBGJKT+7iL8laZfRj+vVRsCc/pndfprAFzes3X/doqc2bSTTr0VDDV
qX3zB+26Ibv0Wn5HY+ZVHZeKwtRteQSf8eTYjyt/IRovCRv03iKyEAhBnKVmqJWS1ErcV6MyB36+
EX48Mq6k+qHG/dYWaPPiS9BJgL/iK5Xsw+HDSL7m0o7uXMEFmxJADOg0glg/Iodqrk0Vhk5NfW2X
1H9epbjnpykmFR6DjPsnkueM+w77HcEaqsvTNRsFZjvEVqBU/joRQFx40fuHDO7OIuGH76Wk/HrL
eiHRM1a5fwJTX8Ofy/6LCE4M0j6PUJytOlItWh5GI3SZoQPcB8gR4rzgFpiPRNyCI5ZrCO95mPkI
RkVMnFbRk0ICwNVq0zSNFtDcqyD6J45IiNxTGePEpClVK6eMaSdm2sw7hLjTTNYV4JMpiKPEGkCk
VzRG5T8+hJao1OSRM/+IWz78+b+2z9BuU1RSq3g1QsWuJwklL3oOHQ9bwuUnV6koB0uV1f92VA9b
OnazLUq9ORqQeR8j23q+hIC/f99VpeSihe6oHJ4zpjevF4aApAPrKBk2Hic29YaP7mO3ygUvjuHq
dgbe7QTjbZ+AIcTqcCYI/mDRZQ6egwWikS2evOm/50vDkVMlkAv+cpHzXeCYCe785ygz8HRdMHWY
m/+hOj+R/LN0ABfF6lFB+d6gJjci7Dv5CGd2dN+LZg10n2AP9qwrIYi7O9PIr9z7hfTXD78RsoYB
R6SCKR3wR7cqR29Cf7szVSH6BHtZTSOyRXXkLq/hY00eZm0Gdx4ERFDQBknHfxQ/5qUxMm6B7RPS
Rf/eCAIxRwYmJigCs45xn9sobQUH4IRbBE/wPzGwARsRjuL1h8IfHNHBHUcdBkSqgZHEru4vkeZT
kdQolG2UfUc1wDsW7TPwaCdLSc6sobHkblkdlNrWKHhxFFvDe3w/nlEG7hgaThXzVqKGgG5HiYKm
chjgrWfStgDo3YxMNuJdrhBviazVMzmRtuvtpNvzWy+aAEIQYtAN3uAEq3k/m4LiiptZaWsThcUJ
6QYjjMLlxx5fQsxwnN11WZVSy/DvOeocDl34TaC/xem6bEBvDFSXYzbVpWn2MdrS2KDAJpuUeRS8
GuM0VRkPpNQQ3UwGB3WdoUPJ8Vvb3QDAp6Yj6idPASTx5mxx0OYtQb/8DpfBiRF+9qw5tRBeMJtJ
JJojs0wXqHXVucLBcSnCLLIicp1VqztlRzn3pRjsTbRdKd9tOYU2cKhcbGK0vogn7F1MJTo7JH6T
OnVNiQzUyqKTWSLB3zaxFVjUwm1tE6ZE7gKX5MlEAFc2ZEoEVIHA058hXGDn08BaeQuSYkGQzzwN
tbXayAmkygBD6BUGG3sMbDfUMA0IyBGKVMAkYwB8mt5plSrao9zjvSUrjZZEMxm00PyxFZU2+F2S
dySe99BHLLcV+S80jD9BfBqVKBkXe4iiPFQbtL1uRNwRAcU6q8AQ6C17b0fElcscQtU8NQpHIzKz
AnDo/9jQb2vUa7RmeP72gYZxXp5u/hPNEza2KI6qXuXtmY0VKgukklNp5y6KlFI9s3ls8dZmqnU2
2HtiEHxoV7kNfus7+QNCPhSTct2r3/i/Fh8BeOGGlGQepl947x1uO/e7DgMJGW/gF4Z7Ja7Vv+vm
69Jp8tM2gphhNJTNPYwaEoBFP+3iJgOuT9rm6k3g7URMsHHxoGHvWVQvH+viltSQtmRV6vDjLA7I
VhTbgziJ2p74vkdTo6iww/l080j0YHiiyaAMLw8RFz0bgshxLleR6VRC/UxmfMFeVvJwr+/qvEQ8
TDIvC9a/boKGTZPEiymOR+DkTB/jX0YioriK8VhJ5fS/w+Cbn0vuF32qVqAEpt85lghOqjI/roJn
ymresZ0o1gsad2u2PQZQJIzC5WAaxfMt8cKuHFu14hVVC9YNqai+XpAzmDgH/6wZMNvK6fZFfAjN
2aAUOmnHl6ISRnXguDEoiyQFkzgHodL0jpgVgf6hFHTyon5t6OxoTvjaUlZNUnTJITJpDhVIhkSq
nuO5/TWcQsVctHlzdocQ9AJJed9FzF5Sz5tDqL5EV8uBez3Ydd8zvmdHERQFg+O0QdQPBd8q4ZT8
Tl5AMyX3a09AiOZqFVu8FiRjcswLKRQ30J8TbtdwmdUAHXHXashgMNZS/2r7x3ZC+0f65OwgB0WS
CZycF7FOCGvajOQyccPywRMIqq4eyUk96IW6iemK4RhjABOpmDqcIUxClTHCoaTDE70qfpCy2qOc
q1dYhwecgBTynFkbSqpTg/n0tP0vRQS2V/bDXwQ1oLAUIszkmPQCXWbJEj5qJfwv95avzCA/T9m1
ozJg09opuZ6zCNdj7No5ehGv924U0WpPithqpt3F5GLnn3/TSpbAfmJNuS9r5Ya+0l9Z50D3Pi11
bPBsIQmtI736dkb6Hx4wZ/5VH8VtKv8mZ/WeOKUNRW8FJedDcEsEf3Rp0fCNTqO4KnB2uKj5R6c6
NIVmGhr6Pwe8JubTcQWfy46tHC79esEVgeTOyoOzyde717GF13lIGrNCXt4bCzd+keIeI9VND7o7
0nvocsqiafASPhdG2aTCqc/gTOTlDdeKXLq2ZnczKpcdQo8NeHUTUi2uS4PCos4KcJ5Al4ZhxHN7
M0h4tjoerRg+TyhPgV3OZS5O0ZDqssgG+/HfyKjI+fmYuAa9pmbsOOLAPoWcy5hGFBOcNq1Hv2zN
5yAKwV2hNZKZIZDVvFWTgJzV/v45kS2ATORyVlCYbv85HQKUYgRaBBC/ipSC5K2bNRi/sU9RftWr
o6P9ctX3QRawR4dZJaetuTFZuac76wwNLQFybpmY8PkJ74PkRsIsMFeC0PIDcANEPUW9JFd76Tp6
KCHMJ1Ov5S3nrJqWiRFzGlhzMe3oqHvwvxR+Gl9Sx/vCDk/HOJLYhwn+2lSs9s4OXh+9FmXidrkb
jsRb4C9XGxSdS4O1keuYVbpozeOsqOqCm4jGXi7MjxwKB2VH2nTT33Ui39cFj5TUr0tdkCAiY+gp
ZIhLrludtmdsx2gQH5TBv4Bsyf51Y/uVFLbn2nM69ezYWGOjEHJ+fH6hjN2arSn3N8J4lFrOSZFY
kKa64nNW++2kXu6MSEDUo1804gghxO8btsCClhF/uNXHL/fDZs09mCQ1hfjQg7TqGJqmajpBI7W+
ZpgHQod27dE1QWqi2lKruiZ9SMInFYrAhwi9dO9eEIT92T1ts2VS1uHwWJOPWdUTyOKO9/zgcTVS
gmbWzpI+dyH6Bu2ejS3prYMNNniFkQNoIc2GuMHVKJxeHYHNtW7qvn+ogaa4Stc9AHhSteW8V6Y7
yLCftsnlJKiEMOj3VBG0OGRq6dksH4z4b21SU2Yc79Pt/yCrW8HEP6NZNxYhd/6cIQ3hKvqwmdYz
OVlCTkEmXQ26DBnkW4kY/wzKcFQWRy4Hc/rvB6XahEe7DPEs5GzwXhR+M6D+60NKEr/Qna0dmo4P
ibBjQbBEx53C2FniQnx8wDCMAF0Lb40cVfDNcEt4ykI7p8qqANWi85llIPi4HSwwff5l27PPop9b
10eiKTOrgo7rHwGu2No1njjfKxPQYKhppBZqLrUXxJ1p63GQVsQqM7O3x2PNChFkvtLUKqN5BH4l
3NUasx92cCr2XVYNdf3AbB0p6oOIceky2qFtDAHOPvpQm2ZYf4//KLvSZBo+wC2SovujUfUOyCF5
ueow7+qjlt3x07JMdnwJkwZR95hF1pzVP2jbic2KN7c7rSj5WSn5M5cvfYUObAAn139yQKjPRrYR
2XFl2Wwj46RMuPa65/Krq/PYkuy9So8igivbem5bjvjYwABLLQmLJMvg4qcjnwt72PYRKC4ir4yZ
aKoC+F3sRAChl/f94nT2jKh6CTY7djLyMJJN2LbfRzOtHEEi8ja4k/0BWpyHXYrRv3ZFlH/Kjlsd
Iarai/ID8w2o6Xvpyr0FG8oytbNOCgKkPn0fmUdl6MPMkgzu81CEJ1BT22a49RK66B58ndXrlLoZ
a4QbwExvDId0liyR9XN/Tgq/r4V6caSAA69s5uXAQAMoekBe4XxtOdzv46k7ADpwOKZAzms1EL1z
lP208/Wp6e3uhfmZya4Ruma7ajQPcgXtXAILHWWNWuqgGaQveuXuwqiDrqp4qoIsPf/1U+EBuP2f
RODr6VWzOLZjPKeEzNviJ6tnmSH4Csn8r9AoQGHmCeqHUJv/95KylqVUWyaG2dmY2dofoGRuawxZ
8sPpxadFlzle+64/SFXbEBPARdpcd51EPkEGanb0Nn/4a4k+Joz2+IOqk9uOand5IPZvvGjDH+gL
ugE7iX4yzO3uD5Hg+cORtiRCIX8pl05I6WIib9jmi+D4aqxwoGw/HGtbiSX45KxWpl8lg/HGhDXY
mMlEGehoUId0jcYFqjh7QYSsYhVmTc0f/QQNX2yul7lFzjqWBHvYIKlp7PB1THij83sCy9geHjiY
pJBGRNDLGFJYznGOuGjw54hw4lmAj3OPaTc8W3yqdrZ8Z/w+WHdD65OsPtG1OQuFJ6ar8vfobqtU
ZtYmU1lY414m8OitLlh6GOXSmmDN4sperdZCM2lfBC7iP+47sHih0ufdvlWmZpvTYB/YOruDKZSE
gTJ6ZV6JN2aYQ22bT6S89dWr/TbdvqmR57u8DUsdu04LQRY5cDxe3ggFo9p+/z1Fz2D7iMB8wC4t
YajI5Qom+Yp293hA8YQKjFtmQB6awQGX8HabwkDNAP4JmFZQTZek7BWw3M8sxe66XK5by/U9jAle
ukgZy0FHp1b4Q5X0bfRe/UsbGC+HpQFEDYaAt/zOZbuc0pEngYnmR5IXqcu7rw4wLE090CS9URoD
laNGvQbz1KUGx1E/y5MjPgKpOjqV+n7QFfq4eelkdIntcHLYX6GjUevBttlGktA3msclBUArCId2
gzzkXrBpFVlnzrgibty2E0cuXAv+NpWz5GXgelJOd9WFluHSMnPw76zuF6LtOV6yG+loFH8UZfGm
/iGZizNadBhBF7p6hIADemhn4E6MlRVwn4p3zRPxFAtR63Jdzlm9KA3I2/IlEf1EamINhlGc9Axz
cZOV3hary8IPUtjBRowRupyy11F2fFdqWhgSO9r2KfCyyC4CbQETjebHaGJhQTBjP4Qz7Vox68gr
E2XlYtQvIJrr1Q/mn3A2h4cebf+u7RsVqLXHUkSKXdtvW3vbteJM93Q4Zs/oa1USvs7QIEqQ6Q/e
SpxMIk1lc2MzF4pdaIDtWhFIFG0bumljwrLA0vNp325wQM6CpOHR+/1cea9gJEJRLweKhIyR58BJ
UIAdiTEMauT7ZcyY1GJI7PHmxthts63Xm6Q+fhiL0CZX3qqu2tY7hLRpmjjOTARjrauosnXZtYUm
qkpACHi9cSJgxCpBHlpUnEYj0dBGApwqKxpY0mu+A9EMO8zZcgMMWCU6opWEPa23jIU1ZjTfwVtG
PFxcWC0IN4FUQnZyI3BRlvmTiDUTRDEnUhXW9f0BHZqESfSAzMI/jcmi4Ov+WZS3NSMy75Usxmrc
JAdZ1C+uqt39EyDT9o1R29qrUrZMXrA24FAcKGIZLd7hDKtgqQ0jj75vLeBWaWTJdm7lldEo80+i
VsgAB214vLbiJCKjIPNV0KroCVs1c82BuEcNZz7dyW3B2PH6y0S7I4tvLgrV2FBq/TinT+5MdTbh
VwOP+ltEnDuUTmEAjvWErjFgyp9BFT69KtrdoWN6rBCbSRlt/wqUaqvF+fU8EMUz0aXeVuVb6Ecl
KXYtX4S3I0BxDdrs2SJuvyBkhY91i9d/djwYMzDkAdQGlGkfvwTz+1+9vO1jIZBZUOua/sQSIEAr
+e3VetakIAHR0qWR8Pl66LULck5+JelmetMgMcA4pzhYGaFJtIPbblOXwjS//Ac8x4r5Pci7sajh
Zfu6vOHKQZpUtGy/fDTlSXWVrJuuR46FgBBQvm1OZuavA4dzyEZGAlfhGkql4xQnkcIipekPwhsq
F3gysqzGxLF8QM1Mp9IMti3BnA7/jKEs9ugSbATQ9Qsm0r/R9TnbGNH0hxp0gxHIGR3rVjQcQiaq
TZIa+HlBepdfNN0WeVvfF4O2BfDzgKvDo07S98GohWmMwQsCR7Csx65qaj01rwVOIiN96s1IzOc3
vP3UXdgCCApPP8LYkDnyTzIuVdffQ7ci5TUvTPtiQeSh7EHByojK33Tgy+isWpX7GBtvC5FCU99i
ioCoe8KJL9VAGKf9V0EnNx4xJ8mmblcQJvODG4J9F394nNecCMDMylBaYhZa9TIjccXDjGqVyDuX
kQrK0VftZ453WcnqUOwEmSldqrLb71QFIoWepTbT4oux7h8SBtH7CSD4/hVdFRbAqvvQpttRIfWY
6NUlU4mjFOaWgVoeWhwbPLdJbS2PuA3MFmOLyEMvo1VirpsgEJqy03iSul6dNn5VL309ymjR6afN
Nfc9U7MwOZkFLG55zMtw835gwgUPAj9G2XyaV+s4tkM+2muzv7/Ugwej0XYYMOFNdU5TdBlhhh58
ZElwkffM6INJAizTwNA5//tI58CnZtHrBK4i7LhBoEy/ewBDK5+e1NG8vOSE+qXUsPn+9RYjG+id
fetzPffYm1yggGKtTj/8l61xf0BVU+ksglknW9F793S0IRcDQlHv8NptgZWMT0s08KGXHIZbbbPh
7/0xkQpzTUNaqwNfxvc9aTvSLTilB5p0njkjO/sQvnmYHY8ZqjhN2+8wZ8KMIbQ04G/YkrMN0UZ3
DFLlTlXkKj/RITesmV0i9tTYkhuF6dNynxTzoVrhvvX5tapvwXiYIXF3KMuXngnNA5QpSGxNGcpW
LQgy7h1PSnL3dpcQm+YUcCdIrYNjqr1EkD3SJixCVxdpggxSdDIKCLE08HF8LW9hWztQEPVzKco9
dLHQL7SWRdBPLaKcEaY19T659Pe5vtENK9e7r7gx/hDWkSC2aQGMadKzuRo3tDtc8y/M9AWTwRlq
3Bzy2/+DMajib04T6JTRSovyrBMnpK7+jCYBH2vMKkpM/uXRNjaqF2Fg64Fphc9Mvd3lVuO8kZe9
GesuTfvsmQIKhJOz8IkjDBjMY25HokwnhgpYNOZaBY0wBxpft3lTbsHBaYDJVF+dRqZ5fAu4OozD
WPxXDUX+HdETaTn/d5JOZ52ipCIhYLlY5H7Mwr+HscN6E3ON05t0Jf92wYV8og3Lmr6CShF3jAvD
GypHjjLI2qTYQXSB6Qeoya5MFuj9z2dSdF2vaHv+r+EhfSKYQR2V0VOfAUVo+7z9c3quf/1VtVZT
5qkrN4EIkJfu2RGizKpWGdUNx+edIcSS22M5QIknbacOlLmkZdX6jhMfEUJceDj0Y2rHvHysJXEO
5EQpomtXtMzKIKn9Tptvhv+PdINHj8cqHo3Mj+INwbQp5Cbk0byBMlqgwq3UMNDH7fk79f0VHNQY
+hSbeW+9HA9FJdLGqn9iTUAzS8uMu7x3ZIGGzdW6bdqQFwD58MZ1SWHBAAu6RVdd+AGcCKZ5VG7J
/N/xva+ERMcil2ORhdBVvz+vfmDYkLSUOp5ptDb551YauxyqFCkunThjXF1BBUE9ipIF6z2y04kU
m5UCnfFVyqpGMJg+BHbQDJKvhWsssmGJbmaQ6TW3UkvOPmb+PMAX4ypLP+hdRvskv5veadAWVvf2
FFeIW+/ZhXYjCmWJFvhxpgFx+3KCDC3cvkOn5aNyn6K1ClYMb/6DbpIftGVZl1DgC4auVAvcQPRf
CE3YNRxghMEeSf4JScDpGS5CfmifIAWXuuQSWgvuxSrlVHd7APsHjiHdQ8dDQoaXmLCPWsJBotER
E3Bbv6HP/Kp9k7c4MFRm53bkYyT55LcQ3xM/sxxn+tCBMC8CUkXyZr2JbKY4F/1kZ+i4QeibZpR0
POXGT8BRDpSmBWB4S6nhG7jEnL/YQT/Wmuv1hqZh4psC9GqpSFYo/LOVFgNWQFKTwtrI69olEiau
WktF+h81482yGAJ51GwKzxWidh2SObeC0uulsN4algUPgreC6MkF57vJpyd04m3+Gv+i6bZ85w4Z
y85X/GT2/PFoyMBcQamM4MgsIGyTFzfrA3jBJpv0q7Z+gW07D9UOPaPAManGzNr2C7jaf8kiy0eG
rp9jcSKfAw4+kVzrQubRXPdQqlj5+YCWOBy8Tfj0N+q1m3u66yWghTbZFCtD6N5POJMplf5p3E20
qeOJt0nMM12EiNYGjxB/IeyhJx/mlc9S8M20zSHGEb0qs3L5JU5NebAK7Ztlku8GoKBuR8I3XZ1h
ddYYE/mJsq+lOuHHdk2AIxUUtFmKrvawIZuWS2XL0cEB6sig3X+p2buWLhF4bb+yf9SvZrgMB3Rh
Q7pfBsRTOklev8bvDsgBtqyGgk+9W9nqehxbIRKi09mfzJb+vx90C8O9BMOt8pwTtOZqpXsJC4LE
44955CNL1PlLf6E5TMQkA/hUhCpT87RlteEVRTvIu2lGVStyxCxuutTaI9l3XZAjnMQkcLL+MBjA
TQWouLeBa9vPQgcCq8S4e6a/pjQH4TSFNTpSD9e3b/PlReTgKoXmkZEMmtGtimEcAW9aP84c2oc/
xfsbgkkCPsVJHhimuI1CiLdTF57e2sgVBAyaJVQasY7xbmV+gxsw+UseyeF5JhKbrQVBoRaexyjN
JlYpT9fe14cOUecXqUmJefl+oFjdzoUNMSAn4nP65D7dlolqqF21sONA2M2du4hqg69dqhAmIvCT
XNjfY/ahhc0x+HzQe1azBGq5b+9RV3JgrEGJp61Q0YerH7Whb7M+KI8XR3+w4VQo9FHPRT/m4F6n
VbTru3Ho7PZVsa6Y5vakDk/LxKaP7eWTLq14c0Q3GIvvAi6Mfg8br2WcEF/Y+0lQdCQY0Y77+yN6
8sS7Ms5PVQTq7IKT+cPz8rYmaZDPhUcDQxgjnR52XCWs2J0tV6l4Ql8M/6xVor0u/MB7CuObd6vt
re2TTAXm8jYfj0m92HHRP666xq85gRvS1D1+s8nAKWqDxcWFE8066YMTB+zAPan62lEuQM3Xmn/a
4BaBALIA+/D8WYBHGTs0DJB2Qf1Pl95+eHQcEU56b6RBzKu3kZzIYzmm/q0igMgOeAVO3bbITrfo
86fHGFH407dY4rXdvTHXzinQPpPBnU8IZDgcuih11tjCeK4X5g7sYhoG32EtgPGugADFKeb6Pres
VwiXNxMtpGNzJcb1aJH3hWNwpQ6/v/qr5T1ocxG/qPOIWNUKA9pkt2JJER6nJf7RSvgaHaa8lsqX
XQxBsrwRyZSssAbozKNMDVpKUKe5WaGvkzAkURbUuZUC7fIMQg/K4Tdj0c4tdiAYWIn9eV6rQDmQ
Nez5Ob3iZ928iZDhKL9ZaPMtlopFT/rXywKlcIYqO4C/QRiohgayJpiaezm0ONfazdx7ZzkHzVPu
bEp/Nho5qA+JHpGM1kTo+KKNOkd0ZvLM4q8Zu8sSJuPEhAN0aVSolA4q/0UDBTwAIoiXnixmReEM
/QYQgO20uYy/jPBBRf13RFfiVqCrqYMuGF/9/fNUHutARh8nE8MIlDS/6T327z0nUQsoh5wZxNE3
6ushvE3CziHzVWMHUuTUz99NbGLIdSokO0s+DqSnSIQJOJLAYGdLFCXtjWgsBf16+Hh2fdcYqbSH
6SY5vZGEg95N70kE1bFePMnzhQ4Rhv69c4CSSbVLmWNkKm3a8y4nZ09F9T2BWZJZm2lAssCy451H
bkS37ZhXdvSpe77amo5acbe229pP7lscXA/X0ISxT4xDgfbTRLHGRsOkJzCXnNM1ZffUPj2PTJ0K
5OaOlCPYkTTrnBHRH+t2RE3LFcoMXZIMfG59Xo20toizKDZONMD1W/v2kEXiQhHUr/Xp9b4T5zLe
6ZLs9L2/d90bUm/7PbrEyJNk+iebTu3ZeYNk1498H/tOJbF2Qt5BlvqrgvTYWSmUlBmYhmPjGizg
ufYjJOUkug3alU77Pk+laQLOICS0wof1GQl1XvdZ3+D7W2p6RePzEktwSvpRHOaHUjN/7GzsVyF3
9X1ftb+IZ/E/K8wMP+RTHKVkHoEn988AEkh6ZiuHElbYl2+DgtZkFiMe0V3dP1xbIZZgsou4rXDB
VsKZqeDH7DCahRxk6WLjQmQtRACJakW/7Ssowcwolh8tbG1V7P5j2Ac75V+eJZGzfxcRc+bA4qOF
4jWQOD502WjSyLzE5LYDIY36uKNy5LjoxnKJ+RMwdxxllVPguz1PwQcy+CWtqy17RbPXVA4Hsb1G
vAe+qpZmYj8loq6b5BFdDAKM7TzgBjY2pNIHyVMBLSQbr/egw4GuRZsiKIsJURj5L19stUp1Vfxm
I6GgqzIa1uG+nXsm5K01uEb+Qv0Sg4uKpBhsWECvWgoe+2qZX5oRVPk4HhjX6tk9sKM1B1uNLx79
l6qoZ9GikGtUuM8EAmg74eFebSGtnITTV+x8FjQnSxD/zjdAvBdEcpNHcq2xkkbBwoPEo1TMvdaG
ECHZFuq6G2OscLVvr+UUWcEi17JAHTlbMvJhmoH3ecVd/CSOOltKw1usOdgRpoyQX+gP+WA0zDfY
abG7pbYXNsx2ro15I8sbYtXsB0RKMxK3VpT5MNshWZtDSN36ygy+FetJYc8r+oCv5lb/S5A59D6A
C5sYOu4hxeqaIjvFnTap9vm051NsWvexNz0huuPvU0V19h2UHtwmpB4ARUxvKe4pzs30lc1cEBdK
0AhwSYaJ3lP7nfrAqV0WZGyMWahGjU7eUjbJtb/4267gd1iYt7syDXkQpK+F19BYYTksPNkv+ftg
peztCyG/F4gun3OO//hZIbSpv7S+DX4BD523o3PyELeMDrnVIoXzZDK4jtZtHO5NwUZ9uPtwdGaZ
yWsOcTb6/xwETNKJMmxyZqMoO1JuJpbnA7F8e7BczkkfVYjY1MIlGF2YNdF17LOVxDhpoh8HoBUw
a9b0o+zwOrTttM0N4BUUIkVFAG+JgxfK/qe2rdWNPn7UdP/bz1tBPkRZc44Tb8HnJeuF8H+keNvA
OqRO9Xc7VOdVh9hwXQN5/PXnF1NLWzfcr3n/CqTm5A0E2pLW2crNjm7Nqxg/ZGZJXaLWqFHhogf5
94bn1BmWUkHkde0+ZEjWf/a9OMJXTglqt+3Lt2ZwIFLLF6T3Y/xpLMlIC0flWkKg3JjY/ZFMow29
ixLV979L72QoCkiQSOMDJ5jUphzkg0KlPgfjYOxJapTuN5ZB2Ca8rFq/0cavYWt26+c471QSkBFy
Kl6575KPPfPm6r0qj9N3kTj8DD4b+x0HobTEKeVDP2rJoRf5n8BKoc+UZH/92ocOFqb3DWZwrfKq
4OgLUlPB+uKsH259Eygw4GO43SRckLiev5LZueMSe0c3Lrb4Zs18NaipPQPKYhb69xBeG2HdpwG+
8B2H5kdk2/x7P+YNHG38pKuBR1KfF5aH6p7yBZKlUioCQn7/B6YMpb/r1lFh++h+47wGtZmlwrMb
Gcz06gWl5WesdjDyARgvI7zeb4uUPeJHJFYoMFwPOvfh+w4s+FcdBX0dHnQMslGM5zTcpPEvJ2rM
KIz96+xuQhK+lJwbdfqJobK549ZP/JGcnVsTHcLefa6qASmuPEU9xhLdA7NlrTDLDbjnBx678kPr
+r2+Q7tV5srx6tUvhqNNVX25o9S/X8EuAC6uNfZSdSIhFj9G71JLFscsS11goZeIHlsqbZI16SNC
AGt6vP0PACo7a+nLbhkS22OCY0Kprh9qXveYBFNbIHo7iXw1vkYAxdqeycDjm6B3wz/FktA8n5VE
NQLeyzS0qjEyShHCwAlIt4b/soQDvuMV/adnTYpz5epZqlzS9U4k+2CXssZo3N6kgcKcaeQuUUFB
1Cfhtuz/TygWWAeIi8X3vMqtPrpmPi71Kmw/H79igYBwZRvvD+iqNl51GQyudTbf1aWcXtQ2AXQc
9Fq4f/jqHwZiVDoeTpcMdAqgTJHWoNfo0ZZ5m+lwyX7VTGmBjc0QAy9pBqnkKd2sYGzB9ndFpaCx
blTpYQFi5ScZ3dzNOTlrfcfcwPo68KfpOUOqfHAISrWZh4UtWNKQHamt/unVSoNSKN/+sDekOyKU
4AGr/gL6n1ob52C6dtMVrN1kY042EA0fnqcVC1prdRliKpgpKSSX6TTzkY+fST3iVXccGHi3ZgUa
h6KrKDeCKixT+DGyUbi3goVlgpz9+lXttZ1izJn9AWyaQkyYqKXC/TXXe9lmee3YQwKLXtbufeZ+
YmLJOKnZ5FVjJcOLrAbEcUeOgzXdxOmTK1z9nBStWlt6qCqQTLzIx9H9ComV9Ozoh0X4KAa8SJ4o
z5QX8Ib91u2PDQ5JuUNMVShPxcWto8tmwYZh6pnGqIZWyvoluYmvEVg9wjxUrCheruZAA9L/rLM3
YKptxbs8ddyog+QsEk7FtYB3gImDJIMuWz4zDCVSg7JtozpiCaQ4xce+QEv+msr1zZqOvioG8vEA
lS6geFBjRldBTYVZN7fv1i/eboCpKijM6vNF07zwtvwldfBpNO5P9CPYoyW9WwNCX8LQuYjJbMxr
ESIC9+mRDZYU1tdqdTOYD7LHWn7TMgK/+nNHXZYAr4URhahHcsHqkGNsZgRQRD0A90n52hgej6Ov
CDk2C1oth9yOmWDYW0X9FUg7G3uBjrDbJdvHj2RUclsLbveK+FYOD6JZjSmU0PPONFrGBmwjpZ8y
MtbDxgdhHzCDn6Z95x4fW7uOPXC6VNeTc13MVjzBzLRHxJVuV2jTKTz4Xnnp8CugjnBhuW3oxvU9
wt7Ptg13YRQ3uS/o/BkZyPHHdPt/y06XoM3dKkLrnDOlDrDmn1VE8e+bILTMCYaVSioIGowF2l7/
6BSIQw5RVlWxl++sFY7Nybakfpm4c5hNIE/cSTmqSPoxDOpMvL7tu0/7EzwgDnQCgV0NqhnFm7sm
rxUD5YGusAKb2PFX64zV4VXQ1cSx1srcxxjwfbwt5HjqqRt/3eNl4QEaCkKBo8+Rw0K/zBav8XYy
SajWM+sciHup/N5OFG5T1b38/xv+3grBq70SFejoCiZY13BT0zsF3qi6dkjUY8wG90jOMX5/I5Xh
Osws/88mvBpLW2bHC6QCmAAdXJ7JYDgv5h9NCNFD9crnSER6K0kwvNCX+5zNu2rarMh8/PCZsoT0
/VYpwSIZG9rPx6Am4yj6INbUtFj0+jlp09YO5ZKC1WhDzjQ19grzZsa8sDRRTFGK+3XJAYCw59a+
xHmm5ui5KMJfUKEI2hw0R8zPbuotIOe99UKgxMaam7tbHfjae4llK9RDEt8eEoNvSmHH9qfzb8EB
eXj5lE+tREsRk8auqy9kxN9DdLEeW7TcVxZLk7vKMhvLZm5cXRtZjAMLtgrbWvEKDhPZ8eEztHbq
XtmgU5LPvi58jrn6SN6EYLPI2eQdjHqxlZCPhQCpfHzNTX8n+TfdGOYf4p1SSKVpM+g/BQnmpyyE
wqqImDnl1gtz1qHHIncGHi0RuEVMJ40Jrqx2gM/N96FP0nqGe3nsuJP9Vgq6m1vBJj8YXpexhO9I
GyD7KXA0mJVBsoNcohD6R0Z5RUDVjL7xYKUyoSbrszv9lEipZ46XOVpBtorJPnfxjJgbHV9l12KT
gTxMFucypJk+N0+DJAreyNvA5J5prI1oXqFK2i/t/ifWcPiZv/tNHAmOALbpepCCXGc4yEH4U2dd
2fgnZi1cRVgUTA6Pu0ivKhwIJtOgwUH7yFRlXk9brquRpxffFXg5G0RxhdmJw6eiX54Y9DotJUOt
WGTuH9525WmVOSq2QVJO0xsGjM0LA0qhurM2sPvmzEGMdQ6VzEyQrCG6BzkvMl+tFPoam5Jhw525
V1PLtzlzcE5e6DKgD1FFxLewVyqEf6lP+3avCCxQrNMPdTQuBJgBsZ1yk/ia5GTc/APvdOnxMrJG
fz4vKvFQ38QBI39MXkyegOkc5v6fbRT0njKxZnC1Zvt0YMoUPdkRkgXLbfDm5gXirnriZauDtVkY
d9XHXLjdV23Pch53S0k7iIkjZWxBJ+hcjetaDJC7YPmnERURNgx1Rfs/yVIvxM/BDt/7E8jElWiO
zVS3C3J6iPkI6XC3aiESnocr/rWv2y3By5gij+Us5vRZNklf8JKRrdoe36Hp4DWXscgREgDxIGPJ
EOdADimSHXks7WxuJs9Zp/r+Z4wv976JJUdJNr8sZfI9t7LLoqOD40vPO2r2krRRHR/yh8oI5vxn
SymrD65JUdarH6z6L3UXpGdIzMtB/kT286x9/btGVOVrTf2+sxlPr+RIowPcqUVlFqiKIQtORWEu
ep5ptg6sdHmnXtmQF1Pd56KrvX96xUYigmGd10kztGsIPZwvhrjkJiSBauqM4p8wgRbWVphWGabf
6NjBFQK7hwnEiZCR/fRJCZCHNmNyfBKFppx7tt4PIO67bl+ONqHaRvCKUwg9CGOAxgLKqXxBpXYD
lVJu8eVnCS9cUKhmFlobhEUg0W3dFkPu6m7RVY0jlAiVYiiu0mCGfwZnuLFt9CA0rSygyKl2wYof
1SkVTwTeTqGusg+1rZX8fCjT3Zjd5W6DvZJQtcAGKsnB8AZIMyTf4vXoYMYOe2diLi9Ts7lrMbr3
Pbol/HdB46+5rBfozVRjyzVrBBGStpXeUSSa7WeCvTQEcm5mywe8O9pp1xM98YHN3T5+kKq00E7+
UEBbmeqh0yzaBjGZE5PVi1HeNxMpWvmM9lLFoHDdbwHi/u5sIDprWPjMwIxIhVOKN/ZTMwSujtLw
TWvIx4aOGJz8j5Nt4XXePGEn8kXit0zHyf7DHS5gteJmWtNhlU8wOW8epJq5PCC4PbOWTM+VSm4w
RqTBpa9arWj1xs/cxWLHTPM4EPWHdHiD/VJ3DGji68Dcw1+SNz+P3WuogQ4nStT1vhFupZ9IzOjE
u3l7t9mgeYguSqIhQZgo4zFxwoJix2LRS1TLAzMOioyOhWuE4NRaCF5vU6gIJRQAsiXJrK/YFV1D
iaDFeAlXvTsLBA3STiEOImdw+0pifO1Rmb20OTAG8jAG+nnff932YPmcp4clI4PgaK1wbl8qCYNB
t53w/2jJuTj300OPiV5hFRMCcnGT8qEixK8+O/tVj13zk4Ht0zKzt7QWEczS5CAA9PaS8QZU3mF+
Wus14VHBR1dnfo1d6DrDajgTU1uF+GuIm/yHhqDJNO7ah5BcRSDe4xbjfk5Y8yo3+ZazG4BnWcNc
0stFithMMcTxjS1FO/GnzORv7o1hHz8RIxIrVMdmrUEUepPjDLis6U/fai/jh8yA3/qN4HfI5ocv
1EtLkQ0utNKEztTsJtt6zW6xu6Oh0kcrieZUGq4tpw/K1LKyOPF5KOQIIqKr9UQcjzSz9CYLQAbs
aBtXZcJt6nWkTkrAFp1ISFh36rKX8N5mVOKX1Ct/BMV5+80kXiu66PRj2oJN76qzryRHqh+s44TF
GddRSLxCfr5L8HJCR0DpdoRDDLlT4r/SU3LS9t0KZ16zO7rWZT+h80tcd8LOPBF9tAyp8auFrsW0
gTNzBWan0C8QZRjQOJO9J9JUCJrjs8idObyVfWtHO2mwZnCMmsDYWr64K9dUVN2O1X4Mdrnua3K3
VFAO6I4E2E1r57vwkL7csg2T67KWNxTHpU16f6DEau3bd85d8YupjkP5fsnXS92JQoKOk258v52l
0KYHyfE9O0Neq8dqXgDLzl7SbRItwR8MOLunC2OeroK05I6xR59xOGT3CPVUbwcmyL8KPdxVt+1/
KRoFuY/Nlo2fixXEDcR4gdP+8vaxM8gWGvaSFlFzOEkUKpY2w/gdU1I/lR8rGO0s2OGBq14q2vUi
WF6qw35mieKEJtj32kK2jfB88ULZWGPxGARNWvD9cpGkEols2j5cFOvNy8DIYF36Snbo52J2aOmS
8RqmcLignwq/NW6aL8Ct1gfXIctO/GIxc5jCVNA5mI/mbi8B4g2SiXJAZdSPhcxfrGJgnDKhL9s7
3E7wH9KT0FAHMp2i8yF2EuiIFyqLwHQNAGztHNvtlGLlPz7oIet6Oi3lBgC00RvyC4CdpdPz9ui/
KKHqlap4J6AUToYp8jKBGzxRdktIy2zDOE3pLblV34CZeJKUy1XbEBTaK6UBP2Zmbw6wpHlvWSS3
n3ucOVqG1mCFztfNWebOeIXltzEZq65fLHNQbUiiYGb+dSfSn35l4ZRQUuYyRhPiJeQwaThoB/0v
BnDVE1Hh0f2DmSvULqPiBjRk6h8mjYOQratAuQ24w9CiP7FUPxMi7xTs/XOPMZ44+W105yif2caJ
6ltzBlrb2ZBGVhwFIcISIyZ5ewtE/a8RQo6sJ8Ijgm5+fempCIuAn+1P+MqSA2TKdLzPChUCd8Dy
RbEBhnCJp6KgEBKNMpigWYU4/oqlWJhRm2DjdXEmeMyrX4LdVCvZ/hDfb6dXKcqh507OhkSEpcAp
gz5w4O/l9kCr20Cg5mD+KCCoUtWIHaW4GJ1R/2NVp9E90xophsPY0O/VqzxdbAEwu0iayzDQ5Kg9
z6IEqv6+r+cUoQYWkvw9ka1BrlkndLMM6BIUU7VJ3GlFLclrK0dPhfbrPVHkuPZ1IachAOk1T/ad
XSwcFjS2SI6jaDN+afUftkJDelxGM3K/49MBVsKqg5S5aT6FZvlBTlOT4MPRSJUH1rI+g9ELuMuR
xt+NY2CTs64Yxvs4sqV1gGgq2iwiUiENzRHSVeJSPv2fRDhuhHcW3gpOgvSAuoXPCMAad6cXRYz3
3VwEHTYUO6TeOixJ3ZgA6huDR2XgudiWoXDG0I8y9WPLwhCS2kUdzcHB0+USY3s/l37yB2OKvg1L
L9DXU//CkIe36k1us6Ltw33Lb5wFt57A6j8u3ypWR9v8AS+loSTH19IUOVfSROnSJVveA0oiELF5
EJ7XydXbYMu0/U+wYrb6EAdSZhEM5YlvgwZk0NlHF201PdJuh0UJ8Y7ihgwoDFZJ0CE9Sff8mpuB
3Bv5AN5uTjOjtF8iHfrtpGH2WYHhH7Z+AODK66/mo2lql7srrfBG4yiJ1YsyHXnElZsqp3lcK8DI
KY1xs81DueQmSpmarfgETLdNkTuGbSL2zZzGN1t1pgLoLN2S4cEmqAVMn6vAxq4nGoAVk92/e+N/
oJiz/C8fVLFtOt3AaLxrEh8O3wRDAMmvV87fVrPKeQo2M+QwXbQsE/tnnFGgYSIatdfeVtH8kTeJ
8TAodUJ9Xd0XAtbV2sx9dXWNoWwRD7r2wxQKa7yKgQj8VJyBkwsmmwrTRczXLpvz8WlV4fNWxpgy
c5RRDah+Solo+Ms6/Iu8+TrpEFIXW94BQz0iEog28n3Bsao/vCLzTdYugktjdntCAcdPUOnwPXYP
hEhaxAYByibeI/DJDcMPIakaf/9S80PEZVFfobsoRfia+Tlb8mFZEwE4SC72KcoEGrdwAM9DAN5z
r+sRApNYr3uBvZJMEQHCQ2KXySCTDqBD6k0wknoRqf93sud2p6VivCIsAKexy3E6Q8ljC99yNCNC
fMFScP2a/TUn9BX3ECeM/v0xCxFPQ1UudbpUO/LKoSFCHAmHfqGkEHxbbsDKuqFIGFQgrTMYK+/v
pKIgoEymLtSoJV3kVYYqb+jIY5LonL3cLwCh2j9UoqIgSYllcCiD+OTlIIjbkRad8xD96Ff19zJ0
K0GSb3xrx+qom2XS8Y4WSomz01qLF2QNl33P5YWyHDBlZoRo+svGILw7nEh0uy/KJtmwXR2eB8Ix
1f0At8MrMQV44etmq9q6hr+c6iltYkIjGRYXl5O5O2V8C6Yhf90IO2FEPStEyH9vCX7FqD9yXRby
bS4dOVJX7dcrnDdUEjnLpbPDlmGR7063SeiP5e/o5sQUj7vExku9IGRNaJh+MXxE0FpQQHH8xvOZ
piASq477F99zlD5OYtx1iETonW0kF0eeprvCYZPRUc7Qym78x0t8ju/MKOKKkqlI3Qy2jldj3clV
uzzmE3NJBj0wbznJDpBFMAPgTslPCO9GmvcHKEj56im+XjzlY/bpNtlTSdrzy/f0ayUpZL7zfsL6
EUcdTs//M9o+c4vS4T1vh/+Q9s2YZGATa5a0Q6c4/95WFPLi1Hf/x7wS1MOdTc8kSq/8COTL8ANM
Y3aTw2FN7i1DRK+uCv5mTC50lyyUFbvjKMliQheUAXzgY4t+M71Os+SSuAlfsHEjvp7pSMAaQnjE
c2vwgir+Thqr/OjbcU5xQH9ptVDG9frClfo9NgJfpMnULL1IMF0IGk0wRBvoi/sQnytVH6KjyRTG
vH/1A7Pq+FWaS+Ww5mhbK+3rAsWY9mNqybl9zQ3s5BWMQYF8dhyoUhfyKjrbkuXaL/KOu8LHyFmE
XXr4y1ZMyydENEZoAntnWBD0baVwDjjZETQcFvmJ//gHxyFuQkiZu2fzTQqct4UDa5oDGxXzGPgP
ibJc8COx02TfaqJ37p0ga0A9ucoOMUoOIn5HWwZfABnNNG5rCXUZhypve06ynK392PY5duiwU3x4
NR704oxlnvlDWG5c+cy9JbS48WS9MgTXY0wVN0taqI8oxQYanGoKUwCigTmqTwJXoDW+5O4LmgLz
1g8pTwmKpAMj7ToRugJLgr+7nxHY3LJQYpOW1kHUP2M5xZBzbmbKziuYlGa/Fzl7THAF4GAG838l
qcT6Tw8Q33T1MDRSiY2s9U0e17n9PHho4fZ3juhBKWWxlIgwilwob6cInrPx2dM/P3k0a0ujRUIz
27L8Omx95IpXC1ovft13gKgQkjLdgFs6jjx3IKCUPThYTeonKwUXzQOSQIV/f9ZSCn5GkyQKt7LR
7yDafFLEaE9/U6y5OEqTfCQcLuAL6+1JRhAxs90UZjRYTMADnYE85mn3XApwXNoddMvOmQ+yWp4y
qKfyzAp+WYx1HpNNQV38a+UMoHjD1J6Ytq0JwSAfofnFdcZ8aK7S5CNiw5LBAiyrUVLkoh/Cvo/c
OxfH1yP1pDXQi0XrqacLDCZ7aGQJpH7oaSR4w63mzoL9F4CY3rcH6slpiuyRPetw/7oxM8ENP77l
8hc7aqmUMqzzAoLJQBy3EELbCrLtPEIQk6lHadJEXgnTtIqSGRW5nLXYPC7JTbiEN+1EA5tOypUJ
D62Z7Bz5WfcAW4Xa0SqtJxQARIe4QVlhb27ePRhbTJISZ7oujFUL3hIDalhxaTugDy8E5Gi1tg9H
86vJZ403qkcN9PQtjxDWLxIcaB/LqwH+dOSiqaaBLU0vaFBnaCHaN8rhWxJijgTZgEgsl6GzhEIR
qSJfgHRUNndQsosZRLsdq/MqHsC9nqQhGq1IadpB8Qc/233VrLyyTNLZpHgnTUGI0Kp4sAr9m8gL
qAQpEVURc2M4lIogrkwTWsJarV1KPng0PxpjTTjHy4+Yk2hU9hl+adgIygIoGNOybhK8msSbvw8E
cvEIwEWzLm6edcgtTVeaeoI77VxLa4dhNxv9MvEonDLpZsEn4S+hjlcnFy7kgFJRySWcU9t2BFAd
rirlDyUhiIcnI9x6aPN7+DwQ9+JngHoz4qHBvBx86ttg0zbt2WhW4gDLYUkmXUcTKnTULkVjKZzZ
lk6dDs21sokQHjmWL6eecqpGBgU8jBNcfo8qA1psqE3SWK5tXr1LfL2UmqIR7ZGg82hxFZVfio2A
IIQOVE7EpZqnzvA5kFF3GpKpruf8rHT8nY8r0eATy9TVdLIoiWKIdnqC/3wI/ojE1E5IH1ZuioX/
ZLmPcdL11sgHp/5BRKoqUNiYDdUbDbkkkRfkBs2ud1L/nIPb+kfCtnwVRTv6VV5dUS9pq6PypdPJ
A2eqfR81fVlkfRH7ipq+ZWyul0mWLZuf0ggtnlNAd0OqM6OxgI9vueYpXrsSGaiKCH2oWkHnjjKx
0/Fc1C1KQuCB9Qd98LTjSTDox2y5x4B3CqjBRGmBu/PcI1gpbWSWwQBkkFa4yD0XzwUAdH2dtFxO
bBX/iG8gERiSEl+p/p+TEJQOMLn6Eox43H0zBOopR7Fw/dC7iJuuWXAr+Xa/HaxJUOtrIpKNCgKL
7VZCAz9y8pXoM/BxRzZuJUgY7wvO8fGDMj0pKlRGI3fotTKNW3nSQ3i9pQUrQ+e4CJ+NqSBHclmo
OKTUxTP2I+KmV84mEQ56UnYDFVfWgP/vx7PyZcDvVfy29X6NjPAPyN7uJzf1fGhTRU4dm1t7rJW9
gdzbTmfLMD/xycZSFv7NWRwhg4RYpp9oJfG2IvGSloI4qx4gz6QaoRfatZSdM+Cmq+zed4I7L4Pp
jIYwsULNmNKDTN/1VBDpCI/Hp3snBipRk8c4YVbpY9bMVCofkjcopuYKkaCAxNfrSz5VOBnsHjk2
j//j2r06qddh+TVV50qzSlUOLwkL52Gau40hfZSw3qLBA9p8kR63FL8QVtAv7ma7v0fFU4cPcED9
g7lb4XoZn5nrEXS0CJicKHHKG9Tc+l8eZ1TQKgJMfdbNjTvnT3R6GvXr2Jze10J1BlEMm1Ter2mb
9zAU8+8M+9GfEcBWLpugAu6LldSojDfEv4k0dypTITC3wrRihtRUvlsjV+Q0VDKTHKHOMPEVOrdt
nCZDJknEHYtl9TA3mk73bWmPBGnwMB/eE6jbGucnDYM0nmAIfxjZxDelHO1RmNwdXbGTP7g1iscA
YMzGZOn85JeRaxL4XGFlwaHOkn8pvTGx6o7vB7gqKK+IVZt9knqeVE3vATSdGdDMqc99iRxaGjwz
ADfgF8TqKg8h7IolloNYREX0XUyjQFF0xOF9duHzb1CcXaR8RQHrMwtiOhHQWWLvEuyJv2BbdL0p
aQjBv/wvptK9/+ZFQ9oNlyNF9jeV5nerUJTUeZsMRZ5iplrnGdEMtLpCs51pWBTLtdJzNNqzcCkN
vLLZAGMYWxIgohIt3434Iqtk4zIBsrP7rn27SIlotu3O7mgFku4z0ZlyAqhQPkra+yUE1NdkpkSY
iMN9NIIrSWR4ivqa5vAoGzZCCkZua4VjhwJiYk8bM44IHY11DPz8dPr3ojzA5aphet8yGeHDUfeU
YnXVVPMzcTxZjUFj/ZUUHUxKxgncs76O7QFWvO+ojEQHHqTI0jMfBcOZ9UnrPKwzFBWnO7Y4qVVu
ZvHYjAYbgj0jdN9heVlargbstFxdahUCSP60qcTKtNlPuO9vYPNb1SfMj4J01XjV5Z+O/BPboQjM
ELTuOB8W6ZLe8pskmpf/al6f33Y/RfcgCL81KgICCjiaIqwTG7cTgeeDgCTwfN5kFzCObmuYPr3G
t/2GqL8Sp3j/WUHi7eTmZocIAmyL5ODxlMorWmVQeHtVRXSsY6Yq8ORo6gc7HiJJt4BO655gwkld
PsGCUT7xWtl2gDjWyIDsZfjtY7qNwnKTG8jxFAcYBm9vsp+hHEaAVl4sapma68Ep8inqw8MytWZR
nvjsaV6yH/Br1g5k5EANkQZgnxsHXrJf81iF66BSGInbn81nUWKyMDjWVzgk7eUIj9NqyMFHn6ib
InDxnIYN1cHmJr/P4OhDJb+0PvxlQGu6r6rV01VxrwUpsNUCECZh0G3pSOxQSi8/91YNuf50R71w
RRhOBUDmBuYMl3BNSFT8n+SjqXKYzlhWB+395O2n174iRTYP3mZC1EMe19CTLK8yBbJmgBpMhTtJ
blq8c3KGv203BNfg97ayi5pkwyTUl6NDvdPI1qC6QoIO6FRJ+p8lxIBAbhqbVUmiPzE2dEYd04Ze
z6zLMHfGBairGeMNS96AeowOjB229xUCuvlkT8PHhM2DiWJEDbVBPfAPsB70WM3rfBXVw71snzA5
rbUY91ihsChntHaif/J2I3fN1TXoUco9os/YuG3Y7tnic2J7r0obQgLl/YvCxnAKi8VCP4ybxcRf
lLwwtcxypX5Jjx6nLyiDKRiGoe5gOWFxUBTaLg1FQaYbCWC+J25JTTVpoy7nhgZ2oSqSTM94wke1
Q7T6zd9+l4XEbT/SE1xCQbrACbdT48uynbFbQuh/dfVu9nyjTgW0VDflgATGxR55U0mqPKK0Vr2R
hsH31cYaT+UtnabenDz726v3+l3I1Pp77vNGZq5+sQBD6YUNmQfkQJ7qtgC54oLfYw1i2x8SiSH6
q0/Ik6gO+JmzKIvped65qHsnE3XDtA0iN0zXBK8DC7BGIQ5v9UiOBY0jdymIqeji7WMK2L0z0rz3
VFC8hxyG5Riga3XVx6KqRv/jIGclGN5R3Ib/C1LfOJtghwzt7t3z7u2FEzPK12eR8njUcdD3adMi
qDAI6BKqGRACe8lXJFM0nCPIjHuBG7AgiUWg+HCwYSr81kQo8EZ2+UBzWf11yBcjHBXSKcHO1ixp
pwN+EBjRTmGAMoOOJFQg6twBMLUvM8msVNGBkrr4zB3asboteYZZXzoiGaNDaYCo1D6Hef9VL9HQ
iBkimhPJJgIdVb7yOv7W7/mvhe5C3TqMJ3WlgojPgFVyuumvS+JMC5h8Nii4PtnddbmwjIsz4hjp
HS24ahguyGgxC/qzH5+950DviaWm8/TqocnQNizfxCCFaD1qThGHVrn85xMC5mf6AgpU/Q2S/27Q
IGcj0NZv7YK6PzHpfwXiDFx45rBzc6asT5pAxK+HPaxbNXfZ0QJU7RKgS4wrWw/Dwqo4YwsnhaD9
Z/i8NrmFWLvkoFOwlhJ+PF+zgjlrRManwT/W5ZShiTv8s1mFeQb04V+5/ywHEdf3Ke1hhTxCGCLe
30zXOpw+/0OdZaNI3HGOJ+TArkvDILBv1yp2L5+mon5ZwNv7LfVmVvIcx0zOaqkC3HIgrSXMEudE
fBuJivlwMR52fBgPuxxLBpoKmWWF5luPXfRa4VR/YWqaaJZeyqcEduXppNgR1Q5/ula5pxbYnUXd
Bl8Hos7oXxRXuTPE82PMNfcoasQ6ryNhZ8NdXjWuvKp7tAQO1n62rKXKDRmP+E702tiUSQcrJMkN
ZOx4SXvzU8QAxSW9d/2rBHcLtbQYMcFExFGbIhqCeuirOed+h/ivV4+1BdAIKlRS8dRqWi56D4cx
7zYWbm+zDWPfOatTS6gU04fjb0CwWVlP50d0g1tUAENND8RyGZzsVsGaW6pf9ihR+A0l8pemYKbw
pTwOEuwW5LVdAZqzFyi9FnuloTS/GQYXfXUIjiZDPCGkN+S3ikd2Vljcxh2tfqc17gcURSe3NL1F
DnUpaJbNROq01IzB/Et0gZyo/UVnz8AKbfC53IDTMJiRIVEIPwJ7fl9vq78eGTUYDpKoBJ7fy+sM
kwwuTl7ZK+lqe80x65hSA+mM3Yg8B6eOZs9ZEL5JD5534jazElNFuSpSfj3wrZWwX4jX0eDA/sTS
NpMBRdED4p3LV4p4l2X1WTSGMHiStSyn6yK+Ea2waZ8By8BSuxoA8h13QjVoSGOGQjMr1+lPDi+F
gGBI94q9HxqK0g/s2Mr8qEYB1WFt6oH4rUH0/Xo57k53zElle9TeDHPJV/7GTiJNXpXzgcwRLTyq
cV0so/SkL/jaSBzm8NJdtyElV9Y4v8G3POGSlz3uLY2SG8JLZl3FEvkDN8S9gN2DfLfht06bImKY
1a+yr6FOp8EPraeYV9s9JPT+NKbRBCCy68ig9xr6TqMvWOu+lQ8XZ04WK8Y05xbeXM33Dsne1puM
d98yrcvTNDTJuv6XMbKP2cQSM8DnjfEGqi/cDxO8KeoaLyHngoFVn4kV60m9Gg3Sm/cBE6MguXIB
5gNdW3laua8rxdBdyo8+jDPPo1oOlo7cOzNXTbRisfqPqYZJzoI0+Kt7KNCydnMxykN9xedFnKPg
qmuvchA7DPZLTe17VgQQ6JZIfPF7BLn0DGFiNLZR2O53Pj4FYFUuLguEQG7JzGnBOGm01EWvPi9a
VCgId6sAqh/D42sT94yZgWY0hb0h+Sn1qCBrAjYA/v3k4d0n1guaL8yPGz8tsgyYQSjCl2on0ia9
ALGxjOxsAaGqGZ+o9V4XtG3WJcOtQ3BDiqOYMxiss/TQxN3SyoDJMZoFa5gKJ/XV97boE//TBlT2
SdAGrwALS6f2wpuab+d3sNYGgt/5Q1ZFhHVSCIjSAdVAK0Yb6cszEN32wov4lnx8bMv3mTqpaDDV
b4xIu+vIlJRmGhmbghBsj4ZRB1jbRNsAWtMtYvcrapZvr1wzjsYaPdLy/6mcZBnnqEyuQ8uNIii8
1QYxxAqaSeMI7kQOE9cRb8AXe0ltR7Ao2vooIpItelLM3ffVMaaNQHFIyAexOrTo4ACU1E30LGcM
BNv/luV25vNmaqHWKdDcWqK5THzSnb0M7DKy8iy+FUDxoVGtABw6rhZbZfw/fDqrLAHiqPGE1O9T
lC2hFNBPv67mTWBzp8+28BbsPEgCIOELoTnvvp0XrAcgSZBtE6q6RsQ5j2isXo1GuzS/F8+maT99
7W94CJRTKjG0yvNYFoOqEqQ2vVs/wdNjMDy3+L42ueC8oarGEoiU0gSy4SLC/YwOqEeOBpvotGGm
uF2vmja+twSxQVTOT4i53a7D/X833IsrNCV3jhcGKIrhJlfsU4QsnlPXW9DyQzaWJliSrzpggyWC
WDI7g6Hti6QZX4NkGwHKwdoRu1wpAYjL3W8j8VeQ8lpZbGK5YXCuefnpWGIp+QBdDniEQ3AgAQ6k
0q3XSaSxsnVsHag6Rkd1QQzC4aegpo3XBSuWEm9rFZ2XerOEe6gpZH7Vj3V9HVrNor371bYpKUYb
Z0Iyvyfwzh4dXwzh3EQ66USeCwOzSuai0qEDmWtjtBwmPE7a3l0GMW3zDJKOc/Fr1gIu5YCp+zcc
xzyePja7tEODS37baJ1XNYXvd/28zbiAdqrWhtFJ2Q8ttYUH2cqCWt006ntOO9e5dwValW0wf8qI
jE7rpga1os5vjLDWWzFS2dR6KVQdvaJSBv/JbU8GN0R5CgAizyarHB36nQVFxZQzbq4WYZZ91PIl
PnhKivdzdINaJoUT+g97og9obuibo1dyCacrjbZO/+PqxPf+EbssYAuvFYIE+w8lLMX5t6ZSIsb5
UFx5tw78DkzpeQuXjFyS28RiZJtRAQiKlh5Q0mdSnewhqEglU3RBcRAPcuWFX0DvinlUFEtuG7OB
a5V7eXz6SqUipXWsiF/6BIPszOGTlazctUcV59IvYtBoefHXfF5Gr+PeTi2KSZKMndQ960Iq/9A0
/MKWQm/uH686q8buvo5isDIB/wJFDTZvKE9EfRVzFPkqkJ8VLOYBIbL7P/SWpAXxgX+V9Qw7BXTR
0dXcFGLfOLtxsXzoWvadKsDt1nc9NP+GJRYThANzq0GXPxgj7/H73L+2J5e+eBhvz14qWSdljuil
2TwpSLzqGGQQglZmnICD+69iDboRSbtZv5Azcc2C/rKTyqrbLRMdkxXDg753sjUShp34Q48ZcB1x
Mp/PreXUMWred3j4jPDrkeajWopa89KRLcdP8Y3+Ro3SLefsbKNhAgZvEuVZlfuCsICNKTwPvPE4
Ie4/+nHc7EmaWL3tMnKI4dwkw+RoLOXbMf7gzi5xk7zkKM9udUAHWxQ7mkxWQT0wZZ/KdxFmOxnv
T1E4IbtjWLU+/6aOozcOZsbUXlnPk2t3kiGale43vs2G7DLk7My1C26uvZV0CBHs+jfjBBAvboOt
ahjB8lgpX0PAdAXlaZFaL5mI0Vxs9htbm5KMecVjhkW1ykFyuSN/NFOjiVzxecGifzKm3nT9UKXs
e2mywTGHw106byNc8CUPizm0y6lZ6tbqi88+TVXA4IdxCfxDIj6h7HJZzS10py9JasYWuNQ5tNw9
F0BppE/6kZSta92jrgiOgRLBjRjNr1kLPeZxVZt3RXUOwSdfr4Z1EiVnq3mcR+LOefCwu73oMEqH
lAgmscY7oMnXETaF46K1TNXjhejL0aHwyQ5ha/O55c5uVcJzBbDFx2EI5yzOBlHfZsXhZjGzCaOD
GcpUsjgAKgjDc95c/wguOwdckkqIZ4XSza7jg1uKqmzmN1/9rTEGUwVw7IS05eGYOKlZdgqG94/G
uXDyZYRcSiGBw/3ste9S7q8XwBH/b6H5aK4ldyI9kNFv+jGJSVxg7SnwjgOvxniKjkwE1Gzu4MnJ
WPPqh51KbTrQur9S+/sNvb8rB3iFZR8BM0agHNpvtnmK2K9djL5vy7chCUVTeMia1L6XdP7I2XZL
g8MZIFvN/G2HNanJEkYLR0QWREEaGe03KiXVkSIm/j0gjilebBkD/WwzcLAMLzJZoZ3P+i+3i4Fi
ulkiGd2TnCcy+Uo16bQOPapANBLPp/vY98avnj5zu2mJVixpC1OaXvi6EmYrBpUP9bOyzWk4DHp6
mMdzsuRTp0dzUZEZfuvnWkvWq0qj0kguBz8dffL+NCz1fmPqQWKNzhVZUD/PMJPPulTp9dQwfCMy
lZdiz0wEnUgTQzPbd8J47sr6++tj+XuqWFtMSLVTb9DjrHKR+QWXKcvg8l2bvFARO8YSTTBc6xTb
WbLBz+6A4U1ugR1a9GQ+FPPs26PTrYLgvB6aUs1d4kg8pUVL85BLhP9ulbl//wttuL5wkdDZaGdT
Nr6tvmueVMaRX7pvi7FDvTNu/fuNnWGDRX1ZzXv04hCOYZYY+KQyf4RWsxutVfLPyxDAYxOeUD7s
vudXaQVa2gdGJRcyj9O7NPCspLW2A2n1pO5QwCFLvXa/4h2Bm1RF4Qbg6lPSj4fzrxpwjFluZqTx
0FcmaoeGpFU4ne5sQA8fv3tNBi/P6LrOgIa+SM4uYngsPRQ7bDL0WOQmEW6QFNyXEEtKiYOCB5qV
yQiLKKJzHP2spISYA75lmcU41lILhTcE2bgWb21akEaHKYc4qjcP+QjbMtW5be8V/eQMnt1jYJwr
SdjTGXfG9SicKnsTbvLs3eDJtQ8UDEZiL72wlNTlVmBC2q7Y/4n0alsUTQGcSPOqnR0nJld3013x
ku0yfH4BQ7D0YKh2SqaHhzNeGFkIU0p/DxHR3TSX6u6Lk+b7+ZBw6PCZkCIo+n9RctYH8BWWC4mh
2gQ7rgerTJHjXnvDtr6YsoHBVeAeoesGFNP9ugU3rZrMVmP7d2klCwNeFW/TucSqSZg8IAhILB2x
FO+6455WP8tYCennSrqUzigc6ATqmkaH3HI0WhplD/Xv7awch7/+Od2WUTIPX4x7D9jLYaAX9nWn
7WFbhEnDAxcqccaVfUuKW34GIpvmP2iEPEDgTu8x3KrR4ZS7ZtAKe4z17W1FTmX9s1aCduSLi8gq
GC3HxWRfgBSzUSYFVU7AINQYoRGrDNLX349tMvuUFN2vWaDp940F0/bjP4nQFmEsXpa2cKnP1wnk
sFB2cc+wZ/s+6MxzwGq+gMMJTFXo+dSiiSAEKvsHTM6XMggcERUUinubOIgyAArufFeMB11TrbWU
b1XR42UeV0mwpyWNd2M33ckC6/Iq0DO8tGSPZs9qo6aYshOWQwKDgGeUyhGphgT7zFAco5l9I87m
9xQcX0GbgyP0x/aUQHYvlKmr3uaYHEjOUfcZbCAql66kk0QGFFggfsdMWHbawiRspZ7ATRB885ed
ZnZ36VM6uqJOs213PwOtTtKKOjHjl+aWhu3WaiKqSdwOX/vSS7QGM3ECEcD9h53Cr/OBVajUzNRp
op4SjVFFi+WIlnj3iKZSPWHxFky0gVkdsn84BzRKBPLg45CE+i+R8UD3Hj1Dlb+dp9dlQB7FiZnd
cEkaSSb3gqnVdyrsnqIfTIAUc0r1InkaX9deN4G59szudSYIh73k3NijaLXuZM0joSPWSLnwYiqr
8cmkjVHPjZ3Nc9wrMr2JKsZ8PtwGGypSZGqGBwGtUpWEz3xkkjjFonuBH+5dbwyk6nQ7iXVFqM7p
MnscHjmhrA0RMQLUnxgTP6RS38mYdGBI8Hs7KC7vuqsuvnaRonpD/cd4qhLZB5wOmF+H7zqBBvXI
Xd2eCMwt61wbDL18WTkTlmObUrOS9iLHbu1X2uvGdEc5VxeA5qIKFtYpGEGBCNP9B14rF+tAbL/k
zhnw0OSyDhYwSoXw9PeOw5P5XNwI2QiUbTLJzDPFK/c0VUpTbyyKfGr3Pqn5hl5Ow9WwET0FASY1
rmehCTkRI1nSBkpKF+SnVdILf+6GE4baGwUmx+e8+7dp/pLKxY4kGcvMoPVvHKtCE7N/inhhP9cG
X63IrwsNPK6pWWvSsNdaObnXexpVs8QTArfSuk8qACI4PaWX9Gnbq7Ir5d2ERmd3CCWBF6nTydPJ
gDtX4tWj8hcazSXnMeZ8NTq29a/tMFbbSnqZKnNVZlo3nUcOGlNS77C8VW9yQvbtfEwnxS8zR8X/
V+R/YbWtTzXm2/mLOo6bV/W+zggga6mszXs/Ln1qzKO1+vKPxMv41anCCoJM/UxD5KfqWsZZchPn
b/m/1+xauz7zXyouZB69WndZ6UG8evF3VS6nTkwXM5TQ5lyRWfOL+q16KTI9wMVWUn7R7Wx/s9qT
WbA+0vbcuJ12o5hfm0Ran3mIyMhxQioIkKvmZvol42EtfWkv+DdgNFLcO2YLG9iS2N3AL0NcVUnT
U3u96SnWj2AVo0KpSN4Xw5PsQ+W2Q5Ob335ITbSZ29+XB4PK2OgieUXTt/uA+0bFqxsyWdHBdAQo
4wJTOfBUaXvebEsUvLNUemMthP927Jyff00wNcrkUySCv+YLVq5Z/4HeW3Fs8cHGXMvneHvnus+M
KvxqmEtDF7ihbdsg4psO0UNPxPH9a3O1ql5i3RXSAhcc9t5LQmv+redZudZiVMOBOiKPyWvBuDUX
O8wWvtnPVzyeH5HmrOcjB0evnGqPog3tOtPTvldQhtH4stprEM75XIIQmmpDE9uifHzbLI+4K2ep
/BLiTGpiFjEsm227JERLjOoCxngCeegau2cEjv7T3Yr39XDMBlXLJiJDWRnsSEQ3TFuhnsa8lx1g
ecPnuulf3UIA39Zwq9PWsppJ/vDrPASseqCzMzbWeVzP6XvAA2PUQj8OZQ4x9XyAhNyXzhZczSIs
2VG898Vn58TgbFPSR1QoRpkdapp71mvZWYYNjU7TVDz2DcEmsn96/jEnv1KCfRUGGxt30Zr4o6zT
dsl75PZ30pHIJ9j7BNAyvM+ng10HPfrhW07aO0fFWuxi+TAeVecIlAh6OaJ9UvIfraYAGfgzZ7du
Knw44oNfG0Fi2VZjOpcZRXqoqrJj+uZB+svgaLmctSLYi45xRnEIB6TeKb/lN12L/a5DiB21QOsW
3QPmyvIbovCoKeoDIy1qd6u8NbnlvokWsdj+IhOYhNzaoijfdljZO4ovYfXn+HoWHhBfoJ2T4NGX
c/UWnmI6GdLkLYiR4Xgm7hj1APSTvMKmb7L6ktjkb/pb/+nWSwRxKWO6yDpVy7oXYuPX+oEH2UBR
Nw7TAfJrp9BXcCJjomhibt9DGsVA+X9+S7q1Blwsd2iyDeBlbcrKe+XjQJnsyHf24H5aDJC4u//9
hObXwUn+2YpGyOl2AEjkDZNYtNmZOJ8xuJUGvhIk3SFH2ga7cK5gGIWE4glBPnWG7LsZrx0rTvPZ
2qwWkDJIUSUghSnafY0fDr0j0At0HYljrH1T25Uh+BXFOEawHDYDePs35+wvldgypLjxuQoYGBh4
NkXR0PKlUiinOfUhw42aRaLlikoswfiL2dcDiZ/766xAoZ3HuTjGSQzuzyJxRgcHGKup0r8MXYtK
cIPX4jqNLsCTm5UhipP8Jx7PztpkyyvSbZnw3UBmvy7DrPqgsYSrKXGpK9xqGFAniSs9cF7UHcXa
Ur0inJlHByZB/22O2VRmoSWbqiiONTXOTLKyg9tZm8MQaIRWce96/lsHggfEnQUlulG2zP5DAH5r
ejNJ0vxUUgxVCGguO5p2bPdbDWlVvfdpAF5LD6h6fhRgMCZg0Mu3E45TQF1Pj1B/OsRy1Mtkndc/
/1+pqJ2zz4dp24vmDfR/inFQKaxsJQ+XydlO8ynwyv1p1huEDajX+WIluHOsB7XPlzSk9CSxvBtl
34uvZdSiittJbq0T37//ts+qVwr3RvZBeQgait6qKGsbv2NTnuwVhx5YK2iHYUkAN2HrG9Zcsm/W
cO3FLEXr0IjeL9oBpb46E/iwt2RqE+6yGxr+R+xd8Q8Dm6asNgr2AncnHX2KjxmCil12xzVj5U1a
DRg6+093aytyIcA66z91QZs4NabX6m8VlN2h3HY1K06ZJK8M4UuGJUpmyrvvv/ta/u5fTrh7V7pB
05u8XWe+6pwsXRuV8AFAozbtDdqm1H+FShpI8DDxgRilN+/IvskFkVwPAKwmCYEOGFPyl30fatTM
YBvUoVP+FzpF0YevgC2a9GzzwYCjn5OmxoequbaaLv9/dxJYaqAgFDKZx5BISY14Ahun5siQty0a
vM3n5UDVra9YBB6scT+Y1fpa+W8cteIiJCfB+V2sR4CFLAzxsyNK8LWPivBcw3wPwi0LoAI1wa8c
j5UYZ8uHP0QKU311PPOzgMoF2GxThVv6F74kOBMHI6jx858Pc+vHmjwoG3cIkYuc3G1hKMz6bld3
iuhl4gLLtkIpyZALLtYjKgPK8EZ2wEzuO/i0/IQK0xY3eqBnpgw6FYwKJTqNQbsZweNwX4yc+FHl
3yJia+JJEQ3JaTdegyWeh1uRxHQ7gYm/0yNEn/NAz+p+DgInRjtFx3vSsoznfRZ/bD2SHOTPGvvZ
1r6/QEmcrnDq+FIpsNjoW+TxMPPd56GST2mwEykugkGxFe8LG/6peFkQuvTMBdBGCWZvRxrgGTro
8J+XIcP4IYhA/YKeKFRlUtEj2A4tRXWKDWaWPFLeEPRThNrr3zab2E4SbUaPCBGi9d8q9Q/rnNtV
2B75xW9+Gtt71c19ItX9IgtIPLn0EAQbHqitKFANImF1JNA1QtV8CESab28mO48aAUld2vNZW6Du
leZGK8sHeB68WVh5J+PPa34a9nLKqqVeFk3Ji9sO0OERvxg34i8RDvsDUAeLnuExuRfQvdZMZahN
1rKDO1M0FN7PDsTkTGr4Q+eSy1hvtEUj6q0sXypHcNht2QlH2sHeWY8k1dDf45mXoP6ZDACEqAII
1EgowdNrvBMICfPZrH0hx+9H+x4Hu6V9QDev7qMEeEQb32caz4B16XGzL9IrYCr7u0m+Tlr2CDaY
kNc81jdjhWHd+54PHm4lmMjBV1sAKReyoiBzZx/wygkdqsHQ7WqqNiQ/6dqDQd3uVG2c4gdB8qJU
wN1LZyIgyFLP7MwrQFm8BBfTuDDPnfKegARXqttf2dJY2enEk8idop3mVoxiKVFvoJ5hYqBkavIJ
3hotI/gV0hgUuk4qOAotFVgTLWTeFe9SnIMRspMS89F7EK1szQtFUBs98jkc7DSCmA6tAvFEi1l9
A23160/WB2noLd/+UmfnbcxW6M9+g6in0M3bKC0aVgAUOea3Al6mSiTOOd0vpIY6HaBa+8nvP9S0
m4JBiWJpAjyC8o9GQA0G5fEleJ8lbUmrs4F1MOieksZHgRZSlQqkOvWa2L7r2+KSsGBX+gaZHHNv
mI85gyROb8Ov5kzVWjF2rAZnQEDL0mZfepnfGoPVr3LnbPflg2LS12U/XJ8HpXPl0RAtO0qPuF0x
sbf/WqbrvyvzWmiwG6BMD8FSJfNk25VCRsOwFOIHkL2x858e0zC9w2/sYmyfd8Bjx2EQKeleqQix
6pgTXB23LuUGIIED/nXQyd18zwa8XFcUCnxXDzMzQrlZkmSwzJa5FPQYV6hB7ACJhRnfAcnjPua4
lg3t9dKkPKMQe7988qYy5i1AKw0PTtux6kDMzc2vKMtLzvDUQUmB7Q1WH5HW7ssV++NFdpgRrOUU
dr5bQ6sGVH77PzCoj8zsmSj1puOkaIiGWUu7+NFaTikEH7KGvUfgEcv7VdthXSRfrjECtMcHX78o
qzA8NtwGgSpxBvbqH9FkNx0vtEAOYZoGV01QB25DjawGDZOy2AMEOfYG2J8iPPwWBfTlmoZhSz3y
mX2dCeTaDYeP+mImeDNw/TJTQfLuCUvisqZkHy6xBOLHcAqv+XXRb0dZrH2buhjY3p5FNFLd+LiP
+ar2dKAlC9UxTLcOxPSD0hWHZapsDJ9wh6+MkercEGJxbInwuN04oQcn93eoWpc70gMHVbF6919l
VWf9odqTLtbDIE3VmplRvKnumTddmuG27BR4M9SYRMs6lIktTw2k6szv37njMpfsbqsUv/VPUvnP
yJ6TZ7nLEMy/thdCFcfiI4+rHjgns2+/I4xE0waw9fT0Y2o/dWMpwqAmwh7WxtAGp369Cy6EMbkn
691fFOdPU8GkS/I7HUC8f8t1iK/xWUJ9zHgQ/nK/9P5w3ZHJBX2Tq7+TRzg74j82hcJNtB9a3ztc
1IJ36k00TY5sR371PfIs8zEOX0vw9QtNHGcgxlzEB939M7EqxaAUBekgSY7wPQ3UTQKZH2Zy2WM8
r0AiJu91zHkiL3ZlTmgGvnIJBrbQcl0kjUw+Nip0XEDAEUhuV2/ScRGUAYePqMJ3ieE1EWAQVStC
m4sO8jQVTJQscUYDOaoK576dr1bXW7q/nVefkPq9PhUG/j1MvaGiBWLeZjoGSuQcn91uLFfpwYbN
0GrhItuy4JXfhMo5/TMZp6HOzZZIBsQE/7/FRqoatUxMRcOJ60S9ZgTAGmBdugYA0nZ7BIoYJ6D+
9ZefHzrR3Xt6p3NgkLH8vN2lohfaYfIyglWKm5Nc7Ukeln+L1pnlbfkYvSDOz61O+ciP9w25BTRh
XQ6Oq5dffyOO2kOglhymugK+S2J6IGBGwoY3eSeyFxfGgAD+0sMyMwKqX6zjv9d+M/eoLDfUEgUr
LMPqiyiPGWn0ZQafASucgCtzkUxSu+mMCCKptmw1T1rfU+jTlhotbIAj7MtseT6Mmkqn1fxUbzvK
DxuC04JL+MCqZ/ADGSfVcxy90lW+pfjyCPxLXQdTO974KKksmU5/i3lFJcicBrI0QNtVztB3OYF4
mDJSW2rFf4KIcyGGrwvbBGAM8mv85nnP59dS57pvQ2ATbMJXjWvfrUa1omFyzdpaUdGWLLWVGD58
uHEqvMweZaSVJUIoUN1B6ovBJxjP4Gzf/1iElVHjq/mYRHmsWndCneUblN+hoq/NZpF/oaD260HA
YS5vhyEY7Q3S78ECMqAU/hQj4bu/IfwawrGvsKwTGYEiFsXV6k/bxHTUWlIDgaGDafVoAuoaSz1G
861NWX3/pz8aS1pDP82wMpy6lNknAZQnchpdsTNTycnSoXZwFlIb6jfESZRNB4QqjRH/1EYRIhYc
rcULjR2nZKL+FHKjKctpJcmYhreAaQqrlJNIRP5r3U5lMH7ywqLzovY7S+ENzSE6702AFdubskJ4
SdJncI4AmhJ+3NfuFTh577G11x0CfpvWw43Ih6XG6kCndYxo+K8EB2rP0gE4aGof0gIc18ukGti0
tCnR+xhTw/+7KEuOs1wIYmBAWz7SFbo7Q0eELcmusKf5P57UWn7lIGwJcasOWUaomDlB5ahLyPZs
zxgjo3FZ8dVik/5NThrBaZLq8hImWbw4TISweYHCk3Eh8h1LiuikMYlgNVrGo1nEcU2BRhUA2/EU
pYIND+xPG8y8wT8SNFU2WIcb8D0bsj0pHx5Dx20fK2/lX4EvB7W+N8aj74Xvvf9MLdibxxA7Km/r
L78UGwOMI1hNMI0HFen7E9DeAsTmndm32A7zvdMOLUAfFiGPpJJUoLCnCg73JUHevj+EZ2Ft2cT3
bg22QlwYttYKYTmJplNzkcA3d6Zx8J2nGaviW2QdBxzg2cuaonDK9Bes8m2hzwOYJgedtOgtYMbD
4hlEL6tY+iG+OoZC3798YYW+hIsmbxPAhMaj2bV/KM412FEjjLfcrHImAehWTFuTThMotlyR5kzj
OsZiO8SgIsMnvloLBsP6U2uAK6c+UlZJ6YYF8wkIpARrIOIB1rlwTQ80xE6pbAVW+ALwziDyNArW
ey09puI8arXzsxFlIFKLOtlCB/gfFP2avpc/CinrNPx6zWNLjEAN0zgU3ZeCvp8qmKIFAo4mHc4C
92FL/C6v87iIO89uuVWMa7/eudjy9QHPfa5W72GzGMRsL+z/cuYpA/88GaOr03PwhXK3+WlOl6X5
vt+iu80nrXKiMoa2GZ1acxaaO7pQNV+VKdRyUk01jAWTlgMbYy12F3vx80G+8wQZDF5zDINK7/w5
N89QLWSdcP6t11KAw5R+GRzVu/UHspth9i8Ip5BDEIJj0EXk1k2e+6+yOxbU3Y6EUWL+2A2CMcvN
9FNLkeVMR3tKVK6josBkxA/4AUWw8e0swzsn8sRSFomEqflem6II8+qsU8vEQD2SQMezPZfb3+DS
ZRWHa+JjUeToxnr0nv/v1ehEzXZg5MelkSRLxSD0TnFjFi1wAbTj5WV35PTFcgO8dGtdbCwSCqfo
Xvg9f5zrKG9Bx+Tl/C6yAk42x1DU5lfiRESgiZCLbQ3daDSBX3ErIctzxktFW2yC9iyF+qJ+nRYL
RiD44qjjFvoCmQGzFS3TW4U5Gf1dm9rv4DXU2PDdQFTxc6ocFrHOkwNCw+MRQb9ytwvbiJe10OUG
ZUklYSRGlcy4mvTPphTIZgRoL0V1EV8ls0inh5270Xt0HGFa/ruw5f5p1rcFv+j7RsouxKUJ7Y9H
DvmsCj3gtfrYWM0Il5sEB8tWnwZNvLfSx++QX2P4U+gbPa4QV0qkrnD6WMy2BY5+qp885IcfYN7a
K/K3pWuf4jQlxpzAZB2tglVfHFcLTt03OTb/riKGVbqmDBPWfTMizKpAbC+WxiXkP1xBUT0T9Kxq
W/VnWnOaWVBuxTB40Cicd+E5rPM5pb5gseAdH/HCXbCWPMZX34notYlH0aCNeISd7QVOH0tPnEx+
OzggQM4pNQqjb6O0fs0OVM1uYYp2XfhecNHXX0w/kn8gbgHiE9dvy2Tf3BhFCwjATcr0KkEYSQ1A
S5lPpwqXIWA6mxIFKY4FLOrxY1DGEXsE2Zcd8EB9th1UsP4ubwADsJ1qek2GXwYZM7LJR1870SUG
aP+F1A8zjiY8Yib4fBlSann9PuMON+Nv95bKQ05adQW7d0fuGlZHoG/mCw8607YYNEvDxr4beSa9
tElLYku/jQo54IAW9Ty4gZpeANezji8uzry6lE89NdeXKiFj9rxfqVlLBliPTFcofCJBiZ6RxB7e
BQXZ+Et3pfTJQthtS956Sen5y88AMtWzxdUI3f0taifTWATXo8jmGoGenDpNucOvbjLTjpnk1O2S
NG2oqv+PHta+2xjR9LYeRjY2MeAjxy3aOafuQHxRNhWvg1t3I0DDzbCipEldlgDZpuvw5M2l3z2z
CcdUAxJziwZ06wO0oXXssLJdMPdl8q2swzl9TwaCaP0brWNiER6fKijePzhD28YUeoWVaH8YZeVe
H4tVluh5ck6VJnkfFiqFBImaB/H3Igw4CsM9HBO0yMRBPBM8yq/Gyhzf54KLVIPviA6ndKDhlE5h
xJO7D4TATvkYGxhlPGBNodEq25TZ1CTvG9agTGkVYA+a6dYxC+WwH/oXcjhReAQ3Dg8WBZSFNH7H
onsttucEJ4It7Q/b1//KoqS5mkiMxdbbbGyjhyvMOZgAERY681Tl/KODNe+dtDeBY09aQdMJOBDj
RE3B6WPSUObjlntO/M7GvnAoWsUQ0p5K/TPBQfEheKD/eVar0zJJSxO1Nf5Ce5AIhEgbOCcq/Vqn
Cnw8bxL9d4d+hux4rYAF5uOcvbfO6NL0cwz025BSLUFcVflxFB7WDszAx4RKjGBSp0IcQA9Ffa2S
qAFYtBQ2YwcBVn+1mFEZRCSR939dhozd2l37vCgNllkB4XNgCFXjnqp61dcKh7RU+tTi9wJkQG8m
Vacz9j2+K/6dppPX2Cp0VxTCO1MxbKFDzvBWSKG/D4s0FHnixKlnZEAi26SC5rIPA4f6S5s2F7Om
D2h/o3IPYaS4BJNao2Hm4zgxzFO0keIC1HOKNtqXqL6X9RQdqQG4RSymTJ3KQ1sX7tf8IzjlXsPi
l9tTv/0g9tyWTMPDlBW0bBwnsuFBrEem9rK1s8oqlKeg0cgBkBKl0Ge4aoDVxfYATy67aXcgFs99
2zCLm2N/xFLgvNpgkYP0Nd2/KMXzHdiRQ/l8ia+mULq/5XSLrCKGM8dreF4UMzKIJndVV+ksbqos
Jo30zOA+ss/Yb6VSkWfiRdTPjFSIq3xL99XS1iTMMdlZHUJtouyOnXFdvGi2qkERpYaQrXrGVkaF
4WuqtguJzY7hVzWAsnEeDhnWqWScvRl9HVlLkb1yMEiptMBDTYgt1uOZrRhzAotlUdX/T9AFAWx3
PxUn15tCzWMTbO2gaen7ON/FSHuO3doWYohLDUAio4NC9FsVgthXBDFBxbrJQd5Tht16at8Z7Iu2
adY59Nr3bx5LRGZFLgq/6Aba+IlHI667FBM8wGqFNnQr1liNY0nze/CmgymzGGGPdKj9XEcJog+5
KcXoqRA078QiwH3opShSMHBlfkqEhMhLnERxxIawnO8RNE/qCCzWV+CkEJoDqyY5m6eeq6xJuvO/
h8ibmmNU5Bysj9VHujrTCQPj4PKUhwg6KX8E7TOuBoEOMF3gwsbu1O9tCDol8QTfIYVAl9RwbNPv
JGJNzk0vNESUuuuiKfvY05pxpk+V6pY6k+v8EPIolFA8sCOD3rcJN4C7iKO8ej41itfAnbidy8V2
hyqkxtG5gv7Q8eV8tuTbjKuzbjzUklIc2mvsOgjhtjP7Zl2/ohkBX088PRjEAmbNzp5aBl9rGaVn
7FyLWfUWtD6rwaTxRVb/72kOLU4pEgl8mM+gPBOFdmDwWxl1dGpxDiWG+KKrXpV9RmJU7MQOT8Ld
Kmf/aIHWMEbyZBg58csYhaHkY27eXTlrp8ARFsZWs/5jfXpERG2Ti4ABAHL6hUJpH2pX5v0i/+zT
hGWzjkP8XzEvcyBcBHOHDipJYt+lHmfQWAdywdeGXE1ylhHqMnXbMwRULuXfLlLBTbwZJkWGpU3/
EkJU4fpPdS74GhiCYcnSLSwty9w6U808hmrHqP6FBCGUeiKiXJ5NFg8H9t5pYSOQGPK0ngRODTB9
i+g7YMEk7zdbZl+QaRYrR/D68VGmquExidaSRys/7QV+86ffBs9eywWBi+EVLDyp8R86fypEpA7f
qY/+LTRwDJmrqQPEGJXkhkEmsbNittMUbyfPyoJq0ujgkHOo027Ma9mdQe8Zj3FukaUfqX4U5Rvo
5F+NGRTt6Q2isnvgAA3iduZ1fVugV8owDgmTRZ1vxWPIWNCYcQfyOsLHsQN5QfgVVdgSsdW86rZQ
tXw4g86/HQupIMYP5mxigFA4r1FwdS5WCLiat0BPpjBZscI7Z1onpIFrJGreEJniQyhQ1svMC04J
0cvtT9qC7UckrzCqJdMzGZfx1Gs01CiMW600Vw9u8ZEwavPQYctNe9/tALIDhNbgfyyFvXEwa5rU
HROZeam7hwZBxiaU/OKQiIDwR2hCbfem/v7ChQ37WaST2z3jkGocJcWynp3Ev0dADyidZ6XDb/ny
nDczX0mEAjyr58U+H7C5hydrxSkdL2nVBU8qvVvTSm1D+obQ5nbf70kqFPm3bIc60RQ+52Nc/2OB
yT4xzK1LNGREYl5ktUfsG6MDeYTWaUbiz4gMphSW2rU/rRMNFyxC0dDKM3pQm3mc/X4R8JkLZu5G
cousVL76ptMJ4x0t3SLJsGg+g92d8CItND2oGFhtWuymddqHmIZ5tOQEZX7Se5/2Y7AFU+ruvW4P
D9AIRFg5aXVZubQajohv7VlZogF542UThIoCs+uHuay5xQfXG5m/acadBXP5PT6yFCmS5n7QXopN
dD+RTBDOUYYyngL3WGDf9F2H8vKtwIz4VAcZlJwGOAnTk0RHwMysmQrMS1Q2pWIKdIyrn3pDYsEm
xZFEDH4mQJyG+9WZY+WqYTu2k8BMnIe9hy32tX9tTVDU1bspkGJb4e4xxkfTIfKOoUOCdW4HFCxG
ppeK+M9k0fzbBgyRhdM5nU7WlkK93aVedAjTZM3ZUAvZkfGaw2UsTvqVkpeRn1KS9gTRazg0a2Pt
fDUEjKgk7Z0KvPxi+gb7WmxdPeY0TFLnjFSJO0ThG6ZpHQbGD2EvEpiwthVWOfZbJJcZfJfuq1yN
749C1e19d6Hz0WF1oMOt2Rle4xVd6zOS1b/UT6N/Cb5l2RA1MlGMvAUjSGCCHlv16W5qwm6oA5fr
V4zk8VVzpLit6BaZ+M8FOtbTwKJ1oU3u0pLie+GlwJLL7QscNpnLv1Pr95czvygKltQ7p3t+heRL
CqCbuISt1hCPff3n3a15K/lP8JxosAJyT1WLwgBxkZj/MGHqesB3R1i8Hf6yznY16rjZpBNr5MSL
ATBDyLwi/Dm0jKHSVb+PjOCKbAIeOS54LrWFgF5fVbbCDtr+mbZY9e7fJZ4T1E0bYdPOa6ijP7hc
2/iATvhuWbxaRio7NzPqyYoU5xxh6U9RO/iuRMfiKnreeVYheVvIIqc9jpJ9H0pdDXxBfX9S/DI7
tIRiESiEdmDMUcZ2DbK/kcMGLZEslWKa9fPAIwSnfg/1dsJT/T58CqFEKIcKlIIBnAazGo23Kajy
v6mReYWxiga8QQq7GmQXMWB+Lk04dIrqzUVi6cb0CrkWmRv/4AW6Fzqiw1eyu9lAuYWQOS6gZE37
EUzt2D9Tz49GVyBZh51HqQwlPhSqljpegP0OS/QjTRE6NUVLGEs4QfSEhMTVp2HakD4yRwrKOV9U
fsDO1YvcXFcJSXTcMkbxoy4hQJ3trik50wrDvku37ukS8W+Sa+IuXP4EP2o/iTq8YvOzSjIZ/gLA
BDmzl25nfesaPB3tYZtw/ZBzogvO6tPMdsiUo0gJsF5TXl3X/mIPSJd9JcFSeUV0MpYh/gwMOeRV
Q9ibshfAZcHbV7geIjAxnZomw8sFu8Hg1IAWARiTupeUBRD9LdJanQ3p4RiRNQMt9FaijykCOKWC
6bYNWkH+4mYc+Ch/slaYhR5HzbIKrnSi4h5algsFivP35cVr+Yj3tCs6RZh7A/59rkFr9oKW+yA4
HHzFC3ds23W1EtgwPvGMi3/hFh6/dbMV0bVT0Vy/8ZyiaJ8wFSuWyZdPPgZga4bTDOEFR7mgE2KG
H4HfiEx5Hqo01eRjLrjWI9KoLWBgI2E/hqYiU5PuZRJ07ncjIMDN4D+4AJCSG5AmtKNeZyhFIHig
X74l7CZyMnSfx8JWoFYm0sC5rg6NGfew1evRxxyR+S1K4iSgiNp4pFqNYlombNuptF8QdcKdBkvk
jwxuOp1GUbYqww4Uhan0gzwxvgb5QWYX+gI1Otzut55bUjZux951FWrmZNz4cT0BYRFmfwQC3CQ8
fTMlbPqqKx1itHHGUCWi6+3TJWwNagNIv7MEsGCVu64uGg/72wYFA2ZJZ5KCtLRtq2867u6OTJej
rG4kQgXBwDNHD+ty5UifmE8abVpzxmD8oKwPwSi2/8OxXCsKz/e/se9LVycezX0Q+nMYUi/vckM3
yKB2coG9LDpLMt4us/acESl8YxWiUJhcZCwh0GE9WM6kftz2XNuuWoMEPm7wSJ665H92ZHxMkYUy
9WqUUGgv2uNIODIgtSKg813WYPjGJ8la+F71snMewANd966EXeUjdmVmzL14juwGwv26SCZhGVFP
l8dl+uJweITFZUlIsrvbYq+XBQ38Bjk1KNQL3yyTeqmQ+KA5XLVaueRG/les2+W3Xsy9hw9LLOIg
74qR0QHjZysuNdBdVyNm2vmJDj1RTA3Clp+GcfJWCUpFuBe17zT4ps3XIwfyFYvO7xW9MFzk2mim
P2//v3g3KtXiAuhYVQsGwTHpkzJiTDyGivsl32oM959fgUjCP6fIgMGqwk+cIY5zoDAvbaTcfCQl
psCqqi/TXBbou9BWAm1UmOemJJMy1xPkqNI5ZlbcYqOpcqFtiMMEgPPnX65bMBZVMW3Mfin0QBjk
19mhN0tN3I5mtZV/UEqtV4oDlWPP7BuztetV5qXRWclklBhklLcfOs05suxZfPf0+cP3YuF65+CM
mYFlTYZFTAiR9asyJkgiEDAieszyCAcVFjCQiNoA71NqLRvBCjRlZTpk/JfN2PUAPfVTNoWvjwiL
J2LlevepASBHtJMAc+jNfkWaYr1ssRkqbM44HU3c+PFBjmtDdSuwfEW5ciq2xbsYrEMEUoOdarYf
bNmY0WPwT5osWPhUA/oUUo2ggh33/NupwoVUjFlNWkkB5OCp/fSgs/XUsDQlnzzUSeNeu1xEhPmm
iwk0C461bsv2+aIOzJPVCEktFm13CPNEK7Qfg63y6h0sKTsXIna9i6n4H2XpX728w/HJ3ADYV3Rq
XHFX/4l1FBTSqknMgZt1IBXATtxva/FJlCkovSKwpXGBMOw79r/BmJZGx964SAoNHTR9PCYrlOY5
NzoD7tKwaWrlIZuqSqjh7ggOB5tVmSpB74czUlXlQf1lU+bxJ+FZIabnwvbwbP5vMQzGywCG8kVp
YLrq1ABriBsmcE22QYURow66dQDgZwd7ISSb+8SPYL0mjmUlc7IFFyTCGVC7DDuliWNA3uRTz457
sjfXYb7nHzn3gRh26rRs1nYVQS7oHrtuyXEc+IEQhwsATH0ylX0/0ChcxMJj+iZZ3muyUYTtV/aN
BAtTj0dNJUVylavzVhGBuJArD5wOaWdW4sFccviV0YuAhqceC9um1rRlhj905ukKsCGVzAGitWMw
1T8TXom3nGhSHjNID8gyOTQYvioq8orZ5EOhJSiXTJRsqWqnWmVwsNyUvGFn3hvgEEb6HeotLWNy
sQ2eEPJMErinbffBNJFOIe1lHpew1vyVl9AKtXS8C6ZNS1VxmZgMk6i36UyNqHiEHHyGtI+LLOpZ
EvYNWR95VAcudHF07VzGt5/0xUjBGlbWR3q8EuAGRmGbHBeesxYj+Giu9AqVYSXPMX8GzlORkexT
G1jQICkY2e4XoIts0PBe/lbb9JfYs/Zlmlj8VCWkMkwebamNNu66JJXL+KWN++mM35k1mzzC1MEd
TAxx6io2tSkma0S0qLgUlaOqShLe7lUq/g+4dOuGfi+6+KAjoo/k1WiTJ6OuaFYkgWCn0I9oxkSe
gHR+ViMnj3qekdARZin1byCKFHGj9ns3MjFc8oQkUHCqCnF5D8fdeq748DnHJzE1ltRtH2yGGiYw
btjJ/tZPYPjoi4sgkaqt48OgdAdbpQQr4Creiwc7cS/e6KxICfrH1Y8+wXKdbd50+XZg34FrqdLH
JReUhXDVSgwaFYM4VM71mdE/lqCg11GjdyvdKhjL7cMN0uSInMJ7hYiOKd9klse0dzKlOal+sE3s
U9epIL/uCEN+DKWs29oyuziq1QA3YKw4I2HjTk6wBg8rIOGLqXr0C7AY7Y58W008FCBPW21iXrcQ
D/3XV4FjCc7EYvegeu5TznFWIm/tjZPNSWHaic8L/cxffhaFjSaOfGRLj49gQanAGMpH7LqYqQa2
l60FigTNm0gpqy/2keK75UfH2hYUu+DYGWQkHR4zhjSSgxWd1LgIOw/gpElZCf6YWinSh9FeSOZU
hu+r3qrfruWoP/Wj5JonyvTe50BYPdYGynVzVo9t8j9lX/FPshimWSci5mCoGU20EBtMIxVr0FUt
xNIhQdrrFtec/jMhxUiN9OX38lMQ+Z/qMOUIQ0S+rrduBsrIW1ugWxamo/+0t/xUBwKCpyNUTVtU
smvT0Nv/P+f4kPgH6s+r3lNrkVeaZLZJDIJaNsmkhtN5vEaGjVLpGsq1l09K2OQh4+j4Ztwpqr+r
94B5vli0ENmDNrm1+69KsSD8Hykn5JIusfGfa5SakMAYb35govgpATqRfgJ7tHJnppYlbcUEqO91
vlZ7sd6iCud/d+W9qSKVLsAep5Fc2hdffbsRHfU/c070wF60/f20Q8nkOhmhWR588xZcrt+3I/MF
33UPkJzEisby46o9yyBfvm76+DrEPAnrFMEtSjYsGkFOtZROjRTIRSxfyIed4C2MZ7DUz6phdOmq
nQl8GZyyMyoI8aBLP/HwxQQqTGhbFCVJ14Rv+Ap+QVTrwDonfQDob9N2M8jd+RjqPyjeLZedzzZz
B9JPlfd4nbKoR8dDL/4Q+ptIv1rJTPx5yL0Vci+BcTRSj1HSST+vOoDaO4nrwlvH1+23itqE+dzh
d2G1O0PbyTgM2armwQb8jiMrcqjJSYY8krwirOxgfXoIckqRDyx2LIV14CY7wD6gF8UmPr7OzlVE
CsRa7E5ZLy0rlCF8y6eSjsbYmxyom3hmPw3hELsmJ/FJrWQ7SRQPGeMTK9/nH7hjCgqeTaKkhrCq
jF6Z0Gr4SHFqNmkjEw270aazj1bHFZScb1h6O5EV6vXWrrxhq8F7+CHmnicPi911xPbZ4D7j7YOW
nt5P5v4W6uaUR1jgK9D7xnpDSzv/ATeTXTCDmUScT63YJzesAZf2tML3AfOxCC6T54hlBK2QBZ1S
cvf/aG/gzThBx3ij5z8BYh7LLG17BYcVbhZa143c6sDHo9NWmd0lHREtWofxqIBbTqb6OX5FKCud
sHLnVWVJtpJvgBQn9WQc2s9ggpmz3lWZ7CVEVf2qTR80VUKNbpN11eieXvr3NddJTuUM7MZUkfQ5
ATy9g7JGgrT8ql2XCz4sVtrpKCIKu/w8I1Izvl/0e0HA7T0n/rxhKdJyARicPy8AOGNaSNcX69Zp
j6d8NwDZ10ki4eQG33t6jzG/jHiYGiz7sx01x9U3QN85tiEuT2wzZvwZmx1XD3qw76KqWGtwA49t
U+rIJ2krQpbnVtACabUymj+Rccm0RFeNe92FJW1kKrHQ5uBYECHOazULDvkca8KgZDXDlclbDgdY
3AK870A/z2eeKojwHZrX9FNxcGatGHyV8KnivrSZefluPoeirsrjZX6HNd/jPRUJeTF8E5u1vCAg
lsZauJ54+EW+PpU/9Rd/cO9OT4K7SPc9gkbIoy7UmDlzKQb5f44FnB2jcP5XlVlpUuBcEHsy97x/
2mIugp6wWFadXGsgscf0ExJYZ1dki1XRYb64CdZy6JistLRJNRiJJs1Cc5RR5ejzSk5zjjXYHDFW
n/4LNGDS8V+OLmfps3oaua2w4tschGM4EUH9F0t+HXfDCjVdvypZEzZnEHxlC+ljIkTpnE9fQ71p
IAdtnD9hAVCMxihDIaJg6ThPAs5U5ZVAOMf+bmbBxmw+xKQMuliJloV4Uh5NqHblxeFoUAWeckrU
P4ER3Z76c2FHbIbe2hqhCr8ut1zU3yQ1TApwsa7x4evtbnXd/oLK8gnS2leqCfbpyZSj3xRQmUSG
e5Fj8Lup+l48XYZ1ybbctRaZPgFD2KOCQrmS3mEFrvnkVAe9SYLVM9fEM7nbKaMlTwwwh3EpP+Tt
qBhVqZAw6eEHnTZm4nfPtnX2ZipO+P/bx9VCRPb0PaAO6oP2Fb8eumH9M2i1BQeB4MGDBLI7+dnf
Bj1+LwDZv20INcDfoDed0D3BIeskwMBnjWapS8BkmHj20R+dpHZ21no8mdTDhWxreeBpFtSeo5Ke
tp9cDZ/a7fdutNWuB/gfo+l+REMuz8d8tTyP2rC0xV+QtMtwbAjZSIWEYy1jK8/wIsZCBlUXFtB3
vM71aSTJTeIZoOCNVQnFLwfSfuUwHfyZ1Ehpfk42NaQedltt6NUAgm/Ol89gbplys8wbWVPwb3Yz
X2epf/GUcCMDcI0wRS2mV4cn2DmNLQcqVnbXxQX4jL2k4OMO/u2Jwr0JnSIWCaVfJ4cwSqOQWvuh
H8PmIFIrjrF4H7P0VYZCnJTrnuZKN+zZZQQ6nvi9a/Z+gkfjs1N1lUo/BtfaDJ4ZcBterTe8cA3F
JCJ1KMuPkPAFSKgSOGXYfaohpkFmc/QPH5mlAodk4nOuvnVRYUA9DGd622LkgHPq3AgVByJWlxhb
6Kr58SQX4wvM+V373ICcOP0N1mJbDkmW/HngD89REmrKMQx1VA1WqmbtZsgjixFhP4R+DNClKbBD
G0VNFJ33WrgokAomBNU/4WowIBLTfdj9UKiSSveJEd1NQtfMD33RlgioMkRSnjhDpcfNOd2WzOA+
ESnycdIbzjLzx2PVXMke1J7lyc+J0tybku0wH4eF4fICD9b5ve2xkW5AvAfybpAQN21Xik5Y8apN
KUlNBWKmoQAF5Yp6HUwQugCiFDExmu29M67aH9H1kXhAtHlD1JKxvFLNDBh8O3p2HC4DcZ9UO/1F
ZXBG8N0EPDUEFaHu2hrLWCVgyBBvsHKImabaqoMNdpmKOaoRK+2MjjvBINaAycPi4QNgwLDT2NJR
Ob819zEOAUdDhxULaQ9jhqQsPkrJbr9eppMPFaiBTlZzdT6qzSKem0LjLT0B3EMJvjPLNSZOTj4o
+ZyhuYEY6g8K0odImSz/H/ZOyofDtMDf4e5JSO1Rmv5EorTEgNOasSMYXpV+RPNdmbnwDX4+VDZj
XBNn8TgiKTBsJCJHIaeUhvNJC+PB1UCYgpVkgkHrbf9Jcu4yj7HXe1Z+ZaiwRKqL6nYoPHLI0olF
j0c3m7AbpX8pBxEawJCM7+mC0wt0rfedV6zahdvOztL9wlbXdtRxKwCuZZeWVBtlBedOsThvdliO
XaXBBWAf6JiCz22g4f2pzSevreqRnnA+d3T2qp9+Me02q7Wqh505lm6OnHKOhiHN5flqdrskyvow
LF+AZqLFTX+XQYJOg/GKnc+EtHC2rnD3W+YIyF5UMZnD7XHOS44YIKYiR0dV847WzOE0N3mAaBEh
9v9qEV4q7QkvA0D0pvkobfh8L52u47Tj/Iric3c8Nr0Z1zcZ4mtnAZj1ykKw06YIQYfyYFZIDQ6w
fwUxDKqKFex9PIHvQTo57QM/eA9E6vcSjTQ7C1lrKzxbXAETwowxEe6WxPS8CH3MWOIUyvMlowEv
MTb0PKUq8giG5u/Z/iVcD+T/SLUeJ2e6EGmguvgyvcD1e5E6tmCdTWyu53khs9vvwuxYa8uxBoB3
5gCmIaQfVhSvyJg081NRMUqfHKHqL1XqhGHz0UEF9SnLmOdBrlpepWaqrSeVMh1kq4wwimn8SBPv
71r6ID8F8sXIAbYWKFKnVL9v3wm7SfmTc8ipcdVqHCXXYepzBGH8d/S7kko76u28emBk7p+H6ADR
xySeewvx5DNSLDtcZOR5JNO9Ia5f1ly7qN1x0FhNojqkUmbhkXv2478Rf7UV3muK9SQj9QXijN24
eCddT8pIg19b38wvwoTF/rgwAxbdyo4JsYDfbnqXiSCCJrkLq2zjkWieo0BERIoIRPo3AZdVZxA5
d0oc1P2gC9s7xw75XvjeHdfeWZyY9kJkH+bqz6LBq7BX4IETnr2F6Kp+CpSaTE1JZq8zNfo4Fhlh
ICUK26NyCpctohVxw8ZeKk8/GCzrKvVfUZY6+r8W6m9M/1C7wr9il+UM/cbbHYY6eLmarJ3rFlmp
X08E97IaY427zU4J1YzRCo9nwSCZxeouD8IMshR6armxhINDPMni65tZuLzy8Rcl3DoSS7fMa5o2
jNt+bUhfRmijXlbQaT63yopH+CjK/WnJnTNncRuC1Vd6uzPd6qBqPF978JIaJreOX4fep5QX5KjR
Hxi6SfBhcRC7E0R/TsReBHp/yNlY0vP2lBqGAi3ii9iFDkh2LHsNwO0PZacx9dn4OaN20e1FaTif
rOFJhaoFeRAB9LnWfOYmP+uhv/Hhivol0wDkKLwb5bFCP5hZrZEaW0nQRxVOerBbgymm1jezi+/4
tRZERl1GxB8266+rUFhdlqOAuOxHRUKpdxWKHSL1ZKNCuj3Lo7GncGO0Wu97IyTDDAbDGNUG1N/F
xD6geUAchD8GV6juQIyALdeVsivIJqvNAapNZYlgkKCMMlbrNL3zHxOI0fPU0UO01iP8Tt/kBmPZ
7+u5ijwVrs4c8FuiL6tJ8etUrTnHN43Ni13oo7HRqKxSxzlFwjs059yeAoTi+p/Ynp0ttA78RwJT
BvvZUDUHRTshnhhtw57eEkqzx63KokvBfoJYRKPWvG5qOZ7fUw/cMK26Xyth16Q7lMiziAIh/3Q/
yI98/MajYflJzoAmi0+w9DYFv1vKNVcLOvi3i9xyGbJx/YTjZX3p8Lcd1JJYr96nuoKWr3hNqNl1
E8KjjOEmvCikTWJa2bp2GMrTulAVR/iVkIvluhc1sAlCZrgN3CG4mkw51tW1zEM8PMHV5Qhik2ex
/ALHE/7nIM1zCTERrjNQYxySzAlMnQ25A5iWhu2A//bP3ntjJVDtXz0+BAE3knInmDDe6IbRZ1ms
Y5qM1ZkQoHYjRbCL3/ZDG7d2fT2XxKQG/3nnSexmShYaZ8tHEZ9YYva9BJ0T3NDtNDXeRjqgrc1a
brPPuQSOZwkINANEP8p4KLa1OuYzFV44g7NpKAI2iwR4qbAlRH/AZxskdiJ8h5NEeL0TVTOp2j2R
TYWLM2HPja8XEI0Bkxr0+55XTS1eWVAya9HbHlOfRxbKafnZgRWP4eP76Sg1p1evgRLXvfwYg/58
Ltt7m41085lNQyY4M8YtBy9wzyJ5CS8BiuHC/C5eSoG2QzK8sXOzUBPQsT+SVsU/Nkq+Ef6mcGLl
Ukb3CSjePiQujwgsENmouyuChSS64Mdc443P7NtcWllvsVIdiHA9N7+zQKf/+Rl5eXwmljBo+/4g
8uDox7eDcW+cg6It3wKZiXmPo0GchGE2PyIcvB6VvuVlKgRIPRXNrwgxxaMJbULGA4BA93Z8Yasi
hHZrC3JNRWD2y6O5iXGp/9AtyHX7pssufju+4VgsVvcLJsin6hx6f1namEOukv+DAxn+ZJ/cUzRl
vMB7Ul2NrN1GbtieefOEXuFUlzz7kwMf6vRXBNf9CqVXZCh317rPCDCN7wuOBSXvZXscuG2o+c8+
EFhaMERR2r6BwTMkZ1/MKqKmmZXxfT/i34FJpAr5P3KL9fkyDDibQsJIKwZ1n48QAjCY0PI2TeKn
L/d7pcKxR6SL9hly+92arxWShD4Uw4kzVEIel5GwFlExvtY8S1cOLYEiFBLg2bPLxw/Qpi9qs2YA
jymoRDWnQq4k0QJehwr7HoGMkWC+7x7gKwL4/wAV7G5Jb352TZuKD7vh0TRs+7i0II8KDwet8zWu
y/Aar9cUDFcucQ0kVHIVeToidn+U3lslr46xcPr2ZEa1aqBjeQKBvZtGN/LbjqSB43/+rnX5QdaO
wqisW0pOASLF9ONa4OTkZqwpyLuoK9OpmZqxTe4Ncw8pN+CZ6YaBKyJ5fkJal2+uJQcHzSGnLFgn
Z/PZZnHpGAMaw/97dbGCv/te4QAgOi9maRwBx5AncdATGmhLgnWyNqg+l3jWEF3z6D0lSg4rR43T
aaJ+uMeQNXN0lcDN4mHh42hjaramy0z0P6Mbs9PXGsyLL8jLGR9DCT3F/VvNdBubEB/Ljg6x3tZq
gf1MM3U8wG6bwa2kFn1n7JGRoO4i2gl43mjnWz4SVPuKn91yR7B094DZFrOouH+vGGxcmlzmA6EX
y5GZEK7xKBcgY/civb1cU99Xxq/bL+zDq2LQYSGDvDpMe6NQPfftXTAjflxd+7nD4MfEioy0VwPi
uz2dfTL+LK3PbIXkwmBi5wXVVokvP2M7N/cMGZRksG2ceELUfYR7uQRF1UPUkHLehTblf76OulsU
R7Q9Op0RxP6MYfQMHMcrR2C0QD1LXzPSrVM1KA5wHR3CqaVY+rn0zPEAlDF4adDI0JAxSNYFpDh6
iwNa9GXbfvNRcIBqbj/AeF3l/JkEJpgRecbZGV0GgRKn7qEYl32z6HET4fgPBzzE8Yv5Gd2btiTH
DHwwdecl2RJn5SiY+mL2teHtYTxPVBm0QxWlS28avnGWFGZoHII1q+XdmuZtMATKpvq0ox8Ymgcs
S2f05UlGNpIdOfIW35cs/F2rQkBpzPXOraelWIsfrQaoBgVd2wxp4AzmPSabJVuLdsZY4UoTxQpD
hcOnVRxvnxki78OZkqUD9RJKW6R5j1EvXMnTmUlw39Ph3bNV788xyEmN70QKAL23LDcKOkWSEHmt
jd46QrinTqdLbkLr+hKsiMle4DmJ1V/iqWD0IwEO8MDWpUFiK7lmQvLpJbS3gu0MjtkeAzMjn0jW
mTnByN4Le82G0ATdgDG1v7WLbFBFtJaurlQ9LX5xKz54r9x/nAGsd3LcinDK9UhdUoXU50qS0S1s
MGrSCJXDnftoYYAWsAZdwkT2sqbXE02nOTSNUm0RjJ+1grleqEood5GGxhQmHGeFpqwGPQATVCk4
pY3rZ4eePqdfLfn6s4Kn4uTwWzfT9pcsN27UmLlgcYA9EV5NbOAlF5ArapB9VxqzGG47hPr8u8zV
QHwD3gK6ZGjxKjIr8hKnFAmaMDSWoC57szWB95g+EEKbHJNAa5Ai1HiC4A4On7hebrSAzDtW15/2
eqwSdk3j5FH+0yN72HQX84NAfqM47uY3Hv2S8N8LZRW1p9hFAg1KRwNna93eCgfH/MkR0BsNj7SJ
1A9147+nNxKWDLpi36ZjS2KuFWqQpyNL13g4uAbTsU/WrUQVaaoeFXlarjvLnW95HmNFnuKhx1ZV
isQm17h8fpLq4wgrhJCKyR21mEd/N0TU4jFI/Odglb5nAZ38wYNRgQsnB0WGjeW9KW+XmJdas+nV
/DeY/WLtWGPQm3xRGq58gjB6EqHTqcRfb3/SZi1cmEGxt1VSovWHOMpTfvOOTBko1axhP8MYj7Yg
QkvZ54LlziCLdwlEvREhdQW2zbdCoYfmVz+Cs3VyE3evUYkaohXEwsyAwO111BaA4EiEDel2lSIu
a2/kYVMwhE39fItl//DBiJAhzweJy9f+n4KytI6SH4bJ3d0A1cYzuS14EHQqbX8lfvvH/oB3f9S6
OBnC8LPhr5M3eJZmjxnb9DbS46c6VNZSQALKCcBLpPFCGpT7GnaXdKv2sfryqa/XVthwlwJ6zaM/
ewQrpnj6ltXIfJWntr9fAQmMXwace1vqigf2jaSE8HNhgF5RKb19jzyfGcf3pFNzhUaf8lzIJtEm
kb6kWyF8P7Cfx6QWD7aHSYO5bY3t+eQtjJh4Xq9GcOwR4m//QK3PnGzxpNyIhPrXdPJtpydmSSZD
lNz1AC6HGw+ZYvHBD7bU47qNCcCVeciOxu0sSd3wnIbwIlR4l6kvrWJuN0KnF9HWwA34xmd+QzHN
MFfRaOGg1P7LODdZNOmtzW7aIYM6X6xKNtLPoxwxeBamsi7CFIl0rtBUlMPyPrIf2QK/0hSoBWZM
i5+1FSlnBc91TWG2Kf8THqzarzW8rOek2DaPBudGUqIuY8vjXg0Y48H1CCSyqj/N5FCMcbHcZ2AN
PKeQdL89FVkcibPCRdtxGoXy7L+LLp5YOEnXfsZmA8S39ABT1cLxIOe41FUcquqTt0BR4tkqah0j
5mwQ5SXApFotLo+uFx19pm0CDiXDwIP9G4n25G6C/DBsBTLraF8PGzgXR8IU+5AHOpXzsKgmXwFr
xGDeSHLzIlWmFwrJqPYulQb5h70RGt+zjW/R66Sv8RNLn3kiyMHUBvE8VccilYvN341OQ9QrAFnp
+PHAln9FUiofciO9++qJQ0WINHCmIU6uvHZK252/eKbZ3AXkzHUZzHVcyd/k5zpoUJTiN5QQHITz
r/7VsXq+MHL43WfwIbN7uabAWRdFmMQx9OO1yU1WaxZOdRidqlQ5BDUbSF8vK42QZvNTgcfaHXRN
FABHQ5C2W58zOChugLxlnYMCSXnwwCxDSVsnZrJHpAB7zh5i6rppWQoay0+HBE6wSwL9yH7xkGQ+
TCX3DpGuKy7AGY71WhRG0oVZjvahcYIHy7GBDW2pGMGmDDbYKScSa21XBGbUBJxHs9HLyVjzN7jm
F0x0fqhlYJen2Zp5QUPerWUr072kkQSadg2IuDjUQKAkhJAqj0O/hQF/9AEYatgCyt4E66tu31ga
ZILcBJPMvlopIBxTGuYkJReXPX1LQfYGry6bFjEymy1w2poZuNlj/w650eFOR7m7Yc/YY+VRQn2H
0EwhaymnOvDH+Rvh4TTP+q08GkkDJ2sXqQXHmUkcl7WMd8tpBMUWBFYwds57GRgDhDWAtDdsTVga
+/sCdxTWnCI3KxDgg8YkONKcG09bBT76ldwnAJZM9PC6hXpQlyvmANWK7wIMtM3Od25yi/OmKs3a
uAkzA6af+3LAPMCy93WHekFhJ7vHlfJ2DYVpkMPMVJRujZda65vlTr8/k1a0Xs0dmGk5jGEwpDwp
mjkoWgG4N3yJYyfxvYLnLGNoGLsyDH7jMARKa20Z391ZvUzw8cYEhDBwKpMnDSwkieLzBJKoP0rw
w3gK3AMhHnw0VyI0VBs9YQYhSV1Z+Bj7gtiFr0x+tK6jg/afq6UTnzECPEY8Jmf4VwEVfTNkbJSu
uZOni0aHnpvziAyGKAo5Z3hUFvPxQXnh5DqoZF/lgLmvN63Yk556v7dehE7ot6KGqQQNEF6azoLx
+AmeF5lj4C95QSfIc1NTv/Q1N3v4YgbnG4ooY0Q8BRfV7zxUP6LHL5zO1K2pj/odmk6B47QpkuBY
pcJ1DzVJni8iERiRhYGfidZvDao7Dg6oh+a0gobOW+L6l3Kya0ifte3nTJdp31KzMAdAR+ogBztC
kcgh+ISOIDzaSOu8TxgCnSfHQWIt9yvT8kA/m0t7nNlLbv1c+Hj0oYZixuCnv5UhLGZ8CPe2H7AN
60Xfyr+9BIhtx2eDOq5zT0ZIv+4zhDg8qe8HdLr3IzcMYsUzZWOsYNvbIdo3SzFbPcJRe1tHr+yC
D5voWjKecwX/saf32XFLW1HvD6Jg7jYaPRNX+KGlqXORA2CkjQuTSXfO0vASFgrB1Wufi/yWF5bj
Demxic1Ew6W6G6nhB2acFBzRmbrAFlKMpG0kgyD+TN0tljosO5guPV3vlN0e7/GvhoX3m91ojUtc
jsmmjJf/xqmEZ171hpYx2UEdT+/93Ok2buleZBqM6CV02X6pEmmQ4QKFDZD2TsPFpPr5AzBVSeKO
svhJVXZRCxLIl6UXTuY4znvYBDPsIxCNamskEjswZyuTq7KY3B2rIx7sMa6/hPVrnnQyYuMMiL1L
+bnAhfXZt3vBBVHw6oIthncDqhcC8XqKx/arwIH5kKgsLZVQZWAeSc5xoitu7pQcjKljgWbs+Ku+
WnNK2HqGZrhZe8OKuHWzOpeptQu7ULBDIMDNIWSmRZYR4iskyDGKg+yVGIMGOAL3L1ztgy/aUqov
UvWQqgRAyekePooUehFVSzbEOFzhezQL5g3Z5dYLHGDfGJTzNlBlZ2p/0259mgaQYLn8K5H+QcN9
m8QkIg3AGAeSLh/lAclsSC97RVHJwIEjQarD/eOVdl926Oj9PKiyuEvAetyVpaXCkxmuV0e8cMUC
371HKepz/9B9w1Rd0pid7uHjqpD2WwfuMpPB4DXNN9XbUZqpm8Q4ooOxGi+uLh10oJ2vurUe8MBF
/+O67HX9bAvKCD0PDKq5HXghX/BQKgX3r62xwZ2p3luHO7TmRvDEtEd8JSEHDKnm3VujQw/b9btN
t8qU9qhpgzzmGDwY7OLWfVPWFHJTy97wCvdPRJbItn4laTK3EqwsEs5Bs6/BfjvKNo7nuR582KQt
qsg3FYeikGLWsIKslGw5Jto5zygE0cHTJEoAk/O87vZkbvz12wvuYTlUMnBvoc/ulKCgBfG6T1Lu
xvK5GPdrT/+qudd3uy2XNasMEx2tCeTIsjL7ApIFBYvAW8HBi61dXr2VDRnvovvR4++jnqOgnj39
FhqraxGlW5Pc565yWLH5HuVeYnv1Slax1zbCbBLceJ7TJ3xBDlkV4dPkVcb2TJSNglNEp/Hxetkp
IG6pF9XhfbJyERoOcYdXk5mHipWTwPq/EhsMk37AC6/m06KQqsG5TwNluYLSziHWcLHvb+CLCLrP
jKjtiXVMlGogIClXkH5cJGxU9wmztU/Hz84Y53BeoFB4AX/hquaGahjjPDR01rOA1Ye8N5gKtLvi
k/v5ccltjqM/ebhHEkmz7QhI4TVEeZY82xcx9rv46LghdnSwVLLOg0q2pB30gPj6RZ3R3sgC3SA+
qfn9RLcK/y1ltlbBRnQ1NO99FBJp46rj7vJZuBZjDHeV2YSKPyyvuEgZ4+EnLnzNiQdD+Ke80Ez6
49F1N/BHI+NCB9W1g0YWivrc5bx3hmY9+sLHJxB+djCPQeOwHk4vthe1hyP1qQVSTFMfnH1fUk16
+QFT9jsirliEZwdakAM7/wedOrBQ6g4mD1bE/Kkwwq8WxkoGohZOVRqEXdYS5uowQlEgXsaBShIB
QYNgKOXJBbZeFHfc3jTvNZhzth12iTt6GiE0CqHM+Xhd/Hmesfw7Y+87ewkJ7wA92me0mgkbmZxC
27P+6depFe6ydcaeJ9Tw/Mi05r7Uqy8ZaWDXQuol6Sl8x+B6NkQAYIR13/phPAvSK+W3JjS/DIJ3
P5w94C+s/syyEynq8AohG53JrNId8BHcfpwluUc0vZli02s37fhjteU4qtBpYbXg2EhozoKO14r8
haKjINdf3wT3WYgxTz36EKnbVdSqz/3ati8V0NfA6KxAyuabPTH47ni6cS1orsPbJJm4fm7dPpl3
ABjhp0J4cQ+l5dShMs7dY5Dy3FFrEuWVrm0IpP4UTDo2HS4rpZ1uSR+B9xk3G04V5sQafOB2MGWh
k6kmioiooYfbHv6WQILncrCq84bs8pRYk4aMM99A3xgtYDlYVPInOSGzkVTsHGdIYN02ViObj/Qh
7UiqKSln+Ap8MqdJ9RFDs6SSwDGKaFQ0nPT0OJAi+S3pgxslurU4Z6iP1ASyY6bU1edG8xO+hmXS
jfludaPAfQAGDCkdC9+yOuZPsMXJFd9H7wszYg1xoIeYBuM+Ev2J879ox9qy7+IKuX/EV4FgC5p+
L9XOf9ObxVQFfKong0bz8tVYWPwIWct+Fm0bL96SNfzuyv2aLJfsF31x6GV1sewE0m5edwlk0TOF
3tQiA67I2CNOEL2sEOTtyPQ2oeCqgqdcFnuzQ/XpFaBhEwo02nov+av+6x0mvYwR2s7T7DofuY3C
SGDXcDxFqNqEWH5birbnJJ3lRwuUSL+q9wXAWbdQVoXDzwSLA0Mw4UjxeDzasnPGpmtYBnyFAvQH
V6z81Go2Dl63S3Hrv25opmJFSeCEvtzKvIb1qjAtBNkxtflSCZKB/Ou24zhtarzqlj/B+Jn/Ue/p
vFFFuZ26bNYDKfFmi28PBCpOigryhzjyCOCS4wtzem5RfAyyxWEnTNa50gBUBopoZvHCy4PrTr32
RFzXFtvPpe8HNmzEpz6Pq0Oi2KShkZNeLO2ItJSa8TlneF+v+v/CwnSc//6gYeas0p90WeV7Tb/Z
Gt0oi7qJ9M+X0QI457Tw9LXwU6awe1fywmUYoUeYgEBXcZrlB/CGMtmkgxazGxeOOIl2jTZ6gD3u
uuUKfAVGF+BRWRhiGgHoN6VKJ6IV6YoEFea8ifTeOAGxK/x/DHwWTgd9nSrMgFP4brOLI909cw3Q
RnmD28rhsJqINETuPKM5ibolXM3Cn6ovRCu+cN5bfyRJHs8OvwbnSchi78NWN0iZjQ6aHtxe9r0g
hBY3NW5xo3w3MaCI12Ogw7bYMZA2qbyvvluAzlhB3q8ah4oecpAjuKBMY6N11ezYOWODw8TEglKW
Yt+bCP8Jx+FSFjDPxM3pHmdgLbxjx/yrs6edZbjud0KXEwdDQTLPlAz1g/RCXR3XG47zm0l3EOmu
Kt6jfddU20BuTNe0JVL8MGT7Jh9tf56OAGa65jm6fPUVDQHDM42ua9w8YQnvNVjjtfx3lzIVnC3/
P7r9qr+ypzcrwXKsvaQo6FLkhWVsQxwgB6VylrWELkLdabjJ+D5QIpJzAWhSCWweiIHxo9OW23RF
N09q+KO8KjxB6mPSYYVpGsLHsZEnWbTSKJOYUH0yZ6wk50GwjsoMwjoaHZHtdHNTEG7WfRxfecIo
BrklKswOYci5Wqzxsc7ap9kDGEu0E9yPhNGes68ewJtF5eoGZ8Ad0A765t76+1KzXFmCSTapBdZG
Sc9GKuGoWAXmEq/BwEbSsnisbPhJoYvz7Bm5oglE9G818xfBsYa2/S+CK85BT/Z3uguG3JQrNn7W
MPEPfz34bDQMCrfq7LoEoiyTsniZprK2sEe9qsCiNW9E4sNnsiSBH6FbBH9e9RJMtgXw+2iMveO3
RgCo7CoTj2vR+14UKHjwYu2nJuVfbrYGLqR0AY4CA+zdy6K2sohAQE+BlTgSI5jgTyqBuBv3obAV
HCUDIm4g3f/G57ZNPl4yF9ZL5lPOooe+ZI2zy8ZosU9MguxIhZgfyh5Akr3firG4yde3jsyugWC1
MIGtQ1evTC+jKAOtHqxAJZmXeqNGPv01idh7397I5FQvuxlDtKHA/e7JZMblijaLAy7OM/y/9FJC
T/ISgKZcRiFwAiHG5XUKHJcATfml0ajz3nQ4HwsppLn/DgqUBaxIDlEI06y4f15ClxknYVH/9jSz
9DIKP1EaM/RUWywt6PbRKHj63Ao7Giqb5+jJ/zsKccGF2+l/Zu4tcc7OH1Oddd84kJPhjSvbPod1
fiVRrQwb+x081Bry4GJNmpuWh5M8fXoYMKt07Zaam0qScBA/hgenk7xXP3GqpEmvyPBPBAvRCjxj
wCMKiVArrQiQDsCywczlIVL89zNds8099/dZoyO6YF8k4DkpNJcSyDxp5hzLPD+829wkFXreh337
7lotTCy0Xo1H7sNmWtBw1HHzqsKfQGJhYjJ6fMxCtX/anBO7OPJdV6Q+egMJF2fejjSJ0XvR179Q
krVZSlgzCgf/EKnXtVcJ5Ftn6X7kVuo+TWI3Rrc/PWEWIHZ1IDrwzHap8O3S0nPlOJ7qsorTyh6D
J5bjzRc4YGpY8c4Fb9t1Dg0Pm6Oymvsvgb7K1XZH8QgJAfqSWZHyPPsd9xjfLvD/yWefkvsVuSci
UmSNSkdSpALyhaW1sW9FInFZRnxJXnRKsWO3m8Zzk67KKQ8CquOiDSgcF3uXboUdm1Fimk/UDlHn
2znOj6++IF86M0xRcpMbDQWvLFNoJUzsONCuGv6cOhKuAATLFJHqbgrIH/NAYfZquoShMH+XpqWn
a/kFRH2b+4hXLTj0rB8tZ7JMcaS798MYJpAMvRCv4MZ8OyU7SxwwPTvSY/MZ0QnDDtGpYHoyo12n
RvqLMdwlEvmO9w7S6AnBr4KGPVimnU8ZeNZ0tSDUEKODDzAHamAGi2qWMqxyc6/Vrd8CHntLGUEU
0PJ5dmamHbzUrs6X1cdagAtC6MbObLYqoGXL1tLYz6E0j7FFuEnjY2boq/yIOezGIdsOfxi66jrg
XlpYbafKv1QC2iXoi2FKuu1gdGMRSSDY9tslBFL9PIciMBObH0J3nAJ5ruMV2LkJZPtBjnZoqNdH
CvAIf5lzKORz1SOkzxjPCFLAO4aVQGzEZRnIKxOIIDU8vy3nWd3642WukAqmtaKmwQgDbAfxB/tl
o72woGkVBp/vFZtB23qitwbJntIx57Q0hjhdflWvXLlj2zkb7drsIogO3jS2J/TuayD04lrwzVwr
wY/+qLefIl2TKXiXQgwNFrFIH80fkY/8855zB1sfCYjE9fN8K4rblu2mEvttBTnC7B/bacqZI0Xa
E/t7gOVGLTi5kW1+NocjooqxQFKf6Jrwv4DO6yeOgghjcBtUjTxHs8EYufnCQONG0TfM3jC2VZ/q
10LAg/CW07SpZNHpu/ABNplKPyE4cXdz9pCTYge1sVzIj9wclKECyk6uwMJL3GeTce1wlTogt6IP
lzYCQAi7nP275Wicuca2IvgbtfckLBuIZ5Cz4bkpb2R76ja7gryJ4bxsRzQNE5POKDFrOvgKwm4B
hpe9lUYvnUplT/SBgRY3w2bZJm1E9ye4BmIPiGz6fDFr2WJitSWSi1OBXdA0zQw77rePcqacdjaI
dc+jd1yQvkxvUct2gGDTwxUMyetd3Npi8D5WPXcGN56K9xTVKT38UxksycYw/EwOe7XYAkc9GuLp
dOBsX5gC4PlAVqPulvQc7ZlQ4YRAI8zRmgTFSGY4APx8+E5ujnaAf3UCU0OwRLKFee0gw9NhKRSI
gL1SLF03nzfsat6S6oReqE/iwNUlgr8XLg47MHVs5f0NVbXwoR40PAKA7jeYkV9T1qC7pQhT/SLz
C72q79OGD0xCdhAOraqoGdNGMB9FKwsCC4EjXrfB3rAKdQrq77GLifulfelQXqOZTgnviK0qPH6c
BkZZTbLkt/oRXtoNAHhgqvslMF9nR5qu2DYgiHphSyHGl73I3UqlmxVJZJg6T/knRK9k3c6zWI0Q
VDcP88h99iXg2P+1aZK+Qzu4qkNcOjtrFlfJDNTqnun7jgTq/AlUQ9Pg2cWdVaDwoCAfXT+eZdHc
q9ipof+HOdDbO3GIwJUCxEKZ4noL3AVD/EBBJB23Dt7eqzEvEs2s7wjMBulDmQkZsF31BeYmhOY0
Z50Vyprb9/FJFA33d/lZR0HdtVQZvx8FIaScIvw3101wRGevoKnm+cCerRCJ/XF/WUQAn2hCjYqA
ojdrE66yHsp/dI63DHkLKSKtsDVZoZonznkBRqbOj5D1S9ZWr8ZqSC2MMsgFkA1N9PbpRXyo2u01
rdIS0QFcS2QFOfmQPGEUQpmj9AsiliX/BSbK+MtGwTAS4MsrIPDAi5PxDZK94Llby0YKOYorpkrC
00S/TwviJWaj4LnttbvnEttYMUM8GMA7u0bZHKo84Kt6wQK4WHepuDqFwTTBJbhlSxY9DOp9g3YK
2330WPPujsFAX5bBU/q0WGqOnd4JYqtNntP2vso89FlVcsncD8tgsXyoc2pRDydb0Djv6/L+4owz
t7LxsY0hF1AfG9ncT8Eq1eMXzWvkQYIXKpJWO3021mSsGB/l921a9NO9jqx2VD+tNmcsSXM3ofy7
80zZ4C/sa7LrawcKZLwbfuQmkdHGROLDiwaVJJb+wVFp79BqTiJYy1KSZYRdwSefXirklJT+JqiI
hzVlwtJnrcW//jFnhhpXu8qzSVech9V84eSLQu2smjKyPd4hRCwiniqXjsE0XP31otmIxTGi7Eug
AlqkcMEZHJomIlvZxPdXVfF4viW8J2/oQOZ4GciuvzakIb85bFpj2a/I4Hx+gHle7ggMoC5FQ+hL
R0Sspdf7SxK7B6/Uib6RSV0glPbOHVsC0U0iAtDNAiKWuM0wzi34727/OFAjEuHiSk+DyAyJyXhs
cQyTow9um9e9C4+LLEUYkJTVzkey7BOmKmI6Jlkeq/ltTJHiMH7Yv0q9VryUZ7sdG4NMVNuTF6zb
h1+cE8R8xtJf3tzzDBTpoC45vNGj7CUjz0kgRO+9YjuNTmprvPoep8o6MHH9qOTFHQdl8A5EI+aQ
EZ91Om2iznt+KNBU0sqB2v9MOQR4MNre1ngapQLCgLQhKbqU/ITTgHhBV2XPd7MmB+cwRadhG0cR
LA3ua8blYhUFtNGLUDO5iH88UH3XVqAOV6QcdTycPTgPF5JRYKzkj3etcpPQ0pr5279JqVD1M9Gf
hlIH7yvps0MfrLHz0Rs4yrrh+pX87l7spQGX9oUzLiDYinM7JDYzxjeCapoYKpQNTMnRzVYJD84Y
6n2BE4psn6vxtqduxOajxhUljZPiX93B1KgTwl2u2k4JpQsBsfmNE3C8KeAyc/whdoQ8X5/dspno
Rbb7tYLdieUSRTctWCZsU3sQbiGPQyCjYTXsbj/FpsV+porXs7or7P+vHBUPI72/XdAhWoDYiXyy
j0crA6+nI4eDgbI2HaCAY1wZ9daUBhi/jS9WKIXhv3q4Bw2uNqU2iVS54MTh6Qv19yFnv64Zbawa
K8QUN2r4tUcBpY0oC+Es/cXw07KuTTTxj8LOF/G6amoM4TwlRdPWUggFrlqSkDBB6MUX1MIEh+Pr
v8h5JZgDE4MT6BxldxClOZICvdmoWVggSx8PIaL0iXvbjXfNysvuzmuEyvJGQKD0O/SOXx3hl1PW
4koGueUq/aw8Sn06OZcyw05nktWX26jRqM2wklIsPAiIC+JsQCqHB89LDDABolIGeOM9ThVORnwS
3e15DcPZM3QM0+u0KrwiYN9xBu50fjNGB6bKhcLUcM2jjkcJ5j+LziMdnzOJXEbHg4+l/kF/ZN7b
rC2/0QuvKpUwE66F4m/7gLl+Q2H4iA6R7FhcWKbQ/BVoeOan8uP9mM7tch5Vz3AtP4bwhzdKPj8A
nYNMqMT9SH9vY4AipTQIKdwf7MissxudoS27mhCRlAfYb/HT9qfovzogDM4atO8KTmLOlbBFz1vX
o/0nZZ5vNPlam1JyVSUs91RXYIYtHdonuuX+cpNhxlk71UCflnEZlSuZ6Fo9pHf7v1b8DjzF9pkC
uwKJ8Oq7MAO1LgK24++V9jYLw0vM4Owi9FD7+B3JiNd7PRp0djMQG89Hbs3di1dhr9/0mAYBMBrQ
DmrqQfXhY0a5ou3NUow0kTYsWgSvOqv1Hl2NmjjUko6gNe4rDl820TkIxJkf+g69diugCYf43ltD
KVLFQeX9QXb++thuRP4EFwteFRVQdqzGuRhjrtoztc7ZSIMs9i7CxMUsJBHGelOZ7RyRYnA5XJrA
1kenbjkZe8WxXtctK4qLbLtT0mAx5zMs2qeZDpfAg8oryMh+QmmEJ5pq0JH0a9WPYwwY41VhywS9
jzuvxezZSXiQpaK3XHmSPNGOEhbgddJuz4q7syu+yEmjSurRGHY5pKTH2+UGU5inOkv9n6Wv5p34
/RDawiykEEr/M9AOXO0N/1ozfbSpUcEelOkvBmWFKbHTEDnleN43ithHvROxdxIIKRQN2cjQBsre
lT5f1J25VrTWf8jZoEDjBxctjtV0YDewKwdl8CpR5GCjneZO2tEVpX8iFSfB1QoW9ZpWnOHSWKOF
VF+NwPf4fR6Adx0fafJgBVjqVSWZZv2YEbRYRCuoXl5qXQNcqSVk1pfuIFvhP4+v6da1IBxkhYP3
ZOxKN1g+NDEFyzfp41uBNIaHPIW7AVZaRq3uObXnEYvDlVQ3eYmUo7CkiDZs1gq76SMEc3g/fM3j
4Pi6604dsNcqcfSLheFCvhlG/FDY9/k3F3O8ZwfIYg05iQ/x+7U2hju2y411O44Lma0b168oHlvN
++j6QxKlODRT5ey7MsULbdx2yjbe0lK+n2R9B11FwcAbm3j5RuVK+0Z1Dd4E+bM5EFlx4DQJ1ssg
A+0lz7UCbs362bp+kR6oZ9T7mq/VQj65lrYUNbiRiIcpQqvTzTYdx60qcxQ5CdC/yJZvGwf90ZuZ
W7gmEoYt9rbiJDsCq2cc3EHXhxJoBhOoE2c4Y12+IJW72B8BAIuG1O/ntKaDrbz5AspwUfV5G4u0
TJ4VyCzdvaBSDjYh4yTmvv43+57Us8AeNXbzB9LR9wNfPD22Dn6X8k1Lgpfi3J45pZb4ueH+u43Z
kebqLeEjmgAAZgpkuBtyfKkLfssk1PLWTR5hIJvZqFisQayCDm43Dm2OMmavfLgkY8UJGMLzKxre
7Dn1fFdH3LwrOaTkkoKpqpnt3D8Wa2i352AuaGfJSDIlUR+DvaFi/zgV1xtSXj9HJ0Se9MLM/QWU
bXFkn5uK2cDtBLplmIP8ipXNQgH+zz+egtjkqcU4q2YkRmnAZGLXVo4vWj0sKTJIDOkobOmJauPV
JmHQQ2n/WJM61dhqAURxPACQjju8ynR2e5C2ld99ZCBiLj1V3wneghGOktFi3/37sveQyg2jb1/h
ZutpolwVNDHBqshTPh453ubnfupTRFqhjGpHdgtj/Y240rXy97F66gm2CFHWkU51DFYRPwQ1Lwsa
xUZ4WWZTQzB9ptl+AsYsx2/9Zr1tcYHSXRb3SjP71uE+EgfqKkYBgRyTQ8DvVu2HcIrhoAfaVtQ5
1A/Oj3G/3GijEHwrJtoyqW323TnwZ/yWeCtL/79ZTbsYQ2/7FWoRmACZ+hEgS1IpTupT2oORgmEA
92SUdsBnIsofMAJAY3ABXt6Uwp+uKJbS4koGqf56mpBlAY5ymr9Il+WJqNM06dlBam6F0Qb+fXiX
K/rAzuSw5hYQRtjm+G4HHZ5fhCAGZ7DnpsXxTcLMsYXdMXYOIcePxahYkcJ3NsGXJkxzLyPNKniQ
LKpsDSL4QCt282Y4hejiVgs46K3JLWpW8Y3h4BGCe7YsqYrHFPbPLE18laAg82C2acSIa3SFT2E1
p5gkZhrgqXKzGNYfj5IE/u5l4z69L9CnPE+NlLLLQywSAt0/VEBdCC6IrIC2APkRDrZUV72SbviY
XYzlDOtezbnGoiHWilyTh0V+mN++303fgSTXGEbFK3hN6xMKF0mU3HW9iRoNFrHpKxfbugf2gYw9
Y1HL6fse75JPAzCFv4Xi9z8Xz0tY4x4KXXdLN5CdFFyKTC7yblAA3lomPKZf0cyNWs4YyX5/GIjO
PgLvkLoKU+Ag1e/ZNXDKZ9uaFECqBHo+VpCqf8L2L1V35K3aiTNTV57c2FTGSPPGjrqcqMZxq2xe
tDfTrtUizubjtuh3a8gjprSdO8DGpgrZWpYdgWC3M9y/+AKowidcawlNv2CGRS0wia1k2FBBhoWa
6BCjhmtWFCk0tvTg19NHyERfuX/xYp9+O6FI5dygFtXl9+IHeghTv/ku/eUBCgES8UE9GN39yMY6
WEfQmMtEp/TxL6aRBJnVQig50+dmoSy1gwlHjos+ueVwM1VR2C3vrn+g57Yx/QHMsITgjzJCToHj
2Of+U/C1wPH1RDggmvc02R6TLXVrLrh/dUgmgogASDDh4ijOwAB63Ww8Vxz08lv2iAmddmOAWZaJ
HoRO9ylidDFiV17YBpRLV32XPiqVU9+r9lPAueifHhB+CPEKLYFr54TEJvKx1XIMkfRwgzJSXQ50
bNCPArqjm1BHBnD1FLoX0VzIrqBdcrFUanh7VW9PIYZY5nJDRdCph0ehmByfp6F/Fj1fn5PhzMIY
a/eY+uZA8hs2dQIaJ38eImGOP915oVwhldyS9PAVVWrAZZT3CislR4hreidkc2HuuOkv0uT6fEnM
Q0GKoFR5ymnyfyZPNhpBMVNjF4UJdsnrVB5qRkBFkDnHQcbbWo0J3TAhG2swyhU8Z780vGWmislH
wyGk0nl9oUzLg5nGyXVDyw9wujb0Q2wQkRvLL9gOjT17sOWB4OppGi+Vm7fUW30ZRzPv4c+yhDf8
z+u1QihRKuUTfBNGjRvKOuvmZgTJx6orxdL7EdRkMNk2tspMB555sfQQWLoywVuVRx/638RIcaAs
ylEBpCnv344wbwphhpRoWhl+eXvvI+WzOGSZu8f1d7Pz3PzbLB2aw+L5B4ygtOD4eRtd1q2Xyju7
MQuntYyDBXf66hr+bBqgXLtkify1sb7sv19S+Krh8MAYrHM38X7b/TPT2JVzPnRa/H6qVMhmklvS
PG1qwv/R+SHeUpf2pZEZohWHdGeFao9L8CkbHc8ecX0jhDqjN1b+usvlKalLesmtqdw3CMYizeX/
8qTixeefgb2BiL26C7LYSMgSMpmqr+tFlZ/iiD+jyumvDP+wM19P6czmcnGcLeuThrR7L/2kU8/p
KqkIsZ4yD+goae4dwHc2UlmlKXX00k5UhqARyhoQTunFjXODidZ7F+DHo15ivm2SZjWQwBOaE97x
piPivi7kH2BJXN6xNJm66ntGBwXnClMlr7/CWtjlmBT+zZD6+mbTNRv2lrRssnsA+kSc8X45b4WJ
/FTXJzfGHSHT7NgYkO9l15RYiMgAlzCskunwLN1DYL/pAKVKr0zHqv80xacya/OoeY8UaCC6kEqS
LlBC22R5YfPsTEeJjdtGsOy6Pka5VRG/fH4S9SB5RukIgSINShioovpk2HT102tz8GjBryOblikx
w2yCgOa/WJOeZXgLlsKWtSf0DlfX4xvs5GoOdDPteIwEDImDffQze4uoMJaLtEPBtBNcP1OMLFar
H+LkGGq/seBipJQrwnstXoqtpd4210b4Be/AJvI7BbYlt2jZAoUTw1o+gfwuxhZGSmJSwZbB0VYx
gR22CQ78n+SN2dWA3thcQ16W/Nbu5Sy/YT6jpbOZvG7Cn0YMvx1424D+LZ3KuG7G+c+SCuAt2Lb0
Gh9VBmfmf9Y9outzjYXqHw7IwdnTul5VN+G5tMhD7lJP5cDYzObEZUQfniBwh0+dyGkCb8wFSjVQ
zEgOxi0/maGaIGGMZr07QjJ2lHTO9plGlyK0hHbPKpDwbbx2xx0/etMKu8L7hMk7k7572hiR7gRc
H/EWSRWIJx+wcDytJgk2fu07Z3AxbpvVQTZQGBALoiEXQBxRJI+8PYBc/JHsgnUN8F5WY7va5pEO
CTDOCLYNdmsIAVPnC++cbbmQ0SMcikpZZ18QildDNvrRBqnEPc6jQ16mlvwAIS7bbeTPbnSg5+7Q
YSLzihWVVzxNqWQ4uIVOydYhsfxzVpzXH5Tg9XMuD6gRbBgciEe5PwrFZAaciyk9Wj8cwYUEcyfm
hmcBKYVDw8WmcpUdyy5hOVTOa5Wz+9j2CZpMlLelAkLNDybxZtrluu/4RtrvZvIwNr4FdMqvwdtc
NDkhv3khKGIG6crWoDOp9K+7fdoRr1WN5lRg8WeFDlv3cfWZwUSwEAw7sdydou312dGY3AYxF7F5
PU59oCbaYACls1qzPmHlsNfEayIFd9bhr5zKTHXF0HcIr5JVRh9ZobpXaD766ySYltSJVAIbQT9H
wgmjfgMGFQPLBAHcUGFmW/ZOrUViB52a4N6MR6PF4x6E54KePt0jRFQjbPkzqD7HLI9pYvab11Rv
MeMq2OKLV7MMisJBTcLTSmrIkLHz8ByJAbubmmt/waYA92un1cCmPw4DpTzIQss1j+hRMmCB9St8
JqOYFRPsFNKBwdWIvAB0pfM5XTR/yO+07mma5S1Wk+H4q7jFJl+hNjUMdltvcMpgk5SKEBwb4P23
rrf8W8Nu3pzXZflc10Z7/eC36MdYBmfStg/4iNbmafOz8fvrI7sV/6pBi82HBnvK7xxebIm+3gRd
ABNW9SR9xsIbTGjIHfcvBtLz50UOXbm7XxwmkIXh5Fz5M8/itmSj3GAdCAxkfTNckfZjWseaAaJ3
mQWrDKqAWDj46+zoUzFPVJj/BX1SJpno642+QGagoTChnvP3LG5CMuMWOL3zV45csJp7vdddSeXC
TJXXMwmAZ7IVNGUz+VUGrF2P5MuGEqQoi6EzBZnaPdyf9Y0w8mpO4qFh2tJXPViAzIdirOtrUlZZ
IJfLMVzGY0VGQw1wb1+oSj5vt+unigaDezv04bWLaZDqsb6bwdSc0bUv8cLFHnOhn4gvooBkQwSW
El2nhdB6dhbicQJH8X2EaTab97E8B2/sDYDc7JNUcUMYzPi+D59fkzTIQr2qUB6VNT9/cokmOY1G
nh2tERiDoq3TKTZGRwh+FvF3cMOAwqYxKGhVPt5n4vvMhUFMow31OVkf9JaDrkkHg0BnP8dkjO+B
FsO0+Io9W/ZgVSO7FL+wfN5TBbC7ulZw2s4PE24/H2eux7gg2rqOCjd0u2oTsHuWILgWVXUm3DcO
9lw1Fr6QFBEzyPPvBbgVD7/zcCkmteAFnlSr0fo8j0HY9PsEVNwKLFcsNqFpAOTppgG1S6jpPUdN
oh9GB9OwqyTKldVJl3vb44lWtrRfHZ6D6jvSY8gtztbeby3PXOKjyHON6efPOlQiKWNaZ6pfP6+x
89SDbruCQKCqX6DmzHkAkjn1IfrACQp04oFa7NFabo7IFtHv8+00UELJIecjYIjukyiM97cwr+ox
p38Y2CkuxIIWgx9aBMLhnon1nSMJRZfUx/mr6ZOPUzbzQXiKgqad31gJfbouK7mcjgCe3O9gls9D
PFmlfO83CYgLlHhp0A7tBwOUTritLbFL0I7n1MZln/aVnElm5wbwE0RE8BsUDuwRvPyfRgfzlNO0
GNiHRPOP9Etq78vhhzPX+EaLST0w59Lou7lcKDTbkDFuVRFrdlEgwGYo/fURemG6W90eZKLEIT/K
GXwwaj3XZnuop9/SqKmpqyM9oomUw68iA8IcRDF7GwUWRqhZHPaSopTSFxf40UOyZuzuwLIpTTNQ
rsHFokC4ssrxXCPBBbe7eImtI+9AsuVuFdVk7QoriIbrRpCkuXjF6KmSXmRSh4N7F2F0zaLAQRZ6
wFc85tVznLtI2oCmgayNb+nwQV5VF8z3rHPBPvETsxEtKgtfUtQAm5YBXWS0jqtFlW3lZFP3/Z57
oV3PmVdpdK+GQSSC0CHQdQqcqpqn1MXCPJzVt+BsepBRlcP3SjuW2gFpe132Soa5Z/C/BnzSBDpv
YRwijU5qGOf2hhbXYN66ZbX8EeODBl8ro/mu3WvHduAfk0AaMUQK7L+qCM+afhrMwGiV/y8eIkNu
zaFatG4UNURZKPPOHnlaHeAjVPFQWCEY1sLzZbyBP7gaExmmVcf8calgeNVIzWzrfCIqeLPNHNXp
ajxxtvF5Zoq4Xx2DV3nStESqQ8VHqOxGZHo+pfAjPt323m+7qhiGkm6nS6yNl5lKOIfqkeEkGAF8
zEaoOYLNh/hiNw3BzrM2dpOIT7TPmMzdjD3DgbRdAk1twUTmJ9kJ8yE0LG+DAUBsP/c5e+x7YPol
VEkVeyagQJ4GCyqfd8xynurZonUlJn3HvmH4+CkqBzr0Li7Q+PJt4JRgoA7BRJwYkhhCdGZw7iHJ
dtJnng62qUh2GgeYnvnNySyzHr4BeD7mR2EL6m5kRIwPlK4SnEx1l/1ULn9aCXEo4S8YJEwB20l/
6w1z1DVX0zKfI+HdNcxZ+akNBhWmFBnQD1K3yUiKqr8BAMIoxKkhOKwFBXrhFAjydXf6D7pS0TBc
ihJ/Fm58+p9Zp8et5/c1/i3g7pYrhmIYH21a2Kh0evEL/uP4NiD6qfOH845tCWwZeuItWK7xo9gb
GKL3Ui6d4MwLC8p8eM1hnaSAxYwmCUVEtaWR16TpOp50fsgMC/MXAL8iMIWyDVL+qafz9RWr4fVD
/amSL2s9ALV/sWm67bNr809v+6/Hcoge6PiaNNhZl0cVu7HuJxekRVFoDRFcwnv5/YU26nmMfrN4
n4fYIvduaOvojojrezS7XpcZUrbS+gSpifsrGVkUvXShobVVl4/0jmhAUySdLTX+3b8csJ3ShPQX
J5OMroo8pocFE9Gb/+rWpxHBrooWfyPX38Epfj5KsW63PsWLmf8HsLTOkQVjgPUJXB9tRJg90peN
ykofX/5yTG1OOr6vfpTJLkYZVon9MN/TNKQAjDyQGDiWNNaZnuHi6LrL2vr+MobQqWqpzb4DG6Y6
ZbvnN5NwH2oT8/zcwBDZFFEFARHwUxsuesBhvxEyPSLx0aQi5fOGo6aMt/E4DocxQiE0KdspBRdq
Uzb7iJTlqcaPpWyhcm/iHHaDi2c6wvIr3NGYYd+E0la1ix8Xq4xmQPbunRzf8ribwSWWJZ1abdwm
rr7XiBgEssHZRyxGKn+Pw+XJgcyq6+lEBK4u52syyVnGBUYrxE/tworRCdH0L0Z5ZodlGztfV7ZG
H74GCqUjPSkfmZyhDankpyOYvGPqorStztTXDogbdu0aoPpvNHkq6BifyoP5IUqjpbWfemJBfnP9
cmCkltgfLaAwHYHR0zmKdNVt4xb6rwTxXXV0gRov16axnQxZdHbIO2xBhKcR5dyA81CJGcZrlFNy
yZbt4wUTu8TDoQDBuEbNpMG4uVwAnfRc0xxyJlTjhLG7Eebhqr6poECeJevfuAl3lcXc6BghDjQn
tMlU5ttzjlmUzEWU6hbJCAwm4JYcmizGyBDmg+nfIWI/NS/YYxbQSo4LYBy24mlGOXng2ajG77uc
ox7HKhEOTu7utmplDgGYxfGSHtMAqf5Qyjd9twE/6gk3epMycWbhssFSUjDw75YbSaFK3yaA0kIn
ToAq/f840S5CxlMrc3vH/2CAOE0Zr4Qr8DqvwvdImNzMnonaPR0tEYLJ4jXxnxDxmL9Y0pr9Hjdf
bKPPy3Gm3Ct/T01sBq1ciFVkONhIhLVoPtRrNLljm7tofTGUW7eDr13x9XjXw21YqmcJ1ZFdiURb
YxNabmbEZUOLujq3LMXvd54Qcl+g6eM6W/cgy/UiNHO9ybTVhcZJyLSrQ36ML2Aip3AiX6vbmnao
07EwQxlJxyG3Xyu75wMDsFxYVD7QidPGZXgBEvEtv200WrYdKdUrL+8bSVFxr6tbr48bvFdQ9Hc4
1AEkLKG71Txo78cKm8R+ZGLK/Mk3eESktQIOz/QEERFnPmpP7l8+Cn03BRPcAlwSYTTGaICnZoMT
G2ky2ZYVsY3Y9kUFTghjkK7xxhmdUAyDJfDbiJ3yWlGgaXH8QhazMQRwXB2ekAMRFfWy+afIBHgQ
xo0UnJboUqlov9ayvyW0CW14UGxY1enMoHm/k4H9cscx4VP2kk/jU1a12V2DEeRA85h6QD/wZFaU
UDcGgjQ0LG1dQ/ChSfhwtFMiI0Q7AGP9PmD2s1wezY/RW2I05UbE5NJiijWPll1hgQrpFFmerq8u
j96C03vx7OPAoUxaFF5jbBsDDUPoPzH/8WRWamabFfeLj2vhU8LUFtBSivLNfTtYdcOsKZtzW0Oy
Pd/BwlQLVVtjr+1HS5Makl9gxPkGzI2ZBEPbPt9vw+dnHyvPRNkfIoc4nNHprRUg369Dtk/IWImD
wNCJv7EdqjL3y3A0Ug+aNh2MTOqrVAiyKPYByebUF6FI9M6kDRvIqKMiaHjMpHhs9oWyyldztq8k
/UULbe4XMTht+hwjCfk6EqaTW/VKsv3vlzJavQTkum9fKAGtwtansaFUxLmCczvu+kBHEjaAqy5C
PSchTZXdWgK9NaTc6Du/Zov/Ga0oKyR0V2IEraqZBNbMadzuBspvgIFzrkNoBcvdkicrP2JpOe/M
saE+CydMrD4T/lhpzR2wVekNu8N6s2SufbOWfExLRscAq1i0+1vW5s6/VNkrBomhrzJ5OH5IVK96
tRmZp24VzhFhrPUd9OlNZconW5Jmg1LiGEa4CQ2X64nRra1OIQXuoViPhAztyXxHJrMuo7EF33a4
lAVEev+ZbTSdAnnidQ/xjkTP04DCus1eVKgFa9rwbJQ5e+Z917nU1FA1NmQi583aPl50cJ592xEZ
c3aGW/QzwfV05VvXoZ0I5cLFD7kfbgt5b7o3QzHINKr5DPXfzxVzxBMNqM7cnqq9sZzoIdJ0V/JN
nUPjn9bB2E4WuT0+YAuHUU0fhbhS1JqSIlRNsvjffzIvdT4F6EPoNr6iqomfb+F7rOvZNnj0faik
UOAbi1Ua9tTnPCSx5fMRycZn5tpeWZbvd/IN6AbBzyoPfPofPvH9IlcqN/VVo0G5Becsf1zXOQqu
XKvAunCbvW2mpDeIEYY8LEPpFqg6pQrrlXnR687FYShHMH2glQcjDA1V1kvgwanPqBr5UI32OeUF
vAmV02AknKLItIIyb1dzyWMXUM57o1ROgE41aK1OI7yI9AR0oOpDPevetDWQA2ReZ2fszvg2SkYU
VOfYnEFbHQc9phHi0jiqDcY2Em8YL0KhjC/GOTgD7TdxoD7E1RlZDZRovqgPmOqcr0+dHR3hViW2
T4CjjfeKv6na4v7Zx8Q+eUZz2yLIvK+DNmMPfRpFlzO4kr3gKVMmN9ZvWO/Qrf20B+sfONkiqfk7
BW7Xx3Rma18LTeZyoe2Yc59RCDcewKASra0nEGYW2TWQm4FuHliABBSvETSqYtJ4cKaW5NT7sJvZ
oLYf70kQeJ6ANbc0Zj72AyryctgOsGz4pnnNAyTgPt9VHsNWnneLtjC5ZgSIDtyQcO+qds2A1MUa
P5t3agmGjq9VAVc3k+zcG5p19km6gJc7mo/nn9+sUke5/fjaxQAMNKFJfdkocOURSJQFZobTKicv
f8GZ5/JgL881rNN30iRmRXGzZzZMXYJNgZzTzx/t30kEhrBP/DXjsL34x0vfRy/EziMVnAVlpAUB
kr82ruIPZ6oyzltRhftMRsucw2TlY7000NWUqplQmuhsFJ2IxgZE8TBUZW9oHYu1B723sGDfDSNC
dIiGLPxYNgEHIS0ly8MsL0lOq1IwV1UeZiV3r684tgDeP+TXOoCty0ZZLC7Kh6wQ9+aPohx3SSll
bBmWmeUA39gdaHhUuyRamBt8TM5vt1GEbfle7lAr9ER0EbhpPl7zJWntqi4rOQX34uG1Q9N+89L7
ui15efd8/EiympIvE69bYfNRteLp1yoCbSeSFFH/9DR+ojYNtxfKtAGLbam+2yo6Ht2w+V/y+FOY
kHB10TcLRTJKp/xWLbs0EKexNq72SqC0PZOwmI87EMH3yQvAXdJ7VWmxO/GwoJAbvFzI0tPZD/Ge
MNs7sNcsDmaBl6rWQjsLQ2VXXgNz4cxJozWN9hdLUSjQW0MxazTiIk9Q9K4TqT+aJUN303e3Owis
5E5HOrYU4GH0ug6lyGFlRTFiSTsuH2Ff/pnxQmyLzd8tC0pAQI2h5MFv3aftpZ0TqKwPeYdMUHgi
aXrReAI8YF5Z3BjibDhqJPZnZrEJYrZiJPR7HkfWU/wSzpxc93+bz9OFjNsJSLF4fBfSU7Y8cgUM
cw/cBV1j5dXNmRHYYwJOk9UT8uQpVfAUcBOaCC/hjTtc9wp9icEKEoogTGO1gRE8Vq0spqhMB8Dh
XafiruAd5d6zLBItmdcoKakVaP5o63XJNNnhiaGo8CDJW3fygoAet2wj6xN5lsCn2b6eAma3jRbu
xdVJurXNTKME7eKhwiHewzGjMEN5dMyctzAIsImoVCb12NKgiLA7RJxk/4lTsVAHfnX7DLs00tZG
zmhjOm2WBtTRsrBvzJEULIeOX3QyrnpxJ6iUXn9nNJI+wM7wT0tcFANuhLQdvzPIO8M7GSUbEhJ9
5IxUiJcxaOBDtsF6GT03ka0iDQTiU2106MRzR2YAsadRFOrvWrZFN4+zBAwkfiu9knEm70nTdeyd
inhdIsiKcqNqgjEcuCnWRDfxMxhXi1LiCHgMeEdhWvAxMeA2AplQUvRSh1pYJcbFn0PcnRTAJWMi
9yaxw1nTw76r8JjpOEUHtOW9aygli6wHLqbL1PJnyRF8aGVoRLiIHgHzrDpdSkcLOmTICmquWFM1
7bF/HEhpMBMMsZVAGgwaXKpj4CgwPQVSaDL2y8WY7MnhYqty8jZvhxZ53P4E4p0kVdYCcluXFWcG
P8sCg35XOE9NIzeC9iKoU4xrZBrjhXYde5OghKY1o3tqq/dcLlQWXiffVcCjzDoBKrezTQcSXJQI
XfIra0kkUVybbTCErS9+S9udJyoS+IUY9vTMnLtHSZJfbbJWXmT1ndQ00YYLJ9JWElX1EbAp2c2C
8keDTz6LmkRsJvlIzw9BU4jOOLL5rxThninzCav2WVYhL3zymTzd1eXXZ2TM/FCENg+1PjzcSrv7
IFbQHStVo//ETddOvh3IFMW3bLxJ/LKliR/xPIGTE/IZ5iPUZFrhzJ4EnwjMGCWB45pIl1OzIiug
Uh1wAIrC39vu0CZBp9w3pZf3ckpEJXBOs+bBQc7IMxTax7rFRNYEuSK6+oB7UgHm3xDKfLgoBdrX
2Q1Mc0SnmJ7LRgwDgZ3u4KrhECOwMChLDeoCz7PvFPPsvzkGKFQ++mSxT8loS7nAQ50NRwKlu+DQ
wcyXZSFLjuDDjVLWBJefqdurSDLgOIsEO1LmrZLtCI3TPEaRL9wB9TBSIqYfgQxNkG/r2JneWMSu
BnGXo7w+yBRDdoLgSramzQjnNs5V+8E9RGIBUYgjINpkHm/BJIg82x/IjSFnCrBMa0282VPfXvs1
rQtVogGtmwq56zoxXk+qhlW9uc9g7NdSdCZ6Uh8Gt3mGw+kREw1ZdPiwCJp4vHKoL4g0wLVGKe4x
1PpncZ/rC1gcVpTTBoi3D3bSFOfYm7bJzylzriF9osmxEeAHrxgXC/+JGD6ZIxwP4XmLfngCqzjs
G1zot3PVn9Tq/XXe6TwP7HmF8VTDybF3gIJjEM2dLKzuFnhbd+yt20uK6690BLlQqjJ15V1a/SCB
jbHQsZW+XhgjrZBpuUPKa4tOmtazVGDaNWUiXTAqCye2Fbogw273SjYWfa6WDJkLy2v4q1NqYckW
2d8K8QQWWod8kVA2xUt6qyQZVrKS/i2M0TuIHKXzBmstBpzkotEERHCR3P71DDv7q5oLsbWngtSf
Hs3MbvZgFtSqD4Q9zmM2XDTqhR+eBkbDr1cTVQ/qH5plemPxe7yEM2e7t1JmUUNHZou3kx60vPE7
5raPuxMVuZsDGsSzetPr52dLPwHsIArGQgG6DER/e8K+pV/NirK8AYwPlVuMcp8MofPTPQAfSuPR
RqdnYsIV2sTrnmnBEIYPWuaoZT5Byl1+cq96+3UPv3wEae758j7hAgthlB6M3oGTI/rHNGlf7TKy
OV+epDmg27thETBFbhLFto4IhZj0d5Cxud1cGDCEJbv3NJ2aG/E1pCk6DIDnDPvWFDrBWVICkevB
kELk172inPTWOxrP5CmgaCwUvMnY4L2YqBvwTJb3EiTvhOWEGxj4s7Z7UvBFZIemWaeUWA67QSq9
2Pm1crf3OKv9YOd6mV6rM4eWeZrKSEddC7Sz+g3lWNfqpqK8PoxZe2DlNy3jh1WXL1S/R6ZzEfWU
MnL1ok2oQD+Uwpb+Et/ckTeyJOLUPnwRoJOItxD0OFZ8kdpfsGwazc0rF1aLY923shw8/daPE+cs
9sKon8atwimk7xmF3YhTOOjligKphnWMlJEYOQc+Q74/xg+XkVecRJqvTz9TBPMYsf2wjjh5Jpgo
tsSwG4dJBARNFd0JE6QNo5u/qNxpZoK/TYL+dGteNdQlErQK1maD2tT2Z/itAICwjGqDgDRj8QB1
VvrWdn/0N7+sw4AxYF9pn6A7CWUq4qKfuLHegYcm5kO3a/cmbJoeTTGWo9ZCKtCPUm+wgj1EgE+O
SKeg7CUpdW/D//q5bpmkJ/6bYUd2PGlqtxoZZTWShVa6f1czkpqx4wWLncgwMhkZGEEku6rPdKO/
oYjUrere6YUkzrtansGz1lbE+/EKWpBzTPffZvFhVe/J4Ug//Yy0sblAFUXWyXQQg2UJOwxaYdaQ
i4FPsuTRHtlB+UaJxhpTgwn8/jGYye7H+4rD+o1DrlflnQSTq/3QKLiKxA8g29vI3Ometceu4okg
bauV44X73YqapDBtjc3JLPrzY5SSQHIKwxyfSVDP/S0iWF3JL3CXcze2nt0Z9Immyxb5737ia5Gg
s17uWkCkvrfBlFu75QKxfenIdn8AKnJc9G8Et9aKVlf1mQYy9F4/rSoBUQdsoIxjrIGbsh5FZWNp
xlSQMBICbWL7TVNzhrwfUPsL/lK7Z9v40clm7b8DiFEBwpHJ6kUcOa3XCkUB37JV1GCVZ6rDz9IG
km0Zh0hr6/kkn4Ng/DE3/GaUrxrzO15SyTlOhSUYDm5PlKrjDHEAfTDCThxSP6L6W3MvIt6ulx4+
SBmF8IqKtdWqEu/7LmXdwDpWust4+M4Gb+secHMl6++O0y8ZZINA8HX2Vg4K3g27qwXe9bC+CKBb
hNSthsKI9tlFrFs6i3FohulNB6ds0Df5ZQNpySv6YCm4052VU6UaCQXv0SB0wqiteSmSa+Y7jpi8
mHl9ITVcaTZ7D7WvMzzKFVzfWcSIvETkEGD65hzA/kyzPA9GTy9a9Cfub2xs8zKRlQs3y3grQ/fk
xa4Fnv7hp/oPKyoMoU8EyPQzVe7Mmc88tXh2QxDuCoFFWyFnC9aRzPH/+uWY07a/0rJQ722AwrtK
nkLFuXXUvC24tqXh5RJGOAduJEvcGvsGWtS+zYuT9gCqyDtYMugYgMun1ir7uhk9h2hh1F/Wrm9C
b1kepFoKWryjpzdKzTsECvXYy+Rs0n/pw4df+himbx+EpY1whk3x6f21f9oA/vKWJxoHwcGRy0fP
ConA+ty70Cq9JRGsztV8/VsPQCUeChPRlQYpWDPWrpra8wc4r+yi4B2BdsHHmxe2+3GC5u7JMBDb
Us3urzvH38bWv702I/w9izip8+FZc0K/CMCmEBZKSLqEbAP0CDjLptWe1h5NQ1ryur9xvu18W5jp
X2U2PiDA5f3UpVLTQYxUz8NW7/t/3vz6pU5T0QUSotCrWrzVeRZZeFEeFIeDb4JTXGbMPkGzjKDQ
pFe5FHzm2cXeSIR5Hh/xaQMFTh7yR0cQuWx2WOwtezd7xjav+mzcqj6k7mhTd5RNGwgVv5ZBlIP7
dtEbFFpwMgthQV6fYeiHP3kRHQ7AODxqn+0RRAP7gBtJ/gYIOudNEekf7721AdnfXwRhTdF1epNc
VnNl3/lN+YuI27ikOR3GB3ycRZSzQP0AJ5cxQ3Xnjfc7YT0aTxmc3W1Q8pZLM0dOd6bK9RBZ1LYv
Ildq5CBvhBAe6nS2MJxCOYpMAh5CZWmrX+Y8m55VHQcxflyOMIN8L7GDk2D9O0leEOYK8XcgJXdz
BrkFGbgRnr3Jgj+DQBb+/a8X/bjliwgKE4iL61+CwSBBgb07wMW1Bz5UgWCkw4OytStwyvkyJiVV
tQf5Y++M02dHlDC2PXEXuuqdz0qDbxMTVD6qJyFRtFhJm8CbPsWjPgZkNOW43Hr3dL35zXEmRP4s
pBFtAIzDHmRfidGNWGHdE6vfA3u4fY8/wxd35LrSBXWUKrXK3A5vsHnP5jNh8DVp9HDUmYnqMBFF
03aLZub/NHBV+PUV8iYdHlKDh++d8TINrDCs0gwlj5xdeLTVZXWR3VSGN7y0BS8Rb6fZVv7v3xrZ
mor11LkBZiareiLUfmJ5+UWd2m0UQhewdiOMJfKJvF39l+eWHmJFtY24DNw5Tpupf6xE0DaGUl7m
rWsVZ/Uh5vZaJwCSr4UHu1138/OK8d/gpaNXeyFcDil/o+7vcp76xC+MtyM3QI6oCfrLLy557tL3
XKuEOT07/z2/8nuOICKZVtUlhs8qvkEKv+2J5sroJXqismNwU9szepDgyf5Fd0M8GDxPaOGFpOEH
EQ+/eFoDP/jFaBVEVL9gjrAf08K48tIZltK7K3eR9mzuLkkw/Xmw8U5zkLaiWtT3BCYe8/KKseZD
qB6KXXq4iofH+uP/wUNjwrTSQ0fRntz9XhQN5CbgMUmLkyxai+t98lVd11c5SRdgVU5af424xDxy
KIwtoTa/DVKl7LR2xm8eMbjjKKgI7YSJnUz/2NHQQex9OInZrtqx9FQNs9DfSjbslSOLJsLpOV7J
YzsHca8AkH14HTvKAu7p65SVklS1y5K+NFIJT1T4WIEto2DcElAbY2EzyBpuJXPL69JJAuNQs36b
S8BhKl8c6VspBw4NKbbOMf1BI7bsmYdWpEDFyEgnh94TDO3P1xtuDLQsGY0f6T4tzMla8PqHtukx
L1ly6HBohmfDj2tIOVn8Xva3JLOH3tyn+ifVkdkKrOVTDENiyNx9KDQi5Byxqhv8tSoIf8ZCHp5Z
iyMG6mcuGOKpnbolvToRRlecXGOhutmcsZP4kO/JFiXl8kC+Z+tgh+o1cMZv/cH+Tkm1LbYciSuR
wax2Po5MpPuseldwKi96GTdl+8IPCVVJ3WLFbqp4YpQtOSgLPqvUW7xhOlRwuTjAvUEXoii/OSyu
uiM1tSMcZfHgl3mMPzmtar12Zmj0VPqpE5jhBsU9BNfEaHIh7XPvPL74kVIT2v2iPlMY5kRXvz+1
67uOz61LaZXSTUp9Bt9RU74aNpxSRDI2UkBhRqSrBEKnw0NCaw6HTm4dkTXnEG8AMxWILLte3jC1
Kq1tJ+Go9X3p5piQohp902p1hILd67thr9BDMOto1slbA/LNdO5oY274dK4jB+OV0GlNW/lLEb9R
8ujhj3Iua5J5bBaVHrj+0FpXobklW6vZuIGdhDTg+InR7VWbhH75bIcgFLOaErR9CJ/mu6/A5phh
9ac0ltLgI+e0JbgSLg/QL2BceSFnaa0mQCidHrhZ6dTNmTpbGFcORpCq+S422t80WIGfjrycge3r
Tm4AYb28kLJNuCmKOGQtF1gDPpQNzVyG3gyFOH7YZqp0nDDajRWlbURsuN1oA3K0Fcx7Y+L40uSZ
JcYgl1cUVHRiBLFX70vAZju6FMCzHct7Yb1xqhVi9FUOnmAQ52ahLAWqrg9I7MPnzNRLd8iLEeij
o+P1sN27v6Nu0R+XIxYaBDjDGb36u+VtTGcSQZx3OrXH/bd/tEKgv9bXSkZkHKYp6s6371BmZDTD
bGaICi6ERl+UE4fbncsxTNy2s7koUadx6mgp3srgAmcH8Crym+VlN7/Krqk41Zm7+ayyhStlJRcB
Jg2NYrcjTJaoXqOlSpuB8qlYrI8KdFvrJlvwJ6v8BxnHSrEiEeQ117OiVPIHDK1FuKkVfGNRoPhe
hbAc2ZkS49LsIdxErtvWscD4yoLyge1vcF428Wt7wHi0x71dv2aD6qc0fp30HpRQL7OlpWFX9PFs
B344dOLt6c0XO3BqAYUk2kI5YNhECM6O6rcC9cYC+6/NqgaNjEFn0W4QlCvakk3lwd5e1Uc8YkE7
33tKlPyGrg2rUoPRdlKA43pNADPyCXV1Wnho1bCHPAS/RcGK0ywhvgCL2ITm83FmEnDVy3RuP1Sf
Zv7hqRbEJCIM86DO9mAyaLmUTAkR2XFej8XwPy2YWIdsv8rzQLU65Jt3/euGVUsrxlrbcS6nHzWw
+b38q9bRAVzkPCRDFNHg1DHbQbs+3eXutMEixoMccVrIwMxh2zJqy9TZaqEu52b4EiD8F7xvfklm
y7yLE/zSsp5ojnWqOjScQLKRigeBEdBoElCvcmYLu6fhwvWv8LYWjX7Xn034kkQgwX/osgt3SIC0
1BdJsEZh+vFRkDkqObMJ+1J2+2xIH/IuHcvlb3dR1fDo4XLrmg2Z1OvwnVttUetL+v1jozRYrZsU
AFOF2znJH7NI+nnqKi5NgnY2dLRldU3FUkQKY1MPlNqmegIGQ+TvAB79S8jmiKByse6h6gMalG0P
qIwEfbOvW0Z5QyxQXmUeV+O3wKBuQQz5somKKhUf7jD6XFG/GK2KLLBTlBpZf/6WEobORWaZmiBU
5zFXUofzgdJYqBRXPfSfSr62Tjfwi32++XQBQi4NPVo/pVDYnsd3UlSDIL5C8EWq1Aa2z7UdXxg8
p8tVsAa/UmLiPtDrYw/LwMw9thGch2wtB6/VOnpJhXJRkg/GFIpoiEQwUgjqRo7LNJ95KLNRcJjM
guJych3LwlGeOmLj1jycK/s2ltrCgSp9l9T60Ph5YqfkCC+dtAWDaJBwbYqphGFRjN4FcIZaStjY
ChFyfUt807lURqWyvzPLUG/qhn+ouNIXtTQw/TmU+3DVJo3k8+5aNR67mYHELm5Kj71Tx6WnT+ak
/BSCwVUE55Um+ZNXZW6P4kQVsKYIziIbFG5pY+iXUwR0JRdDcWj2FaceQSrtuR48m/9ppEirHrpk
1nxtos3/qBsNFmaVxc0cQwYtQWMtsEgIoTb8GnTy1WGbnnqauEo3qaTVoD94YvRWOOm5AkEGeKN7
ibjbe/KcNLpbBKnx370QQvXALUJJewfki7uHDFhegY0O4EbEJDJKNPJ5F2SceR7mwebeqnNGx/eu
maW2hiprL0/0g6hMzenhrWaYJSjnOtTC7UBU4NK+16iR8NPfumKWd69Xvlj7VbKNvglbyw/JH78M
4ybC0UhMcumCdBNoQ60syC1bZROmGwEDkRJ2vCRaUbI6DqFqtIIcIgIDWKdHuOWhq4dHwcULxRil
XPjTbGteyWYj3jmZE2tmASoYuRQ2T8Hl4/HAZOUiKjNz3brm3wc90WUJmQs8E8LLUXRR22OkIiD6
WtBYeQjUB0vHkdjh8eFeggUgGnhUqurDmtnWugE1J91w2EC8HUaq6lbr3HV+H9j1GMGjV3UuSzBe
ZQMMhwj6pgvdY5HfZCbh1pF8Qt2CEVgFDWWqwDW/f1wYhvmVvrdY5HXAVqiJ6AqTd8QFapqzMt0T
GQ/KFE4/4HuepJnODU1j7Eu6a/Dc0KoENpgOGFYwV5mnHlgErWxviEMbw+YrS7sx+8dIhcXBLm2f
zbZNk39w5L76Rn5N5XRCTJCHpa1CDCAoT3hUFNS0TQctYvfZPscqOiXauJLD0bcnbXAR29ayTTlp
IYTy/bx9FO9CpOmwADFiSO5ilclePtMr74JYcoLFArZPQKFDJ7s4ZswKN0kTrDhlwydf9rKtT84H
X41qcl9Kw7NMRP8SYuY/s3ABnJOwU+mUNwzpz6qy2YCPr6Y04IU1h2sSWj3vDSsSSl+nQJxeW0Q/
LgjXOBeKecXtNLcrRTnBCP1rGAypio3sMOBgRvY9PMkTPqHsGv9vSpq0tjpWnJMeEeoIFI9E0WYJ
N154IdsEUKvD19bpqCBcxt7i0WWAti6tNEki21LZ9d0sy/Hw/Vq2PgTyjOEm+QegMfmzajhoo4nX
sKUdF2DTodLUeuq1jkFkGufwMJiOo8ktYPfHL3v3zeVHn8pwUP3oXAKF4qn8AbJ8JUC/b3vfxd4H
FrLF0IeqkDtI4RLIUbjwERxBsB31dBLExSXrdp75IYZR4Xp7sDsYySkSuK0ZJAnU9BQmpRqLy7Du
za+j0od70otQB1u4AiwONhdcJOgHCepVyKaNVPHlIxoop4mUAqboadyRope6zRkINBc3RR7xGIqS
ed+E5mrC7MMk2QLnN+TK7RcLIgWs6i3FO0qYeXchIO8YpXk+i7+PhyPLcfpupW8iYL7Jb6lPdxiy
/VHeNUWPNYVW0fFRJEagHtmhorNe32cOFDLAGKDmxnDwUrT+PEYWYi5tG2lk6Yv6uPZmonfrE1aQ
f4ueuFUJvvDcVAqKeTSF9DXVeU/2KOvVHAs0dsvwNRzECSmwvIKbsxM39M9fYBt3sfX6DEyYcP9Z
EHrr7N1qFJRA+RYg9i5aHHhbPviHXvIguGjOob3YsUNuVzeXwuvGupjKj0kfujcXQp6UGn7Wj3U6
np3jo9sz9PY1LRHXHlAdjBb9oeb1adkPbHUl+u7P+yL4xsqJNCyqX5WMbf7N1ZrDwvGBbovxZk0B
wo/d4kGvnd0YqxP3z+W60gP/hgfFYatzLTk7BUBI+hgfLyea4ZXD7QMldu1GfNgaFxab/gOWPvWm
O8j2Q8M/wbRwk74RAjNDh8J29J5PdvtLDYXCfz5bYOynHqkcnapqg96XeOjqsHGvvleVdsbrjv2z
Nk3thDjnAWx4WiZ0Oiuy42+x92yIDIrVBMH2510tSkZuHuxendVoljRBPlMC6ZSmDmODH3+yIO/s
DOBjLVWSs+vVRFVWD+Ug0n2B/COPvPPm1XyvBawXMiYuAVUQz9R8H3HZV+sM7ORwo9GO1PXYjr72
HGrjgCK25vedun2WR9zbptKoHkv9MeaaBnIPijhUWyDAWWeXdFpzkPYrNz1hAkqjXsNnqpI4dk19
XTSJbqDyPHb5bAO03VqkId4efjSzgKsORqRJnjETWAaGmdJmDy8d9TRCO0Si45aFeTUKKdbXn0qK
VBTVLODFaGHVln+mB19rlQb5tF456EFdgnji56oSkCxqNPvMBadp4EfCuKyRF8elzMsmRaoWLY28
cmyno9h97/40st8TaeOyDn3yGmcFYIWz5PUbE52WkSp5TBdb2X6vFGz0iHs0298QIr4BKb4x1jeC
wi4grBWx7COxJ9BvAciuscrbaY+yUKzNVNNzweTtB8s7mVvj10E4y+LgSYO8rUn8eY1OmsXOA/Rz
nO8puN7rEy7dpXKQ6ugk82fgK5f5tSJTtUm+M+RPS80AJ/fe0T18qlo6ihQDTIwgttpw6ZBYNHmp
hIQ5+kN8v6yyrIkOKwNGL8HEQMxikvMCz5jWd5Vp73FxJ4ASxnD6rbA5NZsfAbIAk2FodeG2mlQN
g6eHnQM2u1Kd8ncxOwzq1brsWswYsAiW5488rFBtTChMA9b98CJGzECpprmeslOHsIxSOiSoGHBO
qObySQUaATTU6uqIxTjiM983iFP8mRDwnnBtncE8PTi8yutsVlTHwBu2px+PQyjawv+zl4v9CVvA
PDnzO9Nm3IfB4dBnoFgmeqhdNGidsVAC4gBKoKpD2ig1exgBiU4JMUMrd6qIe5Q0YXP3a3q09ilv
vSInsCgYKr5hZsKZuuRLb7tiDJ2knxr2fBi/9krUF81UMipgHj5s3dtZlC4gYEkMnusfyezC40EA
1PxPKVy1VrfnduGFakLLrXuY0Hsg1xgQFvg7iNf/DwYSxZbEcoHmVTOE2EXT2LBrgsaKNlPsRAsk
r3y0Tx/ZM6AvKVJgrvvQbLGtgwbm8hL76XOOIq6c+TxUyV30iOg3/TO3zyO5hhtW6UloUEVFurfQ
G9+xRnNDG06SrHDv18l3q0WSaN2N16NnaInSoDtAmwOUfG38MS2XUa9xdwVK1ojV7mYPb/B9p1Qc
xiAfVVaGfQ4rUVVh7pQdI4DHFp2yisshS9ADjqh3hhs1dBhwZGks/rJrvMAADzuubVHI8cU1SZw7
Ruh+Iq6BJ0x8uywWXQGj7OYEDvpVCStDWxtLB6AmbebZ1TKRIabPeaza5lmIawq6mrE7QKoi9JLU
vXYkn4L8jLo+jRNAXOsmRxyz0znUTUXTnELzEBEcxHLhpYvPx8FobGt4+qM56qpVBekdQht8CI/8
VB5UbjZqMVbMoLFPK1PpgwdmSCWhgs3KvZOu+Zy9aJEaqnOgh1WQPk33yRZtXDEnjbx3D0+1tqpx
pYZ84K1dRHba8DTfHD7B3z6peDDWIPpZf2DnNyNTexerXBLHu71j5TXV/nekgJv1/mUG/hjO52C0
AemNjAyHpJ8kFFc1qwhWluZixwc4xPCbZP1T1556/8BhuQK41l0R1fAxmUPD2Hjuz7JF3nO5lQR5
CvGIoLWwFKIypV45Z1B8w3c8axYicR4KWTUBXA9z4XnnudDzrGDlQkMon3kLbDnljachHgJbY4vy
Sedrh/xudgitF030SayOwfQpCenwnZwUF7YrxDFie0nltcMImLLm1AQLGAkptjwlOlcnLlV2Mruv
mAHajfqmbKjUSCb1JgDu9bCz3QUs9yX0H1rFzhCjdLx7bdjKoXOEg0pqwxfGckcl/5nRdpW9wG7Y
rXbcN0ZAH22o7DKO296whGuI0lVKN9uBuhSYl/UWxR8fQA2b3gXeJZ1Ctf7TR8bbW/lhs4EL4aY6
pZBoc59uT04bBMpDbzH+rCM0bbgWKasIbtRsYnfX23uH5XKHhd0uAl4SWTOR02rVrYdm51VLhLhd
npJXDK4i5rOiUGSqRgsrM0R4L4IYb3laSKlzBegWA7CcYFfj8N2+gVap8uUJTE3HZYR3d+8cXe6u
CwM+NZLVqMm7snwcRRFYi8o5JWjMd0pAgkURNquRXNNuJ3FvjktnE1Ogpf9jAW0v5kZ1qvhafO9+
aS3Li0gBEFZvsZbdLrpJ4qC4XZLWLuLri20Fiwp5OaQ9/N4nzfBVFnJNm8MOoM/icivW6MkbJtGQ
PaZEScou1VACdgCVAAPi+Ao7JR+tBz7tksu//WBOfk/SmnLCqN4pNzFY6HtALyIylO9yMSQILJLy
HH5GVoS1rN1r38qH9lZdqgmKC8bLuFtQH9iDlqDuKwAh5MugBX/mqWtusuOcjMJkxwmIwgjaQXKT
jAEAas7kpTrMygE5KFqC6RzjOCFvz/tghAqrGwDyjXiI64eX5N67KiVPAJZpY3Cui7FXZnMva3dI
D8eER2Wo82MTE5aaYWskrXFVSt0sODrSAHwhuc5KZDu1zfYIqxDh37XA4Jp3ByLdX03C89pPkRlB
+Jauf7Y/hjRnsxU9fcY+iabJN7fpGPlpS8n9AaaozEZI78mlrXXdHdkBif7/gxpZnanAlCxNUVc9
eh3Uj8g9TBqSY2omt6NTzaF7vV/PvDuy8nyHMuEe/kPugstZaWlsGAApqQv66svFnFlqk2Ry5MDV
Y0am/bWjGR+Pi/et/VCpJ+2anPzUBkCRknH2etC/qVQV7VsOBH9PJbpFvdAL1rBaxxpDEOElNrwO
Vi7NffN8Pa/B4D4PccNBwPCHYtZkg8tsglAmSFUI2b5ofGIJulT7lT8g2rVW0H0mVfG3gy9hwxjA
uC3Do+VGdrd8177tW4Vs+9IfnIzqHW7yqfUYq+6p1L1rad7O43huYjoxbHsIre1cTJX0jUbtNT+J
hvSjBtVWVdlOeYBj8dIncRtLd3A1iLL6G7qSNa+IllD/9tyRf03Jsy1BzHPSKRuJqUwEVFQ8jA1J
M/vj6qf9EwelFf+qnzxG0LmccjwUJeExfTFfi8fKgg3nyI2FxnzZl9Bhv0jPhehVxRrKu5Nnhqu5
kxPq7c1HDJDCt1B+5yVfgHSwNUZixadRSDt79tYXFkSdhHEnp6VoUHzDrkMDQymrY0lqWZXAadmt
REWyD5qHvmo0LrAbAU2lE3ZlL4Cvx+jr67U8VTIelmo5IgF7Vpd9tTgrozxRztfSu4O65r7fZOmy
tQOtJAEdygN0n50q2dKPDuCaAv7t4hOcE4xX+9rUcf4jYUmeNlFrkM+z4n9T0cOe+rKkL/VF4gPd
IonIMU97fjYUodApUCtsjMFOlejSTFMbQ7AZIwtoSRH3lzwofsnnaIRKXHlt9h/jjJaKDaeOFDcM
xexT/9NIrtzkKyV1CMSjeUYQyX4GjXWDGUpFGJO0ABKc1jtlyslzU4YMhpzNrJr9utJwl8yp92c7
BVjnauTtwyWu15w0uJkIOcX6Qsf+cS2i3ESYXdjO7E1oubvvosupvDzsuOYZ/KiEq/zzLxZbXf7X
PDA0c90B7rnGHEMg31EMulu9qTjqhHrsepI0Yj9+reVKGpzhAB7m0eaT0ovDPS6vcI98PFSGfLej
Uc4VeL4ZaDq2buKsbRr0Z+CoVQ6mPtX+NCb3RzZHSnIAuK1w5sKAXjPdzhr+0rPsd6qZKGsAAJip
d6OhgsL+keE5T7QxBZpFDJwB1KZbhJ4sIOxN2RRYhmAuHKG1ohrKCv2woMY2myM04uvgGGJtFc9z
HfCx55UTMCBjBO1pueq+0Rr/M/60Lp18khPFNMeExhJFgiUuNQ0j8mhKACPdG/mpXTkxDuU2GOvV
QNfJrdWv7C+R37cC6BTYn6xtRCZPqmtY8tloIZtzh7mtbJGkzxTDQIJQFiLGdK2joxqJSW8V5/0N
rlE/GPTnVykFPlyq9WRuwcPHqVeMsnlKcZg/lZ8w6UlBoIZirRww4hpr+zRs0Nda92gAPaesGKDW
ziMgZuVhCG07uFzxnxJkylATYzGCduRe/LQqXZw21aZg3bBbQaUyIKmW+IP81WlSj7m6ps1LstL7
FeTdzlBLn9tl06kwkZC77u3OpSCQx0EYJMrAHEgerGp0QNjg1L69OUMxzfMcjeuwZGeqz1Gn/fbV
+5+EF4ata0tmLdy4dgqhSszqovbF8JRYW7W6Qi5wB/uUP+GAhFUnrXIMWvlJTw9fnjzgnGeP0+tt
JKRw16/7UpceWo+7VLxFbbEWmcOaKXhfj8DzfJhw3R69CBTGUMJTUEazWHCHGrSgNjGnCE9PVih+
0nPRjhO9OhUfDZsYt1GkN9foHGeEoCdOmAKSSek9ezGxei36N4x/pW2BHDCO6R5UnqDA09FSkEbc
IB1wu7ehOFUvm5jaFdZjA4j2ITj/3AAqo5bQ0V/aYDZG5L8Z1oG4K9h2tYsErpv01Na6AdVbp4Xo
TFHpPuSd4fN9yk7d3gkjhCeqK6R2dKH2ou5W2soW68wOdk9WA17JvXibm68R4CX1jXRutL/tOpdQ
FZvRmiahti3LAZHsJBW0uQCIRS/8iwX/5m2A6tf5oaGjyN6Axb6mPk1AYgqhkF/nKv9PdWVROwQm
j1qsQggSpRsYgW7DZGOrAmO+bXaVIP9NC4LSutR7LRTyfJSxyNx2hfkeiX3VAHmUzt1YFMELKPDZ
Ao3aCeHsCyVhTxYQIlRTdkZG3QQYXzM0tGl9NLK5Kb6glJkdIkQMZ3Lg75wwp6ghFKv6foeDxAwC
k5HC9JogjHPtXUp96K63LbK2yiKoMi88v4HCK28Niy19R3btXwENOiQK6eeFcfaTZ8Acmgw2B8oc
UVShci/RpunILYW9QHDu3hu2puNHE4q9rfT6OdJ1v0fEV4z9b/Z3Qj5fDUGl6cwnRTl8sQpjC0GS
rwf/3VWr2dr+ILzOy4ud7OLyfIdQdIm7SYW9d0I4baGv6ivg7hK4M6Fx8rFQ7LT4ffXplCvewv3N
mFzCkxJ7CVE1Tr0KMucfKfW8WuPGhMT4/2rKCKp4UTGg910a8fwoBljKdLtWXgyYDuyalOnkh/ee
9aoeI5lwAwSlXYEy/kLGrFzXxWHKrcksLrGUoXr3icyQnlwaTHl5mswOGI/qBlUDquIy/3n/zVip
u/DLqkzmss1aThI8/+oduWqRTM2nTmZM9Sj4OUqfGWVL6EnG7FeLAmJ52TN80+FD1a1fRKfjxmfg
EQSJszr5sbLa0yo7gRz/apMJwCPdfQAOto6QfwG6p76e+Sej2i1o2SqvQ1YxZotN3gmdZKU/YMNy
DuVnWnLBXedvpnzVAptWl67EgzO5LzLk74bRv33pFIahyK0VCtSaKsbRxathzo3nVZeA725REma2
SuIpCZ8cCqr73kKejOzVO7nXrHbcsaKhApEbWY8Kn+aDXq5C9Z5pS34G9Rw78tz1BTeYuhPBoZS4
BXxj5ec5iI91XyZO9+mZQ4ck3cSYHeQRYDJKjGmz7AjlxCT+s7k4bnJ0n4WKmErtMvYZmkk+S8I8
GWc4EL5xnQOVmAV5ImjjcYb2KtjfRjpiTAEqmftMuDufiws3GHIntaA/ys0oydKBlu68Kab2EH+A
lHl1OaM9jXmceu3Q2p7nPYlmBW77qYB5CXhsiVhXVAGbMmMa/ZeDUFoKzK4z0zKL5PXm1DSPpqPh
0DuT+auKTNHwZH4KhntJZp6QVVgUnaF816a+26BpENEs5uIeZObP3OUGaRETrZvnDWM46+63MMnq
NUfJmuoXwijVtpeCcdWLo3F2F5ar8VG126P6lhGzZcYmu1J1ROX4GlEyWCQGpeliGqRmS54Q8d8D
+wv5ZSMXTjsImuHnymHfhIAmouuFhzBHucQF1Ah3Fn3X0hbarUcxFoXLg0GKXt2Bmz5uXdZZGPf2
fJkDhXff7qAHWtalw87XTBroI4BiDc2F8R7JWM6+Ro4fOfuUaSMis9xuLSp/3u6NrNhrQaKwgKS/
vCxNiZqVmPcA8Nu6zg/J8ikjABdl3kcxGxv8GcY7P247yqD5PQwBP+oqapzCso+1RWIUGX45nv4w
nJhp358hsbjHkr7NA/rtCxGtnuAJC2rjHSpDN4MlvBv3gTGqQxQf4xttDZwxjjJIVr5/naYA50rf
0XFv55GOXCGjndgiFrrReW3FL/l/boRB8lE1Fxvgt5EEV4MEBiPIQu3/JbZ3PdhcLSL1r084ilo4
wYwOg35ewVpFUwFW+fB3XKRN9t+JVb3P8tWY4DoOwO2FEvzT69GtRVljPUVsrRtQcAL1l7V7td5t
RRiQhBcjcySqg/nYc6dPEzZiOCT4o0c0TszZ3w8TFQEaVEjLy0z+IgfzgIJl/orX3hv02ebE3I+z
lv01I4KUlZl0J4Pq0HgYMyE0gRUR5H6sLP5sBbtFzIYGhLoZgkwd4f+3iQ+wIJv8omVNmQzf8dEY
HtoqYe/OWl3Ziw4D8YM36xmOdZ3gDWPrfUdYuQkMjYCH3pC4vGFsV+/cI2QhtZXwoCDF++J0Rlgf
btvWixagnubKg5Of+Q30LcYmvbQWNgtPi+A3SlD+JtURWLTDTpereo1UmjBbFmPsAKHTjQkb9CbV
tED1vhddAplNYKf6VUwKusnRqmfdiw6JJLSCkozD9GPq71QbSrDvlWbAtaXl3+49528Uc7QIPld0
Whb8Mni9jA/tqZSiIC1aW915Ab7AWFfGulSN2zkmHxKPP1p8KOR3uj/qkxK+XtL5JvAp4acge1+4
/ylimvAfbiStRV+mWqfnh2b8ljWL2o4lJjIwsU/XkM67xtrqf4mKsXmQsA8xLUQpBT002ePZVHzk
qlNt7wYwcWamKRuWP1p5On5KIyjqd8dxYgcqJHwLlfip8OCAHmDC45l6WVSL+BLQomUFmdAOwOuS
rkLM0L69wu2wqtO1Vta0UqxNkQLj3+DX3zT1PHOcGFZtVambxvCyitCv6RRD0MpzqxguY6IlFAQ8
wAOq4Z5p+Qs18LqRwyWX5nZGRfpE1pBtjNTv23DMEhTgeLl6xmo5mmpVP/7MP3Rv5xvPmhLGHoF2
fBtt22D7Zmgd0NsSennTwE08qmsH4GPfxwECqMcob8z72uwbhqKMEY40JBiwp9UIswM1enotSzKI
YZO35VGoCtknXm8Hn4WUTEPofIO/AETB1B9s5zxqSe1BNuX0bOmpv8YZjodVMQmcmDa+MdjS9109
BcNbb8QExiA9wbmV/WIMw7LgSXHIutwnGwunASEYVP6SizaPD4pOiX7xNz0xVcaixEkGiAfqiMvQ
u3J3Gco1nNtVp6AjGlz51Q07z0TvZ8D5YokhuS4FNFYV/tzqhOUbt7ZA/Ay3C3a/aZQFkO/gZFJJ
698A83rHcnbSgQR+BikbQrhGNCAPEp1a0Acokqa63TjAFkS3NAv6XGQvJSJgu3aAoFVBglrTVbF1
8DtuhjZefN9I3gYB1NXgPxHyeMiyrxsdomhl42Sj1Z1b9m499HiMZuFgi7BTzdlwzork7BOIchGe
pTumK4Mp67QFnlIGEzRudYFlWvwJVAI7SaQ7Bd2zn5IAovNOc7ndDVQbxwfSAU8qL3ctyAONVVpi
N73MP2sVQPUrQypDXicG5Favw7S49OcXZZMh3GMLwzypv5FQwnibSKDvMr68HvYoB7/CMMvHG5Xs
ogpU7Z5N573P8uad2ySGf5BKsF0jprCNGTGtnA4wpojxzv+eEI3U9WMY0YQ3RWTZpKjw+2X6ehlt
JWHmixDaf2ODxzAo7pVqH1F9IstbS0UWcUmu/kyAXdVlE+x3JaDgX06KDsRkjJoteN3at5M3Zwo8
XSWAhDGwpaaMRvOM6+nUpXX8Rfo8LQWuzULhYgd2E2PMyaKhH5gGAI+klVu3gaQqmniA1U+QwWou
BbSPEJOpneJWcFY91qowLCAe0zSFGlNubGLCaekXWcQAuzcxbhyUGMoCNdEH3louNhYGoWsTtsdD
j/mKwCeYiO3IFIR2UvxQMmvzK4hITzp8OBXPeMoWbKWjBFMcinGEfgYMfFTJC5v9k3Lc4iNb1l+Z
HZrZQdgC/3poNXkokbCBzPC8F/75sNexWX1FHNmPVHTfkk3ahtxb1fOlqpns+zJESfQYB7FrLC+V
XUMkjA58peeGYp5VEasQDctJNIvf6GQrxy0GQh+eUI/L3BbIH9R5KR5Y4Zc8g/1Y1cGzjO/Q650z
1y1bMK765TlFkddGsFwHuO8Jjhtm8Mr8KmC6Jfguwgum4bck6xEMCcj+l74k6lmePTtAXiJMOdFN
hjToXZpPxJN9g/oGjpaG3jT3XEAtmJ9iAAPINFnetkTxDsljS/t/Kmbivxo1faUZAPf3bEfRoUmC
07XYnM+MwMU2GrJcf4uq/NDhNssE4NbyUVLGSpq8TjGbe/Lj8vrFqLwebd8Yr0qKdL8l9YF3wvZy
dEjAofUVui2UbGvxIWcPANehPkEmqQdw99Ybo1MjqOcgeQ+FxxIA7hGcsfbnsFPYILlORWuGG+hm
fIshV/jE7v1eHc7y8KLROqDKavFIcG1fqxuoi44ts7Wsfyg5Lh7m+CmKCrRSpRnUdWsFPAnZvu6W
OBCWieTBE1ihAdpVezljENRvOGaE/yvZqrDh9UIbJU0o7QF6TbOfVzhmEYc2sDleKm1/0Ohvi8th
p1Bj/qxGrf2bI4QlBC5dR2Q+UK0DuUvfYNHRMLCWmcUIBAdZfzcig8IbjqeQyzOpsFOxkDfclpJu
gE6nqsSsybFIR6nC7g0gOQuPE+p2EP6Q2kF4PRsZfGMN7+1GRhPMqHDV26Ck6c6hS5HHh7iL+79l
Z31y7SUFgWE2PbSgtEHct57RsnyRTMuzmXfU7dksgtrdp5O3iAym103i+wnugOZd7OJnNdsMTVmn
DkgkvOS5cN5ZL6bTRoU2yIlXJa/GnszSREGVa8iuu3/uMej54539X5AZM58KNDx4gR1mrzVkRg80
i0Bd3Hqg0F4LAT/FOk7nYfQJW3f/PhM8nggMXODwzfegX0kIVoU/gmdAIU0etckNbzTS+Scrgm89
3I65awLvMJNYVaYip7qbHh6wCUaQIbvlqpOdAZfSwKDj0kKTMGVHO494KTzOlpmTbJBZ0SXc8SVz
SaE/S8Clc2/xTUFeLr+hP3FcHmF8WYav3wRyC6pEpiYDw31TGuJ90sWnT1OqIf14sV0EvSpmSSvj
+vpFY1XTO4Owly/wA++PmDRyh1HUmPM1EL/MUdzjMyFukUKiPqa/iqyZNoxhwNrOdOvblU/F0Cmv
EuYD1FuwrhoG6xAT0oCfQ+hzivQ0HUcTFmgiPuXSLPKPzOt5NzPjqjwYxrkNNsGy1WW4vA2I3vRG
v9uBN3631TaaFhey1OXWbLRejX8fZlOmP1xDh8ErI6IRUZrwd5jEfZfYZjvWbyXtSoP5e/gp3GNp
OTRzUiqRaoZv2E59KBRYn8bcmYGk7nWaAGsI/v/Tn8ejRd2l97MScKfkBI9lrCiWwgg72ae3Y1kt
6bqEAzfSubaEufqkioZsKp9BjX0zAPcUNiHHW2zoPahggGh+mrWpmpY5OVIoQ1Qh8fh33gGmqFWg
52JVXZ+58GFQf11ltxu//92CDe9Wi1VYmAwKJuutouEqyfsjuyLbiNCYVyPt3GWNFRRjtD7SMiyr
r4eKJEFSO0wHPgyFJzooR4PPqILu3AWC8j4LTxjbOr+VIGUHZWKCwvhqXUovjqq8ocmsxMMO0hvH
tiMV3XYLvGczx87kMi012JWTFq80QOywmM0+ImeY3NnqGSKosJOg/PaiOvOjbv3ye1Zjr5d2kaBr
BatHujBygFRswoo0HTDI4WICKoF/lWySaaPsTGuFcnp9jFwY2ipp2xDfcdPt2XfvttOVBwXWaUBR
m9dCeL7XU7ZlMk+LpqvIbFQts14cS6zOYdUnaTWK7qIDpwltnI9C2c02T+VSQ4s442BlGsJVxpUT
ZzcoVE0wdIKYRBg/AtRKO0j/N4QXf+1b+FF1vp+P/inqQD34q2A2X+BeYBsF1TzgY1PKdFLu1yay
Wto+E+umuw80aHn2s8xFYss5/5IuXGDVeZEQHVHQQ950jcE5YxzwNKln6xyN05xZAoLdllfgI79a
nKOH9XTpVn9nb7TV8wChA7j1CM9u8U8UWusQWQ4CgGYTU53goZRtCODtLHeSnnhKBQz/r7Mi8n2d
e19OOr9ahQSJhLZH7oBJv4+jaop7DdOd6CJ2HSuJOq/KrJh7dWy8inXzg3/cASVYPzpum2UReG8j
sVqRQjKEytPGZZZ6+eA35kM2dkOPIbtt11V+Wz68vE4+4P6VIIRbAm5SSsMLwQvUFjyIx/zOfBXv
p+iMYdwUgne8wkWnrzaglg8vl5q/TDLhjWSrmuOXcVjQ/gA8evTsgn95ABsm33HRB/dzIUIiJ+ex
qD02A4MdQdlsGDsK+FgKbIwdnkT5CUnhfn0phc15Z/4nkIweY3szxbO5e40fUz3nCQP+8AyJ7NQ8
X1Jop3tsY2zzVHHN29XXdx986eIaxBY0XWioWC9gGYsUBoWfrpYycmzUAHaCXSxtHoXsjLzYnGve
D0wFI8luXhj8P/GSXwZdxc8jXp2w0Bq6xC3BXwB5ans1i1X+Ksycm73T46X5WrGzInHk0grwe7Ig
WLlb+oLYLD7OJi6vHUmxHhurTQDHtUGuaz+akESGhcoSf/cJ3Dbg54DjFPRC9cNezx31debnmrOM
/9F5yzf6GxJzVLPrCtlnDtyThUCekWuZz3Jqj0SfUIKN9XN/bP25MsuPfAol+0f14DoMvS2bWSL3
w/SxuZhgTpU902yVLE6bYPj7uP0CQBPs2B9bPHNkqviMjx8J6PNdIj7bD8tc0qgEne6AuGRRDsr/
l/+PqvnI8A8A0Xh0wBaaeA0XUMmhB2+PETQhYS7RXEz2ECirF+VFHVl91gX4A3N7MwSCQepFLClw
0wnIe5ZvA10VETsNLL18M9scLGqvu7pTn4NPARCTI7FOZd9XwHFgPUJEBw7WeLhUG/dQLM/AK3Jx
o6hoZ21h+dhvXnH2g6lw5lA5YpmKgvom1JIFxHceMTkO9kVUdm3CpIQUssg0m68U9QNkHyRkav2+
i0leHltvjevtZH9IBKVJZm6WZ+/kqJJFGNjh8Yi92x72MDRHtM//Id1/q0jjUEmafd3jv5TmwMna
9/vHSUgv85uU4LlhpQg6Rfarr6nfUBhl98gjyHISA7+1msxa2t6T2gFLg3wD6HdehGkGmy/BsblH
AWsGzncoOMprIRnqQzHHjquUdX8k8GsCIpqmqGZTaQ3WDqRLlfnckmwofVQflLppFZA9Khx9hXZA
trfBEoc7qnJqfxsV91pA3j/LStk3LA/N2o/7Q50PxjqC23Ds3nubwgCXNZEV/Om4Cl7iqonXI3kV
VtlYjJ3nOjxEcjtB+v+a5jGZZDjO1DqzrX2Zey28nMv1aRv2PTdZTfSiK++0x6Uh/3AGIjp91BsN
2MmOl8UiG0Gyh8jp7NUaHUXhQj7L7Qi+19qqXMh/I2Y7/MoBgKUFts3YrH0cM/kOzI3uCPciItt+
DfPvdoZhRBuJRIhvGcF7uOL7a/J5sxtsjXaydUkiDN2cwhin/WxAmPn7zelIF09csxsNMTCQtHJG
iI6orLjscxy2P38Y9x9CSIouMq5YvNSjQdN+9rF1JmDwf7fRfrg6KhzUjDQrW+wNUhXqbdPr3cki
ALFo63oLZ/0AmmaGwzKrPGnPdZA1H8xR3ilvkEQovKBM7Uc+GdD4+RhKR6AA1v7YpAyrj7jAf3DU
Ui/DCJszjwKiFqlq89A+5ALnFCPDsu/TPQKiXeq5NdUViv4txpD7FEgrdDXDFfD8QLRQA1h7zxiO
26FHHfHc3mlImIW+bjnvYDY6TtqWonRRW3NFsuD4ho+mJ5JgIqI8Tyoipd+ZgZTF+jXRQkpEDlKF
9qd3srPtRLdEfox4Y9k7ZI15o8LITA7fsGhsQWTNu0lS+LJ2cX2Ocl8T53Xx/4U5dncKEOHDQlEz
agLTQGjAb5/Q0Ec26VwqE/tajFs94K0jKQjspfhOf0Gfb6WSJ3izsxZWYr5HT+p8omk/FbWLCD2y
zirmjK5UZxrkThM7tFrwGSXmAZv8VeODB6snsh255LMjX1znaJmFx1DscwRh9HPGjtWGfz9Vepqc
3OXru/tt8fxmEQxxJ64MVh7dOvjZW1lVbYzpt1Iif45JehGdoY5FxiTkUn/Ffo49QtrPcQdIIJ09
aqChA0qxgjFR5ersUwa67AX5IEYO+GJRx+Teg7Wk/fuF1wurAnGFnkGp+/PfYlcAy3EAUyXlduI/
tnebRq31d6AvbbcuaoYF8h0V5rM0W05w+SPB432wkWRi7hWIupx1K5dz8ucduLikxPGQm9EqBoko
/CnyUnK93N3tm1ccGzJUs2SFv5t7Siwoz9av1kF8IIXI9LCcVZkuZj4gWRbR0jUP8dVaOs9nH9UY
KdsAu89vk5+776Y2L/LkLoS3h+VyyFlquNy9osFXKE4Ei3omGTMwBfkCfr6up5ojCfyx+kukzoSv
4wbfh1ByCFTV4hG6dAIYT+qR2wmjsHKLeF68eGGbrX05TbKdzTUbvw5Ig+WRuFx8Gn4yw3RFQZoA
pi8aDX0sKLnVSCiikb1kWJM82O73vmCy5+rqpsiqS6/GuhHerY4RS6s2ckYrindFW7bVGEDuS3Xh
XJP2b8t+HYkpLkM6DIM/NU6uhvYnI9Lp5s0h6+FeqrZTTqC5gVd55Yg145qSq98TWtFscypyziFJ
xm3wKERz7HNbY4nTMWIla6nnRMsSqRKep0eA5uoJ1nhRPr8Pv54wPjUYSCv2+LcENkhu0NXK3mv7
8X6Lxvz86vKi4sZST8TqpUo9BkDWSUkpReV233FmPQbFB9EXbnYBDTkS8Y4d2XfkvNUE7IBiB3oe
tg2VFnWI7ruxu21b6jQlViiTmYmFWgKT+YwZf5/tLmnOxvYbaSTXg1W9o0Q4NG+dKfFRZM3d9dot
Mt5xxLnkFV3uQTgTTbJI8kQOHibrArSRCi8Zy8tXvcL/KpdleeyyhmK5wjGOU9RVYhb/rN5K//JB
G0eWtZEgVB2IqduTWPnvJesMsduH6RkewuFE44jsopwBiNzt4j8JZEwRSE9kvdLcClkZ7d7+CcRv
TEizXvuPZy+KLdpWf5FwfND4d/4KcU248vAWi+EpeqdvLohgJrR4dK2zh7mlk1bTATHwQImsD3zq
lr9CSAmxAWotZD9Ci25GJitLsIvpZ1hJUdXqtdi2tEYZPhLc2ajkHoVYEu/d45z4tc/k8rMMUgyr
U1tUBUGsXJDe7qOIc4tcQhy7lBmDsXmQMulFizxQ7sCw+j3EJexbpbd47L6FU44Db8GCqkvlYMid
m8hLqZWbaGYQHekm9rg24fD4p6V1U9oP7o/KOq2hJRbX8aIRuYpigCT3vOrSX0rdoJfakDpysXSf
zA3JJlb9oL1OH/+5SME/ZcbbJs+b4WPgtaClBIbEj9ealnewtlZkedNwOxX+StbwTej4T+7TZlAr
LOEkJe3qZ+pdS8RuyN2PMd6piKqTa4lfAk+rDnE78wG5kmnSxDiAarp0GRGIydjiC6CnyYHV1u/c
zz4GGgsvaQ3SYDCw3ObrJmROA9RIPzpiYjP3ae8lW1s9lUgVzmeE4J0mLm+CFytMveOTNwiHAEP1
UTMEKpSAKkhRQQDiO3xFPdGeUvRYicdXjFMcJS/3rpAMnDdagXSqREetxe0d/NunTO474WbQiHUv
pz/VYrpBTu/L9ZF+V4ikS5Xhw7JvR/oKquH5hhsNjffZH6oAodp+9+nkI6dxyCyyVHhufcXXmbN7
maN+9Onmot6VUQvsB68EgI0ugyxaLY7RIKUqHTcEMxoQ4HiHqPYBTrt/CQl4CBCFEOpnxql35izq
aCi7ZfdupmbjbjQYnih8fSdugE2gZG/nT9NQh5anjp5ixnS+xMoLsRtrVv0FGgFN55C8KZN9x3lC
bmbrILuVj4aPaBD288I1Byh/4sHJejgXt89UI+b029obyar5BFtYxGZMKSv4xrbcmEXR/LwodQtV
afIXGpF67DIE8nkQ6Ux1zjGjkt5svyq4jvir/U2CeBAiMO8e11T+PXoBMYnp9OblM/5OCRBA/ael
Z45JtZ+p8QahKSXjhSuna33VdBQJbnxBhJzzc+YOpCR+XuUOzC7uv2qHsZSpFxOUEM8SWUZS9Uzk
Kap/KdzL+Mkj0Ik4btczHbjRXOV1VGxM5I/M70i20w2BXg+l2Exr9g1P/rjcSMGLFDrmpW1uF6P8
CnW16SUCTxLvp4kkK42shfktldK34WX37Z8wd4dcye5JaXjhePa9eRlvZXj0CU8rovSGOe34lQVk
pGIEqqR3IJcfxn9w2dlTw6DdjmM7bS5x5BSbKG8mr/MsodMexDjCvzEbWngbbfmezey2WtgUMLvZ
d2LtK72+nNrhwRqjaNwjoLVNcIO0nMSMz+3rc7BctRtKS01i5MNpy2f+NEqrrY7Dts5UUwBiS/Dg
qQXgG8S+upKv2NUMzMgdkM0KN1CpkYlXy/AFJjhBI11egYzquZy/kjWu5eEIuL84Z8Xxbbxa0kHH
YZR7d1PORDqBoNjTyZGVap/RJIqj8SlqXjG7/87RNNlcA80Q+RY8W/S4jq7we1g4MWnSH9B2gauu
eAK/g9xngEGLzUu1BtR8TRnTsFMO2WscgAnjeK2Mqa9HvBVbxbkW9fUnC9xgnfmYHZVYgpWpE79Y
SvPVGY5YQxuEIwXftT72pqKuW7TOM0HLg5GBlqs3XJ+R/+e/7AkYODrNQ2Ph1BSXtst8lxNw3yFf
olMSqx+vx7Mbx6WYYpfJvB5yIe2eK3Pll0z6I0bfTJF7yap9fiFRFMCbuiXPiBV12BGEUkMQRURM
3K2le4mz5FCB3hh/cIPOFjP3L/k6k9yvGOeM81t6NbfWJtM3KjgxNXZ7gtA8Jy9c4PWtTk5wfgSZ
fn7U2QHxWbYnkfX/q9de9+6cBHKwmotVHFekhZ0n2yk9T+nBjn1wN42bvGxr5z8e/EPD+rskipiD
UF4SmWl7f4/gyCzzFPMOsiu3V9AFOIdV78eMoA9O7pfBFoFiqs/NOJQWGXE6KWJYvJxoFBgENUsU
JZZ4qmJOSNZ9O46LHgYtBTvdsr1ucMchRevo3Go8NyK/fqvmU9hCzgT5hXnhOqWzLGE/GvS6+Wk2
gqcNAV1CNVSoGNe8JeB0fpngm0BO+aHIx/eIW0V/YptD8kfgCMSqP46sMnUnyZ0eUT2Ciy9k+COY
nMBia9N3dYeBT+iqAVSg4SjXUVCh/zvulZT5stA+q9xIOT7pTNvCi3DhjjQWh2DEPs/AoW2DDNMf
ojOJYt6FIQmIw14gMq0k+1r5BmCgPmKrA9nhy7bTklQ4z9YEOVKAkS5auUCaDdvRN68qFgy8L6xz
7a2KE1VBydq6meFFKtCSCTGnvy7J3/dO82bw3iooyTjpviXtYdj+crb7U7RkAnZTVkY8esEj0LYA
k/5F1uJCffofUW1U31NdBajtL/KQbjA+ekHyx8FkGXf7XR3Z/qmWH5bB/AtTXqwb4fwoEPBLnH4e
W6ddGjWW7iI97tKoeYFHkKSaQxpRzADnEl8lElUnUE1xtYABqOifejryIbm44HWHlNykXZQCGTvQ
zTQPZBacHmJfzcBauRBC/4/4+SLsUhujfglwPFgUYQnuNaX5VtwEyQn3dmSIEznHP6DG1B27dWHR
EkCj2Ckt+nyBRnsjoo3RSmVQHqQCxDwAAcSelmpS8DNjklqiUORva8c38sOvMjP2r0xl5yF6UbDK
v6MBHM2Etmx72Ax7FMS9prEsKs1k5HfFfc4zKPLDORaZ602efGi58cET8qr/I7nEnk2QGt3vfwHg
L+oiLEpbizhsLLZCC9ZMuohxaocJTc2v0e2MTJW16bS9R9MCg2i22DKQDc/ejzDbuxnz1Hm8bA4f
rN504CGKHujMxw0AnUX+OwBwh/snrZoOKIpx5ypCZhpXLyjIj4cR41tbZ5N+wY1FLN4GE35uemXA
z7pa9Tqzmeott7cPCATqfCdtk1vTIOiAG9MFilsfl+TIODtTRHFpkVvUagPLPsLj3llwl/1Ikx8B
kQceW72rjAbU2IgEBs14cogfWm79RdDfYL9tavqqeGqvjSPlz84S+VSoIFY8mBo/dSpJjFiP+McO
iU5LBd03H2UPaFSYBe+ybFFO79yAsh8SyJ3o9q4sXMS4SN0Z0+6s/rif7JUIClN6j+0w9ITXIbcB
me2MABJnri50G90lH3U9g2LugGRqu9oUl3m/MmtoaUg9NJW+moKlnyrtEVdg60huRdlXRdIgVFnV
f24+8qCDhNmhZgQTPUM6b2LvShmt+e06ZGhntzWtoimzEo605fzMYvVV1sQ2AYyFRkiUtXdtaDUC
F9HTeD+DLY0CIJ43+DYnG40BSvP38MgfV17JzjMq4sWPbE1iSza8YXAnYyMyk17ay5nIASxIXdne
leQEjqOVXHbcoGkwug/PU6Ogfllg0sOyk7kIzOmxvggYJP2t/1NpcDBeXkssca9WsqaP8JLBs+mI
wXGKERilxFwzYrDF/QH2HeEuqISaLz2IAWTAm+J/wZeqZzRmy53qzTQSGnpTtkH0gzT8VIUorn8M
Ko4cGY2GXLTNQ2hQpqr2kPJ0tFJ8EutElKeSMCz2/7qhZbAzheUu4jh3dY0U/H9Dccu2GPe+uGQp
kGM8E2oVopifsR8RSxdBGmV7WpaW0JjlGoseC2udYoiJUG2VqbRVUhrAfbmRk/RY1x9N6HJfvj0/
z6Rd8NAIfrQEM9xfd6cLbbBvJq6H1eboye4Hj3QYtv3sicJVELuLJg1LRM89bN7zXd+3K6/LRkCD
R4gkr07TRRmdC8bxKPPpG1tNeCpkPlETUMKsT5QuL11uo4k+tUPP+hgqOFCxnewVj0OSlf9tSREj
vtkMOhMBg16+C7ag+0i7xSX2DOqE1ICDGnoRbtlOMuqs9xGMP/Xr9OF6dIVlzeshGzsxvlDxLUnK
/puCq7rKUHw4LIYYIDd5jjrfjzjQ8wW9+736oT46C52Q9QtMDtJLf2UKHHsxwWpcYKGh/rlIo1OJ
xLiN/ENmYmeHihLAPES+pMU8tdj8xBX9fffo7oJEZhs4Q9zbWn+eyH9VT1dopRzyvVTXkjYRcPRr
UoV987o61GwnPIYPhtNuGw/kSTbN1I1ZB/ftRlB9PU42ROKH0SDd+3fEC1W0nouVPQ9MAgUuxf5o
gd72fSE4UWGlTd7sBIqHciwVA2ZXoVu8g+r7lrUGckXracnxqRvcxiwGjf3i+gxE4hqdk34Be+wL
JrjTVIfGEVXrb+tU1IQNilq3eV7iFfYY7IR72+PST6MMSOZTfrJjKY8j6y/eBxnb/cv1yuKoHSMY
CuvGrLDRutX++6s47qCJxgO4tEhIlOoI+Sm4pJxCfPBr/CBSwQlGV48rfWkqDSEZ8erb5FkmJd0S
McysHhBPHt9ceTK0lD/6cglMIrInm4ecsb9pah0/c2zojXEzL62/GrZ0Iv0P9VLTrf2OiFVQ4aqQ
NfrDgmTZYZKghs2qSOBoVUg7ImEbyXYLhkx49qOHt2zw3x0tEnf+/9Jm6ytyZbtvYMcQx41Mbgqj
lzgBJzQ2FcADUcuZhdqcq/gWlDmyGJySmiWlODmXz6/Z6RbndOJK73KLYG8LbtvknGm+p23sB4pU
+WURpSTL+SOLL6w2hX0Jcq4AF+3ecfcBVEj9O7uKUZTlxQ7DBscfq70zz0qKGt1GT/kMiNRvqQLl
fnLlq1xmLzQd+pK2h4CJI8Prcn4zQrVP/+prme0DDTdQZND5Fv33M/+RJ8DvWg4AiPG536G9SubD
9QXkx+76PQ6gWyL6lxOR7GiFRbeIeBXp2LL/laVerOghJL9ZozrHdWAU75wOGRNTSDFr1CHR0d9g
9Y1pHCF5iEIgmvfzsvbeyvxhczzcvMt5XZjU2RtPLSeWaGCfVGaDl0kzcdfJUq7H3VCJBu4DWal2
2xNRxhxYbLAd0VtUtguKBM6yZiCXvcVe3vF/u1+znq0xbIjDktUUQIuMX4p374a87KPLQpRk3SE2
aFPHGRL/UXmkl4szkm2qQnoQ/K6ARO4Vr6nhxQjQpgEOCNf75GVlRfU3q3Laax3q+EtbT4gr/9/A
HawkMS40JlGT7S1q4iwSiZuc22r6P/ikND7U5AcfcF+THBFe/ixbFFR35gcI9A14abWu/W+A941t
Pkrsm9CVEg0tgujB1WZu6pUgvq0d0++E4JoB6pGTD68WmSbXNTvCcdLj+IwRtQkaWE3ntFnQS7Xt
ueOp164wrLlM52iOOPiF7UNzll3OdXnhfGt2Svr8MWdbJENONMzWUdE3FpYhrROIdnS46N9zEoA9
HMGw7ONGc5jLux1RuolVs9Oko7fAlkAcJIXEt0wsm3s09q0l2rYhh2x6GScBABSkxt7IB7jPoB2j
ugRdaNYiSKvu1lpllaOTskxsuL5zmuFnJ8SDY70RpbvI3nzUxxSP8HfrM57BkhSKeLrxxuNcsJxc
/RMNGADef5TjhhCsuwvbQyNbx0//jn/z8V+Q5L7xkN0k6usUc3egss22KSALZsBy/rpx6fDSmPNQ
KpVPUZGeOTpi7xkezzqzEF63uTKp1rURsHZjhQktfIU9PDexVTnqy6FpMTOLwDQX4Fn+QRQw8jZG
TE/PCR/bYqXC0sGXCLCSR/L8oTrPZhuT/hCwCI0wkQWbMi/fLUA8rkaPJrnIcAp7cb0YfgTLM6Iu
3P4+AzfSZOXDUBHH0gc1GuHN2B2CnjCmxL6h+SVivTTqrByCu1JqmFacrevyBdujI2w6qgyXgLQu
CR1qjjwRFcRDVHCQeb+bxs4E8pfiLlx3jMDxlsqyniWYuH17vd0tyh+qxuzP/BNybXwp7jDQqvKi
tDFVxiGERje6KMuVXaCDG54SZ5WqnJbC4st7TWzeWUzWEGrB8EOJtmR3wMWUlef3xlZMtbYNEKYa
iGOEhWNSHO/syl8RZoYrkkI34D48WUpqc4+oKl3tUEvnZnTiTO+ymek3vBMDh3GZ/hc9KgADXmzT
j6mlOCm90lNhES6YmirR8mLTVqRy5srfjTUlvBtou0QhY4UY91tH1X1PEdnjDGQUGdfPsdEIjUm0
abyboVWpaWMXHDMQXIy4A8jMAoDlrQSfIW/8q6qk3CE0uR05dUhagt6iP0o8fOs8FyP0rJZabfrW
7oqDfvPIwN7erz2I7EWILLorNHgIZqFOKS5gimrcmF5d20VwU+taqlnjnySUeaj+TD87ox4VzcID
CyexT0BhbVi5ekrHp1hgw6txRv7p8CyIgCBgzYg6b50nfe3omWNUkqDZmFnxGM8s0tdTKjOqzutr
oPw4H4Sos2vXcK+xwdQ7Rt/3yeqohPi+DA7eYRWJ+Jc7VBxEXZiM5EvcMDFhCqUovhxQ8bqycBCK
+GEpZKkryaHvxKd3PKpshZc5Zr9QgnH3TxLZMQiaN+sqreBsiBneeI+DGXulD24revvjm9RN9gfR
ZSKuXCMkIPtqXN6GD839GBuQcz0uhM/rZEv++MMUCDZpc24Vl15TSH/F1YT6WsWtkgE+t4XgOfiw
pY4kmb4Id7TLUaOcXBhVAPVqTqbqwiNMsHitlw6TTuwLohDEfHWCN9s9AaLHPMy6ShaGTxdukNht
sm9k9wg8oBClPgaQxweegfQwCYIvnjSCGfqhJkztwDnDTj17mLaSniUf1thnKXy8DHPBeS0IDNBI
fpjUeckU3qx/nDqXiHXmGd6zGrdCMECVZ/w/CP9zC5SHYblh2p/yHbM0d41UnbRMwE+aMV9keFOu
xnf7p9O0bPe2ByWnKq0dSX+uMScoognbQ9QgGFaKKtAbLjnycWGegaPI3fe8DN2iD3dUTsehdHsG
PmCpX+uLI2ZkqWlnWYl4EQnu+FBbRumtnQL5ZOpiSt8nrQG1zjqnoOMMHav+/jq54TsOwalj/Pif
L1yhu7kkL4eLHc6PJLPc9qpuX8Mrb7D/mUzyaCZWe67ajOFvv9HISnPNlX+f9g1juyofUguKTwfM
9pBnNDPYniNsqTk3M3ySunPrldaNqJSXF0oUwsemkRL0pRN5NYqEN99JEzAw77jqZs6gvE2CuaHh
eNRmNLX/7pSrwLz0nEQBIfusxpvRfRaAWsy5cJa53WTWL8/+8iqLcWs8UsGfTgWZbUaBeXehYo5k
wvO7Y1rJ7xzkVHQ0DlAN+qfjt05J566U+AdevuyoRzVVjjHF+YUdAUuO9D/nbV4m5ODVI913RI90
rreX5+sjp4NfZIbWPO1vnuImaqAY3BP7mjEjUTkLdFZfNlB9vLAdUW8Jt4rMLqJXC3d6MCMDcLhR
dgUljF/48HBHwLHxx+kRY99yIeG70dN9k87uY2C/tIFVDWQ/y06pL6UWcJCrF1bdL9TyJR2tEtgK
ET2J06dXMrMsNT5KhW9Mq3EMLoY/UkyZgeitSc15HizulKHvpEP1uHDfeEzkiK3vl5mCtpF1V6Xd
GgfmpjfK2cVzZdkS7GJPplUAGCjORk4uYov26TXHaSdZVwsTd+Gg5BsmFlQpZZr9hGIT7lnKgyta
dUbBssX/i0PEPu07ZwbQb2mQ9RHoA6E6EcN0dEaEW2LI0V1fxhgwMgp2x5XINnoDAYJIizAd8/rM
Oi2cgAR1Lh2Yve72qcpuv8QjyqtqQsM0BmrfDQPqI90bJQniM8x/l+C+zZX1mQif44lw2q3x+dL/
h537UMDRukpfhRFJjRzJ/iNUaZ4ud09/nJCcxJ0jYXHgds3LFNGbbEfHKggDW1Mc7u4tdVUGKK8n
OHXFfotENvM+Eb9gKBUGDVOXdyUFMhP2O21HBmzGcXHrhMJHyDUWXASd2eQOGDLWCtUBnPeCs8r1
CWvvuMiPWaWlJCgpDgyQmjlccxTnKSu6XvCbwMuMZrLgTGxkPcuWzuo4r1wuNdnEnES+ShvQkJAc
k4u20Ak59N9sII4H/7PZe9rfpl9ljl41O5W6PvCoKl4guegUftufmIuDPJYJ1P/pNn6Im3x8fnzQ
rW9yYBD9qr2tejvKWEIx3SNZJnyRdEV+TzNpoR4XJM1bz8Ouk/DRN3w/5vQRCI7C8UxLYkmHKFzd
9IwZwdvBwM5k/U4UpnQ1ujD5AvbTa2btHoP85vCzjCFT/iUfErFuYCiwWfcLAH1i8vXKpbKLrOt4
h8LFoDpXadZ2MeekwSD8SX5KoTu9EA9g/jN9Cq5MlA8RqrFKT6IQLsZ+W017peCyvzgCsrTcW37y
DPuyJPzsSMLHulo23HMn5NpipCZ/Fc3Z6XdkycYhFJBn3k5YJAtXKXrCi5LKp4ppqpRTfK7uIAai
ckXdcUIMX7SpQ/xeQjZd6zCZFHh0KkzWnqqr3KeWzXqt95uSE7WgzTrWfkUEwhp0bSTinvXWVGXY
/A3dsiflG2OC6dW2zylFdx36k6CDMTUPMKvLEUQXJ5r8y7YZHmfQaWe2+YWA2TTVmtvc+bpHD+n2
ZefKZ7hC1PIow42lL4TbnaV9ARF8PbgWW8Wzz5SNte2mNFflxIWgND4qKAu8rW4j3kIzPS8kL0yG
/n6JPNWYb9LeX1z2ScauqeGGWt4ZbfUtP9J6+Vxq/Jy4IkyD4g0ouhBsRcaXH5Vwp5sfk8ljMokr
uCpK6YlbYnz+lcJEA99G9q1bXpv0TYsOzUNs4zfRS7NkQy3FDmFlHEDIhmWayoyMRvHuZHhcKzYS
0Ict34rbt6Q/01OpqJhMoaHffjJ6i+lFc+5ahdM2wAimV+r8kdjJCN+IXRc6md4FG9w89TcMl7VT
DSCATfaobReoNm7uHTIOojldlSHl1eaJ8XNlaznOflHvg7lgD3spLkQR+xB6WKxmT9EhXNq0g5pp
HOgAy17CV02yL5mrafprFsPGkZMqXmVfuvsG6tfX+l/FTrxDKU2mRcY98ON+5J4bECbS1mlZO654
+L9TgRpplr6glS5OACQLe5gdnz9vHn8q7KaFUg21zujWeh/RKpxwL43aMMda89TiG7TSDhoiRe9R
t2m+nQrKLYpRTEreLHFB9hpIMtW9j9ILRfHepHq/NLajt37JQgZMWvWHZrGmE6tMWo1gru9yfWqp
lAVjv41yKa8YNuZbtvBRABDMbtWhR6rpRL5EP8TGs9YH46BZVdTFwWIHokpLMw5vmhiRjQGdKu6I
gaxERM/urQBidJy6opGCrVgymjNVWV7gOxaarzYtXBE8E09ZAznUqrP2q0GR3KzRiSe7cMQmsWhT
tmr294DmqPS/7oBQSxcE/LF+VhZXSce82/TXs2oI71rflwrFTv1/pXvMCBImSC5TNwY0+4Bp/a8A
ebzvABFKOPZUuc0XObG31gjmllHyNgOkQv2fees8GMqXqgENMWQCBSnvpu8+BDwryHhREAZzx09w
fvoScaphFzLQeDseC9FP/q87i444IMrzszib2d1t1yr9jgMoYDdYxbq7rWKyHS2vDmaRBh7+GaXM
fEkAL3VU6KNT0Nu5ruZ0I5pbH0Pbco53+zYeQtqgdYcl3xbjfhwUgmMy/qJf7z3hyWpjGbMEEZHC
sNnf3OGM/pfg7e75kAv71uH0wrocH4EO1ROxdpl/y/vDZRe00cBfbBqaopfNcq7XdiFJt5SVli05
R/XujDKBiN2vHFnxc73qPhfPsX9mjWWtI8LqkA79fRW7Ex3FdujsoYgIP3VBylSUPQgibpunuBa7
GUklMojDPRe/5KdLQsGC4FJC7nPYgIi/bRpqaCgMKOz3R3RI57IvKfGuUpB9mG5cHzmz4SPzXNBC
WsmBOVP4B1ZoaINRcur5dFW9KaSr8dNYzdSmwj2y/Qp0rLElOQKYjP/1jQSCuqJvNcsFVTLsJXVD
xvb7Nz2m7XMcdQq1Qidybp/vl83sLieJdKaL7GJ7l50mcLuXBuLVyJZ9JPrdtPeVsd7+SAmUfWPS
OxyTyMd1HSSj3510K/FGhre7SD+Ciz2+MD70U+KPf8nFPe7bJ79HzNt86n7gO/apb5gxpd9tvsQz
BwO8vX0mygR7JTT2PIfCu7URyK5VZ0YjLvPHzdhv6RaPQ5DjhFTUq8LqOobKssqVMaxY11t8Uqy2
tc8ASQgV2wQnovkbTcnz/cKtWGBPoVY3MDnChtwnc37Vi3dQmbmh2lzOEj0ChZo65Mo/yCp7guvL
KDLiGvBBkl9Qn81aeaAiuhlkb9eeqNxXYzRFmAMzdt+1uK95HEcx4SpnZkVHGigWjusBCWkB1BRl
iHAFc02AKH0Svn0T6tkrC7/C4l3S3MNsi24slU+sqGJ7eHOSF/9itbUAt8MWPV13SRW9QCaUbknM
FyBpH+9MIR4jI1Kf9MSzd545gCF4zZ+I6UUk+iKtNUTYggTZmxDkA5of7osUlkKN6XZUOyW0qeJQ
pUXrQwAPbtBAfl1A1wzvdctTAayKh6Vc8jQB0/VO4dyrlZ0CpDg2Bf/R0BZpc2Dh9SvQGnyUlRcx
3JNpWETf/sTXSgf8q+SmGFstrZm7kWJE6PV5GgXe1+C6NPADhRAAP47BjhOWqYudAzrIe4Xz/gcg
BEzk3MLC2YgKAGnC5bMjGAReB80n1iKDrnnrbxXsTv80sX95Zt+97VB58M2Z5AoLqogCHfApM391
wRU/OHbmg9NgelXYyHcdHrrP1uIMYg83PYTXx+uUOuKK7nIeeaqwL9G7Zp8WsFDEA1G+2IIQaVex
cS2oiTQpzHr9lrDOGVMUCpQX0X2dtomrzBbku+X4xMkUKU87pkJvx+DYCmPSCYAYXfO9v7tX1t7N
FZPPfOZlb0whxu9YRQkVoq5SRnZHxNDiDcvCPi9n/iFa6p1v2jnquU8R6C15w2bNg1BO43ySy6j0
JGZ423vIL9hrSSCb1I9L8qunMdWJdMO+gF/0bvOYkdc9aKtwShtejQIpBRo17j1X0pF3cWZzt6Jf
vEwL0WPmXVp4hPAscLPeIpCpKloBpANB5ykePfMqR7WDnkixGPGaLM/+Ue/r0J7JdskynppFCjSg
8UbbwyjVhsjZ/V2j5ohJvJ97oWk8xJTbIsrLRTs31Tvvn3T6UHSF/CMjptQdwIfi133vtdIxiFKB
o+5LWv4D35ivcq01fSGnXP8/Y24+XsH0ZBNrCQZvGkeUdBiIun7e7TULProLI0v0AUg4NEURKZAX
wGkGV5bMfcm5fGhUF+gafe9pG6mRwUBQYdF53AmhkPuYDb0x0Ey4LSNBryoslVsL9cy1nWgw5hD0
LVNdXbCG4QfGmSR9CjkY6CgJYWANpdrOJELmVKkzAKIA2rI29ZIm12o92/OOK5lVHL6QsPnkWGk+
S+Mwy5fYXUiycYwH8LuGgZiRdLHyW8JAjU5vAr074ssE63vXKLSE3onGEnQwPNzu7wEr3Sy8/4UQ
wMKNgmUYaP30fwf0ADqgpZgzSa5Amb9dIVVt9UkjJP8Y2VvReIGlGcAnXHJOq3GNP680BgOPKJOc
67rkdG9rXgp3PHshsUdry6Q51+960uHsXPNZmiGkmakNmanVOWwpFgZC5mkIhYOF33HV2ryqU6p7
23epouIgektex6G8JwH+jvqoBeDfCXYQigSfRJbcHvMfhr/Li8BZKFujkpq2rplU31pgTylCS/q/
oWLpN1EK/gp7RVz4nMaJXxUn3eEZPqRLhU5dDCy4min3SfH4W4iUzLbep2K97VmUA2Co8/07gq7B
vVSRxcld5hc6hImA/loIKpXuWuvOuISEDsMgnXjy3t8W/oKTPjk02yXNJzvVjJr922MbzT9DMRgz
CyXHBKhsP+mZgR08SdyELzLzO2bsErtuL0iWjlJB8rnlPU6QTZ+h+F/Af/NxAfJ//Om4rHSUaO1j
Hbp8V5Lq6qrly5NdYlDXkmYjatncw30r3v3TnA+1O+mvStSfXowM4Iu/z7k5WFMgnKjsyQiWgUt4
8lWBGZsApfJwcj28Lumv+lU1hAy+L6jAjpL1JjbbyLC4CVllliLfswugUhaosYsYHYrkmp+vGBme
SuJrkVVSKsL7j50wfs7bkxst2r8C1VeA5MMx2TYWkMYIBBoI2PWKIyIWktvqEVjBehJyWfoozdcT
1k/SPvRRqdlrWwom8kRqxEdGhrvxCJDRuNNGtI4mP1ncQDOZCJ6mIq7iNpyjoZLENCx5uVI3BRMB
U0gkht1NPG/NlWvkIMENKqzUOMatvdm14zSZhiXR2F+fgCupiuPahOKjaByJE0k3n4CVIK1fJ1NO
Q3xcCz3M4YRSUnFJKy27JzEKL0VjfBfBp5Cy3vX5yG5D6CS+woshC6+vRkwoxVdq32e0v87wsFx5
dbgtVbEUMA3eI3p7zEhm1uZITTNmqmJ3mfSqfL8C6XrHyQ+6NL+NWOOcl5k6+c8QSSEKiLes8XX6
CgbtP5DW8FWYheAeFPJwFNEuc9UrXPJhGjOf7L/my5aJuPW3I3UOqwloT/tb9cm3y4f8jRQ20CIu
/ftDMRva9XShpKoTFG29anU7S5dNkBDQQzFrRuvXFNnf7Ecf9vi7z8VCVptw7NtX7pmNyWSWDpJS
yHrSveGi63HgmiHfayflR7fk10KdKLQJQlagod6MaVNG2+cKUAA2DQ1o0Oz3Jh2znIWA1BkvcPEa
H7hkgblFA9foDzDRL8a/dhd0oSHUUW+wUXXWldr2XqcDAUAHcGhIhvRwHKG4T6yGdTp1IiWdJgU1
U3oTa2o8Va7bLXKWOrDAedob2uDv7ON00RwGmzvLiiqbV8tfVDo/0JUhI5pyokPNiwqs/iFMPibA
FUiEuY9JkYvxxH5UDu+jDa/Vz7X0rxFRb3H2gN1SxlL5XfNKtneNvrNpcHgTyI63g9NqRykvcgaw
4RSKFjR/3exU2egm5rzmm1NYEG3PUhA24KfWhVktLX8vn/0xgj8CCCH29Ijx4M3r/sf5/Y9kptYt
Ua4vlN1qatDH0fG8sg2+Nh5BghphsGo7rv5fw7qCeTGvi0wYwXHSUAyNRP1w7TO4DU9EBspMo6wh
NPHlrmNxcFWx0N3TiiX3uPL/JPs0sw5WzFUJ3s93e7Gg7Vsplihq8iIuRqbCSog5zuPu77tzUY1z
gkLXcIqFfrGsp+ejL19AZYl42tzeMtcLPAE6ZhyB2WsUq/+ZREUcYM7DT9YQta+2MztgwRPKBbnp
p3nwjfVZd7seZ+C9zoLlZdfK6fzeH6kN3UIjQkX0acxtlpzEo8ECWDWLax9PYndjXfUdLW7zvuGl
KhNXO1fU9jkPbEHF170T6L/X1wYqjfIRqqDz72RXE3bs+0pSUDpwlElpC3AEGaGA9Pr3ist/B/TQ
ut5amuYj75BY+P/xk8a+ab9B7rCJE8yL3JvBrTZYZ9HRDedBwqOBmwneQoQLXwlFn95IvBSVy3Fr
cnE2fB0q0PMS/uBeSKguo/pdL0EgLV8gwBU1b8if49yHjPQ4q2vFwYzvaLC9+XUzJzrfUEJo3UzF
4cTWCAs/GczC0uG5RZOC5Jty3XKlqUjw1Vh1ONBccY5aGSkuUySh7p4ERjAxs+F0xrTuhBvNLB7H
Z4FXc4x2nRbIGx39YM/OqgW9VJoUa8eYkNaaciH4YrFS2/W6jtMcgehjOt4O4uoXfas31Yjt3g5F
cp1lcPU9xDwQ3iJLxKROBZZhEbZFScxUdEa+42Js9j17i8j/cNaT5TjQUBTMehMVl4zI2+lw45et
Cy04bfPvHr950dY4uEEPFE0swcENgt7KraoVaAJ8fPcPX/NXljfyVFISBz5dT7/ykRsV7pq1spTU
mertyLmxau9SZoJPdb0mDRXmctkrYuMVaeVQo3RK1pAzYTaeEsKcJeR678FOTy/WN8K9Eu62T6Wn
zshnZgFg2EDhzqELmRMDXUmRm8phm22Pl/ZvIRtrSGETms7zpMyUz0PRWazeZK+88dWBZQZMka01
o6G1NgtMgG/tU1DAlN+ABmICnN56EREhKGqpJFzGuV44jXHwrRr8y0ZkYe7CCoKwPzxTTHqbadF7
PLdQh/U0rIXEtXa9r2QsdAF75GVLt/Tlgks/YInBZ3GwsIC1ruWNNeMKbPlgl/zNuqj9iu/feF/O
KZW203G0rYZmb9MFaSq+l4P+/r2ZXc81FXI6IDjnF4JB4tUEz734SqlUW/oPqLC718loQqVS4WgM
WBR/5BlhPYh7dsRMLCjRzVoaOUFntzo6rMxj3W4x4BKjjVEpkImVCXV8U6oSN2sYyB+Z65DZFRus
nVFVN8wXEVysnknYp3pxH+grdIELfab1IJ5rTDwZrXRqqV4+UfHM35laM/XeMChdR21WtROlkCkz
NELsYfYj/yoKbsYyosSQ68q4Uc6NTE37ikbWu5C5K2dHjwLbJ/4iqPd9UxUMnRSaou6W7qu+fuEL
E3aXxTb60FvotaqNO96WGyH5IlpYd3p0iPAIqAyWGbjI7hE+FmqxPZFWwKa+LSOUkU2Mh5J6YleK
2LCT+4YpM8XpUUXpySXGlAnP1vXdX9V+azgDJ3sZEx1QVVNXmy1wqVE9QLP3Wlm2IO6Qg72GCBeQ
QxbdJU1FgsxaG0DB1qcMWm8ucTH+c7hm9Gu1LMmjFGCbTNreUZPjMgVmvI2Sq3zZDH6n3C/kC/MH
lxlrIyl6IXwHtKjflRlpuP3fqwkS93NjHRjevqpqz2te1GlynragOmaePQROMxTZo9Sdof24dNJF
brVM52ItczdH/L3rqy/OLU/DPJMv+coUjAROMSaVbC8R5gNN9SYjrPsSDKwtsvHP3/6beaFx68zr
0yneDzdTkErsaMkBOAkLj6KbiakJnbnusSMxKQb8Y8Bjq6BglmwncEkIOM/fR5qjLgEszfWEEDsU
RnFa3gThV87Bv+Mh6sw1ja+WXPfAvRYAaY1BwKXIQYFco7m5hF9FXL62UP+DF5DZDJu0AG7Fp7ru
9RSFohdmqhj00O/DW5qroJxTg/TNIpi6yMNMSXawmJ6O219S7C4fnMT/ZR/b4anVf7ax+c5cqMwl
ejWGhiUnbhb2TdESW+jiJXEdH/O8Ad40otITSLn44itjGoD4YF1e3H8zMgT2Tz5XYoRNhtPLNqdX
jEt6GNbosZlSyslfY2K9t7s8oQeuIHcb1O7miexVUNo36RaU5AlzomJwe95BcC9y4Z7G2DHeBqnV
j/gnOdVrPPhOhphaA6+3/85qdDYp7hGhCu6yoCCyCClldOD558T3VsD6qgu5GXs5A0PlAaFSvHvK
/kwHwan7OJQEQgf/gm4rhAQR4PEOKXLhjZHqlDeA+0H9ro1SRUKx3NcUfgtP3NzFxUvvfr9OKqAB
daxchK9lfhJ3HjPCEU2YhHKSpf+jVklrUlKi8BCzoAAaLQ999EuzTRIkQayyie4qWBc2UX4ZiD96
aNurh9gojRVf8sXgoCWJSBvmKmGvUVrKOlQL/XQtO8p3CHbbSTv6Tg0HINaHpry6Gj+Ru8W6pb63
bPtxmBbEQGz2mjZ2Ln0bloGZ6Aw9oZklFuNZzJq0wWngbhW8SKEjvt8D0vFJEe0wEBQKAMQLbyYo
OTG5CYSs92O5v7oK9sR7gfrG319atGFwFvdK4/O+i+PCe/FkZCsbmBJn7KlnJ7IRXCHSM3yOpmTm
cBUIaVdNxKYixogc3dKqjDbGjPVJMJ3+OQ870T3lR3s6oTArR8nkmv9dyeuWh9sPewHD+WxO0Sti
sdRC3XaA3VZ8jr6sZZBoFhxWb4xLxROzGD3hWrQCpYr6gOi724HVblhVcUem1ZtS5o1xv+McWI1+
TvLxt6+KlteycpFYDfNpgXU9bIJAEMN0VKQPBaPQL42WY7dUMLzrkCp9xIPSzhcCfyfiGeifS9zx
DeByiidJVrH9/bW7lPtpp/ES7DDVyFm0ZzRG385Rt9uv0ewjkH6O4jsicjb7ncIlqoiZmQpevbTf
Wvr7a5AcmLZk89mmJ1BACJhFe9T46bY5YmQc/dzimeDTQc75HIfTBgevF7niNshwKUP8DLrDXGZa
DgUQI1mfI4O5e3EmdPutCZyo6iiBKKNnxqt3GlIDYOi5TicvKuSpFkmhVh1wcxK2ZpvY0Y6MISME
r8OGB90Fa5rBecabZmfR3BuNBDzqySY6jKVv5F4iFS2sAObSDR9X14UX/kTrU1kocytm/bRaVT3X
ZuQwjb5EgxFyX/XqHYijnwvXq7H4WVA2hMXgZAV8eKIAtLSTHfOcykKDAl/blOIhc1rdH66sCEGT
GUMN2dE5g09IwXuOq9lAPGU/e03eOE4a5W+1JKbvNTSWsjBNIpw2PO5aT4Z0ykD//jlQ0WIvyvlW
/7VlW7lG6osh9OV0tUorKERtPdaBXIdl/IDG9GGHwBXRPhdiZdhemjc9cnRtJFD3X7rmXr0DSLh5
BZnbqazLyL4kBCUiR/TwHmxsobAf+aK3ns+MHHi7sF8t6OQflxvrAPGQN+ES/0QBTctJh5Qmtfi6
6Eerxum+nDFM853bWsNY7neqLi7/NEQqNZX216OuH5aiyN7DnWrYpX/zKCuW8oNS1X8xZsZ34ITs
n58VZIUTd+hGfRPEFcTwFoedguR+sTrK9awdF56tsLOmTdqmOQR3B07cv7qKpF76nyPWZqQQul03
8czHl+Upq9RpRceWZL4KDOzsTq7HrQGB6+N3GNqUVl8+jfdMXorlNTdNwMEDgud64PJ29W7aeogN
VO42x+Mws989AvAMIw2vQQYzLySiY3YgjJdz1Cmy/mJ+mDyfPgOq8edUVWm+KPhT4GvOdu5owQmm
zAm7movX78xqtxrOAHPEYPLpBezBugi6ZvuEkGztJSylHzxw7GIPJNSutpRrPGr0W48zfY5jaTBi
0cJxHalqdlcePJKmR7h+CfxIwzHlQAE4VjSTftZT0Ge63liGU9YHeuuSh0NGo90RYumEKxbrZSey
7Sv2qmgvET0d1noVSceq1es/sb651FA8QGp4q4fzEwgfH1n+7n8F0UmDhMTVqhwd4Q0HVx6LFXdy
Xc3b4NM2+m+bV2Zq/7TCJcnnVe9TwzeBoan5J1OOVAX9bZkA8oDYtrGLcXXcSw6KQQV7nGfT31Wf
YtwAICg7XeWnepg3J678gB1QjXUFjlHchwADcKCGOMby8Qr56NYUVldapZ9OHOzl/RkL4eVgZwJq
ON+LK/ZPPbJGHiYBKoFE/8PJ8arlFYnlsGUDcPkuKbLYFFoxNaISryxJRaYKuQKIauEFptbxLlY8
btlj+E1xdaVeb3+N9UE1jYVgqIG12ta/oh8JlUEYt9fJRWIPw7FxCokCx19VBAQ08OUTCXP8SypZ
r0GNCLLoPd/bM0WOyBf6gK0mYqBcFsbz634kSicVtRRA9iOssXy0GYQQHQYMhrPdqgwBPPu9f+m2
keIzR3ek7G9fOoi0+ZCDl2X1It9YbtUTUqAURJYMRh76JVheIWWEyHs/3tOkjBhl8/QjTra1vOur
o9xW8jmKImGM0KNOCwICLMNcJ9ojnlMApioSrqSld3WUoiX1ctbu3gnI7NvVJ94ShjKWwQzvc4ka
aVZtE+q1VPzCZELPywicdKQKP58yACJFk4ZWzb3/qLGF/CW6aUQiZNTnm1CB1uB/mmOEVOQzN2Y7
GNzlz0hPNB0tEQNOqZnpAbBQLLRxa6SR2cNwrVZAGqq+iDugHl0viNmxNZeV6h2VGtJDkNfBsc0d
DRBX1KoPtQ169iPlmLaiMY844OT+KLJw3mj3nvpUOUdsEns3kYIAVw9HCSlT2Xf5KyeslKulwF/6
CZlHu/QHqP4z1x6PMOlyYnHKt+7oIoUG577fV9rqBOHVv7ZY0C/gX8PlTmeoX+okMd7mcSh7KWJk
uF6EEcHjEZI+n22OjUSgmK7efV8U9bFnSnoDY0zF72dIxtkKjJIwb2rEb8cB4DqVPQ7zbr/oSDRW
j65JLvrfPCMTpe/8o1VljlTMIk+FLM9QavjO+Y1uVBhVEYZZJRYf4gmPfPUMgpBtxcDQj8eOGxBE
sPaMCpyBbX+O0bvb+Pu2DpAbWpMaKXjky9D4HkvIdr6WT2/6wwHK3FWyVifig8lDDdJG9hY9L+CH
0JPZhDt9//88rsSI7HJnrLJHCFfT2Q1C+3qHv0t84Qs0p3SnhlpQNI94whXrdFCg5b731Qgcdk8T
FSck/qvyckUIRMRS5UbCjwDj9p//hYifXjlTn2sbIAq/JycvhgwFQ4X7doLDYcVO3nb2M318UJza
xKvFysJXCiiFmq2zcHiU6USg1SItokG2MMMv5ia3ZKzhqYjyiqjnU573BYFasmdNYH8Zeci9Eg80
GHV9UmteIvUR6L/Inu2hNWUiqTR5y+zkg4KS1QSNcQya0MG6qhe8K+nQtl4zQsURSqolTDBf5guZ
JIzCCWixV3/SCElbyCst4jDANYtwQIO2ORIuy12eguanajiAAGCpH49PNsn8hvXmfimobQGHX3rZ
ig7HorkZFmTNCuYUcZVRQz3KQ70Gi6u++rOS2t4DYtGjeb2eBKdQISyYIjm0cqdKxXGOEMjPIFac
C9xQQudNVd4D33z/lvTLxzCJWi+Nsz8RlocvaeKoTtvdtqHooo6JANcwRwkpmNzQebNR6L/7xxuz
dzzu+wf/jDr8XhHv7+01hVSryT4KYWJ+h1vAXVSvKEFfqfV3iSCQxUwWVGgQ6JQ/4LwJOvydLJgB
Mb9rzs+xD7UuRZSHNyu+8YWpyVCp5gd3KMps3IqyuZ2uBt3Zsos7cISJ4WAsOHrrUlG0xDTWAvR8
Usn00xGfAR4QAAbMWomTzGYDGPP33fcw8cT8GGQuDk6EWxiERGBuRa9zr+Rsekz68qAsvj/L1jxl
ILmdZskrB4CBLEU+j7re7wX3soAmCBFNrMron18/Cx88x3z+ZEtrCRnE8QDqwyi+xdZMNeELv5LP
+w3tm/tQa71VHGAkJahO1Pw9XbBwFPHxewUgtlz223wOEhEZosGk0tgKE6DI6XkJ4/yxZqF6euxm
T7RheOKUPZV+sxZnhiWHotUKziu10QP4Mb2Oflt6fAOsOACRshv32NYDhXMFhbrbKKhWR/uAucip
LvUqA8S9As34pVdaW5Mem29TO8MJEhgrfoc9rrcnXoq+QYxAdoczfOiSANfHT9kRy2Y5ykSjD6iJ
xNOpp43kSsMfJZruhjjvlJsnLYYWTEf2G/2yUODX+yB290OapwlavM5nmAADBBZbA60PMAbh6Ivh
Eml+cTa0e2vxVz74EeeL8sZDQGTMA7cH7TH+h1XE1ayw7S1bG11eKQAEFy9hCSx0YTRo8l3peoh4
JTqDxjVhqXBp+O52bk7AcPBx1NBPeQkXk7yWm7sH7pmwLtntOAOm4UKmKToAgG1gnoOeaPK96mYd
6cb4wXvWWEThbHrLgniTGfe7IiVbssNnaTJ7xjaUoCv3/OHyQqXExvZUSGRTmJY3pCCINYRJw0HO
edNyDobzlnJ5ZZ4KIwmCRybomKOezvFJuRfE4SPq1jtEI4pBcIvLPrHdtz6XUASznK0oMZoCQp3n
TepVUGJSvl+GolkCOuZVs0dMBXu3Mx6npj6v9lpvaWhiZF6DfK562FN6KJLBjQRiH0+JRZQqYk6q
MsRIV1lW7uURmq5fw0YaXhuoekPUfWAbEwSUP7XNpm+TPxAzWRv0uFTfXp2SosynrwKGb/6Ppylj
sAcoLywGGOgMJ8SOFBlScmpX4zoc3sTjsF9wkNuFPbjR9fORiZo/qn9wn5sYIqdzA7FfgHraaSkk
dEvPAXPhTOnA/mUwpGvDS3zcusPgq9FG6466rha11rMjwkcEeHz7I5Nz+xGnXCGyaIrZafcBxzVz
PX680QXkQCA9I77m0POz+odiFRhadYd7p+txOPK+1TXG6nElyVMKolw0Ii2Lg76gbQgYVRLRAWm1
z5Oy/IVOe6X5iDVggQL+90jxhQi1XulrjiNyJ4JUn985wsEd7WC914Ge5jWbOSjoTyuAR4T2JT7G
16Y+cPCbtBU17h6SB59dqHlGydi2qQsoe8ZcYbtofmwTUnrdXzT7RSAJt3NYA52bmv5tYgp3f5fb
UGaRbV3A6Fw7axbyNErVvV7JWrOpkctfq3E27aBi0HZcXBaLrLOgBVqpoSElv+zT0aEbZGZl0O8f
N7QNjebEvrxMTDt91QTETMLzTfLB7oEwKhsclxJUAIXQN1eH5jkdnKdN56BJWI1c0+QibM0CXTIm
vWNjUJs82yGBB+bJ2MDkJgh+cfBT/d4NipTmWs29grr1DhEYcRM6yx1KDM/aNN924ZHXz6t5iWYV
rIAOCaml+diYyKpXJhMCnsWLex+4nkCBllp8OR7iVWzyvZv5b/k5ulh8fAaUhwwUogw2cGTMWKFx
voHxxB4B0NZmvT1B5sWMdWDMX16KLzlbakUHVMU75gSt4+n2598UcfJfUrsq7kRgtUmSElZx/DIz
D84Mmlx80dyBAp09Unz4ehIZg7KsNBqDZ05ji3FL/MdRfBr8s+HGxdg4m9dmMM4szOmMQ18hzzKm
MpUA7WjhCjwuA2sZIYuWIkQO58LetRhSf7GbSdqNbhXoTM2W+ciGSolsmmy1XvJ/drjRC9ImnWdr
3PWZpWqUbkmhGwRK+2FrRwNOshSkOTq1LihXVYMtHkOISvSIHVGxOT7qZdGq8kCNabRmNX8ZPlcb
L+X3BYuAg8MZ5RIMBfR7dOKfgYVq4gXhx4kGhgzx389WlGO3nDgLvZL06tOAdRVRZYFY6KTpTUqM
Sg9yIuJB4d0eSkZXGG1RFuVlgc3q83SnCteK8u8A4REGPxjXiAbmeLbC5KjSHfgSNjTB0z3/DekU
9anbnotVjd2lXxsOfBUEN9Si52/FndsvcCGpAMxWZ7ydDbMRNaIErg65eIbkMHuNdqxRD1yz6QcY
67JyM1HNoRdK3u/Y9qcb6kNKUj6o/QXS2GAxio219MUBBYsj+gfOa8i9U5zrhX7evSdn8g7/8Btm
8P9HOAEuHLUIdM36AGM7ITQwDEDsNvyjsHwJpZyU8+LQsmKw06xmAtuFDB+tM3V6cWqQTH0qMxiE
nD4oo1ucDJGvwJyFV5WAMaITCkWgld2zmpd7tp3fQNKpBpNZVvppsxVqovd3SVz9Qdj18DvSfw+Y
fvRVpnV2nCwUbU/TYVBQBRS/jKip0UEjrjD/VyXzS4irZ1GXEaIutSrb51ZEO6yyiRGbHRENpjsk
FS5Odbn2lKLnsWhG9iC8RR/AtSDhJ8Cqizr5iI3FDqRKKl8RILQv4xylhtVW8liAIKZkq4G3L8+t
vDE891ueVQYhk8VcOdZ2gYViSzqVxpxhkikxIUnOxy4ytRZbWgmm7sknKxMMoZZyBpNWhT9WdP6g
pfChbES4To0e3Vi+527NILFiQx7Kc0j+LiaBpnecbWcT6cLaMEYCYK8rPwSuY14wW8m9LEXk61X4
xI2A2FsUMI2so4Olgv3lpweqYelXlEc/D3wyZP4cSMcLby3cQNXkhPorWKOBX1MZJCYNVqabkLpe
zX5cRt90L8xyTkInXDQpkCssoGepE0eDx6P80qrka67i9E7xv4C1Ieb0yxOqjNyr2TPrkEWi3jk5
pZTBgO/Z/pkX5vyfJMGx1vzAbKWiENemWHjLWEfH4TyaKbiqowpd3oJOKvRK9+51BX+ALjGQwgHk
I+uwHK1sGCOZt9L2/gtPYrtRQ+chOycbPfPrPeUuaHKssncPYYjuLiAZr07m6vxgZikvUhEa0RJx
I0PQZyRPnU6iq9ymttM8WbczUfyNJDevxJFev7RSyTkSVfAV+Ufxo4OeDlLw4LEWONIjL2nnlVKO
3xt6AExg5yuam3vLAicXysb1dIfozyVWfhiFjK9X/3H76+y7RTkrlH+B75AW5aobhBBxjDS1iqa6
EKjd6a7FZD5G0ZbfkSFLlo8Tr47aBCXhoSXpI8GEAsTj0pWwJhV7CsVaWsYtun7DD7rqfcMBvgnd
ATWZwdWsOYY8keYuiDRvOvORDKsBWakBpl6a+LarFTPd+lMxwgJubRJwOFXYaGBpSPYbdXnMGSwW
S962xgXzZwThL+cLz7yQPta8EHatuG81l9JQp8WzB7uZM8z5TzLfX7iJqHq2T9+x7tzY5007G29f
Ki+p9cWS1xP/+oeHdQiPxb/USl4ZiJyLevYfPaBRIhOv5rtTh6IOoHKO5P5yade+czfh2FrniiEf
wmKtZn2D+6q6Ax57blQc0Fq7i5+mvxQ71dIL9ZR4jrpL+smOg0vnM0mD9KpToz2gh/Hh8yrmKCKQ
V9DmeYsz2bmVS9T9/oQMOQlQQT8MsLanMsv1NaFuS5dnNsQQyjQ2sJMx5r6lkQUjiniWylXCL01c
POLq/1YfxStpXsqLVcTBVtV/X2tOhrjS8iTtUIG8NPn/uoX1l1TG1lxZiyCmenCIA1TLNWv+KaXg
YxYC8JZR8q2YPWVpn6EDg6ZTvPvGXlI3C1leB5hFdxFbAnz9Jo/egZgDcXD9Q9X2+oGKiqK/jW8P
DIiaLl8GbEYK470svVgMI5O0mVjoLoabIyqRx+2UwJxKJdrOfYcHfJIiZq7Aeg/dWxJWB/a5Bbsv
BZR3gu/cyHXoPGj6h75o+SJu/eJMI13ORMSfa43FDiqMOauBgXMPO8Sbne5/MFG4MR9hFmYIw+cN
8kH1kpoAuwR8RvZTY49ZWG+wuCENO73R11zaaTVWWZpCQ4x552qsF7H5dcf/UgQ4QiHstTRdQi6/
oxIHVvcwhit/x/KxK5gWCa/W5Wp7MaB1MHaouihpOUVv0QSAlRGqCtUUfLjZMU0O5P/vaADB6KKk
zhTFL9cFTl4WPxP7YLahnl67K6RUUf+Dz599+I2QkLn16J/YPgvYqMRDGyanxhQWa626uQ1ADujF
uy6oVbOajDLdjfPUUeJYOLn+FMEWOCCK28V/0KJoYRsOqLoCOEboA3GkS/SGcchcCnBvHJvUk+WO
Ir4cWWeGvYxUAYsDIk7jWR1yL6BEdFq3TBoFCK7zMR8GtGsTUpB3i3nUDC9V0iUAhwbdcOSP14Uy
nWKeNwadLCX0jw/82HjbWlFouVaWLGFKvCMQbosXTgVdyqemORx2ojVZ60ZNnWhb4n8CqzuPcj6v
aLtzTZGRCQQCh751/1OQzOEsRi7ZLLyRP5MCB9+cFpp/J2OEa+XX1PsUAJUsY7vZuJEg7EpNLF5o
taG6RvM17pwViIYxOorqXTcO2EBEZGk57vwS3RA8mXDBch6fWkovxXS+JvwsrUUXe/iRoEn9yza2
3EqC3/XmT1YFIkoWnyRZyMxz3cq3VlCNwuizT1HPDl1UChDQfCP3rfWGbdYdheVZ+VrqJAMPIvC8
9ydKlGiRzskJp7v+LZDpj0snLbvonfpXpdl/fet7+rNbzBtS/hYrqCsEJaCgpe0JsV12a+qJP0z6
ec17UE7RmFID3zz4yRMbkt5fsRJTSboJANX0Vpy2XtxfnECWjdfLQRRTJiawAnlDHu1srwUsgBQf
oF/apodXASXpk++xMsgFxyRqo4dnaT1I90M2hT87gwJodBx8y9PCXPbFTvcg/d+3zlLiOJx+3SMa
U3BbXIEHHXFCstZj6CLMCDvIzE2cRTwOCW0tSDEbRFw0Sd37sx4RqdDablAf5b+HSKuWiEj35zEH
AmmNqEcaiZDSbD8d9UuKk6GsmNwufk/URwlgqXJw2oPjcBeUjbot+BhV5NO6WfAbaz09uEWh9IZX
vWfZnU8ucmqgQmagIF/6sN7slFVquuPHGiTq+5RA/URlxvxPMaOuUYCd3MMlbw4bZ+enFCftsTrM
roBgVMLfi2iHA0rVN0fQb5lDvkIP6gzdqhIhUsJOX1/1aHiBxsBal2tum1GoBXmAYHYkEJTUh/Wj
Yxcg/62F63IXgJ7r4001TNU7HW/X1KSVk9W/aMAbDYTDrkhJAI251U4Be4EMLHsuLVRkUiOdC47p
TnlmEkir7TUn/+nt3kmuNaEXL5VK0JHW4s8SOlGPUXTewcreGkvZdW4lvfjjy13AlH+7vnodLNAI
fF52tIooYM5D9plLF13K+DOuUuD8jLW5W5FeD9NA6jPUS75ouWUKo5N3BlQHYEzZ3omg/aWqJs9e
rY/jPAMFOAgGh/QoWsgFRb+lw0szFtZRRKZdzFBGd9idIFcdpzJhcH+XzUppQKzr9n7LPWDYu5AF
SevP/48zK4xtL5nJSDeHkTkNdOe1Oh4HKwByutPIJJHQj3y7NlRKXwwQTSu3yY4AAavIvuP3vaIT
2ADvCFHwXhGLglBO1V5ktwZO50WCTK8lpM3JcX9X772d+DipXNBBhEUr8eYgXD37Cl8J9XNaKt4O
9Of/R+pyBDOxdsr18ySZeoZwDBnLHuXedhzRm+21C2O4rfA94WBICIkUw+nj0qdGD3vzWPkfiYyV
3OMg+X3IZn5/HIJIjv8IxkHww1UlSzZzjlulHY0wUG18WTi/eSzoJDzVHnfJDrXxbGAPEBWzi4Y2
U9OrXm8GmqWTnUprCfwg6+hp5aDor1qf/AhpiFRAbqG2rHKa1MGhveq2UyUZH7AoHYSTx4uU3qfH
wFYLYp0PteGr1Fzpp6j7vM9vSA5f9Lq6KHj9VCj+5HR5+Z9EYGrs6WUXhYLtMKwvAxtl7FR1J9iN
8vAkCboOhbvcd6eTO5crEAVfgIM72/5Tv65nwxhbIFit5pvqDLYfLzdqfSTcPruipkXpSJS9AqLv
m4ZVyOOhk2lct0nGD16kMFp9dHQWcKjZgFLTrqGAsfrQRCDbva/LCsoGUDmU+qwyIBXdCZsoMcJZ
EuwxGL88Jn2z/E71Q2Nps1JXqj0Q15xypeR+1u5TuidupWTVICHczZHuUL/tJlbViNDCqQ8wNAWv
3nut9b/4JEz31znRqvA4H3JkBmXBpSW/fByVnfzUkjmFFMZPM3pHGZi9tGo9djYtZtLqHKWLCOa9
ep1FVljGOaz0uGmRZLiZoQt/KaYRwNH2rPdX7Gk6lH/fbVHKpdXXzmNM4GmP/OwtgFRQ84RzT67j
TNBT/C8trphfCISFQfyf3q2ADwBpcRuWyEiDZsRkx6W4GNWz/MvBQvivaKYReAnyeNxPwnp/j2ta
3a1K4IVhUaEE6oQTG6pPqkK6G9Zqtk/y4NgawIMRdfN5TXV/BhysPrI7zO/z+Fs0qTsKa/RYdsBa
5SX7vBeFWfrudXVYLkTHGYEVkNM1ZL2mrgwEM4o6iY+qjPCye4uQdoKsdaG/l40EvwneKxNgvt+C
Fu7vHoilDJQe2izzDyYU1JOpAGuZsSe0Ap+791wjLda8cQHFZvQFFJjJTgPq6uA12cWJ9XDIP2HO
BmWKiYyIs0dD13woy2cJdprd9fUYFNGKx+4ectG7Y5+kRzK0n1igRu0j/xPNFf6TM3dhNCMSB178
jz6Wj688ak2RP3oVYI+L32yze26I8iCltUUuRpZwEHbx/gAlJb15yTLFycQnrAly1UdFautzw/QX
ZlyQt+iHi2yF5ULuEtnLi5/M+6DOiI1XEDBvX/uBeS4pUKOgSifVHoVIUiQn0EamtIah7c0EBYQO
/t6j0lpDbljjvVXZVir31GpbivshdJHtYu2bjeyWoCseAZV6luUwbagiLp85JiM+Yhj0fYgATINs
c6rRXCQmztjbH8UeMbFq/V9Z+198nEWF7UsdaC/n0qz0vxzDgYYRTx4vSZf5NKgPIVJaRemidZ9h
m+xjC4llpZLGX+9XEmev69vGMaW4SlEcHiT9bn1g1LzzY77sL7qHh2YUQFKz82d7I4U2AJkNFD8q
Z8CgSkBuF1EAiLgYFAL3Yb19BviurmWZwUI5YOpgJGAe3RyMhgB+eTeWaOQtPnOKUuS81TO6yLZh
uSNbtm/mEFhsIhuChLe94pCUf8K0LCABJ9zKDeXBWrDqAeRItKVcyyreQfI4B5YwOQp7S1X1cY1N
8w6Kqt8fLCP/MHkppNukxQxYMC0j+J7t9c0S2KEiP4hhkRvuBlcZzAABRopIWDGhQvyZszyGUZ/N
FHWkpNUoorzIh2U0WddcyfB120EojmURLMu2+lbE0/wvG3Mxirn1sCnfIMwdg3LHWdoZI0oXfZIJ
lLIBWQImf74XuI8RJyOWZEbVGjNAAfWQcE8IKqO9qjdQEyJtpOjEfZE5Hgri/gd9JFJDVs8/a4dc
TTjxn8EvUOuQyEeCyMkBbxHxjSREcPThIVVHEsWgyfMIkfm+RrDSVauWfr8AQlRQiVz6KI4Ekmdt
OSvKNGSRqJMc0BtSbTeiXyGcOplzFwPmFUBnOv5IuPxNj1vOmDLlbC+ZKRsvFvvKUPD/dnRfO3RO
o3UV0RFVOe+SXIq373cI82ISnlNz3GXU+5e3oc70otxKa0+SGO9JttK9fBhKutJqAmAvuxtxD4k+
pacajzhYd6+YCq6zblxb9OceaezZ6I4HiwZfW5A1OzWbJHpSObZx4Vrb/+a5EROQSiHb+gNjrlAy
TPc0e48B0mV0oldYyiOIqzobYnPRAgszD+cwi86XMLwT07BHUV/EyxEJ7qp/JYvhQRjvrvHdq1iS
cl8LGVWTs+sD6w+tUKHhKw3BOhKtevmH/Mguf42jzr6UXDsOYFeOVBfxLuzjJB/Xs3m+kP9JShsp
uA1o9hiozVZsvwMB2tV2eNH5VmeYHIHCQpjWPlN0X5POhGD1Q6uFx1YuzHn/njglNGa2r7m4iHx4
YD31LIgj5U+4Kqhn17yWOoHPkLBT5ufWm203Y/ZW3255MEUaQ2C0fARSpujl5mCtNPPVGP/izmn9
qy5zTblDX6eJt7awyn5RCj8DzYmIweSjKxSRWleohZ7nEeK+/mxQTnxbXz3dfnuLbG1Zn9dv/7n4
5LZLJo5yKrSdARf1Kr0AEo6C6FAB/b+/g1oAyd9N+F9P0Dh8y7L9ha9vNsBpx2GZtqasCH6dPZCr
a9r0hi9HGAjADF/XQX3p/JSouGeidGfYXFrxys/8+g1iKkecuPMSofew5AqckZL/RaGAJgHvv61y
3AufbpX7mCz53rrVYTbNSGdiYzDyInjYqLIFUGokwcr2ci7TcltCgsEh+a222HDoCyFg8v+V15f8
+Bf9zto6in4I7pzna2dPjXhB19cr1qOSMGnDU9n9pfVA/eEq3UrKuUQ2UN7y9BhgNtCkDCYR2mgL
HCeYRhDp5XTrfMyS0cnihQN92QygZCLsgGa6MOWQKJ6SJpD1bwi7uBgtVOXIpg+8ELhyZPCjCKSC
7gKQYQTnpORQdaLJmnk9QbA7rHiMl5wTEzg/Wymds19FIoXBlxE5rabYADnKBvwwYH15dGwcdZZx
QYEl5EtHmmXpCxBqBOrmsgghcoda3a4zPbuZDi6daMFcsQEfLlbayMVMoUl9yBMDK8pNsxaTureD
pJvte4mp4Qhpy+5gKB5oes4VybV4CRL3jRhNZkgShtbzHsbCfdA56l7qEkGFIIDW2+pfzsOTvSos
CDKkzdhFhPV4+iYvPsO2Xuz5x3iaRWZ0oITzzj/e12zpATgQL4rfL5b+OHvDIwSLlYv39IS06NV9
anpRzv4D+V4OWDXbKJOBar6AuO2aUMdPoiltrlb1wLF5mmfIZr6c9JqdQ2CoNT8/lzSfJKogy2JK
ZqIIxSNgnugRAUsnVxd0mmGwhOb+M2sOxaBAjrBLC05Pz7ofHvgzP1CqOFqCgiiWHcRXZGcxGLzt
d0hSagHSc6tKtUCTuq1lntQ27bSlvMs4mUbLN29pLifTkfWmzOBAS6/chcws7cZ9l3YETztbHZx6
M/fJYqCMyY5N0ruQKRuFZGrA2V3Qe1JbcNnKnyV/U2KGcwNo10kQ339c9/jm/7xXyyezbpAieuG1
6IZOZvzixfHVmYrlhpbR1bcZRXnqFVtFB/rr5ERMkCdhEe/SX2NlMXDV5J5JZkWmFQ57tsonTpEp
xBJoXmwywhiQ05cKPtWcqNTL/wV55FFSipMKxAr55m2euWq3ywR0WcOnZXo4pOZi5wtlrh0l6lUK
0qXH4RTzhy56SdrRmTuXrtXMPU319z/NED9b6HfAaH62e5jrarkMreKHG5yAPH2Q9JiaZwDO5n9P
MnJwqbRVlImaD8SVJ1M+XbiNfF56o5FKmtqdPlyhqAspUPxGN0f9LVFCpzkq2/NKPbLk7iWzQS/H
LIhwJClVyMoaP40lzfczVkb9V3FxYcnt23hG07BpRIk7IoGCptfP/aZ/6+FOhx+Z8HnLN241GqVw
PbVjyfaTncSalCZyrEiPDdgdnAEKJsRXKeTL+6Mq5mWYc6ArP/OD/ZICipzK2S5rUd6iHLCAPjFS
etbImr/hOseWIyJf6SUxe0Skpag0M7Tw/tnfC1ezZ4CmoEZTVipj62Ek+1udGALBhZRcKn+e2pX9
/hJalZPmXYee6WXai4Lyh3FSOv1gP0SZvJ6VSWqlLm59jlFDWFqJBZCRr0542pf045pM03q4w/f3
IHXSnO+9PochFxbIf466KqQS9c+VphfWAOlld8qqfmxpksCn62aIhGagd1mveu+OP/K/TJOcW4b7
c+opNimLx4ExgSX+cU9wJhWb3J9Z8g+CuZ/V/Z2hsdBpHOuJMGRO9dbrT3QnHz9NAE2zdPtiR6w2
pwVHMBuoDgTyS/I/yMrgSKLsTc1BKcg5pi9D9dPY5J4me/8+mDkKLnoOK9QJQyF+rurhAGFdG+Uj
8tGIFyJ2fBuCxCbsJCBHusEf4dQtOX2S4u6FCW3fY+9Wfr1MB4vR5X6ZJbMIKhP0ONWUJStfmXVY
iFYPkQFE0PecQvjlKbmUMWlLw+slobjoWdZD00rpl2/bc33EqXLf7yXX8O9DuRNuoVQFRM4rx2B2
OfhTmdUioPHm9HgsJGNDy0m2ICAVsM2XKrZJRJNs8WdinMSqd2VOIotrKdO2hVrtOKU9RWp2y5Kv
Cfw9V2cB9OoFBawWdC8d7ShlNIke/zOGrdbHivI/5PazfNpdgGSbKtGPNsHcf3PAdSLQMKAkVZbe
Noo/Xlf1U3ICB5FfW5F7YYhgRo+zqwA4XeHtkbCmgtAzuy0WvEMjyPHd/ru+oPewbm6tF2+uoT9y
j+v5v94AmJdMxpqp6ktEwhMKVI8o9vKhjkdODkRJwr3ss9oq603Yu7DuRE+5ZEB76k+/oV9G92Xr
SzWP1iLeOuUE+pj6BNiU2LpGpm0aqZLxvdk1rit9Z9kek6JtUHwa/q2bfItNsmdKjypof9T85v1R
hux14RMA9W2+HJNJ12LejmUkau/3k82fdzStBLgFlTb2TKZ0YLKr9dP3bnKJt4v34/w1mUgYcis+
JkshS4D+lzAeNgV8MCrg92za9xO7khfJyLy7+S6QEZMbh/qtFOTHoffy0RURMfWcC7yzcKJLy8+F
o7BpCGkuFwvH2sPDbNIx6gqOIIwTOaUNBK1/Wf2x2HQUo8eAbvMepdHheFoU5FyqB8cdpFMeWxpT
nSZl+OE1EGG4f5G5AOirrYK2O0EtpTBo3mP2IVUfHUnqZucoZ3VdcilEyiKFOgih8/ilQt6aCKDp
fA8Gu4cg2/0qzxdGBFuTmELIx5e7wn6ZR8DtflwBFJ4sb1Piqh3dCBHshvn8YaCzWJ1Z8oJhTJ7r
s8ffEqzU1FoEZdiU8jR2ytmSnOcNzfa9BBwlnM7H61yEiciK+oyxeRAITe/WQF1AiS6v2ip5zRLH
dV+rUiEf+1z7oe4w2tqK4wdvmUyE9slx1QWWjoCJXo0nLWq/ZiK7O08RzVm6O69YvDTMH8p+dOb0
HsZRtyQdDml8kbj2QotMRcLVCe1p6PytaoXz90WeMorvXPPjHRhJDHmuPB3t1Bmxht60j7t7t9bg
dcwSnMMxFRlf4inFJiU/MzpqTvOS18JVkg/K4Ik+U/gkPMhSpDlizczpunspJ3QYDM/pA3zHOMZp
M5xpWBR0pSfhIaVOSOskXSIfPjYJTQqCMrGQ9Fe64KoJWoDhgJNo+CY3vVkXZerq/YSdpB6ikv2I
HZtRYHXs0dT6c6FOzFxReWKUOPThC1dLHomUSxfPjrfMetZekQwX8zb88bxBuFLRrG0JsH9ouQr6
d6cZFUTkTt/gMm/9BZHLojsTmwV+8FK9k9SKxTvxdvjIj9FMXNPZ/ZnaeXh2E4rUTuTyqWmOthhT
fgPWVFqPXDpQaftBgED/R97wwSAoQz9nAma5GFAaxSYDKvuyjdX1Smo3RiexDzXD+mUWS0iJcrka
+Fh2n+WopHEyskazt44OTwqHN302nMXJZh58Xau0k+vcDRQxUUBNPvmtAOQ9jcd+Wg4sij0C5Vsq
EYhmSYcmpq6ezTfmCSnZ9x7APT2oLog0D4cKzMYBW7D/Jw/v4jjJvAndZu21edOlh2ppQ5bpF5IT
8hEeIL8uZJjOo5tkdKKdgQnEJh8+wmaIGEhhpN71ZrhRXooqOZ5uOgXiVfsrExyNRcFUeeIN4gkG
3+5yLvwEa6+x7f4JmBP5OT7CXCOXiJhXrAagQi85AAVBlLbV5epCXVuvIvzlDe7PsXYOy9F+LAvk
C4MLvAN+PbbKDG6XDLS3t8Oy1AljefFQlUmmOohCi2BNInoKxLVla6eivnocrQqFXBt8aUqIfRwZ
wSyRKz2ulpEhXaIczZs2fErAAvRgf6rHWlO4seAL4xCaleXgDLgUUQPmg3JnUo+Blml05verTO99
6eYuR88bHuY2ieWBDIdaFE2EoQwfq32ea6CVUpWPujVVaKYXGeeOo7sOT601+1v+iOgiZQ9Nhaft
UQTSAoWtCHBUguul34St7TZLaiLIkuK5fAC6Hy73efZ8lL4Yaie7AZhPVs4eoJIx0eTTLxUrzyuK
ydXuCQu3Ce3alTUhjNOc7GzQ9xaYM6+Zu+42wcPmtcSBwXusZ3VPQDp1IEc9VXOYx2JpsobYQQBb
j0BDhCCL44geIvOvSrs/irT/Lh5PcYNtI3/Tmv2YZ2lmrNbBmkTITR0GMXg+m95V4UlrjCjRA0pA
LjSsEkiT61yodLFNiF+N0tJaa0hznEC/YhHaylX0JD99CSCur2GCNMdYdXXo26Js430/0n97tQqM
cXb2qYMVf7vFv5r+NfJHsnTCc+zrpo7BdjVjupWTYVWlnECBVdnZ9SdXl4Opag4Rr4O1xoWYswB/
c0D7GjBGH0H9sFUKdy/8w7q8GwgNTaRDJcMtCtBSOGd3TcmCXxoC1sI0tfxeJKR0qVDV9OF/s0OG
3A2FFb93b4raLS1W75canf2a8Vq+ZQE4fo51l1+WAaTbVLFY/H7wom40UsAuwJ9xQSI+Iiflb4zO
YHlqeZNGonBuT0ITo+vnImrP4l6x318cLwwMSxZZLRWdeL62H48LFxurkpQDbsg4DN0SDYA7740s
rBvgJGdpYV5comD8p6No6u9i6LCGAIRhlBXlxDP+IKs8l95Gjsf/DMDworHQqCl3g4co8fCJKIPH
AQi9waMk4Lgt6rKCNu6Ba/eORhD3rl5MNcq9chDxuUdmT/Sropu0l9LOkWSn92nU7oAuT8fKAMmk
OmUprkXjDt68fk3wzuv0Z/98aIKhGlKt+cPHhMxCmO9V5i3qF2qZD41tHaRkooJKfrBD2LHV84Im
OiEG5Blr612Z+FErecPDh5gHv8YmMy4Sd7mXIMcOK8aE3r40Z3zHGquQhzsVmg02Ijh6IR3uvNa7
ao7zVhRrAVCzVbHNprOJm0MhGGPY8z15Rsz9JFJ/LlFEwewod8q3kFE0d78rp1L5dr1TMcPoEOO2
6lqR2IMLThrbYN4EU3SCvvPEq9uv742b6X1M1eT5j0GjehC9xeKtFj7aE7H96NHhoaN6uNHIm6I4
jwTdHySaKCyRxkWIQa2a+MGl59Xrcdf8zSITusLrLs/Xj1LzwlU7Mn9PTkbJVxpEF1AK+V/jqLND
h4fhmUKEEMU9H8+s/EMPfSYVF3gUoX2JQA9hmktNjWNexIsG+VbA8Q3APpYilcMBORTugaszw9Yl
2Lm1FIC6ZQK5Ri8qJwq9OeBAbo2sF24mdB8nZKUbcoSy+WG0k5BLcT3/Nd0cg4pAP6q6blj/1hr7
ihkze7K5OXwjOLfCvRyipzc7hSLIyGewhdkVnJnz7o6D/3CHV+5FgsCS6QR7nFAaWgjc8QmHTQ46
KqrhXUw4Xfg2HZ10XnSUwbO1MlvaOLczKyBdb8aNoFonY9zEAwN8+1+brmS31F1EbSQ9jg16CgGw
nlil2cgRH14vViJv7czHAucDTeoO9068X0ikoGBM4GFWjaChXIhoQuMRNvzV9Rg9XDmbFnIs3+0p
+y6NwqPkDVJz9ySrJF/bFVS0DZ1qqDFDCHwuArJ+uE041uj8jGJyKv+nTu76XXwgk0xlRcDZZd4/
cH4Cj3ikSbTVE5Fo+vlUMlf03Wo7shzdUuQKKaCy178iP8Gy1sYfjQAkk+TQD53tKYCkDOGwGdpC
cTahiM7cCbflREYiStXxO1LDdsNBNlqAS5qX6mPeqe5b2Uqx51KfuyauK6PZa1OD10YfdHMX4Thx
+F0JFQXY4U2axDoO/nTmo32b9YwxhSzDpbGffHpDANIPzS450DsNzVt6qhLZV5K2mFZbE3zDexTs
d653ygT7JZ8iicnGH112lgDSaxKG3J0fBmaaD1lcxNc1/ZymDBLdz9s5Ip+14Wv37ncCAl+XblKA
XzjTu3lYnGi/kwMgeVjGz7DUVX+peh6QkYXN1aGCn6nBZn1OPAqUQKO8aXstYWZe3PumZtif7ch0
hHbDDXymLhQnNBEDj2/s+aqtXf5KE9J5BLHTWtpKoNwAyTK6HzDnuqb6WURvP9FL0CwvaYXZUqzN
oTqv8lik3V35iUw1jZsnRKUkw9xndKpnFLoyfBPwvtBUAq/aZjqLaex1A4+daiicRBcrcEdJRaCN
LvG37tRck0YD7Nw5HwMFCYpXBY7I73EgphK7n+ZGAF+CiezeZNtJg0Ho3kyuDX0UYfGXkH8Sk389
VKcuyhuodEZ8v5PfY0NeFcja0jBNjoDAdHRJgLsrSeoLABGfDKw8P1hVVRpfcoJw7/Kn7hQgBNj2
DChvsVsMKJ9ldMFLkM2Qe+9m6qm1imYfZs3vdJKcPfHUJ/Uo0ExBqa49bQxy+F3P6eU9DgBfOLWW
ZcTqz5BwkuBOAK33/ud+TmxisIwe/3A5kXmesRma0XeaM0YYeVwoub3y+BEEm9keJXdYgnKhgdkc
RgHDs0T3C4otIfPXX5Mrm5XqkkuFfSJkdP6oI+siW2c8AG9pRvRmX1lOy3RUAKCxqYoirpxMvkbc
AQVCWXXJyzuYkFo6dg+7ebkrpZ09IsT8Bn/hvclydxleVDb53d3rpIu6BYkfFvKxS7Bclbq2MYJ4
vLyVLIYrhyCRseI+KDlZp7NgbO3hp5LFZLo1kn1caJKz/oep44nGKyFP9VpOd5zMXL6CaHYaYOlk
eJE0unFZyIT1ncgckzzrpXTWjBA8LhO+LhoIVWtrPBbLjV3JnLjjtT4ROD6ZjZOUo3liX+7zRH8M
gLDzpG3q8jX/VFDCOczhD8C5UM737ITrF6oSyzTFmPtiELV7uxFag+/zvC7Poq0qcT+bzRsSQ4hD
SFkc+Ruy6ZgRvKLwPVN4c0SB3AwVPFuELsYGDYyNIKS5LbkSzKhyuwQvq2SNCQKq5RwZbF9iefI3
cc2+mzBgZLPk6uVIglCzTGf5D25oYzP/POVwPapoC+NRQCly3zso796Yw+975D1vaKRJ53QXq4oK
fninOOAdP1enAmBMPJaxNcmCDnp9pnsn6tGb5/O/S9TcDAwTCrCE1cAyQasKdJJ6pm5R+sAiHCBS
uWM4yq0n9ho3ATY2pgumRRPmO4ORo1xBm5ND058Hzq8K9cEsJeki3OH3aTclAO9QEZp5f7SKsbmS
6QCewDFdHDKXa750jMEogyNahziiOtW4ZdpwrSeOx8C1t9FI+ozqI2tODrWpDgQHZgZRagHNjO8X
AgFPM9VqpD+tJMfFFPxZbUQ308TArD0h25rPkgvXWga1eZw2QcRtkw6wEkl43p0LL62KsshKXoXU
ap+ZaQ8gEjjuWRqzkyFl0M8ZJn3rK8jHgwPMKMk1qld2q+mEUqv8paVirPxYldzPnV3VQl7acKLN
zl1kxyk+RLemIeE+PTwBVtCPprRR6/ULVF3LoKpuK6Y9Nug4EaehIhgdGSzLNNxpzZfmxvi/AYk/
I48OiQ5hjcO5BPSlF3kVqYnEI3xR6MFO8d451g/M7u4mhKa+JsU/NQensp1/qAzlI0nT+91xxjDl
2ZjXK73AqU/GCCuygCB6xEasrwy9guv/uWoX9dSsj42WOlvN1fFHo8TkQIgx29Wj3Rf8zEjR5wTt
R/hrYt+wH7DZgJDjMQXWFjzlY8szkwDR1d+GbC8eCTiadZY7TZhfjcBdgr9hwlCRlsakKCt71Nfl
oQ1XfdGkNNu7ZllInVqap7f06EYCnfK2Q0m5TyGvnb809hTGBiHAjpcxsz5o4SsKBPtCcq0jmKB5
31QcF6NDQ8/cLq0s6GA5MV5KJfm8H8ZycE5CvxkoYBQfy0c6RXp9uXHokhQGClzs7ShQNrU6XzPD
9hIMJf47r3BOP63qP2z3F0JksdLZWpNikxjGHyb3YEgWHUgHTccQIdNTAAM48Em00ZsOhc17HjcR
Dq9BAyQbvGGOu+TP5ICf9dj2Nl3+YIUN/6/8QbI52/1k3S0kF4/T66R8+jo5rk8dU7pU+DFBZoFB
rWBY+DtCFpDhgklLhhXdUECOXMGmtB05sMEOpM1pFUBv51d32ecxne6015CkX1vznfIjoB9IHEi0
kN/Ovy+gIYCepOCh+OamnJObMwFaqxR9kf2c9K9WBtN0OnT0J7SvSQZmTHbYtCSl4OH2Iv0ivqKC
a2Y493bNAzeXZPmVV3Qla/rXqblsFYrcVMVBXJJu5oKcU5MY+Ik8N4I7/nR3acq4XoQ2k5bbaR68
B31aASpPr+W0SBkzM6Zln85eomwYwXsUJVdsHSNruvPcSrnnRw7KzqI4TQfHPA4xvzHhjRhydNba
3AVpbJLW6E9pmICGjV3+jdf5bbT2VeQ9h424mwc64ZkyxgDTyI4A+OnRYkkn4G3r3PjSUx0cfuD6
onLAeizCU/jdtJ25RCLjW1nkywiozBWZZhJ/ofT3AG+hZkl2w/tCPdkGxrGO5EXI7l4jUKWFHywn
NwGLPuKVGQnPGhu5QPJlNrb7uqR0IJEowUEh9V01qrxcJaXqaMc7/v/tKN6xm6VReV+gkBQ1zqls
sj5TRAGel84jeJmZe2DZwsSaWrmI5CN7PA3BYdiZPgErtXtZprX1KiEveVX0yRPObHwDRk6hfj5X
+OChLJS2jcfHIpGNdjY6+bvqqd54guiCNImXy8QXQf5KXVEs5LwRkbyEUNSmFjYkbfDW3GM2+mqo
qoDN48X8ZTt2vq8d5ApX+cpWAnzzWZ3bh66nLkp0T8Bgrd5D9beWRvwqtkmqJpGRPTUHc8fRJWKv
lrnWqH7gpCdorXXdn5+gSqHOctmB5XpdDgMiEo6lkKFSkzctAYYg5aA+jXK13RgECLQhaf4c5SBI
xyK5UaWpld21ohCVwfNRrCz1LJIQj5zKpZwOF98hy4+dAr+dqP6lUm3eB/xh5aKf2VFo+LvNr5JC
zH5RAnXllLCDasxb2JopjVNujc4+vsNFs/A3jDJ9Aedr9WuOVxq6euAmU5uIlsm+xQN7tcQEnS87
Z0XEIj6q0Ld71cHI2QgG1uvucDWxVA0HU9CluL/WoyeIYe2Mo5S0wn/awKjXMDDEN7CDEwm29ABz
UIWFAeYwR86GyxX7BwX73FMKIHGx5srLmjA10a2M5PUu5y2GjojDwyMDp/JR4+kSp4dNqMn3GLVz
J0YjnFWjccwQfi+S5PuZMpHYOnvOSsxDb3OtCUZe36cml3gLd9WFcCmDJ1mGKq2WjxYYcaiY+3B3
btjEzVd97CgbrhDxwWLqWLKSVu4gb7msSxfJrrdRH68aOyC0IUiwflMIx45q/3U/EiXmki8OVdtC
bDG/Lx6TpfJ98XxpgOQ8Mb0m2Y4rO28tdJE50L5BQzFdh7Z5W8SQ0ODtD5qCaaA2rAINab3AXaxN
lvtR+t6toXs3aDYsi9VdxqbuYh3MrMuptVv/ViFNmpGtluWAtc453qedn95tFQsMghu1zIcmB4Ee
fK15WgT3Din/j0vGvsIvFllS/A9wSqKZxq8QaTxTY45PVng7cgyVnFU1/zEjB3eaiU/pQtssK4Of
j31eVFmWOY67cJCDNLlWOknjX7EgMa5J+b6mtakY6o/+O8BCwflPYp81BB2qTrgwxv0cIZGpxYJ5
RJVpT/HB64QufiH3x0yBD59EXYKu47EAk0xdkf95V3G2l8fbB6leT+vCaicxQ1B+JPHoi1K0qjAV
zj73LvZtX6EQxEcCKwhEZdyoYNnGqZxJfDfnsTdEOV/HDVWiOisyTbQ1GmnKThZ2qN8nUai9X7xx
vIEbXSxF7HNx5paUegl7RgEEe3A0p2jTkuTXq3w5QYUC1mDzSh3/StHBm2T+1BErDUrMmMK+OLik
2ArWNukoobPKZvH/CXoLnyCe9bhjAeRJ9TwyhZyJmBuY0Vy0rLouMDCldX12rRQBUZdo8FP8fegp
zpa7YAOMjFXl42apHUZcP0Yu0fFYUYz4bqOYVlGHfNYaCyLL6nSWAgLGeXXnhz7HriYKZF6Z3DUg
+7s+h1TcHtcX2HNzxa56ami+th7gN0uu18DJWtuaS0lRmJqNK0tqVlPn7ent8gMkpVTP47ej6ROe
qQJNeSe8gyUNfvxBtVKXxI5I0doKXDzp+64U4GWVvp9T5Xu0OWXuWBDcxRZyy///0nMDzWQ0twUS
kfnmAC1J+O8FNzxylEVxzq9FQdLsfgYSdkSPARepTsw1BZM2+jDcg3Eu/NkjMRNEZK0qfFsEBJ+5
2NH+1MZspjwbQ+wxvmSjOc/gPxH2zI7H83r+m5Ald6nL+EYpWF01Vl/rwKZc5shzBG5zwT9Ay1uT
N1BS0YhsaUAFBxi/Ooedg/uZWNWXy/tD7P8NjTV8xhY3a6Y9oociqhujbJVuIr4WnJDxTpyL4tIq
LjoL+8UvzYrMb5ZnGH6pmGGC/VDMCxzq73KDoGip2UviEGXVpB4lo470DgRO6dobw2o4EF8qjY6Z
JdnFG9qwv1bJLx7l7MKlqyqkLEF1FyZyxeOVqm6nONoUDWKC5F4k8x1bXSe4brtBvxwai1OHjf5I
UMLCwDSgrTGMYxWoFLNEcshBR4OeOnvRiTKQyxg5RjRJ4Upg6SrehW6L7VXdrU9sF0AuiOM4RX74
rselhQgrDTWn6Ummz/xB8xrT0ukOYEDgC+4vJ4noBQxn7TxOjekgMFGFtDVuVopHpVZeyCWFdIS+
5Ju5+VrJsC0UbRSaYfmndwhWlYrfZ/YX3gMeIIxs/AotdTbnpZLWZ2j4iWI8zflTJw8jRrSjkywq
dJVqUuMyGFvvVPRSXbDDxSudlk+mA8Qf+szkbJCOvrLxrCUUvk0+ml1khbcbLYmFdsNGVL6mDFL1
SlbmREMLOzOCiAwTokBSdXHE+BZjUsuvO+Oyt1k3pmImkbNCPn8cZO6vpOAnUPDlJugv11vJ4xKB
mNyH0fDaHKSfUoeb003usTRwX+VvqnMw78Nrd2LDm8Erw5Bym8Nh+sMLMC3lSUT10KjHGs1HSFfe
x/mqEqsYTIq9DxTkyt8YQekYxEKdHCrPf+hOHKstFyFE3KLKRvROuytMDBOzRK8jdI4O+9TOeX/S
3HmsLvNRMv27b8iJrH/TIoLf/5FfKhAIemdwLZZ/o7VO51Os3I85Xcha1fJEvI+gaDKuJKqKPeCg
WMqWvqfxrWI5Yg+0uV2CvwnjWcndzjb9mvY6yARu8NLuuZjYFqC3Hwj1ta1BIIhu1PsOLAWPl4RE
gflu6OohTYywvvWSA7j7yIQYM61oe+mA3NO2h4OLR6D9+GDUXoexWEWMRUWPp2r6AQ3/jSfbKIr4
mdzcExeEbjDaaCMaGPuibc2MCrQX6pLni0J5AU5dPOrJMlY0iyb124889FvMhZ4MZ1qqaYHT0Tkg
EBXWE4qvRgSUcrnaZI/I8zC0IQG3OwCxavoMl/lsQa0+OCwlew8MPfdLa0cHfIfzjY0aeRmT4Dpy
s+xQVoumQQ+u8f7DGu/ennyl4DT/+WzrZvNIlazzbkEQlAQvtt9h5Ak8rLJu3uzwOS9MYaq3cUPM
uDxk8w1SpA0fseCjBJsPzSBATSGQSSRAoPv6XBo7CNLvBM4fCPsCKOUPRoRSSHobqCkRuI4207Q5
uYvcIGeC9BCuuWVX6aro5ameSEDtUU/AOHahXL1MTMAtiBNs23RaWDy+an15xfEQ9xdQSTpe1lQJ
5tdKmED1sLgOewTx7KqZHoa8QomO/bORNPf1NSFiAZY5hN8fXYIqsMUIVeuPcpJ3/hbF15MiYeLj
1QxNL4GFcZdZOSE8JCyN5Qw2D2mDmCi/oUaOZ2ZMHURLxXBmSAKcXYw7dekQ8i3R77+lBu/xun6i
YpYFx9YL6faoULE/p4Cg2+WWLcsHXzrVHfVV1Tf6BGmaGdC5B5IBsIyqiuGl7kKpe/JUs7nvInyu
FEgKQaS6uN5AE7IFgCQApwubDtAiWP4ZQFNbCnjKx5kRxZSHC2FsgNug+WM0i3GZh295QpDDGyUv
NCYb+23aX5hAfkQaUl9BUQv48DdYxchyQU1v2V8c2q2CjXVYBiSpRIB8mdlpCtDRTYywBkPIaah2
UOfHYxaeEJiqUtmlDVZvlGDF3gTEDYlbfNGCtgU1TdB/RyD+e+QcWgQTrAbK4W7b2/w/FJBSGD5D
cAfQY8ORzRB2pKb83etZy9zk1IHYowWfCOOWQ4bm8BgUKv69EQZS0GfbabNGZnJd/v+spzMQ/KL8
azp4JzKuHxfs5rnf1jZ4lKdEDax8OtVyARlwBS8sMeACtQKVFNoFa8D0ECgi//FdBXMmclwd4c1x
fUCdS2X5mOxner7iMxnfZln6efFeQFJ69ybiNgG3LN8KpfbJXuh3Dxh+BbQqpDEcJWkka32OpWuS
B5w+kyJWzjMhAywCcm/S1MfIKvpyQdCZVweovJZSnXf6hyAjWtTF8Q94xdge5uChnNkG5SQPuCUu
sDeF1vGfjso4gCWYSGDqHRovIqXJg2sCzvu7LJAf8lPMWPvrgW8hu2YjtUFmVR6GjpJQ8jxVtxSI
DJC9o3o40BmdMuEuxc3fbG7LaXwceR2VFTWIb8SwfoFv6iATav46zuyhjh1uMLoRCZUTofN8SAXr
laZkqLV7VGejv7Rt7sf6wB5lCJpj8PGLiKAmn4+MV8aUGAKPSgGgbuuAsY5PT1FcjOc1UyFE42zq
7gb6rfq3dEdwAXwk3CnqhdfJFetzXkqD6VJA/vSNzq3xyRTZx2TL42bpobxZqpUkVnPXQo3a2YVH
VAktajtw+blFIBVcq9r1/F2zpQR93rcJdL5Ofpp68q/mKwSBF2vNpv6RoQUJ26I5QQvxxIF2asnj
ptyHufEDtGnf6R29mEup68dtrBgZ5rEL7fd5OSyKub/w8vC2uDLKX4AXMrW255Zki9JzbizDvSor
WlbqIlwLFUqztlDJzB2Gzlj79dSNTSdEHCgvu013MBRtgM4c+avLSj/A7r8T+5X3g9voSPR/iyv+
gmg3qvSS73mXm8qF5L2AeP0zzF5JmBLomrCZBslBzDBkG7GVAO0Ky1PsISY/P+xehA1z/y4zdHdE
GiBmZcA2ntH6dsQ9eRtoqHZT9gVHeNRgEofKucyqf+jpk0uFSVZZZ0+vHHQhcdAN4NGORxv3pS8d
ItGl0uUC8F9TmrACbRKkSLDZv149Cru2/LlxWwF3LdhDTWNtJ49DymeSQDDJRBUt6aWuAexjiTUj
iOrvBmA4MrFV09hahiCHiAl78cZs4hqkez4MK0hy+jQJQYQlTEMhb8iHBIKGzuHsfMBLpH0VMEoF
Mdmc4pYmwBZix/SsskKhtsKdzIN1IstWZqqnGgHlLIpiraW9IwWV67hun6LkTHt7mySOyqLc8Qow
kLRUDYrAfYYdjz9/xq6Q9b6VnU5Ywfl+fLpOK3QpBFCm0FvN4MXmoQkZ6dNr+ek0bRctp7bBsb62
phO1m8CIH/hzzRWc63Fghucl4poKRBBPr8oTEUCOgEZ4GqNnX/SkF54OQtrt8KgpHXfPb1v5VvDz
e3c4A099B4cQvqJKhRMiln+r/JcXBS9SstoHZBT5l/f5pIhngYer+6SvO6bSyAxhqJLx3cLr/xBJ
H0kxFGTZbhTs+I1a6FPcASzr5cdmJwbajRmn5ykKZUv+fal6+VeSuxpHnGV+amz6aO6StViRfsDR
7gA9KI0FA2K1xJB643iffzPGHGbEBtCqvFrDnJmefgYOIYEjWD+iDmqzRIWPm0raqcfxcDCfvTCo
mCYEUvghhkuWmAyU3SACBTHCGc0RGk9hEVJhFkm15AO7F5QXTYELYdMqSwiKSguOrI9IvI0Tjioq
0JYEfguafSO84P1pnnbDah7NA/ppIo3wQPGhVeMvZtdJUpWjslzJipOys/adKrtCmfKWkRt6kpLf
s29BIIRqmWO9YAwTPqxyooiRdErTdZoCsDhs9yyevaKjbogYTePSq5sMEWOdOQtWouNaBrmKuRBL
kFUIwbKdwM+XPNUNQWJjaMk4KxSJQTGMJkmopltflIrqP2A/gWcKS6CMIQc6mMySRci0GTALjsBW
HFsPPkIQHFIN/rloKn7NTPdks5Bi590jeIdd+ujQiOj+QknOFhutrmUAa271x3P7hp7IOEL2TWfW
mNbfhgv96OwCJn3S5FAOE6HxhPg6uN7fn5n0c+lO6qsC74gi4399bTuJ4Sk5XLvsfcCv1Mn1cNNE
eFNBNy6qa6e433Se4nM7PozEZvIeEuQ/Q/BfM9nnAeJkdGHNhtjZmh8pONYlEpvnpG7tY/lBTbFN
hGepimxUxbqvqk31JRublP8vbpcdEalBesh+W2n2QAbX6d8mEkISkDdo9Tw5MoRPwO9dMYdIbM0N
2cwbzXb5TrS6Cta0ZhLH9uLJXNpISTz/2RJHs/Zp68cLLH+Iz5d7fZqwxFbVE5xvGF6XVbbWFZEH
uhFA+1Elw6N8ZvBFtAC6+y6rACBegYvstxdmlj51sYmq5eQ9wxUYhEb/RjodPAAE6MEx9RmUZ7Lk
Ru2+hkiOFtRKVRehtgfbOOm7wMYZQBRPOhHBhq2NGvinrazBTIKbO8G/nZzuUtm/QS4T5YwRe7S4
kEDdNxI+TcHyAo6eyWnHscd8Tn7jTm2FKYOBMANRoZD3RaaTOyStgwpF2ovrJXbdo/XSlorgrFLX
ok3ViyfxKOHY+wnVk2m3kWX93AoHVwmM5X4caaNKK1I69JXAHsH4OCmQA3t/P++eaEtXKLYiZ7R+
L5gY5MUshE2MDMsN9Xu7IgiGzPNaXcrTHD1sjzno1v4pZcTCrB2vDfvgeGNgJQsMfoHr/xLYkaNN
1DGUfzq0ByUE0HQSFHNsvzYn/L3FGTRV4YO396CDQGXDYuX37nCd3oOcB5Cb3T2pvr4+8Q6qIsN3
7/ve+dy4GpGR1XnCVg4KbbZo3eQK0WwqaAZr+drQVYg+Y7yaybM6PSHgG44hcu6dm4+We6x3TY6Y
hnjg8VJ4anHR0SRhc/59HZ9CNthgx8C/Y2m1/RzioDtCEqd7/l3rQJeoVtjFbQlaU03tXZFDSkRE
1JejqimLPqWZw7dwiakxoE0HhNBwZK5u26EXmsB7ZJjVObnBbYKQ7eAzZQZhQFuVdQkCGuf9PCt2
rgu7XCNQOZDJno8OvILVE35v+PGx6040IZmwmOmEv6ixjszggxN954wsol1vGh54LrnvfBcTLWMK
rMcsDMUIQVfMfUT7pu82lij9o/CUMcdRfL/wUgsFAc0w54vIcN3ho6sWIGCtubc47Zes67NOOUNY
BrSKfUIUkYncbLEFgk5qcs/hhldWwfpydZb46pE9c0rj76Km4FD2EjWW/pSV0Djz0nAgTh5KgZyo
yLojFKJlCeae3eoT659zvlhPYlNNLCyb8HV1fQjwHoKmJT1QbCMlVYgrolPTrTt+vkE4kF8HXJmS
ruR7qmAkE4ngOl7I3nB7T2mEV8A2Aex778IkITlOi3TSNRCn4HUwj7gnQtQziUu/DxwGvOdClgJZ
NpBSeecHnCIx1dXxgCICP72ka33FHF0lf3I00tW/TaauYHw8BfubMUcfKYNrKt7AgTtdof1T+Hry
UWHphDZPQ2nnBase3LeR4eDs9rQ9pdJWGpxEwlm/+NwWYg9+bUF01rLitL4QloANawwTq3O+0ZRA
bdR13MZHT+PFN/Dq2MKGYNG88t4+zbrtiFAXwod25jtun2rzn+MK1tnfySDYYGBozk3V2s8orBvO
LIPy8/57SLudV+sTHFsSbLze6IUblJ57p+yCOYh/hg1cZrW4hvvr/5ao/RGR9brCh1og5QHTMOrM
eS+IhhWm3yGkm3ORBsIccankmF8Vp4XwbGp+gE70hpZ3WyPGc/a76F7aHjSbNR6jPqUQtWpUAvC6
XW/wrPEFmURqPb+OWyRb3HIV4YkKiry6vwFd9awPZKKC+kveixVqI6koQ+2RREkETR1hMUlT0kqH
oWnn+un8LiiylUkEgMhNUcn2yBZKpXuL0orItrzQ5owlSqA8duEJtYajXnnjvH+JOsMj6mEZqQ1L
fBFhzD4VDh/XoBWH5pRfAhPxjaNgDobJbKyQkK7J2Zq7WzfHFDvpwVsH2CoKGUBS7vQuPPvWxVHc
IhqL54DiqfaSW8zyLg2zVHoMXWRNn4NUjBtiTbayLPb9SMpcEt94oNsZxAnPfARLYjOzD3TyM765
cNQd6MQVVHEURSv4k7XgdS4tBQCDkBNkZ0Tz258GhBNffyEX94sn6H0D2/p/LKyRkMbM3F3K4QHl
mJuaDkwQHTxCNL1+VeT3bSBrC7KT9pfeBmRw4JLx2nGjn2ug6gxU94hcTjJmNyAhfj7a3IxeWIAv
CqXJGUUevzKVcH93iDgUSi5SDoLX9dQTwwq/OyO3WrXlU6UlkPs1r4TEfLYcVJfHF323lVfopg3k
ONTgvK0j9TZCCQ57fGwnwGeMAqPMtnogG4QEF4NE7hrNmWZfnnLNz/5PUdFvl12HEh54xCbGKwHc
sTXzOvZ2gyUX231CMKIyLioAFPDQjh2mUT0df5fMoQurNIHveSjvW/HisO//e7WXe6AMyTPoDA0l
SgoEuBGuPrIKrx9X3HE1vRvYtbF8dQIe4nC2hztMz5co/4mTppkeYLlxLKSsyQaKPRWp1hdyXbj9
7R1mBrXspEMGMTPrqci40ODJK9zJIWGTk6otNb8Fda/KLGfgpVae90Jwp1vTIFce68Tj/OJevtQr
D+x0D07sSYCXMiXig8fCxzXCfB6/FXKQ1w/IvAkc7xdt6IN6pv4Gcy1izKf/b8uxxWVdb4g4HZVh
/g4kNFAPIPXNwpQjbrY1E4d+00jTGlkuZBmTCc0YeDkt7L+O0UYF0z9+5qvW2QjPf4HXvfIVWbFm
H+NN0gY8bMW+Ak+G8kKpGLqWTdFbUKQ1gp3Ecj5TInWzQE7RsNiwQLJpUqowzW7IqA97deteiG1T
c0W0py+VgXzNmJhemtkR/r15RmdGrr7XFHD57jJF3VMfleJPwOGcYvsakZJ4utqPzMDuKoHHso5g
NrPVhBV/PU7d9FZ1P0IHuhrGe7f57xOewk/fyEJ+3oXuyPO3ZHPB0nsFi/SkCXUrMlujoqbi142h
C0Zx+vx/wXX9ZZb6qCgHt0zmIDyq8Ho5ZFfLBm/XXkz+OBoljyap6TZRoMX0Y4NP4MZmoYvlFzJU
s6Fma2AF5udbhxXu2QXUoqdCTZOPcQxLAcEy9HwJStfak01noL73y8fvl10eB9PzM+Jd+0ffusod
IXHg4gwnvkUp4ycj369bpqGU/nATqMIei6gPPJ18pHGkXpUXlYjInwcEMJW4U14orBArbnyoD8Zn
DgNLhDHrHzn+MEE5uIYJf3bB+++x7LQTXxReaguTMDuLSZLFZFiNhQxeu+QnvzEL9Yhsw02ERteN
NZSm+W6AbM5KY+gPqEh5ueHUkjaVMA/ndpfte7QKAabS5UNmw++5Ny2pjmMeRsiFxKv6xBGjq91l
FN9hg65lvAQKHFC8FCThFUbuQsddhna9qATyjia0hEIfR9uxiH/IufoQy6QfwX0Nqhft70gKDYKd
sDC4afip2BWLOjOXHFrO3B6yq43jXi2UtL9PskrD7kXLw4gSzkGFhEbk+LWhDLpb4Rkdb0HTmiem
k2F+pgouMMgKkCi4pdb/Mp80PjhLxt7syDEf/Sh8/IlRWFW1BH+NYrpxUusq3vDOJjwasIbi32Rs
eAyK6jWJBy+THIUVZ5+SL118reNUMMbgZ6bTJqS3cuG+oz6qzd3Ds7kYn+f5PHKiejkqoLwjvwM9
VWLticSirumqWs5zh3FdPCMRJydMBDksQ26VT1Q3Y9DMwLvo9Mvhy00a/QQcyMm/4Z+WD+Vaxmy2
TJGxf+ZL0botxJL+pAtmNRiCnW0IHKJ8WflgcMO9X+xpugBhJVbNYt4P1tboIay3o/CudG8BhTeL
L1zaBTcaleLSobFOksYIkkj654RajR6Aos4WQimyhKGR56zqTV36VHqy/MVgk8hR3noPJm0FFDiM
o2MgkdL4I1V6s/LxSuQhVYveXqAObG8q3AIJMD+HeX797j0SjZspA4tydb9Z5xcUFSTDFbhmsJVe
I9QHPnyQkEOHcl2tv5JYWFG7Wir+N6s/K59cXxDj34rgII3m5Q0ddi3AAYNgskKOGgiBQk5Q3J7n
uzA/WeWHz/Am0zi8ondmKGv2mVkiMtPnyvDFTIH+y7X/KDLVW7Rwlz5dO7wlEbJKzJA0twou1066
gGQ9k8fQWriMGfY0l8Z3W/NfI2NGm8PeK2QfuAGxCrTTfUdWAi9WBj60BU9Bk5p+R3VAMtTqDKlV
6kTwXwvg2sp96L9enPCMWVpMF6tB0OnBhEGEng50k/bhGKXAddpIjSU93W3orz14Ib7aQp8XEs6y
XQtfaWLgGtozgBwUKfwsE/NLDpyuiTLvqKlm6mScwPeWtUAyrjHbHBzdbbyw/maO6ObDzSoCZDlv
wREF/E63Ckj2pzbAhaosfUfUoxp5X4iZDwm0ixKWGY41R/GJj65gU6SYN8AaYQxg32MQdYgCX4iD
IQs5dWvNC8Y1180lNrZy42jw23jPg0UGebDf5bf0F33GXXurU24WgMZ5bJhYQ0rpj49o87F/pwAA
8QCYB38g0ugfzNPea3XyO78u7AmQvJDr6jj1o8KSjsLaty009wousuuU6GKbxlGgASwOLVgk9m/v
Ol8kwydVdaLW6PPsgktQMO6RSpuwCtRYf7tbJJZEC9trGovdbPl7uyLJSAADR4aFcJ6lM/AM84PE
iU6Osx+wvkG4ChBKIfNrNYIlpoaWVKnN0rRpTScgK7ePE57vxhThl1IFFqmz53ChjUcVOr/hAozn
ssH6ttoW5OSVHHre5NI2k/YLJocs+jjhK6LOVxdaF25Q2F10qUGH2kyAxoCeRwcsb+g3YCkQySdi
O4BwbaBqir+0lH/9JnK2GRG9u4iZKj4BUXa2mXpMihHLzrg77/nCN3i6uZANcFwHbwBx96DUArRf
gFWAIJbjGAw6xz6du/QNK1dFqKy1S0MIKVJl87qlyzEJq9jI1nip+wKvIOzli7z8ad0lZ3W3jSJG
qmA1WFKeZaYnMbyF+BmF42RuylOf9b3Gf/bgDkpbnUK7mM1PjxySgh6rCezO6BF9Wm83mcyuw9MB
zWsCUdAQfYT/gHKFGkkLwtb0gNBWyvYqfWwc+7wv+rTGftAMg5wTikpuLFCXXdQtPA68qg4uO5GF
waSIGIed3ks/mXdOabm9BgDlBVphk4yv8LUbm10IZBr2pkOoDXwQ2v3xJs8XFVyDm8FYHFuXp+OX
evyVB1XyriJsVIyVFeFfmjS5gtyqasXFsiw7NaFSCjaQIMNG8/vmJZtubj2XG9do+iDQf8Ai3DtR
1ZIVOWYyiiFR96g7Fi/G0PcbT5HW00Z0DpaOENmEOI3AalpEymUKzQtSbT35cQsZHofX6PfluoUS
AbmxuTxb1jRW4dJt8dROLY2gTeLUgOGH0Teg7nDEJzr4OI17brHmqUa5paIEU6TMb2G12L0zqr/v
UahoFrg6KD3OcXbdkXi/T1wcxEePscH2ZCF1bRF6bATKSvucxg+yTARRA0Qj6pKqr83/JuhPpQCd
3z5Jo5HXz69+TDnsDzDSxWEH3gdHs5aYxUcinUx0+nrtZJcbzR4/sNhd3TOEFXm53NvXb/oIEOVI
wyZPjwT6tfr/kLMRAY7Jk51wmt7LeUIHj+x9QZJXgEIQlihBcp83R1jzNHrKGjzzQswikUxd8+6W
wzdag+u2s5sdeeBS9Jy0265g2bMdadK8YS64hUzhfgZWoSd0VGrRP5/eGHJfN6eiY4qrfg+n7pw2
pZAAD4RDSN8E4rFQPlud3Y+BoGoKcwCMbCt5QdH96NkgwzvQnUwz+KJauihxYax52+PZ+E6/0s1S
JH2SUYrWViYPgkiWQgOzWWaKcNPMqTQSp2Ip2/XhL9u5MLLvUsb/TEpzAi3MPOT86vi7RcVOtHAF
25cuFZIJ1xiyBTiHSFKe2zo++6NPvkFhG37ZP2LoGovhYm4WGwuZSg43TaxvyAPIulVxkVyW0si1
pyXVJLLpyp2LelDHQOltPJEIjs4btrDktg8M+SkfIGxYMqE4f2bUMEJqMLaHvGWRk9HCQ4l4d2ZM
EyQ14Ui5uI4LS1Fepu7q6xWb7MXYtlUH5V0imvaSbTVnCA+ruWqadHIluTQIpSSJg2mt6ySrop/y
9OTQvhGpfb3Ukl0qhymqiL8EqqSe1vbP6uV3CQdaCnpjXUoKbupqaE+s0bIYhUXPthdsxAMLGTPs
iKPIvNqMEFVQpFsyoo7x4t583mowi86Wo6eAVIHsM/ozibVwL77HaLqTLQ6AWDkwwPY4dbxpm6fq
gQ7TNPFttUxuumtHhf2Ykw6lfj/zVlbfMzADaqxRFmDxzLUlAEoMDVpdY8uqN3+47a3lhvO9Q3HW
nRgmmAmr/SRu7IiwtiE+GDfEQez7Vv3dTM/OY8KtvvXSPQDx2nBTSA92hhhXPFVhUljX7WTXWVyv
odNMyHu+m3O9SRPvrTdepK+uJh0Tcfe0VoJEdC40h2KJfof1m6W2ZAJvPIY5f3wlOGWH4wkRw6F6
ywZuUxHSoGoUDzhYnexmMLd9edvle5hk1pEjc5e/gHJaJJjn/bDZCVz3c0Rdb2slikEBnNoRY47J
EKWvf1kVN0sxzglOBJXPH7fsObHDZEoo7LdKoFzssSi1i5KfM5s+6BCHx0xenV8NKy9SzCwKKH2j
tkfNfKptFHIzIcCT6wWu92crgcwhoehWbfOqnjiDCFeCAupkJT6sOy9vm2/mjv6mDbF6Ma+pHgze
1fIQXnIjW0dCUy/5n8tnhRMltJoJAzdGa4tOuNiS7mapXyYbtUpp4d0JfTHJNMEVBsEpi7KGoZtv
KgPXor3RaNVX3xv+CmfwIcC6je1fWYE4VfdAxh8XWqcQnS37hibqZ4j7MjJzE1QAaFBqZ8v21kCK
EpN1ZgW4jSqD+/XsFXImfLeK3QadjpswkDFQ+2MliWRjCPgaZrerzygP07W8LV+5H/8RRAV7izdQ
fZ97gRDhKnIf9LfUeibX68J6+k0nqaloXnLuP3BiZtuuj+Fn6GOh0/Oz6glOvsryePtYjgNUFFR9
VwhmjgKu+yeh08+fQna+Z7GRENl8+ylY3a6XrnRNs4GfP9SJRI1RlVEUZ5NKUMYiG/7rjygkwGKP
J8rCDm1VQPrqrdM+o+UDkgtP/shFxgUhYfT2UYRR4yuHnmvg/pd9pk7GY9sJn6Uk5nVa1RP3kwGE
8QlV3GaJx/cu2Byti2DddzjWRXQQCkxxlH6z0+3T/1g0o0/1tO+Ld0HghzBbvOqpVKnFK+uhycWD
TPzttTanRAY2iH0JnOYzbGQ/JtGVs9RR0+23N6yIkUlkMSu3C5jGQVuXDmIGIbkWo9YtgaDhbxlI
OI+jPkyNF4sZX+2FzzlN+6eLNRgNMOxyTPEpOnkBlwgc2ouoXvVv4zkKvGPSjVSDNoUlfjmKtSoa
Dg0zQhnI0FqU/0d6Iv7zshGToOIVWB2rjtacJTXd1cyDPnLsKaCUwVTZJZGjqnipZQNMKCk45fLr
9IL9Yah5D0CWv0d4BpivmQ/L56RkF1+50eDlfl8gT+opUAfWm4v+wBdfgvQHCd6sT145OYf3utnJ
LzlI9u2YsUQrFZ70b0WXfJK0KSNIZqKE4o7bR31+ZPDGFKP67EtSLusdOh5qK8FDdKrJBbmtsC1f
XL2fU3KyMHzNTXivx+0S2MUO87L98unJMItX2s8fkYYw8tjn2ctnJumEKavaOnUnjiEPGvrIgcRO
gR5jqEuzOkwLDAIiWXrbQCb7Qrr9MJj40GLtAt5fIYHonkxopd0zS3kPTPJ6DjFoP8zFzeSF6oCr
nB2L5y2ND6pbWNHoEQp/blxswVWHUpODgImJbIXugpkiHwz1nxHmmKuKvLzGO3w1wWCsmXvOurVd
6dM25SiisfPFzGhJcHMrPbXDFmI/e87PwqwfjCJMnvLDo2g/HcYSfYYE9Tl1jb86CPrrnvhuSXj2
4eBpFmOjHXk8jNPoCSfIOLJ9PaBQJlpkWsFi87F28RVzEg7gAD9RI6U3qb7kdn+wm67IlLkU2W+r
JNhDFvvhAFxsC6BJcSHFBSkcl14TPistKRGbHQazq5fEaT8D7+5F4E467UP+OydYEPauUv0RihtA
ggkVlhZvJtxZcYOJrJ6NX0Yd1gpwwI+nwOaCA7zmVampD4eatYVN0LmaSYmXIRyCD4zegna0/hNB
i4P7SUEhr6fOCO79E/DZM6weBTWH+FbY3ZgA9e4MQ/ikgtnvVXd1G4uSV8gjnsOSkpcS7uYPU0WN
488ACg2lIxaXyF+OIsCLsPB/vto/ngszjXmP/VKcal2iJx0F22btBm7xpEcH+11Y9lyBAOsDeZMz
7IqP9uqELRMpOBCZGVpdchSJfNzzij93T89KLXF2DumnN2EvCAbXBscEj0WhIvcJFQyIx3NtefAr
YXQpbA9f4SbiOVJmGA1E2Mg/wIb0VJb8YYR0v1Zapy3Ai6k9typeSA8BOyjS3xVK71/1oAAkQue7
9WjEXjHldgXNyFkMoZZMVIec035jzVXk3k7w5wNA5EH9ScRUtzkFme4MoF8bcYol1B09/NkcdZ2v
7tz6O22gtAJK0B1Io/ck6iqSpqlSKn7MYdJYB7bZlTEYLiMUR5qRA4KNU07dLo45Dy6cGNGsdO7u
GXkr7phq3rUvogfNlUY8rFoa9ZVMzbum23FyMCzW6Uexzub/J1vCxpkmdVUCBqHjT0ktNUaUo7Um
zouEciuQBxp1IsMjU4SRJCfxYD9IANs/9nom7A9pWH02plsB19N334wRZ3TUXGJpaUWDMnFIVCBx
3quj+6ptFX87gF563guqOaeZ5KNsafqKqCIw6WJ5HigB3L/0vytd51hChEMtlg0XiJ2FL3G6kFse
jIkL5GpuQF68jEhHEtO5aKVxyPFjrk0f0HAkWJBQxCZsagSVW/UzsJQhnQafjjEoA85cPuRIv+sr
wdo2Iq9EXSW9jUk8XEymVS0qG/qTHBVZuBTN1+OXixNBuFo3dj/WzmiAonb4UUcjBswtDVwD8I+8
pNw+I/BVPsGAAhxhL+bsufX5RkoVtduMzPIRgTrS1g8MT4zcXXbaaUO9XVbeQ+SK3kC+EXAy6XQZ
h4/mVhKdI2GK/1C8rDM6jM3kgO5MOiGzedv4C0uDq5sc33GT34u49xopoiIFner9yx3w9LmvGQlK
Z4Fwa1JkWVwkPKY32O4/zMoOl1VZ2+EJgyPYHLURLtTeovfmviop5LgiL3wOo/wBFMGEyOT33O1v
x2NjiaeJUpvStiHSr5a4VinK+bikEj+BSLIf7toBg6I5sxat0wFjAhkzQVzIobuyfuYQqZghT4rl
buI6Pqn9w1bngwF68RzqUgjxst7CMSzp4RV3ZjO3LCPVknJh5v+2ZaC4zQUpy7hgVUdo0vFT36yK
WMt5NdTXb/bZiaidN6oGSMmwWW+N9MVcycBTtXb6mp67QBuFyZjvcVR67KmdG7hiRuse04MYtJ7D
OhRinFe9PMipT1UzoGAdzOe5ZkpPr7H7z5eQKr5thXWFTzrflbH7XTO0Z54M65PNHXnbCbbb7L0F
Ah6E+yshCGhLAqRNSqK8hhLs9Zm7EKNgAgeahf5AIgxzHUFmBvMUrH4g1rAtNuNGL0dAzc0oLpfG
l+EtJCOvbzI76/IETNCRjyONZ50UCtEMJNDo21egCflcs5/L7bbStcdOGIcOx5sySASAHAKGFAFJ
EutpKWJsqHtl8Fj8Lgf7+96xLYjfCWAEfsrQZq+t5x+USMdOrrxlooaB4KpE9e4RYPnQjj7MATWy
uvhFe6MzlEa70wAIvwqZNu1yPasTwNn533b8TqpkS431b1wRTP0s0YPbzgCNfVp9jtRPur8Ndf/N
uXw1lDFrYKgdFg0tvETemIdHMnJ+8GoeTTGUU0Ai+hUMGqSO7eHAFSXMpcLr+4efb6CRi+lKW0Vu
Bpz5+C6CyYdLSy4cZ0+9g3FrZ1YBfrAJQuPa0Ck+N5XAD1AIM0dgAvduNUJ0eb6eJwv0fywYDKQb
fp8P2THQDG5yr3RtFnkEIogaC+d+UgDXEe2IIGheyAMi4GQR390qicd1QN4LdRep6pMbYTelhFrh
1ZhkjM9O78RMn2xkDQHt/Nnk3K85/qEDZRFv2+c9kZhAKAz+lRt699hdyFkQxXlh8nOMI+T7F5GE
D53D1nX7wN6t0AgYisibrVmvTsbcif+nMhLH7zQBlWQIZzH0SlISwMJyfHRF0pESQGa6YmOYDdcr
dlmXDjkcLS/4SQ82ZcO2ketoxl+Y/4FgMzw9eFi+iEJNFd1Pp/6ReUKysZ0ACp0PztMTZ4zewyDN
8zof48Ws3MlHcz7Dim5h8ILa5ncP9/QEQgQRjy5A931qEH63JBDI9fRtE+keOdpoj1mClWhKIjcQ
ZZ34vHZYvK3Rvq5afa3i+CasQlk9Ql+9t8LSDmxVQ4uZ6q0NhjHxlv3NK5brPjS4icXud/xhm05e
50epaeKTl+6b0xoeaqqsiTDVZx6Wh/M0dFBBYm660YNsVIAuj7TSxm/YgTr/LeqYJygu+MpfefiC
QBMSX8hE6FtnXnPmwQ9pMZ1WiptVdYypMeJHEbnznMWyT3DDfKwymHjbgo3xXVQ8yX5sDjBjp1Nv
C76jzus8Q2RoFW9bLX8JsLVknBWPV0J9XUovrGMivs1DFaCMVPNns9bNKQrth4Lk3/e2q1Hdxp6t
L27HLe/I0F0BEG21u9kZujiMmX4z5qYdW4/czLcMT6zn2jTiw3oL7DPe5Y0FTMoTVhvu4HXJEEWB
VZ/30gQT4yOwU6vfXFR97w7oDfCCDTjOxPY1LUjXBUnHVzIBMbJBPa3WckLhbpd/fpAMcyQboWG3
FcWv/v3Xxm/3P1XhVQfuySWpLViL4qETxj3m5p4Y9ShJOK1Uk9DclKJapjkJqZIjjjmvvn/PNLIo
DlZ4S4e5XFxoRfyakKNNZsb1Q4TIuAtrUFw7zh1cf8Ytqu6H543BKeQQv6CJUuUKMYCIyuWfUiwr
PdZxaclZDT7FEclZf70uK+Os4z4EdvrQvTH9xP2hGhWlAIP0jTbA6yxzX48X8WmWouB/7U1WhLDI
5Mrb8KlusrBg+v8cc6GDdu0z3mxCzEEUMf/CL+uMl2C6pwymRTnPIj0ClKuCruuBMA+bFnWpAkax
isSU5R5MTQ/0tRoJwYuU00X64Oi+8eIpi790jxPmvdLN6UFDGTWo9fG+rRH9ttvjr7qvuA/kn1e3
XvSN8mi1CYp0K9HLJrDuI6ykDN0vUjeoBeOxDMb5eHpPgB63tQNVs6shfvSCiWRCveCE0Sopvmn8
QBLA0IU32Ap4u/2BUCvRAGApglLcywy0hKSvGgaAMRDXBWj89Wl/bubIZGzWP4YhwYtBQEMlvf0E
OMhhoD4MbZwrvXpw5W5x/8XEUCljEEzbc1n8HO5N5Eg5M8A6cVNR0GruqxU4Y//SjPU4Q3JCyzf0
EHoBzdl3P3ELdM+NUKELSv3tB6ho0Rje/9oON0zDsSIi18PYeOn10+KjgBCxM3QJViM5FpcJHOgl
T2BijCRXoeDp5tfCyRUtDXp+Cqu1Nsqs/idBRUgGCdCZZNk/y657LcJEHK7yaxtBvRb9HcwsQ9gP
cgtPzgHEbOtzsTir1tKGCFOkrJwIONoOdasaxYcdbNAFjhYT7vrpnry+jCvxMpd/Zgsj4WJjmE9r
YIW2SLfCe4Fr3C5A5NMXbgChi/z5macxCMsIfx53tvHdhq7VS1ffRuMrpacZpBdY36e8kxWPpB7V
ePvC0TVOdwGiVjHymwVyztzT4CoyO4fiVBaCFeExLlqzTyqJwPv5+LiMsPYePdh9TGFIzOyqXa/1
lQzseTKnhDPFwS7PNW0vfNy8vD9Rl/LuXhtY969bBw6P1QyHg7ZQWpzjxSI8br3ZaF5iN5Jb64Tv
riOXlVrNAzlhMQbgQNvZUrGVN4zt/tTNGrHBuAViB7LylX5Vhi9fCl/zqrSho9IC9W2BTAtyN4pZ
HWF7aBudE+8gh6mWucr8ZoIwdk8vQdB8G51T5JwbIr8oodqfn8qVwRFHo8BxxLZ+LTozZTN46In9
LwSED0D9zJQ8ikoCCFYTfuQNSAMf1Mmtse/Z6VsI/6o2ht0Cyu86GnfjXdnQwcjNlWYQopADtfSd
v8JQVmAWH2kIXL3yl/EYepVJHYzAkyc4cxwuvMWe9RQx3qAXnTABIgSQ0Z8/KpSwgvnLlCjKTZjL
IZDczA47Ppro14SAZ4UtwpCQc7KIkTY4fjJzuA/GaPu3GOyGVd3hRwLnkRWQ+nunm8eBeJAI5o7X
VRXsHk1xtQaR9RHK068mSiPEpeUkDj4oZrVfFu50HDLXFU8tqFuzgpmOBHHYTyIGX/pXq//ujyuh
fFvfnpZzO1p60NElkVdhsPPKYYGkzI9n5xvg2ZUWqzRKRlxC4iu9Pld+424RrXlCx9LwUhjkWQcG
hRzZ8yoL+cN8qNyoFQf9DhH4xCOEyD+Fee6qLPBcob3j8bL5fjL6S0AgSmYmMJQ7TNE5A2JyWVS0
MsYC1WUTvkxIAckkOTlFiD62nTYJkrjZoueCAynXCVAn2dDNVfJ6Cr92/ayQIRg7vuV5A7YT2uJK
91tCk4+D3hXoFJ2M2Jwf13Rt2/aFY+/GkQqHlR/Dv0sUTuwSOnR2pkgss0VXYBAWWsji3jfkERNn
zq0Cui5hQrdOvAIWWeQTwdUsbA3ClrYclnKQZ0oy8oA+4mqa7q7gvMqUdvJapoo/uPb+gHArz3aj
64+2NsakNSnrZnfdh5V3SqiWYu6TaC305z/mdp2kT/wcI69qDGraPVM8q8eFyp6J9t1VktXo9cl4
IyoVFr3A5RFKtJGNKutacw2ecxrRHREHHIsN85az/ULOkzlO7Tr6BW6Jf57EqS507YwzM6snNMb2
aT3kJkkTVZd+73RcU/GIcld0BYUAFhNZjL/Whgs3RuPSiij0KGveeto1uFp6x9pxK/W/KEcwtKxa
DY027tZGg6FC4VORgui4WEzOJ40cDfzMsBLR+YNPc5kjZus1J+JKiLLSXvjliU9f86Uk0JbT3pMe
xyMS8h+uaFcGnneU3imgSnQX0Z9cO3ga4tKHtfYcqFm8ZZIoyo6cPZausuYnXA3a2CJoCLNh2vfJ
Hfn33+wUwY0/N57q9GFBis+X49wQX3nMt6TXGQ6WJ+vi+vKbIzq4FXYTqucXlMOVfHr5NceLwSeG
WFunCDeZjpjwUUFsNpmVPJ5GyVpvcUjoCSaujUfF+EdxDvy8uZ8S3pOc8d1qvLrk8nG5/quSuY8c
e7e5STOgQ40dL5WnmIEOi7QaT9CDB8DbwPqIDxrmDZSnvb05GhawswnsVhEWhwP+FE5ofBhSdbqY
we2EJovn6MEZirl4bv69p+tyYaaG7WR/bdYf67pPQTy+KTGDfmTTJzOBkuKC1fGwXaUMiuVnXoi3
FmvdVME7dgGPy5+ozp9VRTVvEnIUClE9ny+iL4zAp/fuzo0Bz3n52GLjQ2fbWPMGJeOr0Ynh6OVV
i6GcRus4oahrRL2ZD/v+3/+051P2PM4q5kyAj/xsNwJ+xRytIx86J7L0WhIvIjmPkQecCsdS3IND
r4V0OsEXIWNkFFcTSHLDYb2CznaP7b4YJ45bV/naa4hBjUfD25eTJ5VBW07cNkYiCHaeiN28NvMO
IgX/dMbCz7NysnpPrMONWIiro75KTT2F4huZE1E2BKKTNs8lVVL68nNs9M9NGaNDFRWY4fgzq637
He2HqGjJSxXwGCdfe0SiCzjxbBmEW1XIz/gwqnYdw+FPNrFbE0KS9958GiUtrpgRPwYWh05Fs4qB
aQNNlm6G/WFERyEo/Lbd0NrJOtJNr4RXt/kIgH8K0UOJVfeRYFQBWzw9SEGKhhFIhA+kCDm7gV9F
9yjZ9RHZ17SOUqTv+iFIclygW+lGb22239lLqDLUvyDM4x3J2Nu0dtLo2z1TOFyvq19udvymJnh8
/SAB9SmbgpYKj2LZxCR1ypEDy9x35/eP5ClTqWp+avLbddXbEAQzAgYdrEpPBPcTNsYQshdW3ptF
FdqnTdizu6DKrQh+p6p2M+VVuUnD1hoaR1eimvZ909JlAtrEj3bucG9k/HgMwgGuzv4+SJiYF4Hl
bN0h1lM3yge4e7jvYpvPM75goNjQVdiFwoG83AGTlhLrOJeChjevUuAUizGrhszPkAELhv4Hbiv6
/1j+S5jfz6SPwCP9Ob+0Tp9WtoKvnpxC7Svmu1hgSvl8PIJ4GiDDsS9BbpGv6kGRbOZo87xkdiBM
CplhfSLpKrVwe4wTISY6EFEuHCiUwVoICfMgKg7MIA3Ga8FK4Un6NpItMW5UsMzeQ7Qwv+Jo13VQ
LF7IxX8m4dnUACac2gqCIHyKG2DGvRKOh0gTbRexMf6Yl4cYwg8UDymJi1GTLWsnMG9eXOWJGStk
iqFxiFB/Nbh4LuVJhBdQ17BiT7Ws2QQ2+PajN+E3+eq2d+sfyJt5ykTz0Xpax0WfZkHeGFifzNa+
sEppfFtERbdmgZWqEzyaRMCIm/rTSNY+mY81yDZb5wZLLdqK+7nk+0iup5snbrpj73rFkzYT9XFG
80AnB/QlI5AExi+OSUJhuJTY/Dn/+bXg5cGpFhCE920Jb+8NLMBuV2lg8xmNDiOBBC50Mcnnayhe
DvGhApE4x44ccwxJ0hcJb0VmSF3MM/aptEvj6YiSfNZDDghE+bcpB6oZ/xP3yWFOE2O33W1jReKh
l/KiTaSYSrrOXH54aUaxDEslEd0WMbGM5rVO/3CBrGwbgfmlyTfQSaqnH7vdcJoq+D/+bqUZXojC
Fs15GnHY3jzEynsUyVOJ6wlhV081AmkubDd9Thww4Q49oRXrHS2cm2BLqJApSWWE7HORR9ITmOMg
WhLJQI6PHyY8u8ssqU4yZG3j4HqaN5ErTLAKFBRwiw86e4nKRc9ytl1FiAcQt2aysDc0lALzxMrr
x34QEhPT6fASUOenxoOazJ8ngqywiI1M6wHvEV9FwteSK7PLte5VyJmmuW3X05oWH8i06YrHvLzX
f+qYtT5UVrCGmhp1rGOPBpd+O/98bVmJ8wpMAU1GqljtWrDLOCKfoBbIFFdIGh1qxL9hQ83K5K4B
y8irW9Wu5tYJvwE5t5xBBH1vcJJkW0PlhfPkmOG27rGbks1UNdIYAQNNSd4sQMCeJp5Fe4XJiPch
PCzYtgHRKC+ycdk67c7IQbd5R7Y4tYvWZ237890GewTD3nuAnTSp9qozY6LUD9EHS7s1AtGkbLsG
Z18qbzeKn89FSbC6ov0Jh/leP3YKGSnb48nNTpJZkhNf1cZ+iVpY0At5SlDC3N/sIBNvjltLONSi
FVzhDxl72WfP/6gMGNrbOPOhlxMh8+2g8a5j307gN8eBFUZXyeZVkSw87+yvPUORVxK7blt0TWio
4p6uOsdhi1Q33vDyRdA8WCJJ8vyr7/taj8udoiqibBzACKX8nSZPO9V0VsBoXOWKgglvRsKdXjF6
hUP+H3Qcxet1uUz/lFBVSkpgKHU1XzZn6rxlovw760kTYCNtbTMxpToT+MfsIOIRU3tiAp3vPNSe
zqOkV0IdwI4EMDusoV6VZjz/xxh3hoVkfd5HolOL/Ek1T6oRdckjYLTXnYcUewb18njpNPX0A/d6
JDYK1yQ8XygIA6/KAbmLHCURLU5VWywzrNjBEFAPkwAiPJzkme30P8N23yeUZ/U7mmNHBvekG/lc
vw2ixXYikcWFQP1Ipypg3ANIQBFOvzxcuQ6IluXHQlP1r2kS19xOYLVbXLoS+1ygoyKqdxSCVHj7
VmebQ4qf5neJRAjnt8K9oVjXlcX4QBjITIsaBoPk81giHCZlXuy6NLs4F8AkiJvF+K37mRL/iD2U
Z+y9XoBb9WoWizhO7uD5EK9HjCm+2kpj6wjUmBpqB4Ap3V7mz4ANBSToLnuzNoyRwsJ1nH3ZnCb4
Wg8pruiQWL5qzHLIt6FAV7Q2X8KkBiy/Z3i7arWNVBgcrfnvDaFHtuXEQA8jYy2e14WvHGedrXq9
Eqg8NRszCnQLBwZzpab0Es+K0YGT/GR6xnaV7CvqjhjWBrlfM6yxy7eZctvMM8aZrLXHViHnFCk9
riwLvMkneDQWmnbuqcraOFgy1yT6CsoM/HYoF5N+ogSlRBHfJqXAv/k+QBdyua5hfErcC/+4dCJt
0UH+c3NlmdBqJYgWFygJIw0QKyb5wwU1D1WY2q3RMNMio3wxy879f4k+T0buLmbMqm+nSJ9ukkWM
IxrpZ6edAbcvLlqYiLWrDSBlqQBj5gTYa4TpSpoUZRFfx1cNxHIX5I/qPT1PrcpZlHAbbKlN1gSf
2R+MFz4rAQU/HuAcYndigXZvb9wosq1lHXuQs6rlNzHPf9ZJjJfDLrCuNgLDrGMNDW7cnVu6FG2C
hckk8Iv6KGkfZMWxUZuusOb1ZqixpKV7ubQcZjjIC/nTWUXlx+bsBzVJ/LbOdFoUJp3+H6J670Lx
7hehgk3znjH4yyFd4tuyXyqEUrJaTCUAG/6ljBD9krqh73o0Z03VV1axV2xzwjyCovQhftTX8+Sr
Q/+32HLlTNmaaG94MxNHNHOBYcRQB0+STx/zzrGCalaevQchq4uFPhetjlz7JDIsj0abcB0jV8oP
1SsNd8SBAus4dz9L4jCEtAya4945NXHB3htjCI2/VLyZLg8XypjgwLmb1hn53aUT//PozoHrRCed
+Gewn8gg0mBdtJxiiB3oFQhMPpaPzy1yBdbaoWZjWxpML5mYcaT7Px9nNlFPgs4thWGq9jYPRhV2
VYV3uaiiHNBKLe8ipQ0dWraodS2zksn23g3lz5hHEa9hpEcSDat9OeCn2xPYnaM6YktnyzGk4qXh
1meLwa/eZET+KpewhoCg8pa2HHxussa2thzUz+lOfl+A6UCtJka1MSATN7U9SpIAKq1LuJE3+Kkf
L8R+6ij9VDc8sHfABOhU5aniXCcrTz8G5Mp0Trhx8kbWJzoESJAOh3BQ7aRkpTS9i8NkbJlE+gxQ
SII9EP6cpFFlUuNBGQ9UAEb3nG+fNDjAswlkruaqI0FSpVwRTxKUEPCjnh2nJ1/SKbM47GydiZBT
fgb7tFBu+dTed3rNzjqtAe4XOUv+jwhoF3fj0VikvOCJHRavSZCE3DJLYangJfaXamMCnEEYtRw4
KLAouc1QCUkUJfLIW8xdOIz5QLFGKQFLVj7PYlOkb3IwHPC5oE8ysAUxEl0pgYBo9ph04l+6vGBp
Qs5ddd+pwaY+8XNUwVEubH3S/7RVs0k3ZNhuNXwWhx74ZPXPG3aRMwnL6KqJlqrHjIxcK6kvyTfT
Mxet2nSzvVlcT9DZy1X7dYfHFQuBkXNzVNoQnyTnXHYXhEDFlgH3evAqoCnUeERNEBZu37JH6hUx
DFLeUsjnnXuufOUvOC58CU1yIxGxU4Y3jNFDgPDkqzDaWJeB8G0wSIOIffv0Oa97J5jodqy1RAy2
2beqAyIg4m9FlsrkYW/UCC/g5ZoYXYdxUvY10pdmpuPaSJZk38VAbPX/cwumSuCC/yspB3hddnnI
jC6hzwcFxAT+IgvTkbdhB5LmNOF0/Zwlj4bzLWkX1OZua7PaJX5LkdngcX6Ls2dJEamIYH6OnXp5
W4aYcjH/VV65ioVWdOdKXlBC1a0wta5xLzPs/MUbAR6FdFCrhRmX/R3j2R0IRVbwQKCVNcXSZo+H
deeMe4C254bdPoVeEpImYtJtKmErU5OSBwbc/70WaB6emZO35E5PhAPsZHKuvPgvsPzwPqPY9n9I
29zxzrrIGkkqB20OMYNNYd5RNjJwuMm9s7MWevrlNRVK++Pa8llrWbZhxWA8N6MDYwJmi84Goonm
oLdNFV7Yonr19ZBEX3wXS67q5dqHm3hNgjleOXaJfHZl0Mg/0L9tJYivxyQl7SL8r2B5l9F2Zgdq
eV5ZT7EP9Xe3ewKzWBV7Rlg412OY0v3Sboq9HJj8y59JkfaW0aR8xFfksG5Jsb8A4JG7Xmu8CQRG
dKDJNHjMJYW2hzGlT2RqHihsWsS5hmWwY9DDGZi3SMjPcMxFr4j41YMY0C9LtpwZlmIDqsQGcSON
hiohQCqKQtJghx7W1I2nxN+xLjIL4IP1ejuBUQeloUQSxoK5SmdHTBEdfTcoXSjBen9LDGb8hfPA
brcYVH/AFHg8m6XjKcS9P7r4D42p37kho89OY8QpCJxlWjodRw1tC8t0frPzPI9BFba7bJkDFyJk
2oX9uN5O3h3PsInyBEEDyxAOt99qsawv3CQavEVP1BGB/cInYggNapZV5B/KUSwvHCUKKBifoFTJ
Xe0IaRjzXvtgcYbQfjNgW7SJ+1ZWfaZu3JSP3V3Q5MXQ58OjBDTm1NWCkp4lvEr9ca5l9pk2Bvnk
JnxEOhESLVC30KiU96SXTg1kaIQoIfBWEH5FrRCFdNEKFfQFWWQcDq3g9PoAJrm+zOqDfPiSMjXj
Eek9egQL4gQHIq61JC4ykszm2TkmdZYGOlHikITalqvvvuifJJV8QS1GC054w3W6q2G0Ukh5UmO8
b4WkBZpN+B2HYyRgjWQN8z2QZiMJ9K9I57Hb/b+UTMDRlqy6D2J00f0p1ee3n0qBS9CcfpX00waM
u/jk/R+5xLV+uyGo2wDRbys0CCyY5Ub1xAepXqULbcxJ6apW+VBDv9cWpE4KxGDb0pdcGVx7ETqQ
wvwtJQfSsny35X0eZIsxEZokKjWjaODoJ811QXgL78HKXvYhG6AL2ZV3n4XOWRYQNxQvBr7OIcrm
bNDS93jbb95Iv/XFKVQUEBX3V+AFdUlUCoEN34odHGreK3TKtHNv4ME8LQqDe9/nxhT1AHeoBwDe
yupVo7tbYHqXF1SvpRlx3hmWWpsvDZYR3W8DfLwuC+d2QWFmMrMtYyCOIXQtvvzV5ofGstEvnRou
4dj5aOv0qjO51D80NTOxuz/Q0Zeu1I/a4K/RpFvwVL252F+WAOyHLI1ZnwVzinNAxX6tH9LEm3A9
7rHpApylka5cKfaE5LULCQhkOIFuK4j2clUSlcZZnZR6teBjrQ9EhpsjEYva6YxP6iS2/yKo71m0
LtPiwGvd1gl2+5FZsdnPFYtC8BgirkAK4AgFNVvKOiD1p6PJE12clW75aDYus0HC8JLmOsmH1/GW
26ultW/TmKJqtD0WLdeRKSAp9lpep0LH3v9YxzxIgbpi6IQgMWUTMzyfWtzZIVBPo+QETcO9rLD7
aM851DD8U4//TP3V5e1MaBZT/QOcHJnoiHz6HPW6LRqU/2NnFPvSSj4adl1Hi1Ws7GpXFkh9lOyO
H9efYnjZWvG8JJ35Z7ZkzFIUpsEhC47XcXk5LN4qFFTepXu1pFMiEdZaH83AaxIGSPNuJR2VGNPZ
vsjJhVjVz30jevz3IrYAR1JrzzjJ+YRxR4VSy3mAjmmBbR1nBvGJnodMzB7BmXhQM2vNaZVLT8lf
AJ94rz7wcCIId+amd5w1uJYS666lCf798H9Y9/mkh8lG4B0EoFyQAz9lEaL6DO9ZAi1nrkVPyxvN
Zb9wPtcDE9e5XXfL/kcXwhUdycJJMB5/Is5clWMjYF7rDaLfYINTnuoFvJiEI7DyJ+8EIXE0qXo4
6VvTumFL3qpw8PwvoUGtzQK+biRAqkqNcFUfqnJ/VtYq3CkxZElPx2zSo1ZT4z4m6sKZPIxvkz6N
UCMUtuasQN93njsb2iW8nJ8WJKUeHMUyARFZou13rR6jHicDzg00MKjgkDwW4x2Oy7fG0PbLqkpi
Rs7uGrXZiWIel6hNvi7yKCXPaZg+8gOknj10ynI0UGrNj6r+62fy2Y40z7SzFPOCtCOO7ZeozzQK
SrV1W5oprluuABWcArfzJItxHu1/XwdGgneoET4D3Pe2ZEdmp7yE1bQJfQv06CJsByMTazwcbc4b
3BA0ST4QPLP1uFSb3202soJ7V8ydYLSZ4MFZR2EqCWjAUYP9lPdrf/eGgZ2IjktBaAoWpMqyhk7C
1aIPdF4n0yTpOUmMnU1UaVMXUYV8GnwOaG/IutV7NiiVlXvMn2u7qWW6T8yAz2ja+PNEtygjwvfi
VbpmyI2awAHtEsQzbPR+MER5Q34FM6GcXr6NpcbtkEXsiRy8piHNRqZwATRAYhfVbqBO1LmhBN+b
uyRKEqXT8YmRMZ/M97p1cmlJycZyoLUSzxT8xlon7eJ6rOL7xpZByRdl6TqZDzB/lXDWupQYjcg3
oRdFLZ5PmTalLJl13ySbxbDSgbRj0ZfRa/IAo9GLkqCByvvqdbzQrD/1sCv1N3Lab0Tq3FUgrmBK
ecKOVbjQa8JaSw/peNzpqMvpMBTCpcckWoY6ZPJB5SLUalGWO6lpMPiM2LpfzoIDTmyp+pgWaGCX
no2t80LnFE7U9kP9AHcH4MsoCGfEhO4jvNc064H6MyW+3FAzlNjalHthw9VwExflJi9o3Ok/A8lR
1fZFNzMRAbzdoO9DUpKoTE5dQq2H48O9TY1DUk8QdHxvR0dnfDfEik1whFYUYMcdWJ30l1TMwVrt
u7JAc/eM9IM/4a5lNH8fryG8XoiD0T7DA0gUC+sLfxsm7Wdh4CXr6y9eilSJ6ZUHgyAnIGJ5S4P1
o8thPxXh/HlRffiNlWVn7+iUxAgeS7R7UpTBRCj5KBn2qSF5SHsWVN0MOoKQaengzpBpl4tEqPSk
A9HylcHGERSgM/u1aUwo7pqkFlI/TY2GL+EzeIkwr0eLXc4bY+j5Buzx8U9D1f7eoGXTy1kBJhun
YhjMIhiUrt7Yne3xsiUFARkjl6Bk2Xbd5I6RQNzIl9gXcHWgWGUP5A+G8GMmktz4ielvymZB3E/l
pLuOe3qjDP3P+GLpp+/yfIMHVSXTgFPS3qPAHc8XDM2218tmq1yxNFOlFXViEIR9/RVv9daQE3aY
TZzps4nlxIX+0k1mIQ1c4H6JmBk5wrKccpRP99hRYD6QTrhZYahUWdlKl1F1cglYpDAFGU7+4p+R
BqXF+bSw3Pszgnktg3wMLLu8MUnO223aWMqiN/jEagHDbQDgtc/z/KsWr3JaOSMOFRd1Tb0tVSI0
J8SWljwbwFSJGbJOFD6fVIhetkezENjTj9buPDEYJClymhTDM2+142x4jHFQNrNqLaM3yFBbrWbn
CfSfdpGwIEt45p7f+PAU7jwuIfiHVQ30oKay5E/pX5SqkhEvdaynLgkrTkYumuvf19OWaK5P4V/G
Vb5BLJeb5bMsGk5P6cd+7OHO/dTe8z0RauxATbpsv1vp8tTfb9MpikOfw50MHVmA6Ekw+n/KNvCa
O3/HfW7PenjyBQE1huNuH+wUVeRxuO+WE103Kv5+4v+7U/6IgkYjNYu4WdZ/rwbemR+4Q/ktyQ95
QM5OHpd3kxLGGm8FVDa/toOyn7tP3LFeICL73xKqzy5fPoVjSPvD879tvEVB81itUKSEGRHwg95E
FcY4sRR7ZbQqIWTu9dX87yxqsrYiaBouJ97ZskPZx2G8KymyDxDKBtE0gpvwBpKtt/wuFOQapXCD
/ikthrFWnyjJ82sopybqnakFp2BA43CvzJUjUX3TK1pqgEzPIK+EGxMI3MUt20xtZOSToEpPxdf9
wbHJYECKtuFddqhljOUE1BGgm5JGCZ8gxppJg1xHfCmlqGvDaHaNxFvOh4HhplCrqcFMZZzQjNJo
b0MkhXlSS/uL7DxWiQQNdlZ5coPqyEYE31LOOotnwwaaRxL5sdk3k2/3MzxjNxaAwajPwYFoKviD
NDN8VsB//izIx3lPLpcW1bu88ztYb2pbKBGkEpvc02mzepJDX9ICCH60YtgIhrr2ZzGI0d4Wftjq
FlmbmxaFd/yzQDjZZRF+eomvbsEHUyvMWXjfCxEW8+bxBv/JIWrDcsdZuadN+Zjv2TcMULLnRGgU
ZzMEL+vdPxZtMwj7IVELj6betYjmGO8sUbV6Iu7Igx+68f7gzdE2/kkg6NS3/QyN6P9BOb6R4Xz2
4WGT2tn5R8FjTMkfjEdkUQeKlqD+2KxT6AFE1hhvkZMNzz9pxQ4Ecsfbc7HMUU+K7Q3ddemajs5q
w5bUKToLjawtM/z/swqGXf/kUcSaEiUyXDe2RdxGju9l0eNh1F5K8ueZLRQODlqtsdgqhj+Cj+yF
N2p4UFRJpiY4+cbg4xancyODWYuzQeK9mUgq+PE7+iQY8V7cnGB6E2ZdXG3epKDorV4782cGZWEt
DuCbKzf/JDLkpQtuZmrOADsVDF+JVdQAJ/6bDHVVavS3jo2xAidGgB3ngFppCcLXLOwqwDUufeiA
hC8V4BPryW9Sq9CXUXTnFYnyNKpTiw4t1gAvPD3RN6uuV4nTtwPfekS6Q5059q73qnlndei+aoKL
8aXKy183GMxAXk3EXSUUMpxrmKiO2KfuT9/NS3lvOnvEE8pZz0anD0/lAiOCeoXU2ShmOKIZ/f5u
HbkrhAFZ65aOkdhYjZjU6WzEwfsnub0YJl6BN5cT6FiTPtsfYq9z07i7CnW0LjKDPTcFvlpbwH0u
f/TdFiwWAMzF9pAR6etM6GRQUtWPFPVoJOhg5gcR/s9qApD/+iUKxH6pX77l4fcIBa9jAnCfz5Wl
NPcbBG69XvvZbXz7TU42fSji4FjdzTQvbmTYIWMlkczi74/40HjvDpkP8e13HrF3+ziPj/vpecPm
kkPO/1hdDtCqSuFGnfLsYXfGbxFb9pMa13FZek5/CAY4zsBhroViDEza95QASo6kxy9W5UR2K44h
cjuU2jT0Xvm98EZCRoHv9kdB2OAWIwSUx0Nk+RZwGXhLe1lH5bzg/g6K5F9Ytjak3TNGlOTwzADS
8Qi80/VcwGR9SmbbdO+PoHKDFuJIU2HLBrt5q1uM3jp+EBq9NbqAJ47H31YsiQxgI29ZzbxeQFcT
mkwsddF9+8Yc7YRbzCoB/W6JsZuNH/Ki3/eWteEmHEnxbF+6ceAKBXVFs2bo7zxZHwPXmVf2lgtC
jFVsrB6baMYu+The5kxIcoSsUUcRxgtrBfTYMSiTG0x3Zx0UfkxvAkzYWRR1OmshCqzsAFYQJNqT
2OM/AqjI2V2Q/gPaA9gP9ZsV6bloG5mQj3l7tihImvODUC9Z+mIDG2fl9y8rC4Eyod3/NWzoA8zj
yNI3/7PNpJWG6+K3UEkDIMS1DiC+heuNzqjgJKZdcdBzoezG/rGFBmjY/Nj7LI1WaITN6S/Cnx4K
Hk5wLH2eTpMA3tfNCEHF8j7yjPk1uO/8dUC34INf3lLIbVWAq7z0dap/5OiOnb+Ttckk7tVu+ORF
c1cqpktN6SYxgE0+ene7PnTmfDw0ovjtliwq8Pg+KjFFsrQWTNN9tsXUrBZ9XblL3s0dvB11z5GD
HvQzHIO3/MAST7k0y/ZePppVmB1uh4OpdLFVy7kfj9zgrgSWjy2Gx89G270SNJZ+x9lB+5hgX5i8
0SlMatGElTaWtxtrIU9DnTQLbxHkMZUY3uV/epgbLEDCwe4DXXv3at97i3PCgICFY10SRz6J6wi4
l5sPoM/UNDVQnLfOjp/cSjONGltCvvf2QQCkuemGUWuJYC67xnub1dLfIHV/7MX6hl439ditdnU+
q6POqGNrwmtQVy2HS+TjvXR2T+y41F3QyOYYMY1i8Q7T9eILmI/u0is/lozWy1eZQM1vhG0puCuN
NLJ65ebwG8hs1oRM5PV0U07ZMMnDkxtqVb25OvIsrzdSrOu3x8zT0x5QwI5GkVojPY3VrgXCHnjH
SWij7YN2qOpRoX1WC1nor9O8YMa7ym5vNN8L7MkY6g+gjZBmR+YEsok7rrCZR0sQQUdbKhx9QPuH
680NwKRlWMtAadkZjaIV2yUpldUyKkSCnXw2JPKzXx/ykcHuuznnzLRNzyMHiTn/rmFGdWnTRhkG
MfeKiNahSaI7ug/BCgim7H0wWFzQ9Np/EbRNG1H4DfpwirWHjo1UaT3gbAdNQgnFVjQ+w2qKwnBn
nYaS60inQHO4ferfIv8R64t1FrVGz+c4fIfnkkRMTak+CpiSwR67SJZEyged3ugmtX2DV81HU8Qo
4s6YolpHq97EM5V3C6VBmy7rSY1rJXrRx4jm6Os/svVY/Lgme6t4uablawGnQrz6WFDPnlMjUI4h
NGbj5gpvM8WzfWuDBHyaszTXMkMtKscY1/0bG+FFmgLdPPbZaDZ4xgqLAD6izV4MM6fYdu6QEOXU
4iA4mMyqMiEcsLGvZnXF8U++ox1/sAkBsuayN1uCYy6Jd/IGDAGZ9NXBeUWXgHzEkUj4o5dcGywT
wMm4kBoWmJoRYlCvUjy4odSI8rPjcE8su+bCLr+53DyBVHij1sN5YlGPhJxlEHNE1iFQtHbUi3bS
GDB0p28REbOrabi/cxhH4nLa03WwaWkAtDeHTcwZfeXVCGLqrfUFHLvcilFRxLHbApUvSWJ//7BX
HvARYhvr9oMnJa96fiG/nn983Ir1EgRueDJ4Z8Ebh1K69cd4wnlGIMpzYOZ7eN71yc2ePJGutVrk
DuD9s8fJJh5Ur3eLfIC9hrKEtv2wEh1RW0kfxTyVQX6qSVwpVZsmDzcG4I8rojCWyvPyxgtohncg
lZERpEBFRfgC0L089hbv6xnEOyCLVS4xbR8hgZEUbQSdoO+dT5XRm7fvcUn3q8Yo4hlDtVkJIEg2
DUO7cQT2NjohIQ7giN8cjo9c/k7MFiaJs0SJjXwYzSqjQqhNoqE7mN1b8vPWRyv2T81qmq7B7obb
2oTObT36B5AHWevfrunb4zQLmQ9txRi0PwgDrJEM+WpOymrs5xqEoXjEWX+qQF8lBlNi4TEuXbaM
3noDoqk22JrNSN9dSltxZiUSF9lnJlY9l4/p5MfOituGIXP0m8io7v2vST+f1G0odMQ0Tz7istDi
v3s2Q92KyB3dcBzIBTV18YUxlvgrgvroZNCr1xN3+kuhZJAq12Iw+g3ziFhoXqYkIAS2zFiluuus
snxSI3pd79CcADrNKSSwaSSY/tJXj8JuF1eau4tboBWXZvT8E/VJZG1bpGsn+t7biLjzwjqtWXsC
8gO6WJXzMa6I8p8n2Z8VNITqfTaaV99XA18BIlGXVd1Wr8ng7LZPn2KKsinaeqNtrTy832UJyMke
xgUfNSEGsGcncpqPPOWYup5XYK672VBad9JCxaIQ0OqPYRxZrKw6smz4+Vj0mnAOUx0JJ+yFqu64
wwwi2vn20ke8K95SxK86leerQ+TF0pjGVH4nXcPtdpEfuTyC0p7RAsREwJKMz/aIw/3JPT2PbBhX
+ANijkhB3cbCBL+zwx6iH/ZLDGLto28C5K8ksQNrxIQ4F4PKC9ZTOA4Hgb+8Rpyw3+mNmVtai67g
kXJfx/yxfsYmECob4o7b0hf79l3jXkrC4e4rVPbx7olo6+QrtT6NF4izNSPOIrxBnDWJgc+RihGr
7JDKnX1fUJF2b4pS6YH7A1wn09QRuzM7kvaB5Sg8mNlXzyGMESFYOR7uID+n46ZhhAG+TdxJzzAL
4GSDhpYyg3/pVBF2n9UNvV1pOWTdoHfECUZjTboHaUb4l00ZORZOdRu8VLIXHSkgVCjWqiOMKHda
dORJvZo535SAgeY3Hm6ggeBc/+sv0Jl3NmQum1uGIyK0dlLqX6w/m2Zh4ai5Khb66cLkcI4G5Uhk
5wb9ZiRzp5cdfo01R8zj/mLYyMvKlvXDNUvGKIlEoY4l10ZHOy2PraRJp1qFg+UiSIRx0KZKEnhl
JQ78izlTI2C1asNAZzynpqMJOYi0xdPvCiIz9XIlOsFlBEFfzYWHxJJAfPbz8lliFduLfhNo6wEd
DxMyo0vAM6A4KrqvSWp9gEqN7GhSmz7DF8+Kxlsqsgs6UTatPiOgAYE8dfwm+RIrgg8LuNAgYpKL
DmXCpIyZdrVxAhtNrjAGcDgJ0L50SZeEQmEwz4FNzF2Q9QnkPdYsy9RVMOsR5Oi1twEd9iQ+ZIIP
wCv5N4OO3s5vXoU/WGGpY+EC9swVX9u64b6y0t5d75BnC0n7fL81cNRC+nM+4XdLLSesRrVNW0J2
u0GEJFxfLS5lQsWEZ9SzGTRg5wNF3hzUdFwOLlfkFjqqQtKAZqQZBij+mxCYPPd4+yBTgBMPDBUS
5JTaYhWg+R7rdAf7uiFUZyz3t6srKbgBhaEWGOZKJfQK2txRBgBnIh2rObcY6kSF77Pfq1NYi6ps
AcEgS6GzIFzzwS/KAS1Cyhos1u5Pdp90M/5LBuG8PnsnVsKIjHDicWxuIWNBt5ofBIjAPmXLyzbz
AJzVNMHYgayvXC6JOrkPK6G+4ousj6Ps+A7/3h0lel/C/6Usf6oJ5RGeNR8rf6N3IcGLoAvYPl6z
fSaa488NdxPIySjVFQfFrQGdYtzfh+Z1/2LRbLhmPe8vu0cm5r9rT2z3EtEEM75XsuN9eK6RV0cB
+6UzkQ4UUF75jUbMceIVCCXkBNfpK/lp0A7M9vRCFkxwyHDcxpI0ARHzCtltD7NL8SlmAV1H+5QI
lFhnwh3LIKk47cybY714x8uF4BXCGcFLAf6oUm74nneFXXTjRZIJ2eQu4wdpQiocH61CO8zXNVm3
V8+E+vn+JRsNKhdgDoX/yRgUL3rE1J5aehcu4G4MeBaj9b4FW/5/GAXAp4k3zn86A9JWRzAwDtz4
iJ4pPXrl4hChTsgdC1qvdEhdjFNASoAZM1iyNYvtOOqNVxunck9V0LzWAcJ91wO/kV19KiYikbb5
xJ/DZmDYLeMyO2JvPq3Mtcp2qV7s4fWUrTk01e/0O7SaKSjRKfxlb7xuAiNF5qS0bCpDVuA9lM6u
Qm5sWNq4RgolNgyGYQtoHK15lzdiQfzHov19yUqs5iwjdpSg/AT4RvdOVHcTVqQDvWWYF361Leee
U8OOW58Zbx8TsTbVcw5n00TyfYI5IQIwUDFczcjNY8P8w2eYnfWdyGDVcAqrVBCGkgXAoqgFjZaw
500/a2SQW6PP3IbW8uASvmSv6kTYuE6RrZSDhvJBeR9QvWNit9DwxiIGg2kQmygNaYY+dpnoNBoz
Ipwh9kQdR3rJ4haEVq+7Bu7ZQyNBnTyk0UVJ/x3pPHzTJCdxmZDRjwnBnaj8SqD8OmxGtgRlthpT
Q4uN2oeUQL65LRQOQaeTWxpH/QVDeSFjRVgPmo3b8lddZE5kt1DkCAS3/dUeasvtY9alPRd6WcLd
o2iHqvwICj59quPrOJfhas4XKGSxEErylKQww565f0lp500qMHi45R+Ijogcv0YLUA4RqXtdcvlt
Gy/2hhVuEwyyjAzXLMNSQkU+yp+kZIHY0r5EXOzijFXdk5+JxHH0NqVry35UrJudh6DjVnZYvCYZ
2JlDkVMfWDp38c0VHB0pxl3K+zTYLHDxCZFFT1dORszDn22/vayReK9vv+d8GqzEg1LZoyMtRw7k
HHsUv7xd6RC+S71LhMVTpRzJcIaF2LT3VmxxM4gTzMIDXVlqym6Vz2wc9mzjS/CjY6V6hBTOxQHA
nJLgGpAo5cpAmsP64HontimIrpfLuL9zZaVt5eeMWI1cYeHQO/wccKLQyK8A4f/Gwv95GED/8FZI
psWJEhMk8Siou2VjkGoC+HRPYk9hn6Lx7KjLfZ/xLtXyNUL12xOeoYuEDP2TjBEgCeDxbU0JzV2y
qlBACuN5245YBCnvkSq8EFG0SKC94njWgaMGJESBZMo8xeImrbMEuVPzrmoLOzf/uddV+LJgCmh3
pW+LM4QOY5WhX4LgjwHlr3YeKsD3NwGbm+LdMpgoa4TcR4Crgb2Z1UPNcXqPi6QoFPkCFt2jeLhO
+9yVk6ZjJ4WM9V+Xispg8H+60E0Y+fi7GFcZynwb5QSOCC+eJUR0x5jdRGLH2wxULWpw7KuZRuqH
JcqKrc7GNjrmMUBUmFpeeGTIvXEDx6wS7VzYjdFpHHNwF9IS3eoheyhS3FjxQq+mm7t1M3jjCPXD
JBTyAELQxuk6hZKJBpzO4BXGESdc20DMbhQQB8uOwDciuzg8m13gMj7nfC1pAceJMSIeP9Eeiipe
f3Gllw3NLfhFJwsdUUrgCEvQJvtpxyae5oqnmoHhgGgf70djRUPtxrwszotduGLCEYtvy25xhGnD
DCWLtfFoQd/zU3bXGGbcMZf/FxCGuCxXEUtHgoj/nrN+xwvHou3lFaGer/5Nv8Sqav164mVaqm+t
uxiIegEdZby1q8O7zrtB0i5HEQ95wLmaNT6tWCPYKf9jIzc0ERRuzgHYL8/1z+MzF2H7ybxFWN7m
K+4wEeFE4krM1WW0a1jdSXzOGbMhEif4tab5JK4+Z6aYLpiTJWKuiHU185lY7yaCmsZKo6s3Ah44
fI/OBWSjArvzQU0WTbxQ96KIzV55qcNqG3tKg7QByoqahnpbNIRgKMjqcYRDNl28x4JYBIOQb4Gg
i1wkRPy1hjxeHgOijGEBH9DLpIy1atn3cYqGCUd0i1/FO6owZGTz5aZUF/DoSaF7C9tFbhnyZc0B
eaT7bLLsos+j7MKH7maMeJlTqiwCkdIStvAsVOcEA5tVX6Lnrh9/tQZN0bCaOhxGPje58l7oC/AY
L3AxAf5kOB871xri0QLZooh0uTQE8oyiH7DahI3NlXIxK6in0iQDMQH/2felNyrArLcdh7ZvC2rQ
Iuzy6VcoN/1uoMaxQViVRZPAqjOS6o3HUickWE1GOEntmlC8mnQQFk6W9rHUmq8ofOM00ygKDKky
v/HwOLtUUg2MhkhbwHGz9qaKcFiTvKzo6i19HYW4bbfpDMYKW/U5NE2FrbuBL8b3FXcANnISaWf3
o3+lloA7acGg2kgdCIXxF2wnq7nOA0/BMT2RqEdYpdBZ9/Tbw1zK9/yUpjlxMP5mdNhIB5I1im93
AANaWdL8e5NJtyY72muzwIHO+mstoPwA8RBFSuocdjr8aVc27LXUyWF50TMMlRsHIjGlEBGH5Pwf
wkEPbHiTfCv9+N0Pe5NqE7oNMB85qhjj+nAAPczC6rJxQmQomY/s/mo2EOcDy4C/CewwZh0QNsKD
XWmICeENoy1J//s7NoZmmH7q8hBgEojzif99ojyQlyvDfiZCnHrGgn1Cs1d5A59awrwq3HakX2l2
M2woG5OBoYHUZ/OieAPV/9Nc5/i+Zt2vJsYB2UIx0md0oGTikNsgSaIIKpP6r6N+Fi2XkLhzJA7P
OmEzzDAjujf9pdEOxo18yxFuOsF6uE/PbY57xvnORDZM23Ea5BgYsjS0WlICKNwiXBNoFiX+q01n
PcDDBTkQ6KFX1COMiiL6DOocOBzgZogbga0dnGUcmTY8/sVpTuJ6RAN/p8uE99B30vMNOHVfS6LI
PeAQQQauP/oH74UH1bbFrezEmk3zc9nAafR1QwoP0X6XsBF9cz9rQEcHtBv1SjnGgxUC4jUnGCKZ
klwWrvXu4NBbR7WyW/3J0E94LT1CBirEWzpGimlXanrOpLyV0/hQpMoIZgIKpr434dJ5MGR9fuT1
QlgqQBL82RjS+6c1+p1iGW9zPxtGwxlZXPP+y+UNdetxJ/lZppiPYgjNXQqUYc4sHk140Mn4QLcL
PMQXCM7AGIsCoSIof6oeSWREBmZa2aSzl8RcNr8OUomXkM9vR8FXZ/NyQOPIT82jy2PabddtwOdt
/0Ez8FHJPbZVWMLoP5BPwypMWYk4esujGnN1hVNgWpbaa/dgpO6Lhc2k5TffJTBmoBMUOwPSFOGj
XJsf/odx5ikgMuTnskNXE/e1JPOFp13fDjgLAzWm4+Rl7SPuY2u/+KFW5z8Gpvyhtj1nSDzbtKiV
ii4Nvp4Ac6rT7a7fjqDqrHBJwKcBdk845nPrHxwGSFLLciO/+f9f7oJlYB5Yu/t7PEfRrHErvg6n
VJQzl5dZ7Gib5XLijGrhLVPTvVotlk/w6N9W5YS/x0gwBANMDaimP46JThPCJZi63vgCZt2Q5EbE
AQtbSUX73LUfPIP4/38880Lv8u8uzMGv77X+gmj27on6qc07WRNFrT0fLnYkvJPbYkeTCZxqEy84
KTDeU0558xdZhOl8tQMaGNf/HRKWJvDJfdSq331I1CqGhC7KFrg3kbEW1PDRfm35Wz89/zfcgAx0
SIQxn/bf7FHgX7XeF918Mq+lYNEW7l5dXboP2KY78v6/aZrMr+Xif3O+A8kf2xIM5Er43zC7vLd5
qbFu79gHa1E8RSpm67z2UXTq1OBDMiMLurUIkmr41kR179/w0jF69zmvBg0NBA4ZVwvrrgmoNAWW
v57lmP1vh7RgKs/TUh8i/BOf+uhgoQ7TzPaUclN8smk7DKu7uV5tt/HeRDVoQGTYo9vxi5JpzYrZ
JMbtQTcRAGmrEk3IpyiArknqA58fbQUe7xp3CTQsqCh/su/iDlyt60PL5iYpgg28Wm2XCSPZnabw
u6yIdWojfWJQwq1/YdwP2bTmWSdKSqOL8yoCsjyU+T6EWQJZJQtAtj9J0wWKEu7xu9iSdJFXivdf
fomWPhGLIeGbdQEPtmC73uAtEC0epOiBVE2A8+NBF02OlysuDezo/L9ekD3uq7ql+2tFB04iH0LE
V7tNqKu6GncuCjTCLB95JvX/CBrWAMOoq2rzmMTlAi8VscxFh5IjM7DvDy9p6oQRR4fJMuMeAvYZ
21UylDAVkmUxBhat5rLfpBqGzMvA6aWmFSPO15Qo5OJkF2rFqwTpUE41Ab52rnwvgU58jp+bHmcP
gD9SWLOWc8KWc0IbTfPHMUlNDq5JZOtytxgaxGftFk1jP/+vV1TGn/6wCUK+9JQrizFgLtgvG9Ig
f3bc22v8IJsU2LdHwbyuDsEpLlTFflkRM3cw7RXBM//FNcO6fSk9HDyC5N716Pbb3sCJEGBb3hHQ
uCCUp4mbsQQd3Bt60Bl05rErHR2KEZOJtB50aMZlJOmNa8zuThPTIFeRIrdXI9xzUpH3iZj1Zw07
bJxz55+s+QgIFtg/JtlQOcT+ppyKoz6RetIgYI3tiEuI6h8fbqjJWMqex3A1tGkzFRQxV1SDHsPv
Ql+6514zIDyy+22pR/oMRkSdI9c/QQtg1cf9D4ErvjZ9sidSFfthhcBt0m6PX9IQm3S+r1phK+ZE
3aJY9JI5ifPD01mB3t2QaoOgpyQVy33Pg9lQXzOReIDO8pSSoY5Vw8SKUohGKCGZTpUOX6ogzmWv
HqUH5uLRypNPl0oxkT7q0JEbRwl6mvRzJVTvF6fwbzCx3QlcKwg6MefogHoIg1MM+7UE4e01m9rM
9kb8bjnwydqw631UcUW1dETKGp2ZpZdoJQMJynmXcyBoSgqf/32gAggXGxNoRVhSoHn8HwwtibjC
drpGlc89gZuVgQvnTJ0wzP84DBH9zpN3mMPdMUdZnzJTYFH2qKYKoEVftn2ni25/lWW4Dqr2SgAu
G0Bq9PTCiqtqbJBqkdYCyJLArn6CnckG99RWe4TgToeayVWZVv2MINhefSU9EDEoDLWfs0lIFH6d
RCOebwGa0lyf6VxMIf4jXqAFM0xEwhy7dUFq/LWtXaDJuprDuNaVjAjVUlb3dL5p6qmi7FnNb1mA
LwVpFekCEHfnQni+9iSUH5HuOiZQpty01lTp33+1op8JgC5zgzjH0tu3Mcq9WLzLTwFZBh0TvMuq
QKm5WZD8hvsxnyRYh1b/E3uh0ZF+6+vFjAc8CAtssL++d+X1euYw+VTi1c6i6sCe3wZDVDxITagA
VwaYdjmHxu9tKikRru9SfeIzNRRg1rDwyOQNSjx+1IG0NR531FH7b2JpfLol72RxUTSm9gitzFwS
AQtEFrB9hog8Ab69RbDgYpyoUfKzuiFsqp4K8wNoMmwrlNx///mTilXDNNLd6MdmeqizDhJ6Cnkc
ZofQGisj2Gi0HebffYco49Z/fOZyt2HcEgVTXTJm9zN98Hod3qEureeoVkN/8vfd09ssf95VA2G1
eD0It/hibSOvnCnDtz5XrtN8bXf9uTb9qWi05W1qDzszJhIOJPQPjwAwpuX3XtmzSvYKd4J1+43z
TsepTvqsBquTq879CO9uw95bCpkELFlFHwXPoX+n60wRCE6/d8RG8f+gid6temJTxzAkB8K6bed5
VAJLn8i8Gu+s7DeTw86GNpMHwCehSy1flTCoj2SU+G5pVhYWEbJiiDT50bX7ZrALCb5JcU7ZsZ6U
baCe0lQ5kyHv3kMG475UEk/fJtZ4yctTKRZ/uWW9GGqadfANJQuwudgrK2sVDa9jvPIDRXJB4uO7
8cUQm9wFzqbJHOXaXpBQC+tDtUBGhMo8pCGjkrIHvneKFWT10vHUhh7FFOgvMaLxER9JR979ajz/
xxbKu3MwgNNjgfCDXmfjZNTkYgPV5fb64j4WKM/yufxGBcSBJrBu1mLTJv8NtnxX1JEN97+J63eK
USBgi/bNIO9iGhI8e5vEF7u1r4/MqQtCvK2mja1rTkF0ols+9KIH5oghTFjiziuuyLoquGIHzcTD
XNsoSJDaS73Qby9k0ozg86DQSbR52UB5ovI5MfafX3bdXLbnKqrFI2Yp2KMO5nQYXgTUbn+eNEli
L7UlvagBKH47z2f5WTUQTZlWdz8euGe6YgVuSEG1msDeE2/vk+qUHnBSjHBOmy4706C6VB5o8zp9
Es3w2f0xaouJDOdHrIPx8J2QMsuoig2ZBhhyGeMhtEs03kXQidWFHm+kpwb1v/k0imk30XEwHqMZ
Nl5X0LGOadeX9xR9CdDToiHKyf/cLM7CFvLBy+OBARiX+w2xdaj4KohoXAA901xyPAvN4MtpqvBR
IMQvra9fY/V90zGd9lpA6Ac1bBGfOZrt6E4H4iglsPYboWZ4++MmoV7qXzEUZwpuxNpVI6lYE5a+
EePOCvHP2qaEcTiDRa6wpgh82gjAlohMINEISPe+LMvLyOQboKeNxENK3evi3uaZs4ByxXbbebQW
p2exKvi5rpH+7qEO9CLhedn2VULyNXQIX3AUtf0bew5/PVjujWDIBgwoEoEmySUCurQL1uBAEdZF
n1i8cjDneF5rao1oZT7vKHmBvzFrO0YjlkK2NYswIOlpKiWEM+P91i+3qGSMv44d/3+tw1IuCg5k
wdy/w6nAQdz1LsZUOl0v5xT0DfUMmejYOO6l5wYPsB1qBaOLYU4CA5kPyqXSy+kvTNQu0Ud65tmj
tN/oigQ0g3Fjq6La91Yyo2HENinnSMcZDkB6ATuTg9mz/8TlpNb9xdSjLTvIwIyNCkA1oPuY7Q61
tJudPRWefLJRn6BR1DKMVPi5D+Dv4q7A80cblqOt1D/ds5hWSeRgqfnPX5G5IDsC12FsZnyo6zXI
PwLUWhGedkT/J5+G+nPpIQAxeNLO/0YnLOnwU/LacgmPIxlaupqnNAU8OlqKf9QwHIbbys2IpTLm
dGtn/u8po2b3BMwS1yZK70osJcOF1lXkJRsjXxjTssuuxvvUi9algrgcam+0lgyklp+x1EWNghUq
jyn4mfey53WCy4Tf67ciOA5Btbu9W3XwRwuvvswbQhGK1fApP4IUCaf+j+CwWi2lZAvZiqGXn9py
6CKBSZfD5q3p1/ht/yBs6eCABhgbWE9q+hiY2Ej1722ycBweEY1o33MwILoDsmo8YQnDOj4SIwPp
PyRom/wryBurXMqwjUrFkVL23UdwVvo0jbI6DPbBIRMpX+paEwaPb6V8EkXqkJ5xTdmmSazdJBZg
4Wt8/jKlm2vcWmwiblJ136rIa6jHSchyTSnYrz5WS26CzEdr23PUX35YmdZv4qEY9o2WlpOtdYZc
uvAmiAa6gkflqxE8cMUanXHxykGUfPk7/C+GTzAWCpjCAMTyAisOytGngZERV1SK22J946rPJfN+
DVY9Fld8MUKwJ7omIOdCm9lyYU8Gz+a715Hl5kHlnDVncHOUcQYtawIJNTLGbN7AlAUpk5GulMHU
ssQks47VOMmantJeGyuzejn8WXouLwSSP2O0+gNPBjnXeOrWmKC/8jp11/yJDBL2iEjtRr9wHHos
bku1vW/LpZSYSF4sgecp6Lhdyr5L7862zIWsH5316Dz1bSzhnAJLDVnXxlsJtzpCQtFimVfC4nPl
qhsNSPEu56GXAAVAHy6BPpvPPEWco651sI/PqTzRhNFOl5JsK55nT+vxtMSoCWOSqtLy/ogMTsEq
cCiF9wE3pLGy9VAyIHFt1j2vafMfE846zdrCnHLq9nkluKZSWV0P8tQymkmXwwCO4V1Cd81+IdFH
hTTiubMup5Awwk/hAIM4h8Il4m5hOmGNYiswaV3zq3q+2SwF4d9v43zRvDpO/HOPgBamYi6pqCIt
Jh0MFwBTUYClkDrqnQRMxw3pWevNprzUpxsnoQsOSl9Wih33g3Jt87Z1LG1lwgkFfdGpdsIoFuOM
89kgjMveviW/NOMQgKcm6MihGCPnHROCg1GYMpfzSo7rcTyjEnl+oX8xQ27S3C7DeIRmYok8Dryy
DuxQEjKNB7Wkuzl9rEHPzyWnbXUfxFuOT+aB1xLX3+/e8CK6MKre+aELXER3llLPVHbtVy91jDPx
a1Xmi8WOswGoS+lr1psN9x0OxMeBeLN1+bVO+3v6WLcOs4H4Wx9B6JrGLrFAbiCqDATh7n3pBm22
EwcgeyZH0u+OF/1LMVm1rdCmsXruzu2GmMXq/H6MYRfM/sVFJH7P9ivHPUSlXahn/7W7itwd47vQ
W6DO2GZIeIg88/eEG1h4FebR6VVjbrbuI4eVyAeQvf/8ErYdO70xwbXwMnTZZXrXFpcS5+sdvfdw
yn6leLwk5UAO+enz62rJlJcHFgSegop5/UijV83GJNp3vCk98e65lQ7lYrtp2lphUeUjs8hmlN27
jQYFSz6NIqSkjlawmdIuZ2ADTf7xYTAHEta5nxOZGZtFLWsWmg+AbgqAq5wYsMXSFCnRRT+ypw6A
RscbZ4lyK5Ru1j69UoDMDQfYh4Vqx1C20vBfnKB1lcyScQREVsWiw4mXfHMrx8QSxRcYkhkbfPUz
sANKw5bwYVPCWXG4wl0MUhBVR4Q5fRB3gmjdfUrFQD0PPTp/0VIzYKSCKo75prs08pHr8QvGskXU
1VHmHU/ZOKQ8wmtYsbD6nb4iCgC5zsjdPysg1ERVHxzDU4cXgPtyALJqabYeU1zxZ18mRYd5gj/g
wXQgbC520DUxTbWJQuiHOM4lRyhwN7kXI/GN5oSEtKkcWjPEWFHKvGhUKWskQeCnqdnexXER96Jw
iPa7MnWtDJl+VdGtWRjgm1MSeYUr5gkhnrXSXj+/cInun5EZZCYxlj/g+YKNRKCXrDD0LcJn9fsF
3BGEU4D0Sq0LKeox63ktdrCtLJhmyUth6aDFqWVrYSPaOFZRe6a5MxeybPCg1nB5MqlGhhCdaq+l
hH9pWSW30mt4/wgmNnxTG42Gv/EFzmwJiyr8xY3V+T1iuiV2Sgk8C/UAet2Un8ZMuMJED4PYI4hs
SHrioPeM6CLdTIMMpzGucgOoy5VM7qHJAovmqGDudjnXPhColsHkv6noMTBlr5m8lABGQ8AQWTLv
GjnjsnYCnvNTClCKZlJxBmzkbnE2Qbl5upzZK97IcvCL7z2Emv8NchB+y0KHhFmkj/G3n7Q9D1c0
2+NcCNW2Gmx7ZdzEw1dJUz85tbqlgGpzSoKBlqlS+qe++cbRd698HBXn+7Q2UZoeSMQWQ11UElor
kMw1Dam1x9e2xFAOUvjd6o22MLap5gr0PGcfBJ0QquBtdWJoWKpei5vRb8oRlPBYVn25foDq3rUh
PLw45n4iOjOJ2555BdqlOQWPSAwPVUDRxWf6FOok+ioXKwWGs4De4xtdWkjy2dDC3ZgqZlh6FQt0
FZXzIhICdFsQsbH5u1yiBVTMIhxEhJIqUaQT7ynfHStKqyqefcA8ERsxjwHMIDuzW2mTQf9hUdUu
CocGXXsUPZz4GjlaaY88ct5Hhn6hhmMeH02qVM/5XQcd2boeAnnN4GBtSIRx/ligyIJHqXPKMpyD
TWobYScYldrO2J+AgVH25N8MWpCBtOya8dBoroo+s0GLc9HcMr1z0nQpGEwQ6lKHqytJaSloi/Gf
halPlyrdheGmDxYhcL+6DjfAkJiS5MoClzDfHMKBrbU6CStx+G3TfiW8nupmUtVHQT7xLhgzApsz
h5ltLJTFKOkqieQuwgGRDimOeM1B0YjOR5xYqDYANspn8/8SqaEx0MB6R8B9qL3unmqJTrOnkIu7
/kncwlP5YE6V/SY7ztfoh2SlnNKoJLJ41QKsFI7+RaZTYRQg4PpUbBZhZCyalgcfEZsdBbNbhC5y
ecpJOjhSxcEjwOElT6GW7LpSpKrRk8Ii7KY+ihc8GZHqbiTEK7tPLvhB+IsIagC5GZqqqXfMPNPx
Z7W6RSa/57xzf42uSF7HAPE/iw9WqzW3/CH4HiCGt0bDTk2eejtuRPsxx5c6zklKjRtn8U4Areex
NoCXlpkijSxGR7dJvAWqNfspYHAD8sYBDJ3inCM3WWdARi+6lx3yl7x7Is/26mJE1iPu0oqEdjKS
TtZDHtY4N0Drjcw9pyUw2xaD4EHTwHl3jHiAPW42UrbSZ2hjmmaesSwCGiv/3U4p6x0bXfjDBm9x
e64C9Lq4+XlZAHXLJeo1HvnBVNWlIA0Me5uwrn0ii6Tn9Fy+H0E5J6oFmVTuZBJ4uR8UV3FZr4SZ
g2G27+9ia5Eh64vfh2XLacRVdbs9a4FKsrcnDcVBd5itakezXgYIg1a6iP1nnQbAkmUARMDsls+0
LlA3NVacdohxIrEI6vCkxGFlfwXu0/zritxCiGo5b3CtqNLWyS6IE8GIT2OANN+6ZppPYEblQsJv
vwNHamGpehfQRmdFNY42GNTp0jCgdr0tvJ472vNWQVJr4Dkudj2DbEMcdC8g4MF27MorNwOzdZmZ
izyO38AWzvzEibjRC7nhMiAp3jOIkSGdAZVZSGJvC94aesn8RWBNytw6bUnJxND2UIg4cZ0PbIEe
FrcZMcPR9ttdYui4h6fm+M6Pe94Xln/uMR/GO1mw2crTUkw7sb25JLM2lk2emVuQiMWSgjn3VyXN
8fMgIXEzSudjNr3VNhjgOFGt7gxF2Jbjr07NahSMBUQDsK6FRVOXhNEko8DVy2ozjhuSFzmaowby
h2fgH+f705Dw2WNAMlh3QrCDILKeAhcWjNjxDVSRTzLv019qBSC0Av6v8iUpXer8tjcNl64sYqAw
0QdMoaCyK1Up+rDluT+7Fp+2qH5eDjoHSV33j3g0tPjdnCRg0hEIOVq+Gh95yfUNhakmaE7pqyMO
ZRSp4DPpR51qYZLDwDWLmzp0F2UfUVAXR1ELCGeuydyFsZ9sGKUdOpycw9kG09VGoL/xIhjm1Tzy
aPq6Gt2YGBCuFu3wDYgvLVX49g26OhBNKAcp+Tf86zjeqp63tugeUzNK7jN5csnhMm+RNHqpqm2R
WbXFUC9iPbKHu1j/HZR10bLRNIs1X5WBkyhJDBZiAUJA61uRfj113AvgPiV2QCTXAcSJ+tB7VCqs
TacvShCFnusnv8TIYbmAl2/4NUwDQUivokWMLwLoTXTibYbLVz5eRwL4oVrflFMTP2nWpL4ltaF9
sKFVAme7x25zN9i4pPPeO02cL7s/qXl9LermNr9YNkBanfJd+27+xoBlY9U76fSkT+MAPY27T80P
zq+QqTybccxZLa8=
`protect end_protected
