-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Z6Q2+KSWGyhx3kE/cI5LpVCGpB3tASah84PNrLfEZqpQ1iOjZkYCkGNfPKoleeFv9qle7/yWnb6x
O3jS4AD6dG2VyskBRpk0Fk3G/F9n4BLmzD2yYL9/H5UvA1gtE9EYkPP2FkCD0ZWCnQXZO4e1LD42
BjAAEAX6/0EtekibgVyjYW7KB0eiyfCMIb4wu4VRgxQ71J4LXpNU7piwXy0L1b0l/0Y0j5SlNxG1
3+lWxIQ+4GDFw5tsF8kWE/51HuzgClDv/LyUwUxYVxjTy8QK93z01J4EcsacwjFbwOvtoEDFRh56
VWEq3M+zE2BZP/pI6Ps3mSTk0HrULB+Wj9lfuw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
S10z7bntw4xlc5beWq52Xv9YUnonp2V32XKnKLmysY5JBUGZNkLrYnv+6iFUQ3fC7fA9O+rvqkqN
MjQmvGXJLmGmZAq52IwXi5jHPB78V36MVuZZIGjH8fCr1wiI4TtR0DE/LK+k1hCddzF+awcO6qBh
0zxak0xoeJW/+Zr72J+mHceTOFdISDdPdIo0hrfHFKuOghaMXcGWAMxcYvORaMklU5+n4mGfdP/I
NwCsv3Js3kUsTAnPQ4dMVPw4WK7quCMNyk/xqCXbuJ7/buiA2JCPA8/mMZDJAO7SabEuMw96XEzl
QbFeNYMZbDMh6llpetOeRsxX5Do5/t5bCEl1NugUG59WplyayQ9IThzEjLL8YfEm09jdQVgR6K2z
HH4GzJhy1bmd5h9ZcYwsziZAGQjrxsajAdJByEsieIeI2OFXPWJIEGKRve8m1XY+Agvb5sHa8IsZ
aNZqsSsbJWR9ivleSwAJNvFh0OonnRLWDd9Tu7t57bWcgezHn+LjrANA88POzt4o0f3eYvp6G0YB
h47va5/FV1WB+istyPhylU6mexmdDvzFdLisIsCf0lzdTfYhyQmbtrd1xqXKDO4xEDPy/hjogP/k
sUqGcQMzG4C4ig/NuB1nkfuCijh5HBxw4dvWMzWzu559OHlcKrurerLxZxFa8m7XY5n9ludJjRDZ
KKQGpHc60bAOqOrIwOxS/LQyfJdjwDvbXS8PEFo4mu/vPUmBefvDvE63uPDwvCG6uSeHw1C54XmD
JtYDNpRF3NHjBocA4DMgkgGIXzruzrFDtcq62PHS3YjAWHyMwgCkVqQHfxrmPjEdETQ9XaRVWb+R
k2GQgMR0C+dSJG59gSzLv4Imq0FQ8/k0zxiH7LlAya/O74BS3Iyw6ULfKQJMObYEZXjjNRfzny5m
SttIDkbyUTHvp/ApScyCyzZ07ZSdR87y1pkB0ffk8DaqZzXUvB2s1L/DsVCS5UfiKqqZw/0eN3Fw
WkIMLbvF7rLiIJGZYK7l1jNk3fM1BonFwSSJ1vnR8IEH0SBgV85arKvYdZATfbHd66VLhguqDGid
at09pXj5vhJwh7y+vRzAsTttNVNVqLv7RsCH3vD/lucG+3mc/r+C7VnEDSCZyZYiwUj8hcMv7hVG
M+tkSUT+L6ad1x51GPmAGPKl7WKVm37Me8bQbd/EPygd+u3GhoQcZm+FKW4KXkFc318km/ypSw0J
1ZhzwehTzSWrkWm7BqOPP7EzFLruMETdLOt5qAyOpJ4bD0MeplVBQ6n+zxYCZTpXfGJM9fAWi+A0
gP3esug3mRSBT8wTpxO5AgiSTtAUBkJDNmkxai76gbN7F48ZYL/HFH6pZmpowXgt/549r2/RAoUj
K/l+XUJkBT7C/RRdtaljgcICCgcv04wL1qb9oXCtDheMWiqSfLoy702cr16+B0iPotY8yLAsFIml
k4Zlzk4QPfGein/SLBbes3uaeRPgqSopzqnWH5aOg1gnhF5fXi98NNPPxPVKu4mIOI0RQjdcEt9f
PVAjpv4cFWrfDIcyBWi5KD6uod3D2wcbWbA5PwBjB5y5Y87y4VU15vGYe2/4he9P06JWhvvp3NMk
VAnhCGe7kfPXo9iKiBH1iceqxdsk0vfCOWbY3/sNDko8nJn+bSCfJBAr8XfWU/rtFkOV6JPOEbC1
s+D9gYqdtxfPT9FMnZoslB12imyScAU3trYLvxHpD3Jo1m2uzA41WSaTkaKr+yqBrgvHRmfrj61c
preYu8yMtZ0XrobhNm/ka/Y2IyAniUHEUErXkxxgTxtJ8AgsuRESwriJ8e2Ks0XOULaWuzSC2t5B
0jMvxV8O4JoTk/Jc4m7mzZudQhxyZkGnfXRTQI/ffGuaQLqllAtQWo4Z9C9ovSCCVBBJMqLCxNRt
NVkFoncy6mEOrbWYlNJndqAuPeWCDaVOA8h4fGCfYTX2YWzfY/Ad+T/dYE+a0l97O05ek0laWNx+
PesVo9tbMVUocogP/BrP7PfmuNCBNai843E+Lw1rYw13JL/u5iHD2vQ8mVG2qt5E3n+rkYC5PXbm
nExAUc/uK2DsZVhxNAI+/unxRYw3H/Z8iXgVswYp1hAaUrv6zOUsjBLavkSjWy7rcKZSnC1Ny5o2
mQatSVT2impVqzvavYw0WCoWn0Mz5cH6o29/jgNRTbKtA85gIhc7T8hzf/GZb4sX+MZpYSZawZq2
Bpl2CivQRHUk1yWBssVRs4DulVmvwYf1R4nOlV4YIz/z/yQ9VtSc6tCLFo7iBEM6naMPqn+RCpH6
xvV/NCCjD++vH2UsLclYw/5aT3mTnA0ZHlkga8HkzrNjr0uoB9AuKQS1VKOJ37cJEzvSwcYVavVd
oBpEP26c5z+pSsFXcOrBNGVDXdzVjdRSrI6SScDnVJIAIlD3W3ND1NaNv7ecTgCrjbIygbSbDxEk
jhSbJ7hcDe8u1k2Lf3YLKYKCDHpauezz8cbuVVyGb4zWzvBd3QrG9/Lt6MxOMhRpSrfVsiOJYoav
Q9inImM+sscCOLoTjGnJSIvv4ldLh/0Xlos0zrLr7rUjut9rOECH4s0j7YSEla0HIdHYvoqBGZYp
axo9txTMd8/QqY76w+k6lvLFssrw/Ryqe1CjWstT8YGfAU0c3EKZUvnfgv24iA/j64jkVjyjHp3O
wkpyE7I16RMdYSV0BSgKA5LIjQh7qnIHFZWNnwm0HOUNewMd8sjb4m8OisiL4JFhhPSw8NdqSoDY
Y82E8ixbOqhXGc4LywI+FnUziaD/0XdvgiVOk5JVOLnmvmNqGdcHuqJyteoyi/ewaQeQ5Q3uw5zd
RvzRLzHlbtjNtIA6U11Bv0VhRZ6iC3eLy+5DNQdJuz30Gzo4pjeB1EHJyGXCPl+Ik+0+A/CENDFh
/KGcB58doFK4F9Hm23r6i8G88F3MiV4LZJ3cs880rWM6D0tF1u32WwWWdFza4Wzh74C8kbpQWNA5
hBSHEgRgW3gtpFdYkqCrMeBp6IvuAPOvbEUje8pJndgOnRI8qMfkZB+9WMHGLeyhwc35SC/mvDTM
IHg888AbE+fDKQ+0k0UacyJ7WzsCacaWST3hiticcpTwv80+8b1tyrbbLkdOklAHGyU/yRAZFAEv
b57SoBgb42TAmmbYMLCdndbM7E1/sx4tMTJifmtASZtqS2m32BS9bacf2lks43d9mrBvsF6n+4X/
V5oHuxSPR9+dx+KoJLHdy5EcEOJO7TFdmHMNe6raeFpHY17U9G87LgstmM+dyGyZVZMMxSatsjOb
qoxb9gw870d284qHKnn2sFvS1aHgO39w3ygOeLORMXYtuYBlokl3oW7/ydklsrGT8xrung3dyarp
zmZlFI+Z4hlxT2u9FoPPUPPeqYEbDQrBMy44zkjL6NGgR/3M2x2j6zaBgi+tiNMn1JMxxTFd5IVF
tF187lGJdXtYqc3SHRZlrpDxUxw6YCIlbiC/ptE92gCsMDo+hxwUKPGQi8EvoeEn4E4II3cbfTCW
Z5ebB0DlM8tGa7+6SZZVRCAKU0Q6yI7Lx2SaFJ0ZCXaNM0mZxMdKPZG9TzIV0NU793wNIsCnYMbx
ceqZKVN+kY9D4NWVTTs1YdEvWUtzDyQGmcjHqQ2Nwfpc5qzZvYx1nr+pIORaejMCAjGYGTb/uwvg
+pF/26E7hTlrn3+pgYycRujbODH1/iUFTGEBfwcLswKS264JvGGZJie2wRlvALg1bRKTt6nSji56
jusBG7R8aVhxzlBm1fYE94zuIqS9QkF9TCzVLs96u5FCDrLhrDwFGr1A19eFAkNlK2iAPJuKmw8g
KHi9pFFX6J8YiIEYQ/fvXnx3/eJdt/TxW2uzr94R1mCILVVKNwpHJjAPniPjJO7DuS+8yCr0gHUP
lPPFeaQOglUNm+oQG+9l+B6X5BEnpaAUG+/9P4RwmQ9eo1OCfa9aXimEHQvDnWitSrGR5CeFiSbM
XLsS34uPRcWghEJnlHbMWqYAbZxOi1jV3/jGFfgRfCoLteaApK3soR/ILlD1fMWJMFDY+9xxXwsm
3UfxzNaSI0tHVKhg9/jI6kpYh3dDTY/zqLi0abRpEjwgmaukVqaS8gQZi9UpKSw78xCAmxjK3jWy
LbuDWqQtzTexkzKnT83HTZm7LP1m6vvW7BrB86BISY+jBKhBxyFSM79Jfg9PIQzfJCuGxNdmCBNT
dGRNgYe6p29brdnCO6B6kWsDFkUKwQuCLGWi9UdmOZuBR+a7aAlAoGJOH7o9+U3baDbmUgTAudjd
nIltuN+Hm1YSQgb40nMLucok4kdyBVeClWDx5OXNzF16RBp9ZOx6UkUopnKBGlS1g8hU2FpfQKHe
Cdy+4eBbwgOqiBDtqqsB7YqipL+rTmisytpg9UGnaqRCFj7HDt7aH6s+9c/CN4slHgIIRS7LrVKf
1nYKrAU6f4c9EV8/PAI3Dk5ZGf8lhp0oxlu/oDclh8RI3yXUsi5MmD3FdxgL8TZJpJ48q9GmSdtB
Cc1Mo15Xn/hVy35gGVYLBfWixs/3Hon1s3P7/E7sK0tmipDAbp/62qfDWNiuLZ7hq24xFUk4f1br
5/uvPxs26jc3E7Ptmg6QRKEFnwiL0whELOYAbn+eJPTl5+5I66i9P1Na1AGDYyA87dUWQ4WDUfyA
1KBC0rh/up39qhzysuqtlNXRmFeW4K/sI/Vf94HPEhbjMdbu3wp1A3lLN5WmRxPMU5k8xc9T7Hai
yaa3BC4S18cb9fKtJx9jomcxIdzQjCxGfcqAGwep8tn4vhmOPX7QMEw4LFvigkYviY+b/dPw4Rfc
r+EF9r1x51H5QyX7fltP1oAROxGUrCHCIo6pxXv+OKFPiU9wOuiOKIs9ymY11yaOx5s602uyJC9I
DhAO0eeuf+8f+O6NYYY5rO+hG/5kI6SyBuKNfRyiqmJSrySJX6KPZshqSHFg0zZo5PhN7wQKKSjA
nKF81moe5CRu8AHJMB04qyFCGfsm5m0gNZRdSdJKcNiMQXeC5Oez9Yt3wc0emm1VZCOR6KiDXn9g
TsF1BRGjgDtpciN1azVyyikCj0rIK+pMcof+4VWJpB0GmDw+baKgHQ2eSfZaY49lNUFiiiM9kpK4
qWmsSnqf3GsYKhtHQH5wTowGlszENN8Fb7jcF6qpSwxatx8gUe9GcLgZJqji3mv3CxQWf0TK3OZ5
QzOm086PWiroRaow/be1YOSWHbkw8etoUO9AB9YJen14odNhcJ+Sdn4gtTv6bRkoitYGfDK0/Al3
bXu+qwBil+lEjz2Bziqx5e+Q9PI7o4OFarkNiVHIxFu6WpQ2kn9LeeT2X7M/GVATcAA/o6mlGEmx
/cjEsDmrY8BrKsSar1gcHVvHsxEb5WSNDkXndg97jFhCY/lNr0dBU+3n1acnujslI8aaEI7QG1Zm
K5u6EWn4DywZ1UqK9DIFfk4pG6l6MvbxyVEh9AcTa4ZSj7+bOK6jrKuyj86m6nz0Kq4xs4klbr4d
iT2QqFAvygwS9dfyD5CzDNN+NPrvHRFW+R/JdFt5X32dXoaWpRNHNtBcQNBUD8oQiqqHJgrOh+5c
FcddmEHAxuxI4t7yZllPoRxCopP915ZLHS0sENJ20FEJM0Km6sCi0GI5t6bPUKNt/xJxDKIvyf7S
4v5nDeCIrv2Jut0WrXxPO60zMUOG5AYdZ4V2dOCwrm2pdjy6IVWv96M9E5ugbwj/qKBLWMNVrSrE
oigLgF2536R5PX6T/pJ6MHutH27EHuhnu5xPdmqYIZRUhd2SUxjkAU/xXCakliLxiL3oSxWINzzu
Dr3VN2L0kXYk93KxkA3UpfJKxrS7rSAL5h+oGKSh40TR/FLjdX8Di2q9Qf2rmK6LloWl6sa8Wt5H
xqo69kZ69wPpUHpJUTv8SKaW8SXoJQv7Y6CIIfZU7Y2oRouvQzdUYgjYBFiULY4/Sfn4kzeLhl0u
iqxP5Q5fKR5bavGepkhdu7UhJfUkfEu2quQ/COgggKqQMoags0MGDpvJKkum9i73n8LCbXsxxVrv
2W4Ys9Hc3pc0dpwD4+ppWR11FTAOzlPXlNzfmMEfC17u4D51pCuUXzU/RXOoFpHKOj4VCa9G7Zlf
d10yFHlVZuPfgCYueJG2jcYbRpC6QgrH8LKuLlNKQsKZs1rhA/AsPr5TfzNtPNQJaZFwII9DYzXl
LGmUA4JXN+qxM2c23vWwvP3FtlLHGmdftArdz67EpRiQLRob5oU5eo3eVQ1Gbp0SmaxazE22F0a4
Hiyw3m7e+LDenkEEA4usC5bgpv5SZ0LAeDBPfRkNuvJ+qlGg5qhGiA+vA4MwHsv0wH7EFdaNy/Hh
y+ntmk7cgSiGYPWP3tcK+6rs/9AG7Wbvz5mS/r3rhCkUYwM5Da8zdBhdVEmWWYNeHyo5IeROfSsp
IQT2Ppt3DWsuJOiMEqrdx7vgo18o8uhUntkiI+j3LF9+/eICJRu3C1XwcB7DRm1MBH9yISFastuO
KcGEeulISuiL6WJEhzEnFz0E08IVJWtl33dndhkdsjgG84luTH+f9RZ2SWKayGESs7I3+svTRgs1
Hrz5wjgyr+zPOVtNBbzei2WU2zneddGZO93LT6KwZgfwdkkDqptjKuYuTHBUay9ET5VdZ353sL0I
2Sh9rcfZWHBQ6uA4d5X6b16fZT3ieN+HP07SMwHewn9V1oRvRe7l8A4oGsGjEXeH5mef3UjB4n5f
POvVuAYzplpR0oDZrDkZJSa6hiM3P6N49Z8vb0bpJHGo+3O40nT+plVsy5xKaqaLiTr8TBzsgZcm
wHSrGJAR9O04+7sAGNcnN7IU8vXoSrsC9SeC3E7JyHnUYSsXh+0Hfw8G0HhvfA47xugZZder8V+O
iqtdP3VZijbm8fENyPYRwoctp+6chGuCQ5uvy3rdqMcYBf4pzGU6V8NFRRUxC4L2IuuBIIiElk6W
qF305oyy5iZAuoAvkD3/qxjxZ/VCWNQdj4DeGgQ6P/Hwrph/R292JEAIdLQocwcFAMAHJS4lHLCF
3Cu8b0H1dB/feh+Bs3nC8c3/YQFaeNFeD1Ummadn4q4n0lBl53Rb3YTaCN93JIfgwdR87yikrdPF
xNH2blnCAJPw+j87BinFVu9ZibKqAJHXkEW0CtQMJYO6Om0H9sX42TFzdNd7tbZN8ahItUZ+9ymk
9xXlxi5iZQ47i6Pdg/fsxii38a0BlBPewPKwbF3D8zxK02TVkQKwNNXlcLbOSkfmheOFfICIIfn4
zx8sH1omdH1wmGlsqpkATPOtX60SRlVYNgoxrCG+sKeemxfJN9NihqSXglLrlvIqDBQQih3iICpN
FGVXop3nj4JIGqv3R4oRt+iQJ/rfJntBymsQ+NZ+9uxxf05p8u/FY7VfqW1Hge0PNGXC9S5rZyK3
pGoeLIQezAUSHH3nkGggdElSlKNPK2epX8ntMF5u6/RChyP1POYadtfXIZk7Mah+qmtW96Yr05uE
ZvxEWZI5s8FCJya+VAZ6wnseDb67R4a1dx0iUysftEDjZU5yukjKcw0Xx8MjA/hDRTLjd9qy3dBV
tan2NzlsEwWpJQALdKy7u9KLHf/+iCXmpxk8hOIpnC1kXyP31RBKI/xuce4jZ4VIkTofOddYiqdq
G9/YN4zCuxrLXTtssTxJOjBwT1sAztveBEX7QXGxEOsj0jSHeQ5jgqh2pOsVcd5v5qdEI8TNQpWi
+XVQH4ShSDgRXxTd+zIJhElRu6igdlSkCgHF6eDvUL6EjePpYbTbvJSoUUi1vdVe2WroVWfhGZCt
iHhsgGf3lr7cqW3ojNhtBU73wDjnQNbEaP+P+mGzn0a1IZdztqj3VBxq84v1FZYEIh+gT+9X1FYG
07qsETcanM5SHqK+DcIKQ60fspb4wNMzZteVfYCPKkwhhV61zIB7LW69XKYvgZJVe05e0z+dHraY
uK3lDyoDaMHUOM4ARmWBWfKfLHN378VbEGrpqjJn4pvopOl0rzT6AHwosIJsWQAB+NblW94ajHA+
L1nO7WUT1QanP0Y5hxWEVpYthfc8SKwF/p4Y+QjkTFneJSf4U4UatMqugeGDmngGmvZyVOxbFf0m
DsSwNz4syAfVR14+Lm9wKB4xu8iJq4bnZ/M7htuUQnaTYoK+hYZTvYiHKdt5l+78/bN/GUSJl7Z8
vvwNM3ois+Fvj8g9ZCEYGRQU24frFQNX7zpunyMqGY+vpDRhRtZ9H8bYdu+FwDSjkE40GpRvPYp3
46ITo8mFs+SQuG/3cTEli6l/ti57X8J/wmF8e0quOsZ8ngycinrvzTNfX+jmuICK0eSYsScJucVu
uHNc/Haij3f3iG1EVJgqifFUzjKWkLYq23BCZkuJ2a25pMHCWrsWGVmm/7O1k31k0eTRB0XQwm7b
1Xy8Vkd85fLb+pSM1WtERCzG/15c3T1DS9BpGUAs056wj4/ylSDVblCji5TVYxdFpicNyYvsVfEv
Tm6sWxsl/aqo+A0CNAid0cv+eqOmNMcWFr+o12S1Wlc79BPwJjvz7iCIhccjKsA4eGkeOwRUbePn
aEHAXNyWfykb5pttvu18aKkXMxZtuVqWVHHb86LWJSBEqo53Dj0xsWRh4sAMwJ1Uv4WN865jyRwk
4gXAYHmnDRbeghZEWOJ8QVcrsCA2YpQObzhNka8KuoemJ/bJB5unzTM2cJbC4mF3pWRwL0iRJI7F
jBudHIPtUqpEXAE0l7DReTh4TaJoGrK5ZyGzbcR+1CmSAh9LlPGtS/AnmbkP/UeJdbX+4L08RdDG
BN9l+RGZ5FYyyqP4wrCnVhlzDIq5MLbtQX8AQGv38fdTLxhII7ASWwMtMGCZiVl21/ZN0cIdBAXb
pZFF6aY1aMPjgKIWXH1//IJBsWPoENg2PTn7es8D4cTpXP4ZUXTr6xVPmOjlwMq5sLFHmtRcZRzW
kVw7LZ6ufaLzVlYmiYPPlmMcpM1eL45pcYx34/3iVAzEWZPv+r/ZQuUwkH5g9WW/3jBqHIG6ddI6
xvjf/MeKVcAF0tmYRisa6M7uGueSganDvADangelY3hDWVwhTSOCuuw11ufMQhT5lAa1SJmBJBty
8WxgOS9ARqwALV3DyxG29xWC3Phng3+8PW0Vorb6TFGKOHDgjXLfOW2+sPN8GmbSNfDolrMh5liV
Xhiknktma1FvSEdUxtYjgBDqWvDv8cAapesaM6vuoHU9OkbqIe8T1USBY6F2YYrYocXacX+LJlUT
hjtDXvfXQNLzclI7VxP3EzxJETzhyv6raU9QDaUzDMwFd+yC96U5fMqs83KJi3R2d/5VKCns6aCi
NXrpLVxMmp7PXxbGxEyn0y25hHuA7jgIQy3kl5/HKUV/K9EnbSsLjW/bEh7weS2MX77Elvt0KGSA
ijBYWLkfiN6OAygukUz/gDF7cHY97LQd9ONUFIcXHYSYHTVR3GcPSf/QXYubRt5R5rDberaq3N4J
+yozOfkBF/6PMT6gyjbgsO55NgHrYsy3+YvkZJZo57WGGAEwduy7k5XHCSMY+VDTlPOMoUA/c3Ew
z6pk+FBEK7EMSMEske8cWEGZX/GVOjadyaGLJOHhUYnT1lobkQjLJseQvAoI8aWizHW7sWr7kcMY
KubTnXMMmoL42N03onwxXRldiyddE6qk/55tzUdDhieWQeHTnbHc/DUFXev6tJRiul2CRSuB0eUi
/wXz7V8SdA8N3OqTIskF24wQwaUGz7hdz77vazqqvWrLbKQAZFFrW30uhJh2Dah0wyHLYMzl1T9A
VmPj1KuvVbrdEtM5h7bUqRA4rhYCjtZ3C39K1pLkKfwOeUrc5xm5vkkzx/0+HQzI6CgHwvNCuKX4
EIrNSa/lNONi4IR3zWkq4l0s/MNGNtaZ9VIFy0ExLGcVapOsmaGYlgpUukY3tRcvcf41WK97wTAo
IyCIhExZFf7E4n07fuZ+xsMYT8kH05DDgNS1XCYBFf+Nqr+01kVovgL/SFtKLij5WbwU3B5mU2Rd
hzQuGzTjtK+kbJ8ttUOjf+o2an1Dsc6KdaD1vH4RflClo/r+qMdLS2jhwsROq+kydtjRkITJWvZb
UCksLax+BQQpNL0aECiXuJu2rRwJJhNDxCu/NP/2MFmQJuPnM0Ti08cZdwNflP8x6dSGocgr4Vb0
cjpqGhe9ndZi8wrTsgC1F5w1pbiJpbOXKLRSHdNAFi5ItxhJ+R0YroP6kbljgA7Fsd/BKcVJcKtw
wHrkw/ljC6vWUD9ReHLz2y5lzb2fpahYX/xWRSc/h3AoZFBr84NaHj0750MuNYp/d/QEHLEcQKIF
n7CxEiLnIqrBplS9YMLlgl2DETNfUfhIwvTyMpq3bFZ3RysOPd5on9TcDyt9F8LbwZrbXFyRshtR
Sw8343VOyvhe51CUZyqLOnig8Agc4pb0NML3F+d2CrxBrb47fxcl3QDdrVaf7DW3LI81+CE2c8Xk
LA0nQTKBwPhVh6jwR+8m78XierBPbz0y8teR2bXhNmeeW11bj3xv1rVNOalybvszzXQ4dAfginVx
t7PAE5g/EJbWcOit67wTwSGiojT1FJ3nOuDgexY7rWbxyLVsFlckiaTltMUx2sUzhZSlA3iImX6L
YQUW/YOaljUj3fugdxOhMAsC3SnWm6M/U6L0p1NGkwDqpMfnjEQh1L3TOV3lMD+CQIQoKZxKCoMm
6/13t72HPFQO2uRFoaOVZCFaptItPhghf6D8ceHnebHVBLkEUwhELSM97Kf8hhXJ20srWTgfypmG
yKfHL0Wr5naOU3LtoXielM4UXl4a1DpkZU8NzHsJEnjEu1H3AKLJTRAyjto6xBraOEuVacRmD2By
ZroGuiHodRTgzeoctyWs1lL7hpLeBurIfChNdB3oxHuPdoJ1y+DEFbw+XntPwgtm1RTgtDbyRHlq
ZVznvJBHOdd38J5l9J8mVTRwUZDWPwZEtZh4lN2nl5K54ygVl8R2JdBXlMhYKNCelmJrmL6kB7NH
v2MTw0qYxwUnBWoL+FBpqBxWPt7IFaB1FJDA92trHU9a2NdpDu80yg0lwOr+isa3P9/kGsccfy39
GWsE0bTf07JNb4FfGcFI1xRjEkSLFEWUSUOOthlwYKL7LRQnP15SZfeWLohBSoIduMOFOUnsdmSn
2CUlBfQBnJGE8fLeCrYMvdVrmVFJfmVBi+9ttHU/AWoN+Fk81kBb51XdK+f8SKCOe5a5C5jwL96w
SLF3qfLaoZ5cXmTHq3k/owM8KlN1+pQi5WeRS/N+wx2Vgi2vbK6FpHsrpTBEANJkksziM/uY4QzT
g2y6IOm6t89SPSWk5xIDfJkcf0i3zLj7lt4BmEkPm+IFgNRbxA5W/TGcVE2xFaSGKTyoCz6LVu90
KnY9FEk66vCFsRjaBJHXAbYU9hmymXr33ZThu+MtvWpePnSiE8qOrO5Aery7y+X+uCBc8lZvpxb1
ep4MkRpexpaxogAwvxNd1UPAq0CvIuysWq48dP0HLfCZbQZIJ0bWvlp2GlooZLD29ENnf5w6Xk6w
Aiamzsx8qF3hksA45hD9qqsd1XOk3TyXFCXv5q811saKAxX38WD8R4DMhRNlVNrW0OgTYKNO0+wF
/mAXoltC6EWAdYEXF+pbctf5pkCtNNOdMhqImMb50reUT7l+QpPq8280eLpyIVe9+Ae7/xIX/WRn
uD02cFv/W0viguSlaDyafcKJLq7yXUxZEwhB8/d55C6iA+tCpiO7sB00Bk6MOx5fEB6rx20+FLv1
d4kO0kPp1hgLckRzT2g4pE+AzJ3aLPk4aCIUX7py/lzqKZl1LsjET6dEgRaeCMslrMVJOjegaNje
C51OtWdd/BE4tlWnofNJw82Zs1ACDJ1pVegn15wgKBxgaR4HeAB5tgtN2EWP7ItRDnWeYUpNcGip
IJDkpX/gn9dgbrkNsZsh5DaWl+QVGiJhK2BLGIeqmzF1biWUuo3v/PM9/kTgl7WqBcHS3fvHiNXS
+tYQrrX3WVYXzQNxrzffD8n5wYN8IcURhOZuYb0ypG3myd4qwxbD1vevoQLSuzLdIMdgg2xkY1FF
K2obDK+Uo4R2iq0ZzrS3oRkB6QR/C7lBBXlyzFH/b9XT1cz1jCuCESSsXO+LJgWXGpNAJaVkg5eF
iBu17pZQpgr5ZszvH6F5m++rKc7OCY5Jtuz10dO6jJXYA55nKzoRCGXFBiqbjVxogiz5nsp7dlvw
ZIpR7q6nFGV9Q7NHyZy6pqiTaku1adFAkt/KEMetNlP1e42Ve6hrSzqfwQ4G0JZ6+iL+prqpKngr
yCrBFG6JjuYN4KQ1EQCCqujh04yiWpxAnNX7QdxvsgOdO8puS3Ol+g74ESjjwDKNBp4l43nJNfk/
Q7PdzVDdEPyhKW44CJvvVSwQ57LQElPIszCR3IdK5uFjGLY/zhCtq3x/qr2SLCreVlX5knzcssfK
Po9FWOK6n6W4IauyLZsJyxb00kWylpN6CioaQCNg4nboNiv8hwGyajuI9Tn8ZGzwRHFnnwdYUcNt
HxcjXDwCtIwI0pY4NKKvFWlWIS+HZFh+kFukuKnldlQVtRYQgoXvUyELbO5DrD4Cz/SnmBD2N5fr
UuvCeuKFVtwX6K0O4YAyqP2XTDmvwl43mjRYHXlk68/oqrg/Z0o8tJ64iTpFbKUTTIA6c5Nj79Bz
lOrJnAwk6R6ZoZuSH1VcS0yFEHOcbTTWFkbBsOO05HkoqVjMStJX7tnk2oslAKnqwVW6YqS+cMhJ
VUt7XidUR9JypC3pne0nf+reWuH+jmVBPwwN0rrggRE08UHg46wGu64XsS3cP5Gdfn/ao0kHbya8
K3tMOv7yEKlnWohOQVgeet+zE9dYtLVNN3K2OhXUUSGezPjKSBDJgF8ynKPEaV2TNeZsJXfh++k5
HZXhX26YKyIleknWIaalovQuyVtJ1O8h+EajLZnQCAeZ9/VqQSGQtjEpUgGC6AnEQGEIr/lGQylW
VkBe39QrpRWl+XXp9vNIW54pX+ocjByRXYQJ+uVPJ4DDJ4lqkfBrZYpMG5WTZh0Jq2Q47ADRcsOq
/z7oda7YZZUHfa8mkf3qRJLmBjmUc6Wm2rnJWww7ghNR6uwIyfhf1Kapc+fBYDcom6bhtcjFoBnQ
n8BRANkRv2/JJYQK3Xb9gpgNB5Es8ttSHH5sl9Jw1+jxMCLwRfsS+0/pJ6IJQLbFtV7SSrOMb3np
Jo35nfiG4E/dtTiLhuiKh4ULDMl+h5JdiHwJfNwUUFRO2lLIuC2rgzB4mhSTuAm/FCL6xxjETo7Q
KiPYACGlPbVDk+sTOI0Vc5sF0U+fP4QeX7BJ9kMzG6QRA9tAuiMvcVH9vPPm+BVysnUwbWdCcusW
UBdMrwhY+zKxgSCJm0bzeEPJt2x3Ts4Myd7fnDW7Wy8/2g5SGzHGy5K7XuIv+f/CiSQXl1xzlBFd
vnjDB1+2OAs4IrLRmbSj+lE9U1nscSoJyB1Gockf3zwEhZ+LbsWjsHqPojh0eD69LK3IEMpCaUoD
emhN/KD090ebApCgFS//0m2odZw7/kd94heqqM1lq8wjwrqAvO/sj78BgCRJnnIBb+KbVQYb3tR8
c6jiCANew/iw4hnCrXdvcSZ5jRgv2yYlEyues3WJp5QEcg7+qHrlaLuE6UE9pX9S4cqi61ZQ1zNG
yIia1GjEV1qL9ZpUDgSArSGLjOeUZYpKUZSwahc+OXlqZdDri1Ik/no32Hh8TYYQ9rfIdMwzbdoM
TpqLpSPUb989+aDNgKzoG1fTKxLD31yYv4QBEhQmm6MAAUuVBmLsfV1BlQmP9cwFHtIKG/f4kqAK
R4bXqNXY0kBARvNIpA0SkIQKDwnC5MIG6ingAuU6AaIxqoaOwMcTGakrmHYbNGTGeWfeL9P7Nc4h
UODcqtbrIrd8aXiuSFqDJuTsi204aVpbG2DXkOlu43hWuXAYOJ4zxXR4ShLkt6O3fcsn/AfwQR1L
JiQY5oJusWmlSGtzXBBgiQdY5oeRfL0EZY+uKwyiRV7gMrlqolTrYvtypRpc85CzB6N5TBMe42WW
f2k4MSBKnr/CGmbRSluNQU3znM4ZpC4/+XqKvgeQZtLHj8EVDK4RyPBfmD7t2JbBUPK8l7KYmh8/
kmR8+NV+De5GdlUiX1H20Ire7ZCOG5mygxkoNPzbFT9SyQiOej4CZn4+D8Ubm0SDX3d2sAFjqN3d
QlfEB7nrTA/tb8Tih/q+fMNvJq8+fmK5txnURkZvo+nFDK1uzW/hhaeM4W69MR04Vq6V/9HjFwZy
aHqnQQjoWI9c1lA5OchgQ8Ww1dT+ddqSqnBCxYkXwdTStc3VUfAoK26bEmxDDffqcalgtm7wBesc
3FZJuG1baNIya4aOT7W7MyQhMEaXhT3ctX9PB3ZXfpRReRls8onlP70UxpYV5TNGU3tZnaMIesPY
H00QjT+xQ7VzxnnhK8EavFHs/aO8dD4N9eWM8+ueS+5Knt2Dk0QuXowGy7kPVVN6CAIkcUMGauz7
oYdPzCJrd9nyYG3LajnWl2es1LOey6IJhmPdcLLVcJywoSNLw5Ra3erAZxow7eoT0cjhrRFFNRYK
UgqWHqy86aeCmva/REEPNNr2X5wlA6hjpLJQkQ/bcqPwjcOPtB9Xow7fLkpRXHEvQjYr+4DEIcE8
Jg7jDlOwF4e+aqFVGBxcHffOMtBu8XlHBw75gfaM0NsmtywLIefbHbPKq+RtQVMxacuZODUOE81I
3jGAM5gyYwntNrfJ1P0tykoElpa50B0HWfb0h4IAHTnS8sKDUf47tTHAr6q6vJL0fsvpS7ExkMqx
AeldoO8GdokPa7Zfu2Brz32VrgEyLxZQDpizEV2EuawLN8uXvO0EXYyjlaf5NAwYXtAw3L1mx+JD
aZYC6RhTgDDYOHfvvNRyfU5Jr9v8ObRSlk/mmJw8E/uJ+N0bDz8udpxmfd5Q8MLYftU08LeW8k2C
tTyz+RB6pRYREXYjQzK7IShB8Y26XEltebeYMAu4+WvwoZ7SpYlXo3JLV4Ow7+ID1kDCRsWrkItB
Dmi6uAiYsCggvSLuefsivfLudB1fQPK+zruPvytt+U7q2pcsvKXazxwUKGNzseGRo7WxrxZiflQ7
utqwnjP5lcoRKKEnIOBwwflhBwYDsfSxg2Ivzj1evHKerT+dY5JW/b9rpepsZck9y8jysFwRU+wI
SVQP+emUYS29FmdeXgQa3atCKbwU4f2S6AbquqqxKWBylLbV/M6Cj9UwGUnM2+lY0A0QnQnE754v
ZSluKtw1bCGrsveO8VC9sv/XApVt5hfNOnWB4tQDkddZB6OrscgdV2fh2g1aeXfmKi4fT1emZOkg
q0rWn0dSu9mIO13sLrO8c8lu2vfEnziGbPzhj4WKcUpK2ViWOhZLlxUAwRgEeUunUswBvVW0h0DB
mqjg/W02waqeTeZ2LLO2fhA33AHwza6s+/HubEd9OBV0CMvubGxAwlQ00gboOQj2Acyg45C7STbJ
Ouin1vtW2DB4Br39w9qC6NqEHqSL7aGjmUO0V2zrP7G6qlPLIaOkrS9mJVLn7HBpvNu3gnWBPc2w
Fd4Ctx5Tg1k5D8wvlTH6Og5C60d5bmC2hyi3T8DjprUJeEOK9U+7Q15ckZoeoYIZwOMbaVvf90qJ
kMuH4yGMWcfWl+gHEA/7hT1T2JZNmtvDJ6K8Qkg0KkdNBkzqbBVnf5ajzPXWnkbTx1S6di+scwZc
UROnkgOHoNY0CUdTQLh5NesAXZV++HXQkngz6dKEdM/+6hc2972xzb9mOVi2XsCCQ+xkucUqK/bb
C8+Q80dm+hymXnzn7r+NVawhDYWRwO1H8lgSopatcOdiLn4pQ3kHouaE3SWBHYirj3Sw8sDHScMa
8lwvJOcSI6MHQ2+HUFCmiZc9qQVf3fz/3qTbsiNwZ5Dmh+hZTFA828Tr5OyTSI+IaMeV5zvLf5jH
VIg8Vu+lK1zwsf9fzQGGdXY5glJTFZ6nkA+/GS8PsBT8V0anrqtI1birCMH74b5zX54OBz4lXj4C
jCpxIPQMEcP3S5Yz5IoxNVjNEgaSoFA+5f/cMpE1Xcc+iwqMixzv4Vkx3sCsKRhHvBS6xdC7tknz
9c/WSnxZ4Dh7DGuHWOudAFeGUCsczLzyaR79pd2upA0rVqxP/8pbszBksS5yVADc1d4aoUSL8Kxd
hw90/ExHtQAIYgWxEKMVGB1KeFjkZzbCKI5V29IjQU04CDPEzuJWXGlEjzWLQiIbJNkRUrWmPJcq
Zk03ZF93cii5XAA/4Z2ZkOHua9FG7NtQfwDtnQLUf2gnyneGe6JEqkfBOkLZqzu5Y+roY4wNzGwO
/fH3M/P/06/GlfQY84LqKZsFh5R5SD6ZQLk+eHoi/bk4loHjDjN7KdTUkiZpV5PivCON34e9hq2i
hHcAfG0zVxR75WLWyFBF+aF4xtQhot6ANsHnBIrvxiB2DyQbW5Ti3ix18tDNjN08Qw2VChIk9Kid
ioLmWaNQQ2S79VaYbzdennrX1HLxNj7wK3b+cIVbGZ4Yfl0LF6+442fyJ6lwk5TMM3ljg+4B3wzq
y53e/dlZcfVd+d6NshtepuZF27oUHdBCcvCt/a4+jHdMcjj/CEGFnT2HJlFrCe7XDBwZ2zK+isbp
0L5g5c9W+P0QaZGQ9rsgiPJtTKaYOQJrWeEZAwaQDyPRe5IF41vyrxoK5cDqWEbxKoJBAp4hnDpN
eX2cwKw39yAqjhuFwYMX0BD57TktamERIaPvoQWp5qiKYcRtqBHPBugyt7wS6d9YHW0g/zUbWVWB
XXo9Mu0Zd5BcmAt2l6IUoNTHJfBrpYev2d4giv5VouoWNL+xsyqFaCR21EpBGbn/rZg6BkeJTgMK
73BAuIyIGOAF1Z3I4EryO3vh12gbMmySZUzmFWcZP5bFkIg8bNRhm8TVV4wSgjtvkY5foraEUCTM
SdfTLbN9aEVl5FerFvGG4agf677lbM35EAq/zVenAjM/nDA3/5yrkbH5k04rky1mY3VssSr075D8
eg8ECQ10dmtyORNHuM1z+0lPk/KaCp4R277cG+cOHtNgYLo0Jv21laV4J+rgzuilVRZ7CjyOLYYN
dJkEkGxrBiMCn2S6NKjqUeJWSQgpAIUe0+f2+qjvopyGLnIX4er+6ZLQisxfXAJR1svNTTtfVmbG
YYS8P4t/yX/RTFGbw85wQtxAZ2iQ7OHXRZ/fkvD6iBQCj+c3I3exn7uRd1FAK3EeiRzM9FGSSWoG
Lk6pS10lsg3y6gTNHTtPo+5SMNhYEkLLnjc7nVGEignRjI+EI36Yb63ga9qBzpfPGVDKxY2qFv/x
0yZLBs2/2HzIgAeOtthxmaRTNoYM3J/gmXMlgtYJFGCxnhcm0GIvY6vbiJ4F689EituYmqXj93iJ
JpykBJVEXDSUv45b6GSlcRty9D74wzABfTQcaVB/jZxZhKilUfdbX1hTGu0cpI9nCDr10jP9Rur2
nuRQ/OdyIRVecPiRSxIXakOKJh9CmWcRzU2UQO680LiVM3HWFfyq0ieyLIiWBdicRTSmEZ7ixzmu
MSMyldSunTEE8V/fqKwayUZY9V4Q0BUztheHM/Qseu/y8IId5x2e3R6f8TjoVd6yG8fpJ7l7gV6I
IREdBFonpFhzAzpD0rFb9Y7y16Ge5bePrWhDViAkAiteTeVUOMsAVWanH857YB7H2yAWAA6zKtIE
gia+kH4dZZ834LTFfiqRoXiX+rxZnv8QQqpqq3jdwF8F57LGOo5KPs1+yKNyPxgnyQ8grQZZgZtI
KQJatowfpHc24g1tF74w
`protect end_protected
