-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EIMcuPbWJG6b6g7vBHclMfZ+ddCvYzFfsYIcaQoPday5OXFDLOAwclCXL0z6JgANNKizj7mL0EMS
2bqt3JI5j+SKvMSQdmOSiE3Vz0fprGhqQ9Zr82XtrZa+oORtBvmpMUjD7FTF78cpgqFXOwfXKI3+
frwB85RlBWKVL8JDAUHbsZQCPR7SOhytFa8lSgpLZeGdMRZp99hawXDoguSbrYu/SCaKbLavCmvy
eClKa5FeysVnl0qQrxSBRpiQYgj7DjYEsFeiIH3Fb4E6ysoK3V8v0BRnupeslBCZ1HwnzHDhIv3f
Vtla39OkmDD0TbseyKIIDUDwnIFS0S85KELuHA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
sj19AJhY1rzbi6jAI9qL1U1Xw6usVx1puVmUy7Pzd3oGqIV2Q8fUcsrd8TewUav42fWkj52r/CUs
6SyX+B3cSmWz+ImJcUYlo0tuvr4T76UQjxw3FrlpdDIyLylRq9oVkZTKbRbWIl8ahi9KhlblAl+D
4UOBfbOpjOXoY8UTCYv3AWJEMt8HjoLoNMelM5WCEMihpQBAGyiSeJaWHFmJyXyBV17ABXOUqR+f
RUImJWQejVVeF/w20D5o8mOdNRakidrsAG7TVD9iOYhDOZk/64syo4vyElYHnC5JLYLTdmaREoDX
e3hhkc6gBWbipoONcEBGjYPT5JACEWCK/MxFkohqwUZ9ipeZ8/tXd9A1dUcwV+NtOTcCbuSt+o+s
i2UrFi1YUkJXRp7oeq+kt4yAUnOsNsnENunutHaqV1mszOZxGU8U54wQ914Uuya6vpZQzAx2aZu/
6P4FwqG7bc0eVSwgutkwkm9Xzmq/IAanYTpxKhlbUeN7AnjprH9/vnbfLeoY/tCxIYG5NmIa6xgR
jFoyFfIsxQR3D5uN9WO8ejCMLbMWh/LKpXTDNGPdLnoYvr/QfNP5klXhQB30jQp9k2aUtTEOnNJ4
14IKe9YilnbYYBtkWgRz347sW/Gbib3sm4fnPB5+BNNB9Y2AKGblfBqGbaViEwndzOEMSObWTBi3
6qmrGVUWN1kxlXpjd/Hnv9pj7NNkqDW2hKu6cz4D2v/bhmHnMVVZEO0UALZKuh/+p2BQCZy3YWQQ
6uTioIiL2mo3K9Z3fVPNZt9U6w6fyZPIbvbjq1mtzigSvmCkx73+k9NWBliZRsmMoCa5q1zXWXWV
86UL09RYcXbiCzVK0KUFlL9WuteNMsgm1Alc9p8fk5DAzcJRbRG6+PAKf6iiMSmvPyEjtiWPrg2e
XXfeWQZz8OxsMFwIVJr4Ke5+8ldmdZYAKlOH3wn0r9F9K6tWJ2B4edrvQkIWxxvpgH588DxlgNtf
BlgBZIIBLr+Bz++lkwuQEBzMJFBro1jYn+dz7GkeCGuvt19afZifYAb+UinubzAqbg1j9+dgFDKD
Pl6bnMHSqC1dc1nlPmBD0udrDNwCssFkMdytg8yyXbJb3zum3tIxuX0jQQGzJUjhLVSBSrvUYoQn
phGbvwVfvRRufDZdjREgLeE1WuU6PoprKgY0RFtcPcU4+Ir+1EEx5e3AQpqpNq7L71QiYyIybNYq
fM2EDkoD0tmuwcMWFpGuwf3Z3qseevgOj5Nn4MWhDQLxDVx1Y07W7YmZmCChX6PQXcNnluymu5I4
GC7wqyOmOejdM0NVkWLOMKZHIbiRk0lscrVZWC0LSPiFtQ44NmfrwzJXJOZ9jDHv7/cgI+gebARU
rNVCImEB6DPiBiTQNZCeEpZ44+Ke3hjJxvoXJsopBlGDdeHTKJvtNFF5/hbXjvpUNCvOuD1wOkS7
F/J07Ne/aPYc0S9SSfAl7J4vuPSOQCeI4bvja1MYSkofCyavHdpxJb/i+a5uyd73dr1JrVAGp3oN
kLgTCB+1d3S2RC3D65OPu6Pk+7HDTEC20LRw7acAkSDRhHiRH5UIVaHb9/QpHlMzorPY2Oxhokhm
BqKGg9MxTRrnmYi4PAri9LrPYsgzZspSkVWrtVzm5VKq/8TlXE6GluouFEAUZNlDJc8PkcmD7dw7
MiMB+W6UMlJzp1b7OKb0WHPM+VrQ9ME0LoirRAG5X5UETmfbndvG8Q/+HKBXS9iFiGTj5LCdxO9d
TG2yEGFW0cCvbqKqwtjdP48rMzbYkXaa7fDJzkKQJzZ24M5LsCz9EOBlLW9w6yrpLoDTHg/Mg/7r
0BGM+GvRg0mPua/CJ9ZbHBCoQCtfKIVTYmLyDSEzt7pVDdQ3QawMEYgg5jP8Q7LfQq+MOrjfXxjJ
SjWyQXWG6osjUggcEoWhOWugZwUkCWyLQ9PC60RngNWf4fx8Bs3jku2VoLmmYKYl8bNgS0wGAB4H
j0H1ILEXSstSgpbONSEwSglQ2cD4+/y09cVMSkCiDr3x1OwvbGf/6UFuzE6+SZF3sja0GQxqw7eU
vgFrpgtg/TlG2iLX0641mQ46T7NzO4sjhqAqhuUS+YDixRIhK942njDPz2Ox34y2GSMmnyWub6Tt
WGJGoZV9tElfWoU24yacAfgkKhfxPsQlppqEw7WOjtD+TMa4LCAqJU0bAo88+Kplq8T+j0yco0t5
iiNaiGh6UY+MLL1jHokZjUgb4P6Sot6JGsLQygSCqPwKb70GTJ4yTX4ffrS4NqxUS+2CrN/b1H+F
MSr8ZFBorI+Ayl6ch6Or7jXALlihKAAo90uYc1SvBH0aLovRJG3/X0QVAvbDzyw2oSnnKED7sGop
3WwgkP3EkNGekV5NLYIDB/DuXwV59lphrVucA1nKn9Qw1xYEMkKt1wcC79H6q8vwJ+2LMiH1P37P
aDk6f631SCpWtab/p3k7rY0jrAaFdLpWzTYUD0koUktp+witfPPd1soj/X2RBi8cK61Vkw9bEvSG
/AUXmQTUTKBmUPH5Dif/S2aXhTBvRdUn+cbZE7yMHRUen6B+Ocz3D1cLWPsTXjXWPJHQ9fprzi2s
qtD3aLX9T+X1RWfuXifEGAtC58T2gLoI8Ybayj15nJfbp2YbsCuE7epaY43e7TwErBOcnRiI7mZg
LgYnvtoC1dpaZtsG40afR4LGYGzwN1Y4mdlc1j3i2Yx1v6yv9jXX4iTAi9/nL0DhiYGY4wLJALpB
50glzzkN1CKBRprpBPga6Re8g6U5dt8c4HyROzZkEnDFPGEao9fwzZG4yi19dqRMyOA3kl85LzwV
Dk61rmopMIYBNDdHLNf5BeTvVl+GnvuW/gYeUD14OzOL7opO2EwOlaBVnHQ3n+0Pzp2yS0SuCP5h
82Bch35wTtec48kKWf+Lz7KcHrBGCYfhO2uObnwxKAxKJuvRNiTZJtJ70598DXMyAQrGedYXyNYe
JJY7v6Jueh3Csr6uoINlefsVTo5yBVs1fQaESHyOuTZq8yLniOhJSVCet9iSZf2U7TUl02O32IQ2
BPVYCQPg+3wdSU82Ejhn8/fAuLPsH08Cq6dfcWSrhUQqcPwJBzyKRgANiLusT733WAQze4SriOUM
Jdy/oLIvVFo44IqoQ2mbYLSe1UEgI16lkK0iEYB73tqUaKG6XJgTCAqvF0DVbCjROMxgdtAWcmXc
M6ZVPIV10YdtBGU+KCJF+jBOjJwyViFmswyCsNM/4N0Q0d+uUUDGcqFEsyvTT5fiqCsq7kPevDS1
fO1gJyVkhibysFzF/z089UclfD82ABo+QTzuM34mXUoi5/raA3U6vxDucLWkwjz62hmbYRIQ90SD
1ARqiFKhG6xMvBnmvuaU5SKEWBiy+6qoU+8Vs3ryUATBLchtUqkZ8OpkFu5B8iLFj023hOl2E7DB
L+hVtbc7lIwDoht6/6LyTQWbIOeK3ebHI6OPq/fPnfzb0Zp94a0RAA5bQja1OAsH5SMK6ftRLEJt
ez+2F0E0caEm5SqOG3R/k8D1uf3a81Ncs72UhZMJuilATWDNtDWp0qN09kaSbP3mvBf7llucp/fY
jwi1LQjkjTyw/LwYhGtLK9d1EOfSus2WOWlFfK+wKkvAkivghQoB1mPu58oZ/JSd4L05JR0Z2obE
dslznMZ6jbqa3SDU3+1eySnoUziUEY6Bth2TrgPd4iQINO/iojrcv58QrTn5bVtS+FD7cVdV76ZK
2WA51MGzKVrpndHNLXZ8GKU8i1CLpm3DIMWIVp3l5eH/3FXwcnX7o5Nw0EArgt6a0iGPWy9PimeV
f6dCladb1xuaewhFYwjBCnl/WhQMd5B+wR/fAm9MuEP+GP+l+yeVGJ2x/ifffzoaEYeBD7uR7kuq
QzDND8PVnmLoZ10jN6eHicUr9Q6yRGXCkdEf7mz3fYuACAPlW7wauuS6XwwWNp+/PDXBllg5rEIC
08WIu7VFy7Z5afaoVrV17Tw6fha542MJKKW6mlnbGEOPL6ahNvUERZc52/jrAHHuuUTdzTqLkyGV
lKJazr+kerzae9EhMdSECZh01uLGpqowB4ZuGK5GEtyh6M/1mBIR/oRuW4KCw3qR/hLLDonO47/K
Z3K18CTW20t/2M4eoh7MXKqDCWfnfZNyLZMPxl/x8x+elhl6Uf1a0X7Ay0NwdSd0hJ/9DasCSlUz
h4gq76XJnVpWJzUdqOcPjssrDrLZNhN/G9hfSgqra4baKRh0Rgpqo7MVrhIMEdEKTw0hNZUfD+Yi
UbhRKhdowIymcDZLlwYKFOn5zkVc9UfUPqAwU/0ok+btcUPKkbWtbJas/5qIOKM5m4Y1atzBS/2Q
36gbCNLIkuSFKZyiTmTQ5neOfmI3jO0GbbijI01rX3aZlhq4kWdD/Qjo0Lf+Gj/rXWlftj0T2YWn
PuZhRawfhidV/93d+GdbMfIbNmlszhCT8CFFcynvCF7rBzRmLzQXwC9dfwa2SjKuUGd0yN1dptN4
RD7a4j6rlkJ8B6snTk3vVUFl2vghxe90+g6+N1ENytXnu0t+wkTPJza0Pe1IV8CesiPRf0q7APvX
DOfITjNIus24UFKeSCGf+UdAjJ/XJpICSd8NqkcJExqVp8w3vN8RO5OeYvm4OhmNi1m/KqQyNWnp
k5nBcYtIpPlQYXYMpMX97n7Z/cUaMN/NI+DHBqumcuIWpW0XkJxZ0ge2KlFlZui066gl5tcyl0KJ
cUP57xun5xpzusmS7c2LgfqcBZCFDOTK47H17PUGY2lH77yAix/27/fAC7XOeK3WS5tBBeAefhod
CL9b2WUUGx0JbR8qYIdI0siWkNJFcUItXLInzQKCJts1lkqFhM1dqaIxIRz8yg/+Cn0oVhwWCQ9G
U2NJ0hcx7AtcG11ctaCSYxbH5CNI5gZjVddK1nHelhwPv83xN9CXk2TjsojQYjG9vZH5LIolQwab
l1vMD484/YvAXd34d8FrR6/Bgugw6NcxERkeql+qKO4bB2mfk87SgRGYTECkyU0QjS+KcuJHjslO
VcEbEkALc9JHMqrRteD/xrBLPkMvt9eMfY053dLKUSU410qu7x+i0Owm+WAlOfhwM/yqGAH4Ee/W
xtHFmUtZwARJF3CRNKqPOS11/qk05jT84AV4Zhxo49hseznMHycXeQ4URgTc4fZ5aqQaT6/F/sam
a9iBSV9eWGx5kPL6iP4Lgvuqy9cCDPI8QkL5N+ReOQ+Veg3/bImGAk8dutdf3WWDZiIoGv/MVEyI
pablXr08zeVXn90Ed414YR5nHu5GwjbKh+MDL/KOS2tVIMx8F6sb2jxcLT6R1n7HxgIdwTbztGZ3
zfc5xR4RGzdmWa+0ehw5lxHLRmkh8u+OLGEWfTWTiJDoTdmumInQPPskRXSP+U6uF+s9H7aVxWsi
Pa2VYNo8Urk5QZEUiNdmsjFkwUtdthuN/Sc4rhjXu8p52yl9Ha0lcGPzRluVJcH3i3wJO/8U4Huu
zLIW2vtP9jUrdXluo2coMoEgo7MofI4DrDsWKqxkpKX6UwqrJ7d/E/tZCuemRFW8HLP07SPvT8yf
U46uS7TaRxjXasO2j8Rxl6zHajbguKinv0kC/17jEpr6Byds6HisnrxVQgrAKIj2nNKhz9M0i/Wn
QC+JcWbE6nxYrKfETH8FiT6oJ71WJtEYAuayVW414iX1ho4ZvFFxmk5wRNoylROraU3Bcx2UwV1o
G2bPN3SQI9NiGYgGN6/rzBZILfeWoiO5FY0ENKLnmL2X8brUNqCyjW22Wg9uk0Qf8x7SYiCbFwhk
FOcoJRqVYe0Ctw1uiHlo7Fy4ezlyRnpkeVkaU1R4sC+rU6GJxoEFzfxGH48t7gY8c58gKlmgmoT/
a/NucTZWWNN/O5OgoIAjNCnt3TzIUp8zbkgY5nTUHvkx4C00yW4QZBlDPT6GjVAqF73w2PypRlsE
vpeUF0EkTapJmRZohAwovWzjk5rOVvD52BqZcZB3FJVWwk+jTbZlhvxe/BdzhqWoYz+eXPJlRfLM
Yz2k6XKXW4FAj+/8nTfUGSp/ufYjB7B6NbySi5NYBEtz08864S034oSUJmX/kqpdw0/L+UiHIc0y
0rBlNPJoWsB9A6jaQ1iBP2uKhEld1SWHex38QkG5x3nfFk1UkMRR3jcDHSAQIib3nVkM9ukB3VWa
bezwmiyPde3VZjP71E3R1uKqiXpu8mOepW7LPWD7Hf7cK/88+nO4eX9A0m6LFejEgm9dNgaUAYtR
bgRipWuEQ9k/Sv6YZKp6qB9oQmh4Oy4VIVUTO8EUn4sYZw3w8xhnCFdbKokDLMSTM1bvZvIbN791
BxOzev0cPIoVrCV7hG3mU0LehJHbvwXlujEIinzfoO3Ee3bW5qAsSz+o80/v1D1wyd3e0TDYKDGG
3zWWN3Bh3dbKdh0HWOfPOT3g4An+ViweOvIbpmmMBQw+6TUl+T4SvXp3TmPd00KvdjIBfz1cJ8u4
VS6oqZnTE/zILJHWaUnnPeG0pdORBGYtDuF8d2QF7oQX7lAByefQmVJdoIyGlkcec6NDRN3NCFpE
CLlYZWk8O4rl+tUgBdvzoOoOzvOMYhyFeEBBsMaO1R7dYHFRG85knmyiPMPcHx+FIvBTqjaExiNk
GAvAABtt8PiLJmVupMwqIQVT/vN47K1rM9dsd3mw5PVq6aykxmNCate2c2zaZbyaKIfV8JQzx8Vs
fMiG6ycQtsWTjrzEwhio6xWZODvfqAzeeco11CIliGr6g1x2zMwSvPRZtZvyDaKAwq7lTbyL7Aey
MBDNI6gBIiZqiv7BNm8srZFYwlk91MXJuvJWEDF3qMJ8TIYhulScA577ewoYW+UBNLZJmmBoyblE
Lw6+s5+HcVbfDKmAe/fsrVs9yLq/XCRP9fQ6ow/CH+MVCUoqsPKl7qhop6pTO8yHF8/H+ipyTOuG
kDLGKfpMJpheFO++1ZHFmguEZ/mtoamUiLwiOkm3UQ3WiLQPtZmSS1vplWY+nuVDoPdLllYOf99c
udRwpzfZejIqPz2dWpb4wVvg+k9L+wfWD2rk6MdFHVV1tzpuogv3QeA077yMbs6zSaqJ/wDyL3Rk
jhlzeoeh5iQpkhrjdZGMfoi2GgFJ/0hiff09AZ6bivVuRQld3ALNOYyKLIQWvdIFiXK+/b4S3jVF
wzHQBZzePuT489a33gCZINjCDgH+OOIHHMspbPPu5F0XKH6kyWui4sGW5szX4jDzmIotVRcx7O66
/qzfdylsJR83P5UU5Y5ZCcKd34Y1Yaw3vUBGoy5brr6y1dMfYMQf6y1+cr7hlProJXYECH1kpVaM
JhRXjsYVGrBGwIzF1GEyuEga0aqvc66ED5bbC9MGOhp1IFjRDWyutC2y9UbDzbO/J721jZ1Hh3d9
YsNqfI8CpT6HxkqpAA6BUC3X/q/W47NW6adcyvHpRLjRPdSuTD6SL6OUToGxgm5Gdftgk9+5riw4
fSIHjx/wgL6D/CNoZ+XTpQzQMmQF6Quw/Ei/FXO8iEibpSHtwjKg8G6NTgwl/yQd4TLSc6Colj/5
gv1DFHdubUtnmqB5ohngC/WEvP+vvn14MVg4mtsCSUXZ+hUm4DEayK7nXcQ/cGKrsBmfeY2EIQtd
acQFjYc6TiX2+Up253Alz73Y45VKtJzzqi9bRiWVMjX+tAnSWnK8v7r1RZ0aIoHaxaaordwKvakE
IcjRyj2FjbJZi3iFCdAyHXvDhddOASZN/jeiSGl5DcCsFpSQfptTrWrVm6dEDejQiJ1UYrpDcCLh
lhK35MXEWXY1IQM2abx6eXkZTrGtGo9u0NfmW4Ze631WcBP0rUGH1uWXxnEh7biq7HLjYZehbnah
o1jfmKkN9Su2kNcYDbsw3abwAGmAaTRxKvVMPTpdRqXpR//FRrJM86qlEeCi3JZK74WuHMaBsBzc
t1DaTdjeKo08zmjvRaPEWw171Ce7WJf5uPQnGAblrAiSN6HgZ5WzfEhrHPwxLtHiU1WmDU8ivKuX
d2fo/k9BO3HeHwELKs0gtJ++51oJ2x932+5vyQjyJ9RM10Y67zRcYaim81THqMprxKXPDPZp1E47
Ie4vxAxurF79tcmVqH+4aYmopBZPnZmG/UtBTXKAFBanLoCMMX/bz6QwbQUWZG0koQpOOAhi5DJz
ehxG6QZ7njyRXui2+BhpwMOSaJ7FSM/i/prSKF+gwPON+EO+h1KbyONshCx6iY9GRj4q+Fb8+Hoi
GWNdoCa0bA05l3T/BzS6kan+iXVjZhDP/GEGNX4eh7kOpaXfsIjGShNfjBtMGt81HmSb7yZiPfXp
WkhbO2xuw4D3ZR13vV9eSWrHwi6axCKpyxE0N3cP+4hFyEJNTbILFgsMCnd9Pb5trI6ffMDKJHXT
0DPvpFrnovV1WAM60/s14wVIYIFkkUIvIkymZl0ih0gJh8wqQb+p/9RTm/waNMUD+rpipIL9jVga
drzeWBbVH4OJdWVdTfFdJtGKQzsyDSiZFBZY7X8HSaPGlxFjLH+UmfKvTWENHwYw4SJCs1f8l/rn
/DcB75dlDVzY5efD/vqrHd8NNpV/R0cJy8JbWjfH0/6sEvmIzfAxhGoLGwO2TVp6JaXqfwXFIoBx
simeflY2xS9uwB/W969orKF06dSyEdvvMfcekhnKVVGGxWn+s35eHusnzOj7yuR0g38hxrAhmXfb
rV+a6tHRHHaOkkdRKmCA1ZB/UaA1g2mykpjMSl+mW1Btv2bu+QZYDd1C3GjR8EuPnBUjHndo1ukm
8yt/3o6cjLywgocTFBt2iYTUS9wAo/5TQWeuQaRL1Rsjt1Ee+LYdy2kXxLCo5kdCSEDK7lGiTeCS
1O9A72+1oOp3BlqrXEfb+buiyhRR7k0OKBzsop5IiwhIxJEutMHPOS76KLq4sT1mSgOvTPvih4qF
1jIezLckNIpEeeOULYRLiy39QozoxrvkM32VyiNfBKi5zI6IUK5sT8SW4RF8iuPrSOl62c4lGDQ6
43imX9UMnX796as7vn9xSHS+0dNpqO7umA6y6fHVP6A6r0SPjys0feoajC1Dp50na8QQsmCQb7xh
5ploiCwQny2AU91oup/H/59W0t6gCB6gwtlRGUQGg/U1IJO6YJYFCvrpmHZk2xj4sVvkystCPnOo
JKaXtJ8i8QtakuS7sCc0iG6JnAXjhBqKXwUwq0rH2hnbqthsoPRr84jX1j8in3s7Dyoop6EFPUFB
TxQcIivYYzDlg/H+VlXNhtF3RzKDkC2ok+hIgjOzAc52uyMxESleV0KRZcSB9Pj8yKA2XGcGuVxD
P6yNg7eKdd8u6WMlXmXk2FnAxccj69MAwtGPYvCSUaDiwb/XpNamdTnJutT5+GNSNKjl8outfw4r
sX0Em0kjSyF4vW2ibbS2MExPXqs27WmrNgXLOGCxDzEO0mIvXQa9eYv6LEG4lJsmUETlEHy9TMD5
dOtgrb6tLpqBXNfjlAZNVX7OycWpf0v9emshN1yWD2UmJMBFrlS2StCqZLI2U3Kohoxkt25mYBgW
xLIW+WHVkRZmfcP98GmTZkBFaD8kesqgvKqYcYq8WyQX3NMVco07NJTV/ym5G+WjtuvMXSvBasOG
Fit+lIeDUIwTXKVkGFLVhGgjcM6MHzVtbJnFAVyYda01oFznNhRBFDnXNyXW5wfz6xZnDhjvN+AT
mJsehFDZQDjBurEAh+63YzNQUz4O379M9SNbzOMQ9Sfy0p+v76HEB32lUbTOMejbtgX+ombdSPrj
08UCgnr0dZMIgAWHc1U7n0c7IH5cU3x9AKTSKd8bUJxdfvyeQejMGLWwPs9Wx73RZgEYkJrG/L9N
GnBRqwgc5gFGI4L88OFgC1g9DUhrVaaMB2xaRd/EcvAKyYVJnaDjqRvbH8bNvA/TO/+7qyXCKulH
i4Kn0/L+aJ2cKxOlMiScNSlpxdKerpQD+Mn3p0uLCmasKiBhhwaVPcQXUX/nANly+3XvyCFCNo8B
eXsdzvcZASV1ty3p8a3AQy9ZWyM6CHNhF4/j3NbbI7g6VJQ0Rh0Gtw2xHbTN7+BKLf+Bs2xGpCqi
k1OV6ATmR1PupMeaqtyDmA+YWQoVygpzWVHxe9Gnqh9NOOtDxOy6oL/2PNkki2bLCWNXLjuTdpQx
12UmOONLcE7sp7AC6fo3yiUuJDvL8HnnhKOngJExlHwAC3CKRF8QzqLWd/KHyt9hzb/TWOE2kJjo
64f9PE8xccZilEfgt85MxqDulO/b4XbI43/NE2TULUUtAQUpzw2Puzc41qj9Ipvr6FWM8lQ4pHQY
8r6+ntMo43bRjqV8itCxWqrbPMf9NKBSmUy4YmpBFjQInvmhFRO2y5s9Khw47CyZeIezWIOXa12e
ge6GbKiNwP+Ld7U0lZ8xsbSG97vYhzzdYsqIczNmkLytwFtc9lOmscCMf5Dz1azqFWk/LBui3Jet
CRji/7a7OtB3GTvXWX6yQJFFC+aiNaY1wMGnPj7r0yndmlMZbfKrQSrPxB5VK7T1XgtVxn3vYi/2
rEno4tOKEP7n5zNCyiGsZ9/xt5Vpnzlgfmph0naD/HMONfShECcCFSuTY6ZiUOOD2BShG3HhFgkJ
96WMXK76pFsLxkW5gtvIRCp45WJ7fMe633cBx2Hisr4hAiRF0lkIT9Tqytq/fCd8UH6b6NoHASD+
Baa5C27tdxRneNIv9pC0hEqdo4IfwneCXTinr8fpKZQuYbVnnYeKwQUkUAwDU/GmWoQGY1bh8q2+
xCyATb9UeggVT6D4RO3CiY67yukfi1Cmwgk2E/Kt0j21rBIOK4DbFf1Hd2+rJDLEAVb3H94dHEbx
dFnwWUjCHwkMf2tfCMbaebV58bEEoC6XKVmNBWeq+R3zuGs0v4LJwXioOdoxhnqL9lU6fZzYVEgp
uPKuT6fixUOB57+49UAsO2fnFrS3sHQHUDQgncheJ+H26QKEgaLCSEm5Irsx25Rfh9bYY3sXpcoL
+LW4wWQZs+fxb2EIky5NJ8e0oLNP95ZJ4B87hcLlp5S+itdWxkQCMoK9gznxizgYkPE6Bg2hOHIY
z5WfTCIFoB6gytm9nV8P3WvW27u9s6UtewsGxKeMwhnasbud5TEO2CJn6LKAItqB8fs74cBd7xwQ
FvNlKUCl9RdNp5iCCcfSiSBhaKFurX3ZYOKhtqtjEzOBE0PRIFkh3poU9SnTpkgF+wIgfjcXHBhH
+pARW11FWL1QnqNTw9IzlwTnsRQRLpQOHLq5RUlc4sRpToQbXS9dZNrRpSryzcC3VB2u9fh2aoYX
2tL9s3s/suhoslgIrvG4v7pLEeyYYm93LMMpy4gWeD26X8IFtZOjRhOqOjVuO8y6UQpWzo00hhd0
Aity2eDIb+V/nYa83CKoQDYXLfLGGwUtxsV4VInBo/fNFHaV4rpxPrhas0gAthHnXOJ6c4X8Kb5c
FVyCYp8ozBf7VkNuZFdpIKwzpwUERquoqTn4BcFqQnHyNkyJTTTfnfL6CyqDzCXEtLzLR7xgEjO/
1803YIawxacNmv/lNFwjxxLZAcLA0gTz19h73LpkOrL4kcI2ZhT5HSGgaRW5sLXsvH5sNqhPYUKz
dtAjTAulfaxiJc87hVqc2CCkX+LZlcVxSJZoxr6ywuT13x/qEHjwRUd6gUkS+KHTazYekHYagUzG
VHXYAXpVjJY+URRaNAsyARWkDfW2yxTBZ1A5zNBAP6HyEtyRzjchsbCVNar34DYvn8JKQjzsmYzS
yo1AKqjb83eJZ9RMDahj23uo+ooXYtwsHHQfiOERMTCK4/rzaTOW9l2E3vFY6Qw+cO2zbF59t8I8
zJeMkf7FG0thm+K3s07B4a3QjGwmdb+mkew5jwQGL6Oi8rjhgc+OLy5FezaT1G3oZkP5tFFttuKR
3Qk9H3SWhEd/1opm0TbCD6rX1zJGp4CZL8dt1mlcfBKsR2qy7mOqWr3mvAuTAZlDCfSl7zxgL5Nz
Ep8ag1KNluwaZFm/psCAOkYFRLd/TE5+ur2G5Hy8HDYFPsKx2fortKm/uQ6qFNdlfYAePqKP3FFQ
Jfm0N8MW2ja0AEKYu+KCOGKGJ4VFbPMu4CAlE414+t2ACu/KRLV3oQvNCcXrNH26NsUSxucLVEjE
UzBMO3jdYgBlWpx/hJ3sS7IoTxTI8S1F6BYk3NXIUR9r4rmSdoyRRGlZ/EBnkeiuNbzS7AHESEGd
QL0C49z7swS1HFkYzBnzcXS8N7T8vSroElyAmROaNyyX0loqpM2DFXGhMOFXYmSwOjYGguD/7pte
8fkCqEO8OLANJWZADgFZpUicbMEQDBnIJlrAeS5JmPGOGvK7tQto0APPSZLRsX7ycJt1gALRUAhc
qe1wqPkh7ffUiGE0wZeH6acEmZVi08K8R67uA6UZ933DLLo4TVxhZ7H7h/asDs1DeIwARIU7ykV8
ZyOE9z7NVnJuhqU4dFYOee6MybyRStW0IZrWfKB/ZAselKbzWX7nX8jw7cI1o/tBNTzBh1rFDU4P
UqUTDhJ4Ap5sAsLWGx5aOtJdP4wU0R4GEH9pgahSlfBoSsM9a78u3FVufpTAINtmm/2DP+9KLBz8
FoU6mMatzBKLf+Rv23ORRowX98CnRQY9Msduje/GiUx5p0CWxwvfOs73fTfqggAZt6zCiMZinurk
1TLDHtOkt66zZ4cmCxfXQ81WE11QSi2JZh4leodv65hmK/7gntV5BG7tGHGBb+xDZ+egi0db7D/S
r+ZtNUmcfMHCa5kawWl+NrI4Wpe1v9UMef4uIcNpL0XfhBJChhrcH8Mh7Z2L/Urw+q/ROxsBdG8M
G0xWWBPNpD+uBPRRdDpGyWG4z7PD4ghWviNKsm+duerMY1J7zwtYPpQDwXulLuOs7zECT5hy8xLM
0EdEaN+To1EjAHN/mQUQPyVxakVzrhG5sWpolAkuyPIYiwaOdDJr4pqycKBhy3xerzpSOwd4w+RI
iN+ORf4o4AEDFUR8FbCfda3Q/XerI7uCxgS1fr4VHM9lM86H3QWsvQ4xWFDJF65hRuD/hFUM4mwp
9Zu3cse8cJF+McUh67UosiiMQFnSuyrmAAYphoJD6QBnjiRpR+tNZjskq/BVCMBQ4UqvOv1e1eCm
1diVVFaeAhgIzLNycUIEtHMIG2uR4AplHQ6g6uQmPVG4+t6By9jyq6yG0D8cpdWQbCVPVQsNuCPT
lUs//Wlutt26bnzZsWp1n2R2IvCA8xT1xKetkd40o9LTG/4z7/o33BeR8p92a0GKgDBzh8ZfEo3Q
GB7yKpUDlA040M3xON7nvHNlpeY0W1B3XTIEo2XPi0j+fqPk1F+5V+BqqaO2l1/sI4HVvVPWeFWH
/uyMx4h2xVaLC3u8nWhAaXhjncJyIddurHmHf2fVFOaKVQUtejmOduB/4V/L62n+Wpxtt/8amaQA
1zskVvanh3fK3hdAgY2RYktbTJ/O43LDfVQT19CkfAwnh12pUReiyxPC7yNdWhljnHxfL0H7XVPW
lyXuGBWiAsVTcnbGNpeIDnchL5M6BnREEaUKHbRM0n+5HeEwbDLVy0ksmuRz5AxhFET5CLGLDWZH
jp7cIoxPoKq6KZQlxEbCw/JLNNsNCZmPrbsghombJlmH7RE7bwo+DLthtd5cjFx3HZiwE5sVw87w
7kZNLPL5B5iKxv9E8TLeaV1/7dXk9WqetwLpuqvm34nG1kkZ0eYP+GHSxEhi8jW7jqhxpFrA7hev
xrEu8RkB90YM1Rli8gD/2AgDWGWSVJrstGRX17j3mu6QvKM7o+m1Z5CChzzlLPm+a0J5+uK9zq2u
k66xC34HO3ClVP7WSPGpuI72ceKS9wDhpKnZoXbc/wgO94tHecMGAXk2KXKNxywv+wimm3lSgz4M
U9w6vVgruiKdEDmL6resdBLvkInI6ftGPM6KWihKsjtjgH3r38KEivx+DIWmvxBRcEeLwKGn1dRM
n5BK1w7ogozI9EjyDNxAEnF25qMGYrjEX3nrPyTcAAulShKeLyrKJpPUias4TqoSO3jDHHzbMVFx
e7QDPNF7zcTwHbJN5FzYgolbgcLBHN+dea5Uv1Ww18U9YYe8odKLrlrqa7w5meWY+oWkrcdxX6KP
WT09bhHdsJTBp16AxZ6DshW6eiWNmigCXY4BLhYJoehyT8ISfLrcMVQZjPwWrZ3z0oFQWh5ryJFC
6ru0Yak3iRy2GPBXURsNZHNO0bvPWsXdrFcCdKxMaqPF6CQjSyU5UFnrwfjh8dY9A4CjjKUHOu3A
tEmTeb19xA9a3jHw1UDdpy+UVBkC8Ki5NTPeeG5LxLrJHv2TgsLdJdCswLsLs3rNjJbQgB4wNjKK
JBAZu8sJzxmpHyK80Ql/plPqz06qXvJqjTi+ZVGE7HGicHUNhjFXuZQ8wppnSlt5cc7FqeLiU4ed
IlfFuetSHR199vSPLBX6oyYkIheJZ9Xi7kGsneR5HwnUBZBZHx5/N2A//oycXTKDMthhM+PldO1D
lbsnRw1l3k6Imr67aGfDdoHG9VPGgYnUGXdkPMHV/YwN9VKn40H6G4c3fCfCJBG4vaCnE3dH1Baz
b6/r7h9cAqdpZzWWoobw7pnq1rDrwiVbduaIgcuRXsPiaxIrwDv/zubdMM776iU926CxHVnQz5j+
xZgKtKp7fTpZIQRK0BLdVY9ZBiJ8wma5broPeSzakMhYsOwqSz8xApsSNixmxCxTSI0MdTWQ+81z
SqjXmudagckUVRf6WQUoVAc6/0v/b+03Eh28ClM97CPbn3ttDwa7hsc7b6QnFqPuEjkDncs4sCt+
29Yo9w/c1XNv1CCypiciJ28q8x2LcBJ5cHAtAekPMaAXDL2Pnd9KjshH7WImxHeiakFjZdZX7vBb
lTIouvTVoj7zcRlVgqqf0+zk4KWt788FbWNFlHFzHazoSQhDXMESoFGduLp8NxyVtCTg68ks72Mg
u3Zzx6TdJo2QbF+jNch6IUtVHtUHiZS5RND/lUykOuOfEpr9RDijQ09fHn35YDTljVGGOEYU+bwU
ZkFu64aqKIut/wfRD7VMSsUEEZGPdzh5sgO5Pb89KcjFcu9n8/TtMKiaKQnj8je5fhPuETpsoEb0
1qAPKxavRKiLEpVV7NidD0eMvVM9M/87K0G/yl/ydeSaYhm5GB4wpMGrEaTSdDOSXcZpYsdX57bP
FxYAl5lNqS5MlSF/tb/aR2tSY45jszSDdZiYkbWsuZ/iAJmkiAC6xPj/Z+Nskr6T3wnoFB8Vmcb4
HzPas0+71CIT+JwrVMaUuehaDxyI84TsP7g4V/M8S0FViupJ+C6gHcTa0J999utn7POY89kebIcV
C9YOht1soplSagfTF/Gos7BSGx0FDLiPXMM1KkzqipqV48pVxBMsxnFW989ukjsuLjLAynscw3zT
XC/j5LFBwVY+vVouFRLRWnyKFzqWoSynrzAgyK3/UzACYtG/w8DflzvM22H/1X/6piRv9Q2Kyjzr
BgZsd78JZfuOvKlTpPkS9bZel8k9gG2RpGuBQgrfTWUtmR6jFuEvFhGJ6Cjtj+Wtb45qLOABxusA
iaoJXpU9LUkr49bK9LnaE25hwbm9XCIpHmF45R7GRhU/NFM+0NIomjy4ZVWUQrrdHu/LZdKqLNFI
zzxjGtsQjHQ2+H91P6zut2UpcVsauWtMpZKgmkjjzNfnpVB25VTTf3N3I9DYBngXTcgmJ46dJQBC
3IVR6oxzEh0om6PKlmMdRg7fDTW2mYs13HLnyAup3NVwc3kmaRaZeYy4QeCdBAEgJlePJC/e7lqW
WDabpNkI78eBWkrmDh9kL3+raxN20CYI9Aoor5q+LSZ237UbmhdbFZb7UX2jyNsls/I5Ihzj+bVA
yIlAnkD9QHfp7zIGlPZnBOcWYHORleSYKlG2/RHo96akgsWnZYRhf+p/uEqHNAG2Gv/WH0Hz27C9
qquZrkFkPGA2/n/Ds2MHiTMrKBDEU57uzSxvjf9trExa7QyPKhSYq89KjAq39QWh7ZiH8zdbrg+K
RM7rT4KEx8Nh2Jw/mr0WgeD7hjgZtAR3BOZW0Ar5AlS2aZHWozX1ZEUpkJ7PuBVVrdOex0BYhQ62
njO6+EkOHp87HE43VM5cvEDGcNSmsYUc+W8wi9PhZahbyA8douuVfpyHamubQgwNT7DVp8tKBm13
UJOmz2qL/DgeFe+LkcMElcCa/JsclNShPjimTgWcPIU9gTnciA5MfLjpx17eouowZ/1+7Yd3of/I
NBtanOv5kUefHulrR5pr7a5G7CL1nMFULnEh7p27kCJDpblxz3X3CajDB+w/36cg8aN8D8dMFjTS
07uFgpZEYdTomEzOZGZj0tyaiTAr7He/IU4FVHx5LQpXwSrejnmsPKveR84NBn76Q6+fs1pM4YGw
Ge/sXUsJRi77CqebAqqoS4gz0I91te/PejOoIOd4vwAfiz8nmfBsXtAwBigUAVN6fd7b34j5+L9y
voSmjuouy1dhqJ+6gHFNNz9skXNGOu3Pc1olnMYl3gxsQk80istfhvk8cKdXPuv4DBPYZeN91LCI
GbiUR13yVv72VM5rEOir0gjsMhdpgLbyNIECGO6uIP0oC0gzdSqjLCfaBDbo9IreaP64oIgWfIA1
UYWHLKCqpNxd6mwDXYe0vP2hbKISmY1EDzgDY6eyMjpxgRdP7Op+VYM8WzBYE0HLguA5/zF8x9yz
xMYnjw/5Wlxcp7+C+eKI7ENlD7XJo0zuYQtfz0SnZapvomyYp0JI8X7prj5J47KOy6YCe6MG2r12
CTy+ABbqq+UhNokUBjG0k+B5db3/slhm0FUb07XgA9An8KlXE5s+L+dVp2y//2blaz9RP2bnN4Cx
keTFomyChOTGYEp2UHW4zcI+7XFYOw4Hn+UEZnpx3lsLSwY/2AZGbWN0VWAccRqt6CdKp8D6zaTn
5ZFoR+GdzU258ceVXjgmel7MLZpMkrNAjyDdntyL/EEIS8zhx9De6LPbWLdsoI/Np/CTilihlRCs
ycgT7FNCIVUt6Dghgo92DDrLW6BTtjUcecbrFdELxxMeU/7CQdUQKloqsGKZHWzfWA/n43V8eNoJ
1BQcIUBpTW4XnJ1aj30hgbROVo+8TPlDYq7ZCfWwSbNWfF5xw1WPFDlh1uS4Ckwb5MCB8iaU4euw
/TyPM/XK4DRwSOFRh6bLhPzOdaSTUVUdPMkg5swoRlg8S79UyP6e/TPirJulNcIrjiwsDd0Glg5q
usqCikANUL6HME6rZMcSBX0REtZKjZ6juBlZMqifS2qZvv4C9JOSk/xbRch6JfGYfdZq5fc7TT0d
03O8kXUQQ5Xe9tKCBpK8QXXOuX5H
`protect end_protected
