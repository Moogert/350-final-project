-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oDidLDgvMelDl4zTMxg6VXh7mhCMpG/CPrTZONNBvzaR4dhGZORNYx84gtEoUUOwVztqHaYHe3nv
FnCPUlsTN8DzljyPc7VFw/yvIiJz/EGfWNU+TG6I1xp7+oqinC+6batOFPfL1R9KUJFR8+e2lAMS
gL76XakBQDVbfbz/sQquRLL29Y/KlDfhlKuyppeFAuBXnugHwVthlXwQM5ONdSdkhzwxXgqF1EWL
Ff6VTgqhudfUMyzWVDWWtefyCmQaCVZGYWOfUashMsEeXOE4M8hiGzAm+0picAUGLnmodEhhWhex
uQcs2i4EESxqcItPYkp2W7m8Vp1hnYLjmoKBIQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
JN/rz0xsTaLEyZp+p5bz3T9PSctmkSTSI0TmPtbpifT+9m0tUmbsEqzG/F+3JdberOwK++3hDYLq
U7XfiMWLgARtIxHXyGWEhoQsxt0hL2TiQ6txi5v2v96WUig94xKUMRGQ/+fXQ7ssepE7YiH+qm+3
dBTCDimHImEgzFC5u6jFXnUdUzJZH4tBGP+BTbaLZOj1nyeSwlC0Q1Wm6JNw9DXmU499LhDIPTRN
xIW4Spm/3quz7Y1/C1leaMCXX3u/mD8zw+0szcWcwUwWcg8EMsNANQXaoLsNKR416N3k5t8eQH2X
yVfDoWxrSY4bDuSJNvvGr1/MyBcde+Bc/V92JXIqnh+RR1dCx280R9cHAvkTKItjo/n2VH7LN36g
MAd9srBvyGtbcc1A0qDeqYMcceblBcNvBvUssUGtg4hbqoa6CoDYSTcuocLO8CMcwy7haCafKt+i
bLY0vTHgaQiiJW/HcIW3ZvFuDptWlOwDLaKUc3S0/WCalKAJFrTqiiO9whhHerU5XGQAsKt0FdVJ
cj9csXJgzTZMEhEGVNJROo4tb0ZEsSraoW7EaB3SsntrSPnk0MLJnJQbBllJcwDxiewwQQZ9wSY2
5AK+DnWA83MDTWndSu3FiRyGKuTmZCv76tibSNA3OCRIlgA5i7n0EK+PQBKlBRokekT8nFsRN/Pb
ddV+1VrZF3m0GHbxap19c6cTgJoPhZC2EqABWB5mDNs02vy3fpA4cb0u9CQUCyhA+70c5T+gmEHY
gLr65nbHMjpVbMQvScePha/2Ds562qT79PiszjOu4vHwirXfv8a7fCak3gkmcaJ+qdNhNl08V5UD
ccye9+cUf4XWYRo8UgydHNv58pUDnVHksi7qbYwOC/B8sZudMBn648bFsVhQBcRDTqjb87WCM6SN
9e+qOoENDQlGKzcQubv6t1NU8DwR8vVmYPZVadnS/Dfx9hNEEzGyjRgb7O56fkQdsDawyo32oNsf
ez1dQ/BqTlCICNBHYvvTczgoTmF9kY3tcCFicr0q/G+WOfLQejJ+wKylgAPFICC5XmCOyRT5AaJl
loE11jsxj7PjjYHpC3fWRt+WF9kN3BGTBsCvNZWflyc3aIds0+r4H+ariyXKeHl/2q1rJyLCKt8v
XwRHSXXGH3K/2UnGL8WDlf+IE6Tge5ZW7UCH4g71XN2ue4sFm2dmOkLuOtCNee/p6kl6/rY+syET
jVnXUjmGB6w9CdYDIbHvJazBM6wsT/XeLIRMzB0z3T/SBd/DevXE/+ZMDc/mgYYgOmG2E4fo75PK
QkT9tVZjNaF0zWUSFsMXnKD2zEmpQ2pMjjS5Zjigz+beVD2W8zV2s2zVH7T1oBtFx2MdXAD+39S8
S/qecGmVpmfu8CrJh4zKsn66Uvqsnj+GSdcRdsSQCW1j3w9gCm0o22gQdHfVzgambpUaL/QvU9fr
jirGPrPz8ENKaA0Fj5i9ZGAMZwGSz2PI8QFmEtSc1FlJ0/9HMqxcK+eOyEq2XQGJxhBMeYLFjOOe
oS8JLchS0spy8ISdOfXoBhM8AwhgjWuqAAJSN8JJkOiBgVj7GWl6Fg3XoF8OqFDmLRLjJNCY+ceg
ZM0l8mkIk0NtVCZ/5dtZgkPw8POQ4pt+HXYXv9Tzlo3ltukRfPeHYvaVQsrBQMR+fN/u+SXkbRhb
IZpZU1eezw/kt6PsI2/v5DGAody3PxsaBH8R+piOayp5LhwtlteDEZqCGLcXtxoFj3xuUQcjOwmg
ZIe2u3bkEIgP3SXBCJ8X7DMr1CkxIY7jqv4T4Pik9PMnZQGSfjVrVEq+vlEP9KQ8K30jARpETOjx
w73TMvuqDutnVXto6pskqL2wxUGdUuZPalWkTqZuWCKQ/WCwF0iDFqMrHFIkPbihvm1rCWJ/ao8S
U2sbW9Z33b/36VI+t7UQF2a3fogGPIh3WdRZNSprTZO9hKy/CQmh5fr5gqQOUOpMR2roy3TW7e01
FXsZTi4M6/HfU8dQbeOtdPsHdEEusP97PB8ycxDJezZUla75B2W98pOlL2HRQIotx98Gwl1vULXc
2O3lTHypUDoVq82qcI9/4nTTgCc7+oanWSdw+WJZ8G4fRIhXcQLY/NxSnYtO2iK4M3eEmtcx+8lr
cbSUMi2cHa3swF/QmIvWdiLwuCGRKnGfhhIGJe5Ez16aZzJVsKhUUdNeBrqUrieyZaEYX47uhCR9
LwtXKeHe/Re7RItTQPXReEbJMDixkhbd7LWXK6ssJUk4r0ln/RsDPCq1kpH9A2MXhxbnk9WTaZIY
HSZLhEgF8zWZp9ScJ9i12MMqQbqKytZ3PQ6L0e4PHihE8bfxpCETGTlEKGVfem/6MCitGoBfMWEM
eLLQTQ8rTtozJBeUNyZoApPZHqbkGlWUCPteXYlgfsTlpbmkQpYfo7ajdZTzLrOAXvUBWq8Oy3/h
BDu35uSU3WNir4OVeJa0bT0XnYZdXMmZm6clTSzy0/qfKX+MkpmGqoUAt6aTu6LxmV46qJJ7URvV
rTbxR3bOMi2q0V/P72Xk3dmkJBEVNdf+/4lH6Uqgg1hG4xvjPcTmx6JAxSJJDutT+kJGeNEXkShP
0ia/iLQV7zsOkLc4OuXN1ZljucxHs/mnwLIPJxrfrgIyATc1gjYCsmu3jnGK7IuIcvWLjnxt5QWa
UWga57HSWndgmrf8pvGlLvgWTXr54I8kfnig8QftcJFWrQX5upVnJDee/GrI2WBA3Tkv8+xL4MRD
egUCaIczKv8LLCpkRAD8zHrdS2C6Jm0tP6BSFC16NFybuJaQjmi1R+e+rmkb4GV0+/RLBF5h8Co5
t47rXRRclK7A8djUvLDmVoPi3TXETrEj+QT0YBmOmsE5KRu2pcUoP2+PdrMHZIWlsy7HZjRR/b5I
QwuU+St6AhZMQHoYN+V2MR+nlSNWbou2cycJg4O2/6zwq7SuAzFj/ytEg8/YNDZzC5PxSKl6c4zw
PFSDJNH1jsA2bK0vdg6+d47BokmHu4pDuhxZ/xT8u4yVnoO2nWmwbS85hERRShcynWCWhZ42bJ8D
tgRY8bmAUn7MDJVjLB1xwWznvW32e5FDEyqMyRGU5EEQrnyGco2q9ZBOZhK3CZw7y2vKXtct0B28
UIiTaMD1UOrQ9UG9EaPzzI5yc0P+h93kdR31rZlydlJOedshl/pPS1E+L7k5ITvl1Z12OrTLkpWS
BOwX17Im6YLKzxTca5Hy3KXYIyZVVc5URd2PD8+tMw1NfBlf10at5SFhY9BBoJNKLNfBkMB9C9lj
sFHe3Poab+dBzwTaipkjT9+/78YdUFXhBN7W8nh52bTQ6DUWbxNW/R2eh2PE8zUyeqX6Ck5fB3QN
RBIWVWWeXD1NSVKfq88f75cc4BJ6FOmg39dVibFenDJuxD1gGIRityB9aVCVEV2wbu6dXy6fjgpp
P5GA2XBR26Cllvk8esTvMY8UFLDlvd/9n8lHN2EGuPhF/IW7Pq0YsE68EKTVj1wNFVKmXWajQGjg
GTT+N5XM9Xepd1itCgUN7TU262ocZDBZjkX1Ah0Jpr3hUSBod0QH5FsUTstzsLHr+h5pyQ+72fVp
AzQXedbfKTr5UXF20aIOHGDttJkoiDDJogFUnDvMrjJis4pxtjjFmZF6r6Kkk+o6JhP6fgcbsIvd
Gyh+69234lgjdBqxFn0p8fKmDPwA88vhfDCslBKYuSW4JC4vclhCAc47JfR3ocw0yaJO1/oF/zOo
Bh9YTB4Of3U/PqvqjHgH1MncJTmtPwT25q3jpbg11Z5iMVjmt22XhcENOpf/0CjiYCa5/1p92IdT
bomLVVyycoE55YDDFcuA6NHX/FSJ/4a6UZnLNv5gI9JSLFlcWHZfOihxtNdwxFXmX1FA+vZqHDL/
1+p4TRGRDGTYHbAPJ3tMdq8YYdq8xg7Ypf81jO6LcpJjiS4Z7jZG8y6R4pr4nrtm72h1RwShICWN
62vORFeXUVLxuWsHm0k28qa/Omrv7Ckt1efu2cJmlJN0fmNBsMy7ktByOWDrby2oa0BBrPsMxYAj
opffDQpkdCnr4RblWGCB8HGUJ5XdOvcUerERjGZhHHMYOx08V+6gsraVy9Y/n4CEa3aSphk+zbAn
+2NpZ7HI7gFuRTVc/5mIzp7Rv85Cflq3/lVsTGMpYt396kEM6bN4FK9aXOdPcLj5ebSANtNiF88M
SlJkLFL/W8QvOv/clbPO4q2NYdvv4dGdZdFetvVGvd1BJpRBDSqV5nbGAouHS4rhe8UgTN/qFpkc
bQVCYr7tAKjIsCYVff34r5D73+z7xJiVDCIu51Mtny7y4/ub10/Em1v3ABc9/PngMHIP1NvBa3Hl
xBDzSnZLB2OBprPwQLZ7FXaKdEQMyuJeqQL7GdDQPMMqltOnI7EXdv1wGysWQKaojPbj8L+lQWpP
YKau0w4Slg8siZ5+9jm9yqfCwrMpBLhtH7/FMeBDoh9/ch4QAaBJFhGWjWH2op3G1RFAi99wyRKu
uh0V2e69MwahoUF0km2mbLwD+amDdkkaJNLg8W1sVI+Jnoj0yqrx/VcxzHD29mkh6UncoFphU5U+
NVXeH0RdxY/cQ+FOZK2jYCiJloRnKyv9/5X9ZOEHapojmcbBidlYVnWoIHlIk+WNvhPDUFQN0PCY
RqYDC+xF5hhUq+b0/5NR/nliI4eBfxW91jrmmTIPGyzN6zWZ9u9nqM2V5Mwrz/N/CoXEe5XtBuVX
pGGPKdVD9W3y3ev6LwRYFblssX8Pp3uNkjNZOaINRQO3dOwiuyt8MhlFF1RdEV3dDV73KC3LfiWF
AJ3i4cbOpTu+VRcTgVbMUDgrCaiUIuaGfbFw8YJb1V7rNVE2d/uvtOUiFrhBxX0FZbTeeEhuL6Em
zF5gtGROb64IxkxpfD9PfqQEyv3i0x0YBKgtWaI+koz+FZlrsEMwnHB5ykEjRzgT5lasmovpvGQ7
s2yrg6Bz+pbNAqYVL9XR00nd8ae63Q3Ko//ThxeJ7lvbJSY6GJ9/1Xppo3VQ6p0E64G7oRJGr0WT
paGc3tHE0rslbAGhfY8Ffscp2xZgiCFxDG3sjYo5/9i/lcFJ02wo6K+HGxxqfi74qbiki/FXk33S
BD0HY17Gr2hGwtI1AzzOxnp1x+r2Z/6MtHoa/xw3j8InQqSscJIFaFDaPFT3YnP4U6HXRdmACTnZ
CncLGFgXIQQbaQhqGiBJy/kuotkoRa2brnFLN0SYbFe0CjUrdWx1c5DQOyjbuU25dfbWDnLSwOcV
1Xsp9B1/R4By2BD5fl+8vqSRZkIQeIXjplBOeUiPiWPlhexyN3iyA/RX1gBQaTuMkGkVvkKCuDGy
fubly7Be05UYxt+KlHNpIrvyj8gYACVqhx2X3C4D86ontoSpnziKSyL2tMsvA0c/l1S6KlhIs17u
T/ZQsKZs+a30iMNKAvbnYViuZF5H1HGa+cQwuekc+MQdN3DC8DIJ9ly+p1miLKI2fXuZ6fKfQWai
2TMd9e0ICcZ8IjZ9w5/wzuX9DL415LGpfJSaKJTzUwGZBMIugsFFqfFkvpF/6Ut8PRK+mYOfXPch
p4vcOZsi0fKwdRxY9BRich0q3udFij6ZxICAcGyn4O+uDSKNwtr6Z7OkHxg7XXOmV4Kciu6ylMuE
uD6sU7fd2po3HxpnSByaezboAVVRtUb9S4pB4OY8yxSNo194r2306ncJ/rPV217yb/HRWtU1wyFw
Ct01TmMRxfXcqd5j4IhZqUxiza2/y6G3/5dtBlBU4h2eVOnvx0+4UO/FVSsjNeXzzjq6wmwIqHtf
CVwDVMGkpOsvCxcz4hP0A5Su7XuZzC20ESUbwYgttbfpKX948jIpjaOQJ4JQ9+0SVgfHF6Q/TJFS
t7SmJnCs6tY3FD7ZT1J9z/IJQT199uEZq51pKLSidxHA8XUped6wweq7o8Mk2JJQQWeUIhb+vO/d
19hpRt22h6tAaB/KCnOWiu1GyRgOdnRhJT74oAVS7vqFvnvwQDCRwqzGSzTBPF6qNFfGA1m37SfM
YUOIDdIXJhhEgJi0+ukNMD32F0LI9vuVeT3iVauU4fQ9+v0hx9uzM5xOp04KWkDYtvXutSFJ59/R
CrQnsRGxfz8JE6A4iPp8GoTeSzQ2EmmTRx/lVxc5voZIggj6d/KOXwXdzP83y3dWS/FswaTA0P/W
7YQWDn+Opj28x8ClEjLq6hLEgZDXJ83kaHu0sWGcRbtCSFFym9eCP3Y5EVSb13xtSJ8Cv3wF2ay1
roDoyzQu98cyQvl3+IGzzs+nUSuasHiENip9GM/jcrpTa+KSIg8qWBPoDkwC6gDOHRpBA5fuH74o
VfClHckZKB10vWZfBGjZdo2TPNOQA0KmSIFms5p13DNnKNeAWy4bdTZY78WFNSnPhBnRdPXV+p9B
DfbmYEaqJY5SmiOr1cZFStlgavqkyPF3jNFNkcn+MZVaHlDCRM22XYnVN5o2qY2u0Z3NxEJ3chnG
BqAgCIonNRgmV6V2lj+HjUGu7IA5FLjbZemtHMoa9h+/u9Hw7y3MoeyZyx/Qca0Bat9Ew1SZXiqo
mzNuRP4SfnVByDYnoYEva+6YZYmnbzicz/DTCdLPL2YNlT3aIJLIWD/v0wDCzAzur0UX5IX5/Q/o
nZ8TFLSIYMwHoag3H0rom66ZLlXpIAiS3qTiPDLqpoIB8C9zS4Mi2QYuPIPT2D4Ma36ye7s29osn
OwVKUU4pspOv5HeJrySpMJ+b8T1gaJ5iS5LICQv379hVUNHJZ0+mA5DYFTNByC2IF1EO4wAzJ5qa
gwQs+x3juCOYyBT2DoKWhUmT4oOq9ojepNSr5cxC3DB6RP5BniiiDSCR0+18exNydjZO3jMKurAA
84eJeYA59PD3EaSLJfCzjfpkyITExp3eL5yq9YXPiKQsLWaPOtiDX4IOEpr0fzHwKRpcM1q/Xxsh
Rq+ZI6ZHkSpyiOxHIUpLw6wQiXLSuqIudbaA+AQ8oAYQG9109CeYUX8fjrF2ry1JF0SoS/SjZqr3
n34GK+R7pyD/Ud094v+DDBm+gzc/phR/NEllV//mgb9Vh9AAK1yRtw+E7+Mhd3/s738Pxd2CuAll
bbvayR1GQ4e5xONFEAAdf5sfxy5T4KhasyVx3AhXt3fYDW6qdamtik+TvbzbkbljtmV/UG40hVpE
ksdcIeLoMHqGh0m6J4W0CFzsxk2kaAZs4yRipRb2iTQdtCAmgoGhzXFTBlM8iMejyiIMgJcOy5Ut
kIcdpGNgrSnpEzlVbNQbOPwzQXgnWYYMSSZEJZD/JkmLDb6b/4QluoA874AywRRd0T7aOrv8svHw
IYGm62apr+SXaChkCKOQyEBqFm9cpiJhO0RRYZ0cDxCjJcOfe7HVidzHxzDgOxt+V9SOnsqpHp/q
6kRRlRykNDLZ6ViFGxH6Pd1cACx1aIF8bxq9kDJYyg0kyEnVZ3yHDmZ3lgkNmev2JB8NX1D7wxQM
/VmugCUfUBvvQy5E99B41tXk9cNdSr6tHInbVJfm9pfv8zvMjNksaEZOeMJ0L5t+FpfXpBuxnYiZ
azTd4wMC/2sBAemA7jTZAiuW7/gwpYF2AtQ4WNMFAieeQyIPKsNMefPa69IPXsYurFFGDgz9XK5w
+AkvxLsCfPkrFHTN/82d50eRl+ey3cFg2tjt54guWSdNPmOqvoK+l06yNyUjwl683gF/lqanOjJZ
koqMGZpbr7fPSHhPu/52jELZHGD4XYqloPRKtygB7yWtq+sJa9jwD4Z/+iRwkVYz6emHVc5PkFsw
toFFe717TlGKGtGFMHxdE0Yng/QzzWivKFtuxZjubbfbAoKL+iw3L9y2ruvS3ndzmUG5Iluhh2Kh
mL/qHG/DsBoacH35UwkQOmy7trFIy6sueFcIhOp8addDPNLkQDeniSjYJ7h1Mq5EUWjVwlijiVi3
eRkD68yvwGIo6xx2BdTZPmTA9lF1R8P0V5N9ID4yREfoqq46pIsD/tSbpw7az6ZTgjKWcEeaHCJa
xd6PyUQTU52/VOLGEvTtoxwuD6IshjLAbQ5VQaLP+UINAcYxC4Niv2zb8YTHssU5QUGIaxTtZRCY
glUjJvJqX79k14iHTvlKrfXBwwOkHLSZItiqPzsjUHnoQ1xrhabrPPN44uwofJOB8eqTtMMGzDwP
y2LKE73KvEqIJxFScd0qAskg8P5woj99RkCFKHdytHlzcjUNmpMCK57waChU29V8O8MxlWNNUpgW
8h9GNVti7xXoDeo1/uOlZTgFJ9BvCWWs+Sgh3HPuafsRE1uoZ7fF1Fgv3JtyVpKcQxfoXNCdtikz
llpwTSM/WxlkQ5ANlgf2f1Sg+iiputlFQWJPbm1eIJ2PpESYy0YHVyRW5gfTT/NhWlpCtvJxJSqg
JuX8ppSyeDgnj3RTxQQ2Tu20FfLFVqG7SwjszUjX0R1Pp+8A96IQnUUesODILCMl8hjy6ZDVYFI4
kiZePTDFE1B0Uokd8eJrapnU/Gvzv+R888E4j5PoJdkrX0q1pLZtk5S1m3Tspxol/O6Ykb9GU9YR
4Nkmy+kp6nxX+Jm7iupnh2+o6b3/K0lXqe8Zp8G/aQ9onJHa9BeD9JlXRT++NRM39wd5JZGUe+ys
B7CxGNTRTB1inp9hfOJ3wfVz1e/EDoqNaoy2u8kGmojTI41zDvSvQrhAJsUKu9MRibqsaEevRe6D
cE+rzHgSnKY2QZ55HNxZ5uBYzZ/8cqA48tfPB+1La3bVNHvVeIxSSXXhGZbwi1D854sImbo5h1KX
SE/vsLrgIQpKWnUuNuIZUviklHX+8kwgxbMTff3Cznka4WMz9zgYHwYUl8IVBOLTKvBU+RxwnOKs
S8e57n7qO9iVYIShcUwd/yXXwvT4LWXmsL90eAdDSUpA/gZ4D+vNxGG6ddMxr11u/Nh8AJ9uQKFL
yAaEkJlYq3myx7oYTNElRUhdZbsghxRlXPgr8YIGx5rP0A6R/+bIJvnPQwBvVjaYBvZ93T3T7CSF
EdFjTQr0EyO3W42ElGzSKrb/af4ymhmmgQwul13d/iamazdB7BCd4kIUmBPs8vXtRLyBUZzBhhwq
shcQoHmvH9Jzg4sHDq3PG8ZZHjpTMKayFjpQ2GX4eJnTfSCpjjfqXSV5qEs/uli0wa2ME2oZEDvi
TTsfw0+2YJra6/KAXy4qyZppr16EhHwyIaLb2pAnXMNjo8kHfiJafrUZRpZjO3FVbdS9LpjSnbC6
1b36Wi0HhTzQ11uXneaid5LknCuXwP50PaVJerLYuGU+d2vGwTprLi4K7DQQ2k2mcunNUUPONFm8
dr9E/gf/tQ+aPd+GhHDU29oDBKYG/5Z6UaortpVYZN/Y42oGqtJFvEOQQxSEnynBqOfS+ZCDGeFQ
p8jYc03XZxtfuYwbHyyBFpXAdI0NxQKXG3YLARnWujCBPTNMnmCm6+5crSLRmk65opdUTcTEY634
dHbWcZrwAkP/b1pcSKZIB7U5C0iZCP7jwtMKWB9AXEUOLnhGLDEVze3rAfb13yxMackM1u0e8C7R
a1OkQzfQIMynoBVVimrmUoXcNTGHeVZJhkx55CUbxhs4ul2wqF3ks0myE3vz6a15WtwhaNpTYdZk
44+nqnikyNxP/WBWMZQMYFKSSEziV82GgFeeblj7SVRQ4cgBYbjqbooEi8lGfUzk8p/yuKnhTdMV
YXoPJNO0mKySZXEsvu9DHAdj/s5HB/eUnOLI9G2YTasQusi9ANkM7w3tqbitXY0ZM4EV++3g+l+o
NSt6GLiKcso+qtUrGizWbgCWgXQdcmudGKFQscPJk9wg7XOUpLxiS0S9Dg9Rr442h66SvRODcrDz
JqJOjznjVirpOjD+5bgKVGjE83xyXBjWWufOv8TP0aU7fkSo0JIVarKpIMwpmIY6PgLgmG7UFyop
mJd1ir43iVEv7wpoI51j+8Nmuf1d8O88Hk8tBpi9J0jzPSGzBcjKvNd9KV3LQiIPFgwuIbHHo+tV
nc7/zBUpsbIFBXIMOHfS2kNsSyftrEFBSih+2aSBWC8Sm9nCWj9hAHBFGEmzfNSh5qxufAckV6Lg
MAIAzPdM5sJF0lEWnPKnWqe0ntCID+gPNC8qXHryeR40Go3urbRPolnBX0FqK1B7FMgkBwcNoXeF
LsADoGFpdeqrdLy0Lm9pym9cpfvUnTbsmIykhi035EfXWkY83eoJRCGn3VBeCLeUOejcnMHp0xyQ
GNC+7ALlpllzQpuRgyVGkF+LDIEQcbvW27K0rawCSKp/15c1j4n4RGA7xg6dzoZJzWrYTudx+V45
4OZfwojshBQjjfoCM6YzJoxkR3pKH7KKnfy1X7nxRkRsWkIoAwloJce0Lx/pvkhv4RqWwJOXC6Z2
J/juwg1oBXGDtcDVw7g6536Uz0Ecxd+sLAW/WkmEHu+chZfhGsmodQopGmrdEOdMSHhos5L6uW9h
Gdjk7cfHQ+0+ToXfOIUtWxVKj0tvycfHCAqB/LSYklsuu30KFLUmapMIRdWPEFdNAtzjdjS7EWhq
2j7NMJdp22MDq9oaOwYG3vs+EsWcZa+kZfwc1TNB7bzG8ywYZ8LQF/epT/IP9WMHdjVLD7qGoSje
E+1xpL6scbI3BhJng/2m4NGaFn60zd43nN8/4MQhohDVZRIY24q/YzBkBip8hOoXVr6FsNDf0zH0
ftZZ2WAOyySVW/tq9gHZZjcVef5wmDR6BoNtS5kbeH4rnffGBxb/lgMxnFb8PAtTD9eQqg3w2s6N
fwSZciOKQU/XMGtFgvHUNmbo9t73owRFwDJgdWoq1NsW2MhZKKiFt2RwcNfnsa94Sxzw6ZMo9GLK
LLA2iq0TGFr2TNwbpLZVZkE+zhXCf6Q1UR4N3Wlbh3iNQYsT24nSmzfRFPiCCqRM8/7TMA3WaT9l
RIqbwSNKIf6rUFUf0/03A0OA0EDXBZr9QOWGEvW+NmDQpgUerMPcnEGQxmp3xlb1Qp3rjbmdvLV1
5Zd9AwWWlGSjjY7YeHLR0J0tqP1/pMhRvG8CMKmT5nHnD+mA36SZvAj6K0571PJ856T48PmenDa5
UuyiUqdRGqGyEtRw23SkiOvE/KL9CEZEyOB6h2FrrY61hyrCDYo/7YqZUpKJg/Dk4wz5lqaTTBX9
3br05UO0rRR7ouyDC8igN/dRZcOVunfd8WxytahvIXqVHvP/Sqw36Iy5ozly3Y4Q4NL8C9Teyp3J
lRDdwrRdGywh2S85pC2SfRMErna1y46Wjy5ZF6TybOQoqtX9ZHaTxvUHD75NibJE/1P073cn8bRK
L6WWWg5IH7STIqNOYqnkfmTscHABeYb0IYtshjY9ZsT5M8UeS+zCSKGCCmq8SG/oSTKrKPg2bAHi
9q6j0NesEFGeEqQ2TEBL9zR3KZAJieaojNKpaH6RVcmDVPhZJEMHIVd+KqCXUE1pfxZJWhxkx5Tc
zy3koV5GH0elQSMIVCNdGUPJ8ZpUIKlXdsstZheEyvLY9piWCcMj9fghBM/gm/pITqonDaI0oARl
BE0GorC3qgbgcjaTxlJttAi5B/g3LVX2OdzL9jZ/eZOokqK+qeHfHdE/dzKH5BGyBeYTzRtxmHsS
Px7ANg7tMbZ0yXFAhQ28dGsRU1pgNL23deYP7SfSuOI4Vcteo+NiD9IanXlNt+O+G29+HZGRnIOO
TZ+NwAtzYp7QmLlJqu8sd3hecP211wwGd7/WKeOylglkqgFRTPRkY+Lqnwel4qhVSRjOX0kTNxw7
Hm3/ix0rmRpjZ3lF6AR+6zfEF3Wnf4Pkam7Z6Ugixwjl+SYmq7ZHSGHFgUoxP/O+gNuCnNSYdkh/
opaJ8Q5pyTlX+O7kwJAdCTPd49mLA11/7kzj99biIaa0x2ZLI5i431mAtWndslY1xJ8Udvo/hj8V
d49KAbdgsYgtWZanaTLU7ptv6I9RBmQKCn6KFwJF1gNODO+dWiTzhjxLdSQJgjAaK5YEbEcL57BY
y40ro2vvX5R5c7OYVWj7cLFBD/rr7Vk0tw5E8hZtjQfJeUIkDOzdK6lzkzwc/8QPnaqunDLBnNbN
RWKR8L8w1UQ0h/9lCHs+T12WViezaMdD3edRcEGMFVTqKVNRX4ZkQ1AJICOy6hjnnkHPyRygpoHk
XvX3nRV4fMhjVRuY0hIsyfGusyCqlwE+gfMQfjlTNyIBvU7C22XbXakZR2uWWwsyWgq2N0t54Zkg
soSVT1tijK+3Y1WUJtjZVAbR3CsobbF7T3mJJc7YBtMTse3h2Dbf2gtGUNPrL3QpwKMg8aU6UvDE
6D99MQgpK/WQJqeKBlLvAv4MhvKrIqNdK56IMt5g0bOqADB4Qalo15rSDjEhwIP/YTURH9pDpE7H
GrkYiwbLn/KxCdDlOO0J6W9cMlc+RqAzA66PPygfELYnSUITpiLJgJ4rmSh8EZAqBEaGWyWsOyEY
xja9XlEYUkuQ+k0gr4orXhj0KOnpuG/W+awWmzXD17l50XP1yrxfqTbf1oiWE4FzSbeuhi+aF9fp
ZT4Ezwr+wv6rR7NBCNYmCmnQ0JPEW/WGYTngIOq8jSbAIFqbboF5z2Wn0kZ0jCkOi+D/Ca8cIIhv
NZ/H7OuCrgVgG9lChVZOerLxPimaNnpAkdGyzy4Ua6qfWiCMTDAIYZqw3MNaCFO8Ir0OHSFT6ftR
yj/kG9NuSKIYYcPhQRi6l9/KnTDaj8PJn32YAZQT62k/KCYy6+5prZBhbd5WbFEq2c4LfzsapHfe
LSWFyUT9tb7+ZxEUU/vWDXXe5RaUzjgmJ2CcNwXdq3x/UtRPKv144A//u+mZX6WOeAB/DVZHGRCq
dg61dQQDo75bxqztKl5FVdZaqRWm9CIw+Em85nn+1DufdUkKcZz7GYVd4tKOqqW2zlQuzYsbz/c5
rAvnRpUh9EDPvnR8TEb29IAJtWrHQoxF4WyaanIgGCKCkoYDsaS6J0t9OWPkBuf733DjvyIZAgMv
R2/gOuIvAT3r8ggqLfZmTcUAQ9JL+rBYAebGayTyQ8oNJKV0EVUUX9/9w1Nv4ii8xjlRgP1A+ioa
RYNDEft/smtfEQOwfT4nxhYJ/LqF5Mw5oE10waW9WFy+QErEEDVZLGbgqUvu23gFjFu2AHOvVsjt
ojSrPXE0j58BmN6n4weOd/d+vjWUCLVIMk1r08oAACVoEssHK3ne3bATsNki8VBWOdpJ1s/9/EQH
Nb4fX516N1znoeMhDiY03zIqxzd+bLrhlHG+DSHR8iy7dINPJxCcxhjeHymH05Ue1b4nGq07n/bt
VgJ+Or5iLmMl+46fPRxMLTBafKoDmXiKGa91wzJSVpmzvmmjifa4GyzLRpH3ZPyixViZnYfzp7cy
895CNEWFOYxqi/kE38CXQvrMZ6TrLAFyZxuFeLdXNbn6BF1EMANRIVKrM/7nuVQfLjP98HgiQogb
y/FNuqIAaaS9vBPBi6SGaxT43JsmCoC2W+j4bk9tbNGGQUA/qRyKhhWV+5FI7eMHtzbptDsaURPg
TkRdRognMyLRiUaitLZ+5Np22uuhsYWGKJuCUI7M5Ayw6NKVZrsFXCAZrI6JSCt24pGMvjc9Ufi1
3U44kTfBtmrBwtNKyhot2iWjMGzqhO5J4tZfIliLgMNBnCUjGnm++2YszPVzSZlamaWgQGb9/xnw
FWNOU+4AIqeN9uzViMAob1c4AlutH28nZS5VnZbhDKULmtF63BBpEl+p9juFX3xr/H2zlrzIP+XU
mhVs3u8kXbyW1zLdUm1/bTx652yni/I5csweh7diHbXAPeHKf2JIBmur5FXaJrap/85zHIctQLYW
ISr455RD+/eoM/9FmnsuZV51M5xXfnxnk+UXHKfiu5jR2Mj5NxyMh0yfY2ToZe6FCnBt1JaVSsyy
TleUyRHQEaEn8v7M444ihgJNQQHlmiFbYf7U36fEgAgFIfoi6uV//eepeA9toiG3r4IxF7ayWVG9
Ix4VC5YbvGjGi8i+U9PDLRNWgY6kpMzPaG3TNQI4yXF4d0G1rBIozkCBav8dfsVhS8klF+26pVnF
LDY1WXMrUIHQD2MlNEI2DLHG+I6RCbvKOxFrn0xSZxA49Iqd1Pcq1teRNbpLE7TpE4+lLfzmPp0w
9G1oRKJCc+tkB957MRqSWRPKRe1yfKKrUU7yjB1YdMnqwnYnPLb6ErS30OhgHftGJL8nzmqFU8ey
j8nt6LAkyB8lzG2Sht8uQMBfhNjN4XNV+w5k94obEJTdeLZgChnuIiw5p2MZpyKK+AZmZbhAQA1o
y9trcKx1rnCIDBZKGreJLl5yA40w2ZhL9O2I/pe9irP8GBOTSSj8YUxIUqWE5cNKCoz/YEeAc0PC
sa86ZV3ZJHOACwXEVz1/QSibED+Wc0d64wHh1aO9370RV2hIjglsk8xB56BVGIAJ0o94IqJCZiW+
yIm+LevsmPddttE/sWH+XxzoyJLOb4x2cCoBtJ3bhJNzn19hhgMdfFPZuY4eqDKD20r5K4DlNfqb
vC5Qjie+8D51kstok5P549FzSg8+UogVzSK25mNR5v6+VQrcuA0+vnuEpoYwsXc40MYpr0PspFFT
QoBjlzWXH/jA6E/FgJVQXfC5Tmgn4k5SoGCVZ90TxsoFlE8utA11OJ927pJQKeqN1b5nt2Lr0hZg
uKFHK+syyOz62Id6JfdO1wUpW/BQqHYvhLnCMciBMOVOAVWp6i9Vylq3oh0YkiSjvwXbRDx5aoCv
TmnqZlPULlcswOOkgAKsAxhsiIrYQEYzTMXCZsxGCHmLvshjrw4AtflrMpxampsqc9WQ+lMtLPny
sdZXdRPhT1MFn7wm5o4tPGv6299jFdNyau0BxPyV7wGy14cUIFNhqda9Z6ZFRGmlIiGav2gpIVf5
3zwrw4S58Yqf/IAwBZSiVkbLg4XDY64tdwf9QzW9iEFhOBc8lbqLeB0kxHr0j8Z1fc9qk4HobjXQ
UQOO1kgXNBmdbe6zCPbpMsqtiaYQxKHlm7L2cQQZuThcoVJl8GBtPs5zfXQSCXG88z50+aCMXdGB
wNr0klqzxLrAfnh962CnHqdQjsANzGbAiXMrdO1rxFFuESJMcZl7nehooEqOU9gjuVxdaywjP6aF
vx28Fro+CWKfDDcBphMm1Vy8AiHcukXE8BpXNLmFzuLSbuzZF0BzSailxCi4Uq8BZlIhumd+jZMj
LCrJJLffV5xQtIHlTMxYI+5GP7sPd2zG783c9FwGdr8ZPgTzcc6JchGC7XLa9qX+qvoZAvPjdH/x
A0dikOCXga3t+C7JgMhM237vXhVqo0FDjLF4bkhs3BBgozjvYWkYO3lCn0eg8ROeGYMff8eZoJe4
xa6sjKZLNmA968sLhD9ukp03nuy5TU2VVW5l9qb1zRCHl6ReFsKOn/fCstXFQMwu2XtByepR8GL2
xcxuvvVEeESNaD9K9b1Z/8EuG0saS/Hr9nxV9ESvPi5LHEqOSXEfNSwMYjFz4W9W7kNFNu/isJ4A
AQE9qZXAjWEOe11O5+LL/4v2vuS4yajkx0t7pVuUsudWs5DCPzk7xp4i4TwNKLwgBixz3AH9kvy3
HRzc1WO/fUhzOZ5ykktNhQ0nO5ip4QmlywlySmSAU3WljU2WkNwVNrpPIo7jNj0W4Ww63ifUcW2X
giTp5nVoIDGGcRK3FPIzpFnmWHu7QT8AX7k1zZEQcnjwxiixpJVJhNu0ZaIGdzWv2lgKntwaYKGl
NHOLofjx0VepeYaxtZ5PSve4klJtO4K6m0yY/GBKdDZmLM9aRUTbI8v57VOIBe1vNw7S8JbsKibQ
6KKmdO5YD9DQH3TTG7jzXd9XU6XjT2j5M6l9Zjd9M8qYOTN/9U/P9Oa+Y4eopscdwNuR6HA6h0gH
2PNfFIVaTuf2xGCV9nv9R1DmGLz9FYfjI/lRFXJX1Op3BN9Mg1yYpAm6GV82MPypL64ABX/0zxIQ
+sYuuZ3/NMuaLFKa4Cbz6rOXkECAPylsTokPrJzsQJexposVWYomi4nMv7A0WEcaktx4b6row0Z7
8MR+H/MHjEnNNniUL7vu/zeQNYgCRfWouGUNhWj5OJyhwj010OXNySZXglo8svMyIhJMRKp1/fhU
EWiPU/OhJLngJy51kc0pHzw4xq0vZ+AjlZHRehh+Yr/+HpJhCxpmbIg0X3Vw0prxEp5mFbhSHTep
WnG0kbqL5T8FmiszQmeMIoQEpTOSIM31HVmQT3Sa76D0Pt/dEn3P3mX5NFir4XyxO8Nnt322koul
1FYoh07tnhnr/vAu8qhkpl3ol2PG6k9J2lIArCtPYUOopOeOyOm/C6V+UQNelbsM4npXY3nR2Ayg
uXL2zjrrufsjz3hF6eAMZneqagKx9bz/GEByOHzkxAHy3IzIdbuHqzxQzDRquhE3XrM/3xvYF/14
a5BgI8kYVE9uuq7OLwDsiIHth3I40mDs0Q30eRfk+rwQH5+4ZdK0LoIPU+b/isGy2FAzpNEnazeS
zutCpozsuoUZDeMmP3u1AmDt5BBltG+ujj2CQeYTsgALtT8WMfFLHJYEJpVOLo9KKIf6vkn7u1yS
gsqcIbfiA0B0PFk2j7alyRlUJ7BsC2fILupyAE/d9y3ucouz7lsfmH1f3DGgTPUbQD+Mg8M+cShS
9jwaXAvyyg3eHvFFw+nMLiYtzYBdDEwjdJVulVZsI0df2EIam3nwxkQFxP7781hD95eVnaxxoPkH
wI4CTN/QB//de17/R+KERlAwoqKryuCLzbSYooGiD7RSoVGlorb/FByMWaJT4m/eU+bSTR4FdPcb
QXscAPzOhyOtWfr3xiWM2z8R9SHYnQDHzRqtgITXvlz/7Cz4xSIF4fVw1pK3kTpq3XmiVMF/BYNE
P5ydU2QhxlaY6yl/6O+ZT0ImgyltFXqfWrSf4bYratZCDZbG9FVclc3tgSFmNWkAYuIh8kwBJMv6
XdgyjuLufTpS5iLZW37TqlJboJu0HbYPDhrJv+lds05MNAk2uzj6d8X4qFB7vDwGmENUb99MKghV
ZJMNcru9QFPIAyrVr1iEU0TLDkdwbolKy+/CIawb3E7g+4ghf0P6BsK3HfaB4D0djqDyNIO1qWCO
BrdglQJpFqGe9cC7n17BZCHl8v/1wDWQPxWQ+rTaySSzPuy5wjwcMYMKCmuRQRr9UO7gavlvl4Q2
9wKTsdVvKWeOWIoF71WfPVIplbReOtD7V4WFrDyPhI2WptCUKpLz7a4Ne7qQtx5vdOmRrh5e8v5d
McSBtXMbcabDRp1rtG93wuZyAe0+zbY34GbZTtmAEHB00q+/5+QD0Czyiv4b9CZUeFUJUnu3Puxb
l+bhgju4yzyai9yqBjMsBP/ptiISLHYSDMiEmDgww77mPuwhhOr0kNd4VhM1QZB47XOCbp77uzP1
fd7KmgRaWlXewghr72xJXFte29lmzAvvxqQLD8/R6UYPAwUf19/M0CyUyo0WlQ82n9kagdrXr/px
Onyt34V5WOz6/IFKeKWdUEkzPYfBxbeOQrWJjymQ7J3PAvuTZzEzM8SRxs0JjzjKU693knLf91Lu
hh0FfEmMaG3Zj433eok4+Bdzfp1Gw0yy0QHeP6EE9v10nZ7xHPBku8nvNRfaztcRxDA+S47hYLZ4
BJmD3gDM8XmUIDMG/EZ3Ut7Bx+f++XmU6Ejnk6G/YbtKVZoLhf9VAPMwrfGLoBKtksooDIStfQWf
VqkToJ8udbkwczyyw6xoTFov/1jTVEvrJ7tDxwfBMWaHFhWXwgoRaxs1EO2aG+Oo0AOIzYq9q8ha
WPBo/cp4tq+0JIZZZg9rK77c+DFMGC0ESfW0tYxYaPQ2U/UVF4vooLPfmjn3y/0d36SGluQZ1FBR
Ad6QBYhRYyyMdZ6yG/L0F8htDRKaYoXFZOF6S34PpmyWeZWW/s9hE26KV8KzwEIuIfndSTgZeBnw
N5PAl/EPWR/zeEuZaE8E5bKGGMeW2uLCtrp7RjuSO7ole8OIjoUCc1T+besZgoEZMZpHYBVQuU7k
jZIeSrMXW+kbeALY4769pK1+MBtqXVUJzPCDqGuyuRYVR9Trgp+8NHLA8foLYgvc3iOJGo8Ks6I3
dwCU1Q8RK45Hx67u9d417sksT+qNYtXEs9Z+aiajCIsf5cLNcWEVt5TUK+5YHZqrn9u8onv1n+yO
4KaptpKS1B+FcrlBNm7tZd52uJ+Z82t4dZ3dUiQbt/ex7A5FzCZdLMGQSE3pPB3CWEFCd7xvq8xn
5u8ss+eHGz1cG9fM6bKYj8C5VMZdemuaO0jQRpL73M8G7I+jWZkBrdhTzqe25Grz6BB8mU/4ZhHm
YMLAut1+vCDLt0M7lIRs5Nj6mxeS6L2epYHG4f17vh1LP7u8rW9hWQ+rkO0iMF0aY0zAN1Gkz9hz
7TFcldK3DYCP1e2ktGsHnQno8TOZevxgzITe90gQq+vPMzOR6rkrL2kK8f/EgqLM1yiyncfvMbGD
IDXh4npMtfTPbBUvUe8FG3KlMcs3bNh9XExwBqPYbGe4lMWjmeHsK7m+7iVHVsl8CF4Yd4aVWFFc
BX6viKFZ+Ba8a4/hVbJ3reFnFe4ASA3Xy0DRb22Jf9vZOfOyQOvdW6SA9T/Q6t87Zr9x9VkTHQtx
x0IZvawsIdMC14cJpRGn58HqUqirsY/ZaMExxfKqLBMguAwMp1rLmyTMicffE5oho6eBD2EsWuQ4
AUYc1eTXldTlzNHSA86r9STFu4nD8enF5eAcT1SaUQnLlFqd/H+o2rS28H2J6fx6iRO7lrJ7y9I8
B3lMCYWlms/BNEDKuMdFi2hzmIZarWqDs6z+EMY6npPHC/r8ukXTuVHX+/FBy+Hl//jbAJyJCizP
JqoLnmQryUAWKmxf5huhAbzxFE5NZ+nTw09WKmPbC2Gi7AlB+Ww3kX9puSbPrUCR3Kn+POujDRVM
J6s+am2/Z/EUoBQjSCXtXoCU5Vkj2K9MBA9cA0Nt8KcgtZ+NWslXhiWNO+hWOwdoiyDhkFzWDDcD
bxS016CMUOGubcBKWlHAvMM8m77MXtKv3Vty5k32HFaPFuZ7+X+mp2o1VRuXAbVZiRIWTLpFlPsw
xR8cKK5pe8bImS22+2F5HAu8C47X2nBjyLHsOSr2/NX1ZVyPDkbDArJehV0ALh7LtQYJ3bJvyHY2
JxkeT4Apl/gyFwPhEeFDUOFraGCzZraNEUd+zEb+rWTB0ivUfLn/+6RgOS79+k55g054+osODX1e
IRdnpJtjftH3ixvOvh3W+Xr40g7sbG/C1GMteb7hAw6+ulpdtOIBT+TSyP1KOPh55x3RsB80uCw/
GfqO7fiF10aYX7pE10e0l/uZV3J8KxEJZyWR1xU5MJhuQb6ay19tyxQiCcTRVjNy1UUAzKrwQ3Es
PYqF13Ifj4gf6APiNYlEIjPkcpKYKqdMlsyAdMaDeM8LO0bsiozIZKoyEuVuC8z+hE+Q2IhvyMpU
0z1siRJriCTB9Bf3QTA6AngmDhYx1N1AOwDWIkUy/8Qf8caTbmR1AwcIu7SOnEHxmr4l7FRAjDlI
DPP/3S295CooKhbYgvUc+AxlRMgMVXhBXJOzfOmx2gZXpXUcgdKquhveHUsochPMDjn4uBSo9OAN
7gWOdhXxlGWSiWx96dTW8oYAnHqqOaF+f+HWJ5O5fKm5aL4V5vOq2cX0fGZTJY2YubX/vhMGD9Ib
rOkeVDUCjsnaDWxUcPz2BCCRMwiJKuCBwVJvkOg+lupCTiYMheuJ8+HxxhGVsmHqwNC4QxXnXMph
bDPCJ9dfXRKExfDTrbeomB1kXEoIGlJiniWke0+YHgH0ukFtBRNwC9L6DxjT37CteKMUQAn1dvQX
bTe3bbmQPln4bdys5vUaXPfGGxc31q9PWaMeK8ALME2NRC0OMxnGO4TmHE8X6Oc7Wsg7UhBxhhtt
Kj+ic9nS19BIKK1IxmexkVS66Tk1zw8US+M+mKT+GUV0t/KMVFZJn6QJ2vYkeKyPe7oiWLWMtIna
fWszVWaJbKRUQ1ua/p6jGiQdi+CiGrTQvHVd9hQo/JGkw/r5S82C0UUNai+RklUUp/a7yqXo//l5
2aHO0j8d47kh4ld01bO1DUV/VT5qZFxvqJId5ItHKdBtb2ThOez9n5yWCR+lP6IAb9MqLb1zXIJ8
g0SM6GmMn/tbTN2G0IKeNJdR8tg5w0j5VAKVwKlYXxNfdRKfeoTAZgaPCXAkoiGQFeoeg4icK4q0
sENIiKgrdE96wfZhRHOXqiYnT0vDwoD89MZv4037Da8z8kJqLVnitt/ZteRRNLnkm5ykUWuv9jJI
o0jkjvWZ+Gm9ZfrRg9X+Q9+P3UTD+i0qLntAP9uV/KFeiWJLYdnS9So5yI28j3vi8FjcgRHBsBlU
QoLBg9R6QWE8Vs2uSPDT6Th0A/bJowehZe7KLXgPwRd4cM6PY0oj1LUTMm5ayqF73SzMa6K93Fso
T4mH/PCNAWbX4jzP7I9WqXOzWl9FOYF5/OF3kyJWLgPKyPO78elfty9Lt4pP/x47qf74KppXEDIs
hVZVulgG/YJOFlGocuKmP/Gm4hDgXcmyOxy5ebOjrrTDdoq0+PdxvFUD5YqZSBtZAKeL2YCPISBu
yYAD7uP/iRgUEGCN9+WxPU3lVGzqaZYUE6gG6Ai66UeH4SKavWQXr+ZSKf+wXpMEdyNODHgpzUBV
PXOGW+a6zjlHRNBZYuHgPhANNd6ls+q+pehLmPJVytVyykCZ6A0QBXfdGRZFSZonZvZlVQX7TPq1
baxNydywnWkKV6jW6FtNrABpxEdBE+X/3VAbifVMr3eyqMNFLIYK4pmLqAfeKG5yNGEIQNCJ8MH5
G/DvncHdo7CBLRCqsYmpZUILER8SeFrmnh8Cj+hN7JLxcpK8mdyPOdPqmdZS7Yv08na9NYjHYJdO
VbodKmP3I5Rbja3Gl3lrxBEclt9Ivk0vfeR4mIulOb2Mx4ojWK4RPnV8q8HmpqPMu8OCRnFxk7FY
t/txENk9hmoypKzfBE4UIBjW4s4khw1kozWfn8ujwF5VGJ65LrpQ7Udv4cAHCuGJ5bICWuVDSdMk
iicZD9fSSzFzDmYUQFA5xL8GAyMOVDeg7YnWE+iITpgdP0sQo53SiYt8YHMq6c2Pv8EPBQChW4pc
FudrCIy+F+E5yoi19zrQaGPVTs1hjIjxGqYF1bcRYd5aBA+w/M8jH2nYm7pAQPCtpy/MvDchYFrI
yNi+N+lCVrV144CaBkTlS/0frVMIjpQqZjeIBcRAKqDlrB5mT/oKfqUVOU+NCQvulBgXui4/95EI
qNo0kkJxveEpkGtg0bkoh9RwBE+3juIC+BD04BknmbHIraR5TEJYR88FVJtNq/DuLdX0udpxA9fH
qsq25NtGiLi6gi4Iv+L0elzKpqPs5s6iMhDE9Yy35Nr86qeQXWCCx7/9TJIi4tc2TSHfcHbUcK2X
GB7zgbyhoGn72GRCc7YErgkclTUnpppXcNjTK2yBgvqRmujtKkA6wyZIfj8H2K+r1rAI35qk/kHt
E6OONdIibXFES48uYqz/HPkDULSuiwtD7rmMuKQhBcKBvA9Jjh38TWMF95b2oFL/baZI1rhyNYSW
wCXIF/N7DAIJP0fJ2x8vGVWi/zNWwoMA+vgB61nDLScv/1B85xYMzPCwp8SyMradAFyaZmfsHrWl
FBKs69UAaTjy3maV5GwhQ0DPIRBL/p4xQTXeiuINkbuT2YWxN0pax/PwJrZ/Hd0gAHsglBJCbIq0
WI4mGe9+nBHzXSsE0IOVld0XAQNX0F+uQHKpB/L4bJQRpnlr6ypVnMJZT4zZ1daLaym9vyH28TVf
E6hNR+11j4z+MAPrZn93mWH9NFa46yLWXxnMgWb6cD6/OMRnV6nvIWBAulfsM9v0Y2t9bPywqI06
rRX5NlAVfeU8YTECfsgPSF3RYYbN7lEsmo/8Nf+7r6feiw1HIvYbu/qz+S0Rf2teuTEn4jfX8FY1
1P++Umc/2/US8WV7uQ5QNT4qGkuqmXHehpAWZBcr5ecrU0m9ZGJF+3cdKEe18AHwsrYe0EoSUxHE
ewaZI7SFj0NvWlJwHd++LcQQhCpIakZMHIoJ8b9d+VyXtsH3TaTDamOcotHtUpm9hrLL8ZXKJQGU
xF+XQNFPdnnd/3PxI5tgE+rJOFE8r8bvAEQE62FMRb4WdB8OpK3e43akXO8Efsc7dbR3YiuGg0QL
o1MKqK0XHK2n8u0gvn2fi/w9N4ogVvWrnmnVamKmOw/mSEQBHXUHfGCXmL28lc+DhzbXE2cpryke
wDdVXQdaYyAIHl1rm1/Jnw4asFG5GGUb34yEeqljTITnMm8vEbhYVKNY/ZztLzEykcBPlKBqgwhE
tQSaI76fUzZfQ4WhFeLzMUZ5RIIE3xTrRWp9ZbyPaKhRnkyl/bjR8+OD6lknE/r39BpIjm+PMeq9
AbtN0cKKKh9iDx0HRYFjwPW/qmByxMjbfp9MNQXrCiMdAgw0zJpwZIwPUOw09JpNT2/qHlXdkU9f
Oxg3ZSNkYZncxabkhXMwKrtOc/s+HVf8NIc9tgoohGLJImANUyqnar0EwFEYX6AXD0CKyNQUypSN
yGD/F3Jd6f8JUyW+24DggZQtIqI8LGzArdidtm15yYrt6Fo3+Ns77ZkQwoCr1J/hId1v5qxR4Enk
EHFYaTnc8OuQgFHLFMPQ+7iHAWyvPtyKG3YoKIqqP+kg2U4XbrpRPYYskQOWZJSbhBoaQxO7lhNG
9/RutAu9rPX2dhlQifTRYn4eLt9tBYEsfvr7TuQ5Bmz8SActPE3nqiWbTbfyDO9Y9RWHF1px5aE3
mc4tw5xlY2o76QUA9nbscm50iK5JTDKO0NUPTSYTCuAi8Ylmge2+UWpJaaykvFwmQlTbboIgfr9i
cOPH9eEC5A1t667J7WvwdtBg+uxlhM41yf/ZFLrtPTn9IbGcbSmDfyAbrGC9qU3qHMlwZ9yZ6y+J
PP7+IhD1PAk5kvG0KNt+RDchCjh7KQil+BK+fZyrKjbMI5qBniwx3WuKQ4ZIfj+BCfrlpBK3JTQp
/Qi55IIBswTY+Xgpe7xgl7rNJyU/fBHTlU/+zUvQOQjSnHiz3vK5RmLyNGBOOSDzCzySd38ZAMio
wfDdvbd8lA8wsUhPeDKLMWd61uMsCaJUCxDiFTFP9VkTfKiEJw07X5MVLIWp1mG05BqiKh6IUCkR
v1KBVgYe4PsUaR6iQUvbJeWXZ+L13Vb6tLwyoPxfqJY9F5pk/AroNolatj0ulZm+OGR/F7OzW2+z
77oNwH1ktetR8Hp1VYfHldbWXmcnTCh/nyS7xMg8S3MeGWwr3xVlc9Ts4C+IsRx+mh1vLAGiDe/8
6jngPEqu7dFSzlMDjZUj7GCWz7GB+isv1OisZ7ZsjdBn/iq1dILUVnkzZPCDrsT0BT9hVOO99GNl
kIRu4HIHASLqgWCVQ8RlmNF6WdGIbfzKheuu8VV5yb27vDOjfKOLWS01AzH36Au4+b/6U1/Z8JyW
bfo4IeSTtk+L36jY9gbsxMtbvMZXJyysrGop5VHZoInjfL/c6XQ6ASh3NlA+DwUxPOeBKOdKBI/B
isrLgK11WyYWxVmtz4M6YzySC+AYpG2nticLZFE+08CglHEXoTD7WebrN/mkz9gcsVvoImWknWfF
DCkWiAFcY6Ro5z7t7WEGRPm/3bVgxan0w9+eQxffNvf13k1ZFkmgTguxtZ9299zqPNt32ogKzxrY
bPxdxoVRf+uUUvZS3yJo5z/mDqPJIucK2TqE7s/cj3UhD9VnDI8+s9l/jKVhL92OlZzHxCH4E72l
X5TZ72a1lCjQV4A6cIbNp/ZB84hbAPs21Suuy+6OZPbtOnSprjCsmxHsCzugtS3n1epztus4PArU
oRclbMZKw9zBg3bxLT3tIx571+XwPNcQMSUZfYIqj4+x6bZeX33oBNh3seumV9oE3NTPShsghitB
qCAJoh6kNK9u63fkw/fetuRtyiHbifShVy55GH2BQOaDSRs/IrKlAKxAVX2vSSaKj/SNuZWKyIiV
Hf+eyvKEoL1rNi6h5uIG6bz3VlbCao5bjEqQidjNKwH8KqN3UmEGFM0a5kOnx4p1BvOQAFb2sejZ
eoWQpTR+RGlJas7xskzIuNdU75s+SH3zaXNvBi29uG8/InGr6rnoyDz448Xf9pI7BQZ3w4CR2yTg
x+SqSXhVFd0UKvObdS+FLjzhNKWOONTc8n5s8OwBpaOp19ARuQxMEhVk8PaaSNFF3P0/7cSfEdX3
Z9PcPx9Eyb1uNqxa2DZN+h0PAd9X7u6vuURRyMIS+odA2DcLutxl+K1FznOn4GT7PJCKWOWJfw82
BRihEf83CrdAy195w7tjWQ7l3Zj4v61L6EP8K0uRsmmix0f0meBA5iOkKH9CuRPpCGGncZS9FOez
jIe2ygUgaBNDaQLpGwM4xmrqZIRQfgStF8CODUr1CBsKEOSTXayysjjL2sCQ3+neM9XY5pHVS+Tc
wCjX9ZxXuqJ4y5h51Rvy3WoV9hzPnMyB4xHv/JJle/XzL7GNjHZjikPJyJhH4dIhOwM1+DIdKeP6
agSd/acGWDKeVk7UIy4P6mROVXYltQzfB8Dv9casoo2rLaWxocc/acNPMxsZ2xdivRlW+CB/08/Y
Wy2Oz2zjgMMhIzzzWhwLrqhhBwtPBx1xogrLbRXoeftQgvNXfX/wMPdry3h4spEtLkYynR3XHgkk
rHAsQd0NTaKyKSDqVvPiw+gPSa/EV5OWnQCFZT393hy5Zqcqh2Sa0CLjPWL35wI6K2V4M3cgoAkA
LrN+3DZ5co0PZDAgD2MjHilk0lPoc5PmhTJrKQgT/GLLYsTQZ59wLtoE8LeOwQ6PFSqY3er/PV2A
kezWJyiBq8TMTlwnC6o6iDJU53/uYgH8schicA7geGRvP8LewR2RexY/8uILsOMTufvK4Gl4pWa5
ZoGU4xy4xek0Jsy1eK4yqtEhL8N0TscDd33mCoH2kHsSD7PfTEJ/zm19ku8ewDg9xjVywjN3H+5y
NZ0ofX9J0IqeXcsn8L6qpDgBQrHcgNs1OQBThdavP8wjx9h9/8+HqAIL97ApLHaidiislEvTVED/
CCaSLelJ/8ZhyD/u0wp8Ijv/EuHvukqNmp2ufPMe2wkdN4yWE1xW2dwWhb+ZxwCyjVhQFFhqY0gx
17Y7+ZO2jlGnoiQv1s2wSfAmQ+JN4HLyWvsTG1avbL9I02bEimkOafPYUDNBynEi18sFBXCnWijK
0PcVqBY/ahRxzsP1/dqkR6WBA7cUXIA+CFF0aO/OZTT8GoO/7NePejkzAM1//KJTEv9vP7M2yfSC
k6CAUzlPld+lRTe4/gV8j1pXvJJd79WMi2GVyectrId55ts0Ec4JvWP2FK9AEkrGiAFFyBHvDDbV
lqLpb64OPonrbOnRFXsfI7gDnazDDrylsB2NVE1cVyyjh3VFFh5kdjofctJ/wJ2dLcJatizw4ti9
ESi2HbVdph9eidZe8vawOQqRPZ0KZR5vuDQmRQihqbZGrP1rL34OANJ2vGxzUmz4GCroQhGN/50Z
lorp2uQUqTl2TZ6MT2loVC0MX2SAWwwzfZaNh8qkZtELV6lrnqvWQwP70YVxIkRJlyzCBSD9ovX6
1ZNWWuqeId6azDG+fbcjtra3YMX8+xiExYFH3LjWCLfc0exdARLMgWG0pMrYiYnv6D1CD66+SjwM
jQSsauVqPcmNZjeakBaKywHBJr8Keiiicix2FIKLxH1u16dTwwX0Emv+eGL2BPcQ1oWJFx6m8sil
ZXciyhSM5+7vmgywUWnT/zKQpLtcy9ySnx2XoWccRIhL/J5lXKGa6jEEhqI4yVCDkxA3Vq/WNJZV
b62APXnOqd+Oyrvfj49H/PIeW7OvdNOAmIh+6KAsqP1F1c8mapc6NebRr8pIql9RQPMEt+s86RiA
NYi3+W2SqqctKncArRy1v6QIPdqBrVZHiGJRc8iTYdzepLAr2IKJzamfMqIsMN8VzE0qGLKHqufm
3IgNROm17h2FAlOA1TThjJvVzVk5ZGrTe9gCOErixRQICaJb3YFlEVnn/BStREH098W54um8nlzt
dAsSBC9cEqJCiuyAdwB49G82Ru58xfSf3yOQ101aM7lHIWEuwjOMmdbHkzFP5UFhoI85Xf6TZ7Wq
mpBSkP6XzhxkZYeXV0KcL538Jzow9o+x6CMe6F08GYYPKW1dBpiR4b4PXJgRZuuMibHn5A7/QYwe
duRrmiwvPjso3IzFYQpVyZ/DFocVPtys/osG2STPG2x52FmMGmr905B7PkdMNACuXna6UsyOvA3h
MFcUWXPZNdmnWs7yLnLj7AYs65Kmy2HQT4iCd7EzbZ5lxnIK5AfU2RyVQ/+XEok+dvSVCDKGvDu6
qOvhdd+VjeAkYjo2k0mZYw6JXEfD9r/rLZX7rT077A+2PO+ECWAdnguSPYrZtvBKBa5vyYyFgyh0
1LjmK8GxOaxB/9XzpLpu+pDlP5f+jmDePA1cSeDawnJpEiFSj2lJsuNTp+tCWjhF4ARHnOoNPCO2
+6GkCZkS7Ro3vYPQ0YiO4Cb8PqesgUA5NEdv0UmNlNUydPba/wAbb8JZ/Mdq02ThoA9wOPoRR2YH
4W6I6dO1IoZfVn4Asu9KwTHzoshKQ0L7egSbEYpjEbfxCWa1RWZZN/poXs/cezmQ6oBEcZeulTbV
ytIWlaPKuuuQOs92q3fgcWbWY7p9XHIz5cVAufGpgyJ/R1iLdnWboprSNBYO/K/fhX8BK3NuFMEp
7VDy0J9Qgc4sFVYX67/X5nupPToxWGm3jleioJ2EhMcgz8cI4IPBIgFdHx2Cx8ZXD094+3ZWX1dQ
R5COJ4TEL7C4+AMVrh/UZbe8gOyr+gyio4CddG0B7NrsX7xsRz4GoDvTe2ShqWot3a9zqt5delCH
oH1ZRhtsx8KWl0lGTT3p4pqrxH3PVUNSGiOJ8+ALXBxD39aDmr/WzfnzhW5g8YO8dUj2FigWamzk
sivb2XZTtJU5USBT8f0VGbPalz1IYNl9rRTrl3FelXlRUUdnGm6YsKaMuRmewHwOzuGs9bFqGkoX
J8X+UGNp1YDVL7EoT/T4Hh3XTjJwwvEaUp2Bc734GUNWknTWafSAuQBnuuSqdtg+RCORluWdOpZ7
FpJF8FX+mRkqCH13ukMKfWAqfr4cN8QjsyRrZZN29xxcKrE67tLOlrJ0apoBd6hhFKylzrTmC9dJ
xr3jVT5rm6sMYy4v14oa5gtR86JF+YJKpnx6FJsf9a8ujblu0O4sCpT0dztal4MVOYQ94PRzGJHy
S2YCu20QqRHaPhFuU3x1u8YD7ceObbhAW3tSYdyj/1IRgfxm9ptnwrKQLZjFtntrJrFoLBl1WN1m
21QnlfHxNMfu3zJb/HZ0QoVAKr+6SIjD88OtAFseeg/YtLaB4cnylOwz6MF5Kb/VOMspuvpsl9Q9
3cWTTFor3tc75Qs1Gewovo/EkNGJb+3rWRMxErcImfUej5DMgIG8n6VH3x+dWZaZdPho3rHilwDN
q1LWNqI1hu2W1V0y3TwdQ6vkkkvcnhffsKrPOvMqk+8M9esiWw9OevtMlOP/NqtzzqIJn4Oi2sxE
xteS/ey68AaW5Phk5Zc5gNLfe0za/QRdBYxEG+JsqMBohzfBzt7MnHi915MN+bgBiut1hyKOYPI0
g/ykJGaxbTIkJHi5MPYbz9dMetX5008hB+5xAkFbgRCx9gYdXnt2eHGvkiBXpnMGeN56dWVdQ3Xb
9uI+tZp3d5F2ywitpDNW7lSn9Wd6A9BefPTIYjbsZ7zUwNWIZ4uhdPBgu4pk/UuSkp2259HbKpKv
SM89WGw+0d9YScCl9w3fNzufTq+JV0IWFcMD0LJfP+LEqSxYHWHerG13cpUots0VEnVbDXXG48cE
ex40g8GAXtegG+mx8GZP6pJIK7sk2MS8xHMkOfyz1UzsntIKtYNDM9v+NT6LNKWYKr+q1F7L7vdU
OdUJsr0QOsEvek4fX5BmmxugEZxUOyI5HEMfMuu+ag3dwRGwTsdDy7AuyASdJyLN5ZEjmYZL5OeK
rmPPZA4HhM4Hw98F3Qdp27DBbAErK6HUkDlArQM8uXuJ9r9Hktv22exFqxMMVnXSqiZMr/0/C+US
rSSfESyyTUhy1WQNqxqpKRs1PJ8bEcZtqgi9f6OWxYl9DZwD7JS8A0ARnibgvF2bj/pIvbupQ5Wx
PxkFrkKBMn66oIqb6ft0XTT2zx6EvEfxiAf53nE37JeBvjVWIt9hh68flHKyAiKSfMfu7jZfsu5q
edN60snFkhcg/pe2RfcVClRDACQra96Vqp5KRu5NarQzLeL7SjkYF9uPI8vSf8JRuVulWYQzLTnb
XWdgtT8WEHqD+bf5XsK4S8TbTIXUbutiu5L9+HvPQM11jyvuipQZ7KQvnwf/bGtrQ9vtOlSVECIp
u5XffR5I9oB70UyP+Cr57ZaOFMklcSP33SEM+W5QBQKTszY5QuKsubi3Z3GCqWNoXjCK28wM7ebj
iFSwmwYXXeUAxIOHxZViJqZ/4sHJCXeVdEA1f+e1Fnm1N26vDbzXyAoFwCPx903TkKlJFCEoXKoS
hQb13IOTzgcUL6eRA4HucZgqNNhdDiU2F5N0h7zSybh/A7bk0KTQ+WCJtHhsk4Q783A4LVpb1los
fyVuQ8zA49ZiJB5I0ix5URdqG706Y0mo5FpamJ2UHhMWQ8EwnlEWggMR2C+YKZBcxLUxzV1XQsye
/Ouwg5aHyi8vf7V4WQevVb40gzGMUIW4LeePuR5G/Fll0jdybLj5rXXBoagAQzjtknosLY7+PiSY
IKUAC5SCAvLBq99PcuxMF5bV25Vv3H1DHeErhqqEsUH5f1apl87OYSdJRlMI9jvke+seosCtZbcH
xUba1Pl6R7BFliAnRKvYSKlXdblxJ0SgM1iXCCguyEwdYNJ0OnD8FhQ//OxGfTG0W/t4fzOHSbKJ
zMGS32xtaw1MhotARlgRkBNxfpZwgV9jWnPzam1gD2T3lcfTZaWmwt4QvNfbLdkGqNlo9D/4A+9x
HFxP8q/Xkp6WtAIkF53uApl3pEct8KtFJZHNr0G/3rnm1K+AygGz0Iu8BT+Au31gKOdAsllbT9NG
vmxbnsvGYOlYRDKC6UxoHXxA53P37CJQkrqsO+du3bNG8SOcovTxE+MsZUmsACkPPzrxsuOrjWWX
N/0Dp6W6Md2fCw3arY4U8zCWHdm4KaUF2ku/TA/WUyXshsktfKKIKWT92KL8WotErxEJzZf4yP5W
eaLcIbM3BOJkh6NObx5VZvglIzsVvHB2GR3sJFT+vhnDaUQAtF8QgdiVcKgc2yU295UWNKw9JPdh
EnuP2jySjEqYgyMYCaid2PnI7Kr86AggNpPOFx+CIHFoPPsjOMadiE7TvCtFo/DkUASXmHHt6Ox6
swuBuK4jWa8zmJHNsoPM+mRh5gk3yi9zv+B8FCSsOAPQkucadxu1LrISd0hd9v2K0NbjP+mlq5CC
bI6dIInkFIyIuMkljubkahb/M1nTd7g8VRMu4uVPEv6+mgU/S3maMGw/MZwy5EizMXTJMxXs0pG+
HcRGZuJLpBHMGmo1x5BaUXZy9dJJW9K6izgq1X91cdXueE95kQIqC4UgWd8bbWRsuy7Ysf5bgnbo
P4msc7aijHe+iEfPQPsQChbK2PFySt2meIqksJz1gxHCh6RNXWMhv/raieMHKC9JGTK6v5eyf5Dc
em/PCyzRzzndXEOtELBLF3zBDkoMcv9/tSKRKb/zbmd4sRyWmaHcbHlPDUfmwh7SxIJsekFuyFZ3
tjsois2aMWwpl8XMeaiyP6OaeB0kvpLPXzBEHDjFVOU28OpIMS7Y+AP5AYy2jR1wQio6loyGSsnM
OsKf/tBBaU7DCdUpieQadFLNCtZw0DOwW8HDU1xAMLzUb+YU25AQgwRSZkAdHuJu1UXMioIxUAkY
01zSg1Eko9/bvVAXh/e0NcLIj+ET54OZid3GJc/qZULZnRGNUVbGqTRNZKlGpTA5LjnlHU8FWZEi
oZdq7RvTrOvKj/A+EYrpzPw5jRGlVohmc3wqlCtCRSfnvALuuLcE865fsvJxEtbNFMpvVTJm8QPp
mUIR+a3fgraA7p/W2wYU3ACQFkiO1jM5dnkEuaTebbk6yGwNvHwP2kPgB7iEpJAVMK4+hNOHAnqu
HktgTmoL4RrSQ97IjzQim76XMgMc8gfOjy2JZF6NmywCexCEBTperMpAZxirNZfCGV2qaGTDpEIT
wmWkVUGFHvAKqN7M3Vl8NSmusVnQ17JN5TA3+bgN3qjsIM7cOleSh+J/wBzTU8g+tukjfqsWf5Bv
VFl/tUeNTCBHABAJkR9w6p+f0iIIBIrlp49IwLEFLtYDxA/qJL47d+2cWc+Pob1zx6W22nXu3LO8
n7tAQQHlyFdRhyNXUwHXYDr5jmG04SuP+FummZpG4o27UF+lxDU6HvTkYRKydQqjT1YgOoteQkjR
JqIShRX6t5VwoFyNvavxjhfzvN05zbFjQhYUVUTog33oeBMAuwQZR1aP4d8tJ749m2IL92gFnJJ+
8kFxGH2CwmFkqpoXIRF5MN6tyge2qUFgABTFq2efvPf6S889Z1A23LVJ+rTCpofykmTIhd3sPMEa
2xRXIzKS5vz98G3yxQFZn1WqvPKDEjeww/FTt3NNdJmQqst79/iDoiaO0uD7T8x64Z6nyCV2leP5
mHT8UYy9sHquA03ymn+dt8PZ/+6lLBlOy8TAzXLc/OoTW69vn3fb9h8CYEtm0ldu55fDRu1ghVT3
eK/7EheMyqhyn3pkD5Qq0pTTp87e2DbS/40lf4+RJYH571Ei8/LN/pQEkaZ+pjXk3qznsEwkDDfq
bZj9xLHzmOmlESaWspIPLiDktcPdEkfCtlEV3NpGbbYtUud71Kf4xctl4Xl+cX/kIEAeCrZ6Owv1
M9GjBMCSc20kIutq6ZQ9z17wBPlzulflvTS8My4hY3ABgNSalgbPtHQXgk7nxJQPjmcQWB9GW+dF
m2X6gzxJ/Wxl6fKCwqVpIMprYhS55Hfx9NWCdgR/uQY+oq7tF9okBEZQdsUz1uXAOCu58oLPfX0a
avQaxa8Lwe22cSdTJB+NOOdpk8MQUxqztId9PkrxAX2gaNbLEPuWrntDKcPGPMSRr5S17z3zlvBB
eKXf4S8dAwDeq9PJlgttnfuSfhxcEpgO64S86usOkqFZsAtdtMcrEeeelkGmRCFEO4rcIq4N7FlB
+1sGiRISlQwb0BGj7gzC9neR3gjGH6lXL1cjGVX9JTDq+p3qzODykgiiOg7KPZopNZ4TDTOVJ4oY
4vKxlXp4ghL4gT8ZKzflFTb7gFp2pg/RW0iPKLQoIFAv3QR/EPyF3Klz+9vwlYjkTXrcYbEWqzmp
m2gMVQ27B4F17sTppKFYOvbB5QNm46RUpaF3YWM0moNXW717lwyX0o1ufj1vCnKht0sEfWO2bVN7
TNPbCzBP3RtOTNQwvXjIDdNwQT2uNqF1dptpoH9sYHin4v6omIXiIhoa2NYkagGl2a6DYha/lmEh
Hg/ThArKaLegQWLPUbnu/IWRB/SvTFUS928a+X/vxoSxqdraILMlWv1reEq9kGGQkcigysZ8ATRl
fl1BMaRcGVKYnPLBgAnLtvOsWM+CGMChRbHnachVH/KND3FGzdR5J2ui3VqVMrV9KyE5wluB5DVI
aiOyZunu85Yd3d1nnR0isdxk2s5dhTn4VkbErhI9QJmoGnlkF9Mo72iRzyk8tNKrMNJcoVCl70L/
9aGd93qio5Bxkpbkw2o6Q45Au7ALuXw47GLCPcxzMIc+VMBDtQ0Kk/2IZZU7S99D0BL+SGLP+pzF
aw/fJoEjZ1BZkgjXHCI9NyGczuySgImmt/UO25C5UkfSMF/JIFCECB7OhwCSaHhHxLLWNEeUWYHT
wQB8+TPB58p5GriWUHX5gzw66vq5rNtmqef7K4bf0VEMDEG73GZrLw7u06RE7FsJLn22eeZH1Tlz
rRyEF9YPqkhz2+Zc7jZIVZpUgm2kvQYcb6JwwKKvrgU1JI7yk0pqsxQNyrNTM/iXOzRo8vVBZtcO
fIrofKLgxnNLu564fr1K1+PEZe5tlbHZW5slQKrhpwo+xUqIYVle2HE2DZ5bpQ+L8f0Z+Z3UHROK
mvFJ2i+Bjx2tBXzN1VIMqfrt3FcFcnWKTZod+zeO3dTewhcrbtzm+b6nwQFMNB4gh9MGTRiTWJ5X
4tBYo7e6gkmpV2RV9PCfwI1SFPWbYcz1pfNb5zsTCawPt2LE4TaDln+YYDak3JgCX6CXMp5P0QnS
pcAEZo9EJI4KbufH6kx0t8JKcaq0M8HVcB5TSnU+yxXPCOsKpOJ1p3wuktlb6niBQgKmIz4sDVzu
rmJxlq/jcW/5MBBVDhFDmaeXeFlcIlVGcG9YKv2Fjez7epI/Lvik5yIDR/0Ujrpzu1PYulIs2kZ/
A6oy6BBEIOkhRa6Y0IQYo4efwv0x0GCYcBAmBmPKkCWC5QLxT23euRFmUW7FQIyrGgvAF4TJIKnw
y9enCDbq43xwRSJ90fG37HqJ68K91HspbEp1K1CGx+/XoEbmNQjkuN5tBwgWik81/T9AX4JV9oG0
fi9mKXr+cUVvJcBDBPB9FYAuALuAN/RKvdIkQgbRLzqYjcpxVJbuVL/UdjLLVOBhTsgr59M42Vec
v6OyrNgHWJhdRr8k7aSjtuRA2ZH83M9FXJ2AcVU6io55ujrjXvNq+fluDMRxkTGY8K4fFBMe3KBg
JR6ZqvbKU07EKI5Jwf3Xh7Du8w3p7woBmdziqtfQ2RhkD6Jefuk+KVibXP6QEmOTj+nm7xwrH9ow
OTfNifixJsht8mUOOi5IFqD5/AfKdwoHyFmqB5noT+Yhp7MG2pnu0LTzeayVg6bAMuj3iSlLJCCT
nd+w7UV87yJ7lfzwa+5HCwasugEFdQz+90khMJk25yqxyLvto5vsmEzr8zze+2lKhna6MveHL0iv
i1xs+AToRZ4tWvppxvYMlpjvMTXO81/KorIbvTxDYv2l90QySBJYC2xaU9gg446VlTHjx2CNMk3b
IEiV7CV2+XVDJGyylhCIkv2v1g9OVCuIkHlp92R5ikztvTHVoZnZvvR5lf3GO7Ff6wQcJOyu828e
r/atFc5zIEsmEWzEEQ2P/bMm6Sqpz7pZi6zMTYDxiFIOXQ+JGky5yr/3c0b7JH9Z6pAetZ4SlsKw
qMBUhQBAfiBp3hoY3vbW2HurZKp4ZCu9fKpgaBbwS/nmpI5LX+8R4olG1NzmMSgh+xj51tbiZGvr
s55RJgqe2EUsWqiHMRcHCzYFhQaGypJj/nKWx+89pPEhYIBClFDSUkftHju5kgq8pFDojhLOQZGb
VJ3yHhsx64GCQfC0AzacoMrmPkkFmtWrtzkQIv+Ppfwgp7ikhYqD6T84jOVJAEe1oPnVMzn6YRob
EvJDC58BphH1xChEBm6wrg+GApQeYQ2gv2A4UJg2Fi175V5cMNwbaHUtaFDnWYahWVa2uxusDNF1
CpKHpMWeNpzNMmwICUoDgMuGGheLE1wYzFOH9IOt/8012iXt9J5tOJuiWasSfF8QbkSmSp34gymv
753uqWwfcI4wWHS6pXRDygeGbIGLyTzPRNkI0KI6kRJgtXcJ0h7JkDCdF4MvDtFnQEdGvh0ZjrPL
jO1pTrk9yq9vHpFHB1ebjuQ2/pLIYH47tk0Jf4oh+6MPWqdauqbgAvWLmrclt8R5aaGTWuEZMNkf
BNmDzRY0UlmctZPkY5czsOIDALTEYqTbkpHiYj3v6xWG+MOzJJeqLTVolAwgElVG722Pmt+m/1Cw
zEh+Rin+BClqbTMf9bb0ht1dIGOhlrkKluW7WXvH4bV1Zvr0nbRByFGxBS8gEdNUiuyoZlz5wUuS
GV2+0d7bwzQpTRaj6MEve+Nz1QyHnbVys6+auFumP6DZxRt7jnBCwzt5K3is6pkeoHYB2pLdsC1S
ucK9ZawFWc+46bdIg6LfYJEefojvECgqHVJR+RHjI4TzbezZp3IUdL+staOnRwAdVnPZWq4s5ORk
vUGoaMgh4jPUXH4gaRQbjrtSl/cDzC2es5hk5u+BI/mh1khppwUL5V/+m2FMSmIHKkrj7MAhZ9Zt
Mo2IqsjRfERjE19Ade8jHjFpiKPd3bPp+zJChhhuISGCEozVvBUuawZQMWHx+xdhkcF+57NQzM+g
+XjE+c0nALuEBvnlUuxfSwOXQLiYcx9wu9sQUhxmuDaUOUWp4BQMnTbUJdbWd6Qk7KE4gs9cXLgl
9yG+xq4SwdTEDuSfUMPVa1HE1rmHE3hWbxPHKym9d8sU7A6A3+cExZ+yEWs2woYcx4K01F+zHdwi
z/y5WSB1ADciPcwdCYfT8hSCNH4Qk7hqAEErRVTyfe8TQRTs5Fn80FrgN4ywAsSvsvlKYXHpjOWp
Xhc9VgNhiUZt6qhETmrHm89P+N4UEyoZeJkKBStzep00mTdYWgSkzEWFxjI2BSlQQJKYeYqpyewo
KBm/tKIDd7jGKz5pFQsSXHyD5fFTr85X9+zMlI6BXzJ8O4aRZNL9QMyaFrW3bJj62nu7zClvWPcs
C9OzaNr8mXTi4LetIEAzPeFqG7bCAt5y7mMARcB0Lq8nOUmmbEktZtQpjKs8RjoXgqOOvUgyrLBN
TjDHLndEx0bz0KJ8esWSS1oKQTZFfTOooUAwuGCdPq4x1E0pHkB9AjyMyHUBhnFdvPbTUnkvQHtS
speVAhmOSmNrVCbBf+re/1DztEEa7H7lgZyolNz9L3bx/vtmVA8F6Vj7i9S7G/FbMaYUfsgE82dB
Fu8UR5aFyF+NUt8vlnQYe5h9YPgIeFc4vFl4IZxOb5put40bEM0qy7/0lo/6xOrbzR+6FvGHTxFo
9uADbbaJ89/ILRzQqOwbROsuNHWFXbURp3GZ2edNI7B2UTuH+F094FjUbtBFTI3Lnh3kJMZei27c
QcZEOi72YAtCj3CIRDv5FG+aiYo7d/31sc/T9ZeEt/jccsJQiznTwk2esBF9BzwS3pXfnpK+eVP+
7piLEJ2j45lHYFoYH0dZvtprtiC+CSz+JPpLeEEf5yhtkgLQ3E68kNg4dIt4M3GZq6h99LqEXzAF
uIsc0WrkfjFkpoDZq7L66stRdtHwNgBXYPTBQb7kA0c0Cwvpx0evZLxFwT6lPTr5y0LApJa9CYgW
nbveqmcQlRalVHCjiuzf/uEJzeA+EghLSbqA8hv9OqSE0BjDUhcJvTmQYVHSLaQ+BaONwL9ZuFrc
tqHXcOgQt54yY/VzTaAtM2r/OIkaqW4y4YiQQBWBhTCLtp8CZfX6S4cuHCZDM6D0RPluSfdTOk97
7jGMZ2rv+IvOi85m4lqIDcX/ai5Rhj5e2iZRoWFpPYKW39dbUiLRvH034WeiCZUyQQdZdHBBmGl7
bBBb52ACNChWIvbw9s1hiFZVMjXTv2Uulo+y/hASAiZ2P+waMR0Y44/S0myzjZ47fGh6ZDuLvAVu
z3wPoMzj0uOVgVIHywwFPIJBEXtkhcFllf19vgrgALrHHVRVZzc6m4LI5P3TgzrtnWIX5j00PIEX
BZzg44f9KkFMqt5F1XOBspUcClVKG1xxHsh1NWAo4WIAM+r1vWpP76uYNybfaEOZtg+RwAilKr6B
ydJVgpwxx9UfTy1J4cSsXIxrqoS/kgrCCv6khVhY1a3A1hrkqq0fHGP21wSnmHX6KLn4p/Fs3QcW
5n5oJgwSU2sbKvU5LScReF4jRHEcvMhUxCTZHPAy+eGe0Xd4ivp49Cz7SQdZO6LLY6tbPSedTzvO
K50n+T+waroUEz07+pko0rENI/RyNziwPVhG1WojNZdDcTIpvbxcZ+hCI096ARUMd7nHS+4IBsQJ
WDWmKzO+O5GHEb23j96RiDpdWLZNaN0uSxU4cIrTTrHIgsusjQe9p85JQSjla9T3qT6pTYJS5/dT
ZjTZhWZHRokgVDL04htjJ66a7D39c35P6RsblmIVEum1/+6LfwyRQrg0dzVtH1j9b0JbQjjjw1Ct
EVmCXlvG+F6lChufz2XANggYEtCYD18mWxbWLF54UtyJX4mG1b96LLg4rDaFQFNEGMcM0S0caetK
LVyLDrGz4J4YMLooNrIs0mnER7idjv6VrwhRxb/AlsONWEP/nEnMve/Mx2vhtqPcyUmUBzV4lTEV
83QSoZuQ+E+aQroi3Ejw68AeWd0A19gR94h4UZYBiMr6tgOG8cauafTzCrZUHLuZ7bBaXbgSiEzt
jHk1eIg/Z7wEROdCqTbXgaeHEoUqCL4DPuCJewnoDmjrJythHHmYN7u33+OXim+JuC5y0BvKGXI5
9754ueswPJsijwFKkwi163a6sIlxsHb+ARnZWpfIAmSKbhZuAAyEoOxd2szmprhRTLXU8zOSb0fn
x8o6+m6weopC3LivThJgop8ORr81rsvM0et7+o4o/0ZrQzoUG4W0bv1EEZnogbAdlpCPoLSVobZg
1+x/2di9Vf5FQi6v2K+RDvVyrgaN7rOtokyfB3kDvn3CnWscWlbL8TKfkX4WhjoBXAnxz1zLQ33K
n3S2fJ8x3h/Hne2t89wcs2SUALJBcl1wKrVgL34kQblNWaXLdVlz0Wq6EC3N6YF04TK9YuPfEP97
ApfJoxzUlMGy+q8iREFoYH5AtKsYsGXSBdTxIalUj3gd4meElNApEYffwrpg8BkNYEdAaCkYcXYj
YNkYwbceGBojKJyCH0LUqdkEilf1eal5qInAaMQ9g5hjS1LpybTIkqvj6GlF2Sbv/CsVX52bcrsg
R8vKKpFgEvWtlioHWkFrgbS8vpYugzZVumH2dDB/ow2Dj1h16JvHpkCsdEwCEM9J+CIE2delvm63
fq9qzlcl+Brb9OKto6rNcHa/13MclqoERiRVnRqO4KWkvEwPbLmWLvjAli1gS/pdVgjNAHhFweCY
p5q5Rv40UGofLbwKsXG8ePr+mIuT4sef1d2cwvqIM3XHUe8xskH+uZUGqHzEp28ayB8mRbo5T7GJ
fntuk16/ld+68fsGtXRNHNrLKEP3Py0M9lIQh7tdkIw+dff8YCSVvPVzjwfuTPUKLVc0CPvB6uKg
c6riEORS6YJpQ68mypmL+meGaigYws5dJZadVRDwQcu4V7tWoAvq8CKvV13zriiqEFeopO2ay25L
Kms5ZfbTOhR98KBbc90l0knu/ynJGz17qgQ3fYpIv8rqPVZcqy2jaAamS5YCHaf474KDpQ0mm694
X51ioxW2ddYcHYNXC+7m7a6+q2WFLXsP89E8nIPItnjBdSclupyPyrYiyKnuEflTPyfdI7yOa2hV
BKMq43D758RTiInJjk/Uo6WJzC8SLTgC55FgJKjJSkUdppedRcwEWvCwFRmJH13Ro8Da/owShUNW
3TfYECvOb1WNAyPkvSTD7i5eHHOwfYk9gbHqGRSFU+z4yGkjZU2RL2ENyab5ptJTYFQKzUQJ5auM
FQ0/JuyLYhjQbs0y0Xoa9r4ZdjEkS4Sj/SeS1EG5VAHiH+2W/MU2EqJcMUX17HmEUh6XKp33dxUc
JfjziS1P4kNbi2Hjjp7a8Drf+B8juj1pv2QpoLUeuWc4UxeUMj59xZwW8HzegSEfATQpCn1S1v0a
MMosPVUzvRbLyhqwKKfjc3MlkJDmT/NqUfjPBMgbkF/vdpMIybEcYdGqE6KTrX96uR2jpSDya+Os
L0c2DjxIXu0MHwErHhO43ziWkfJYE+lvo9bB6ny2cHkOfGcF1M6XHquMeMpyt8i/qthiwIagGCK/
DgkyVaZmKmShy0YIKf9bGxs/1cS4hadoxB5z2t9tV82NFRdnxl4dK+XPyIQqHF4seuhDusHHeLs4
uxtq1XRSr7yZHKxXAYYvmApFZ6u2z8gfqIO/3eZoS6ehabtuc19hBYla6lTSz+dKOnlQFsajxEqN
cgdCdSwJrTzOcB2999tnvWiMYAJ+306ethmbMqWRfyjn6k5+8TQ+iepDI7/gKa3txTn2WyPCq7rr
Ar/kn0i7COK3NLPVy3P7e6Ryq25JJcl41gQD4wiUXBXJIPCK81TFwC9TvEzFXQdhQUHuali5i0aV
AZKpPpRZQXHq/P4Ok3zlJLHGXVZN08SPjqrx8LooF2BE0M9aDlOEjYJMoLmPfzHbPVktrvA6HbMh
q6skqCSAk4sb8pGrvz6DLCsUBonJlgk5oE8MEHrluypXlOkcQx3B3by2KXfwxHsgtYurWF3E8B1n
fJMQrNxx6sOvGLBT9btLSyJLTfOaJbcGXYqPNtgkX7Nz7fJo1jGctmNjmM0BcpetbQaW4K/K0ruk
Led9sE9naDwSmfbBIg4Gy72WP0tgOHtTKQnX2IvInXAAlBK1FHarOWUudtwHo46o8YmkEO62b5/S
WhqUugPY5WhErWmLrKaU3ppFOmLE/o48OF72hTYsSesciAqY1SKHV1v+R2TDxtzz7bakUqGR14bY
8dOI61rh7fLbMREsWb66A3mmZV7GRYvtpYB9qLMUg9dtq4Pz+O4evDUKOatZFLGlg5WKWDwNgcLf
69CsNaGr/Or/0TdUnralescqmGmADRzcY4Vl+hRNjFikp0i+k0oGl60tD3ZGSJVALRQDLV5awlpN
40TUHu+hwyva/Crm7ZXvNmuMDSAWaWfG6A3bHbS1q2Lcuz2cN1065UgfkbztdwQOS8+rJx88qxMG
Uu9lJJbQWaxp85G5jC6CwUH5syXbPXMZ3+qtTe8QhcKjaEQGv8JKA6RqpYNgD8YOYjJ4r77oK2fO
Bd7jLtOZIOzA+gDwJ6GsAA+DC+2DiHFN8jWFlVKROgLUIcNL/EGo9sOASrLjDnt1+8rb57NZxsuY
d1T8bEvr5hbq5rMq2aOvguGhDbvddNYAQVgKmPPLG9KiFHrQ/eGTF2AgPSby4bfrIZT++7sg54mK
cPE+Ylip1iaWXHEtmIVjhX6dP4hNIrHgvIhvHFLbnKhAAR0CQe+mO4S6fNIzmbLT1UAHZGyAbMEs
h8dwbZylOJipimi0m44Bh7XHxFt7+OFofRDewbwFja6ZlZkZmAwfnnH4jksCRvDeDXLisS7L7Yp+
6aEBcw270fN+n1EiDf46EM0dfZlQA3j9gqGL/Ry9XquQrP9Y9NE8lpS8oQpahFVXLiC3+NPr7FoD
WfSoEZ0d7D1cL0xJ/BMV+pQe95o59TZpHbmw+FQRATPeIHJxjXRgVb3Qy3FjNYhoNkJi+C8/eGIJ
nAHczggELezKdUGkr9n1bCVVdhuV1xJquuErNdCbdIwQ7J6ozf2WT7hWPqUpsIQZ1Ng2S4svEMvt
qRCJoAClLDmYCj153Q0z/Ng5i0NJlYFcJMlYtC37EYkUnluBwdLbMKCk6fly4/oHdRjM17LNp/35
f6ZEtHGaCkxDVd0/2PBnWF3SeKQfyLP9o2dlOja0Ml0qPi7PW8P6OHVTwp3PLh8AXddMZ/11n+az
XQubESsmdq7lvY2Upq/jrFmiWkaxe3WJaolHPCf26H0S0y3eKKbuIpFYeyx2I9vUJA94rqpL30OE
imUng5bWGtKlrztd8jPY3B5twM6yH5JyPbOVJ79bueCusctxxdBjBevoAEn1kIU9G/EobTVAnVCy
I0KOG8dSjh00lkszyVde4hVP0UvZqWb55gBYuHAbLvJmyWRnemzSGI5Y1Ll0ROpynpqf8/Y12fzs
mPIByT54W+Mfz0F9Pb/Ub5WEXK7HD1wjYHYw4u8geMdQDKyaAAAZVwgoc2BdPlnon8l/kaIYUMHl
jTWUTv5XnnHHc4Bucq4flUusqcmrbBhK8q2sARG0WcsgiKd7X42zpALCf9I5VqpvpYG7e+kQy9aI
u9uQuFD/f+hEH5mnvMUYhbxP7v8XQp6nNAKpaXsf/N+Y4vhex2Vl7Il3+vCziHeYETYM4goXUzJ3
MX9X58p908mGwxU9vvoSftJOk2uK3ggWEHRE1CTEFY75/15j6Xiukx7v50dvpwUWzGF4ACxjjleH
AoKwAr0QSNcNzeWosCSLMGpWY4lkHJQW7QJtiWBDATuqaurtcDw+chDUdLeiDs8BDsijQRhZvdhK
XHPsyl7Sr4WN/J7Bo1IWzCmhu3Kp1+O1JBrJYetZxI9lCBBPEkxyN5f/yGZmFcMsKegGW5gaJudg
SaDGef3lVrINcrJCMKad4dwi93bFaVFoXZxdHhezIYiuyoA3OUP1OcGu2qm54/agO7CKF8f2higt
WFJ2jyyZYUDIg+Zgm2GbaSK3yuHtkp1F19LsE1LM++n15fuYzvCNRQCM69WJQR0LmJ47lLvmx3bY
auq9PlYkdpRU2kH6pd7W4zfQzrOp/eVhnFw4yMso+vodXn3XRc0s1/RgWmUza9TeZRBmhsklLSIL
/YqRWYb6ssW2EEsxhVzVbpEKYXT2eloH5UJW/2srB1HQmxlTOvDwnT9IrkubtNEb5uLl6fx1xpaf
B1xDm1XwHl5w8MopHl/0EVhaodEoPeyVX3uFnYkGpKJUu6ZhvIND2KgJjhHWLeFZ82zSZDXzmoTI
N4L3RktDK8On8mKvqRJFTcXrzS5dkjUD3nTdJqft0OWhqKaPya32jYQxKRr2kGsJ3HnaEic1juP1
CswKBDAMVWzQsadD+6sngc+OXPpBzPPLZhYze8lcRFM/Yk/dQt26xpARTDn7JhQJ1tV2thwfhy5R
ndOr0JvQmrByC3Q3OcYda36E+NCCQeED13MeyNC2BQ0IHN+8ngMT/+KOyeEObzy4Ymgva0o/nEbq
IkscVqlPiNeTFX7VsC75D5z3Ph3yIDbcloqAVy/IIoAW3oWf39srOQX5r2AzBfBep/Yi5pS9rnFi
nLvOlDthRTFP2wY1NXbsdnlzBXoBIF0gzwf6v9fGNIfsWWMvbPR89fHXFQPROMKWn5Q6ewZBT0s6
KrC5AjVDn3HRwTvhhVbC78haWadJrS1CQyN+Q2kPffgiTjG0iGlAnjlkgkVDEFzsjU98mkzxTJi3
ipPlnryt1vv62qnt3/mwCsla9vASB5vOmh+1EFebmlSVOf+J3U8ilFCKYYwHVX2zDbYK1SZmN1g7
Z4fPcVQ/iS3qwtatWsqbwBhDp2ZrQhP025P66SK6BpVPexqZ1XYMlb4GQ7WYBx02iDL/+WgBCc/j
7udOmRzkiloPgRX1Xb1pFwjbMO7G1yztaOMt0ucd6RUBfU6ZAR6bvpgqUefbAYmbr+qxBJjsfW2m
Qe08/U4sHa/WzLuRIclEs9ELhhiWPWQyOcn+4obC/bejhwFcDj7YTciEtcRAq0LZaPddYZWZJuWH
1Mc2tPZJYBthOfMA+ypdXn+mZjuj4+W/kdsWJ08RMFjrOE1j2Wh9V0e+gcAepyXsrun+IC/Kr+aB
8+hE2bdSLhx+jpT5tcwFcsGdUMFAqP1B9tgORpVmwcTxa/7/Co0ggg2Ew+L0m2MqZ5sWIZ4uiwrp
G+phxkeXQhuQWpYeyZOgYfoHgTc/gS3PwQ/K7YGiIDjZE+eqr6XvRxbTtdWfGz89h1H2go6nwnmW
/rZxYahdGURduq+7VWXUtYJ2tggUELUOq3G4VNB+TLPDPNrNMIuzOiqH1J5YeozRdglIpe4cdAbR
Hdupdi+Q0gHBKEPSUHN50nk0pG6JsnS2awfEO+lHIoqBr/K9A5Q9ouJDWhLWzlow8lLSaGRR4nfr
99JdvV1fvTB01i6EoA3a8R/4UMbo2dF3xaFf6wW6UIuAV3i59knkcHNLdeAi2n3mi6+ZOxZcQo5E
yZ6FxIt31LK/Mh7HoJxhDhJNGAThXhFm9k8kjO8N4vvmDo/H5VozrhIG+qIZ8u89xxf1KoneA9WK
eypX3iduxXbKvvxkdIZmxNq045WZHLqjzRdhA9iL7ixvGF6/rTKQbCZRBgTfcQwxpZPD9oTARtjR
Vka4M0dB3Plk0oe3SwWM+c1Egl/LRhv0E7/Ti/QidOhKbWbQRO9bU0WSy8veQvKm7q1llDBB69nK
nZjN+CPlmGXEdWHBoKMNKmbURPSh3vjRdq2RysfRJCUZIiayj4rSdhYBaUYnJeDAvm/EFZsLzsxg
3PUHwH907K+obJZoQajCLQc7hHLMEa8R6JEs0vejOtTyPgNJUMHP10oQjuG/8j7m5mM49h3g/djI
6u75h5bPO4ruvxGJD9ZCWrGH5lF8z4v7kEJUd/qF0V4PvUQl+EP8WCfHPEF7joxfFHhQh1YoZUd/
ajIx0E2VkGqOyJ7mC3HHFW4wG65g2AfVH4Wu3lwnbMi0j+bapC3WhwlvdnOIuStV5oQphrzZFWo+
VfU0+bRUnFZYG0bDa4NgPODjmbbVXVZDjz37W3Zu8z/XWJgN1NtMoiQpnfekvIUBsvps0tG7gG/z
AfnjbkJxFkysNaw4v7pvoE4mVL2lk3J0pAfh1ZDSZRYtcOuCc4xxUeJR1gQBhCLnk84vhl07aMeH
ZekKyqnk/QmszEBRsK5U+1oOSIcb9T45wdAm5Tv7NMk3WbnNDEnHEtPwaoGFqPAS/jqazPuvqjRm
vVEAnjZ4M38mVi+v3iaPb87Kn42p0A9riQAfP9ocET99fZKDUMhQi1XqsBAlW9RPvd/XTLplUdTk
pj/a9Hfn05ckAOuKvU15xTrak97GzMjtDX39QQZjKSwFnmfPTHowROCEIVJxL7ixcuVqlvfHZooI
/kUOeDh73J56zC6Q2ciUHcRLOuPi5JfFO6RG1PUMGdrhj+iZ298JXdBjvyhYndabRtsb3IruEHiX
H/1lP+bTAsWj0wz2w1D9XPFix9hj/w3ptfntdmLRDQ1q1Oit83P3znCmbuoZWOWdEg+rWW0kmUJ1
OZCVqmqCjT+Kbt4b4Sjnkk5N6aGqZt9+5BR4gN/fFoykzIn1fWktYh+WzJTMvKirTqOdBydl8MYf
d8EY+x8pWoJgHMS8GLVEalpX3JmhntepVyQoupExl00Umz9KEmKIaXp8PlJpb9S6hD4h9bYd6H+u
GGR38lk+eKtOhRSMwUt9EqUmggkinf5D+c8lwFM8n6gKTLjWJlCMketeyga7QFlmymwau35940q9
p5afjtQn0kRupN92JG3f8XDAB9W1CZBVuBFuEVAYldfe8u1BYs6tmUFw4DLR5LWIvs/5Ko058c9K
t8lIUtUsZ7PqLhbL5h91+oZPZE63ve7RqgwmKJZT0bBn+X1PYX+WmA59Duc1xgIzYn/txaBoyQgk
FqYG/Yr8edsD4e1g/8DdliF2oifV+2ep3+J/92B2xTQ55FE19N63QdycGAFZT+KwWw64Yp5aGYGE
oV2kv8b4KylgOJn4KFKgOaLr5UW4P0SnfxgEHcuvdru3LQtm/Wvu4yECh0aZGTQfqGhoSaydDzOl
i82jyvBvzNS3YXH0sdqXOXVoUyzzxkwXEDOSnn4S5J8q1rikNyTG6Wa3MiDI3p97yqxmeYlPoOdw
Z03dITyVWXlwzacH1ile8Tu8vSH+Dhu6pWn/lb/dcn5GT1Tmbalr0T09y8EB5WA3cIfnr3yNb6rW
OxhKaSbr9VzjP+yGVCI4zmOggbh6518uDQ6PiVuLFFBRPniA0LCTxAoGYPd3x0a+wcMjkGxavzYf
jU+vRg08AUOA6boHADQ9Cqh84elWm2+YcEnIcRT27UQTaUdJ8of2MSUS3O9YXdsuHHNwJPMcFmyE
cmlpJpnWVa39of8Yve+UfG/L/xpX5LWOqJ2dFpbFSgXbUdnEwZXwbrqjs0Mf1nqhK3SnZx7JY1BD
yvA1xcUbDUSS/YokqAv3pwoe161MEkourlqdeeQLEPVKLGxgRDQ40hWJkqhe75dTh69cpGBjo1Kh
wh1rd+/qqHDds/EDjYZ/GPepHlV7MZiPaiw6zJ9tgWMDbW8n+Uj0VyezmG/MxjzltKyt1ZoRNVEC
S/1Lr3CSvUmfub7Z0kehqGr7Jc9g3180RFu+5k3l4ik6JA66mZgQ2NkwjzRaZuujS+1KqIRYsyYY
uQ4JtBIaEodvBzMzZiI0bh4GdEA2xFitap72PiM7tvErkctEjeOTeq+G/Fx0k5ShYtzjxMnZkeEE
7xkRrgtoEPbfBoRv+IkfUq+M0VMGHqIzYrk/aqRDOOpEQEYx++64kX4ZcvZiyllX0HcIJlYFNCm7
JLf3RzexPnMSbByXvWs4R5gqB2VBY22C49izWBfh9VShsBX+0TKlCmXqkikWNRz+CmYKmy7HBWv7
j6pv4MbjbI0XKiVLb9rtrqxzI3xp+q5G2Yt/Czz66/9CZIqktw9d8h9i2NmwEXqEvzDLis8vD8zy
fk0GE//sFHPTTqM6uJEbA7oHLxUQTBuyw3cQUuJVT+/fZcUv0jBSoFbn21D+5M+3aZCgXyvX94cf
eofS3zQsVXXeeCldHgV7Br8KU2g22OUYCJoP/SYI0dO0jln7JmPNYoY5mkxAUobPiYiEld1MewZt
qyiyUJc9x+f51s2zfqw3f6W0h9jaJ+/74XI8PGaMClEpltwD23C1ZMrbyh0Y44de1MomnajOcTod
ZJoRYRqzxxDnA6/QD03WsOzFZetvq9MVKiqa5EUcCj5WBtXbiEJ1GCNYx90NF8OvByZ/zOUIqVJJ
K7Wq9HhlgKXU+KXGMV7OjrxdO16aItwqvgdJTFvfDz45F3SG+Ai18eHC+4EHp4xrEsUyKAeL53ek
Q0XKuA7xNa/yb1zWk8tjJ+MKfWxqexE8AwSIzhxOLwJVhhukTvXenvLqZtYD0HvZiFEQDmX3tSIE
DqjoX7cZe1UQ1QU/pU1yJaCaN4UBmOIdpLtUSE4a1apn5gUFNvzzdLy+uzyPny/1ClOmyzd0PRc7
3ZZ2srx1qMmh8BpOXV2b+4mbuekvjT/UIATFMYFDNAJmtp5FL48W1oh/K/TpaecIpiDP64yiDTln
+BguHC5Z6P8HLhlZDTohjFy7OUV4fmqW1xDZ9w1C9tYWSI/EmZ4qh6j/dBCltiAy5Syjh4S1nyhN
QqlHizSY2gEWlLQ93G2JLczFjumZztmzEfMpjgJ8KHiCaelAx3VYMVbc3Sqy/TUASfCryzwypiua
CEhLQVpq6snOjrGEtz1wDzf3aGmcjpXGG5CouqFAeAt+VUr8iMMJ+TbATYwo0nffUQXwoFxp24hA
3L2JMTKrhHZKJid7R7dELKrMvh4lA+SVcKOHEK0MsdCy11Iy+wzPjwCHhbgcsbaAea4KA4lwcdLf
niKuL4ldBtKIJdWlOmcGUy11OEs8K5Hkbf2QRjDKPmaocANKvfQGTLgE1jCreIC/iehfUSvs6ag3
ZCjHRJ6Kz27wHuI3LbVnakoRtcEdS3vWZtbFq7q4iBBxC7QmoSm1ekWLe6q6rv9baoWyM3QvPcJ8
y4ngIK9/PP6bWh7Zi/qHUSvCJScoq3T1I4HWkbO+W+iPYYWr7I1+vOD/6/jHcOU4I5j7MPIh65Kt
lC1zJhaFGpw2ljrf3duzo50B0umT5pFDcaXRlg3lXvN3tJxRUU7YkDYoR8QFH3bv1eRR564Ls8l4
Yo9cpWe3zYZVLTCYdfv9TMny8XSCj1SS4/BSt+YzK+nlj/G+9yUS13R9bimm5SRaHVoPmfy1n7jv
1ShkoP1E7+vMHUQ2GkQ+tSo9SikJlBQeQzeyzKywG5HH8/gsdE/IxV6QrwRBDnSIIz7slT6lQMHG
2FK8vzgzKt6xYL2POrYhVGu5qD+NkWdo+qpAwmZ77im1OkGUHr+mJ0GdTkz0Q9QfOeqSVpHlfYzC
/LH1BNT7i7VCkEtUmY9quR9krVvgh8Jo0IIxFVeE1Sa7IlcYidaIr+CprGV0vB87TD1meO4chudN
VDnOmIz/YT9sR+SEfO7LZe8wggfPpY9j/214I2N6s1ApfsYpwcCrGMcwqoc2DMqMd4y6lKbFptf3
jrrGkzt7vgtLniIOYlbCur+cvAsaKcnpPi4NQiZGHjjuLzlQ3VblkWiP5rZzbbwpGIT0AFEyxTWz
kmc2WLlZNKVKHwuV7SXxv+nASVvwktrYh7jqsSrDv8I+uU9Vfzqfu8J9Z8dIfn5EnUni5NcKLO0q
SNKefw/dG6DcUhc2bWcadyZ43AHcw8Yx9qTUOaHsyG7K0ngn+yx1POWESYM0UIyFTjju1ujJG1mx
NPsikCjpMcNisOuNmzKkrD8GChZh8Cg6JNdlmSMOImxIk3rovXoQnTuj3OqtYtPa8AZjlYZH/AA2
i7eOJjsJ0Wyt3WOW9CPAIH0CP43t6pTC5CvNxaRamGVi15G8OeLa5zw2tULE72vWoPJAz/ArVceP
iB/D2BAepXVJRp2zOcv8xuq1stsoYX5sYoAu4JkM3inSLWy5KQIii8c142+rCOFV8UX1LKb0jffq
PhF5MsXRcHSgs1FIlpFEALRjaV94DjvD8Xr6qx+aBa3BWIy8xfRRSwpEfy/W6v1azAKtVGYVoI9c
catJ4R8goZVZoLqS9M0+0lFwYeT2Pdt3rchMAc5XsaMK9EW6QlSck2zzCrJmzcYJNyoiM5KSnnft
5cGWJQSaoaN5q/IAKPlo13oc4qMYaPPpfxMExGXgTw6cZ9BNI+P/pgFPnGNtwNJSwi2nIHbPoygP
IoE53hwC1U0/sHIqijWIg8J7dMMqFNmO5GFbmFzGRjdmyVpc2xFtYLDrILcpOJVJZ0Lek66BIGHM
E6jELdAglygDYx7hJvgd0bUo36pCaxWLg9y7IjW39JgnRNjTzYkQWCef3wbwqj4qoyg4SeEUf8yN
Muw5VbawdTKvqriEWHzutMR/QBkU4iZdd+CBcP5UkkG32It32T/hz+y6mFk6EOrnUsOOxNGVwQVl
uiZDDh8WJSCi/B402bcD/12IJqfOWI8JEdpWTTIJ8HWvkrYCX1ltgvRMoI0FDfTwLV4AzRkOwDH2
5AnSKDcn8yI2TIlIlhzDAy2LLSuu4iuCRx63JJXnfUF9Yh1cRkxR6+XjKzk+0yg5rvd3ILpFh31W
cbzTEZqRs6IIg/mh6jLmaVhjEyGbndZrmz3XHD6TXBez5aq637VRMtDzJBexJmys0/pVyIvrGlXi
15eHMk4q4hoHxvCEGVBAOyPJIXtBrT/2kX+VYuKUzrhonBoGqZ4kSBzyLptkTfK3x/dSKvgTeN94
25/2oIFeRJqTBVJAn61Z4qXSik91FywcvoMDcJd6oqmL8M+Crk7LfvAqp7ad9RCI7GT/NOno2IJ4
uchHbk5H4UtvlmoN1Km2Gbu9zYgJoJ8m8/6MkDueDfN+cJmfJg9IDcdaFq3FCXEQOpF4AVEQtmAW
h3hHbNW1lppW0wT0lcLtkj75PGRUWv8MkN6ytXGx8YtoND0MkJJ6XVV35io25+9OHViOdRuNHgtG
5/AI8bgU24DtqoTDkX6IDHyBzICyyVsZQ/og38drB6WRPgXL3KtZ3WObUcpRK2Xa2jPP02v4HDuw
ZwKviuy9354eRo4D6cwNIMQSpn7JBlX3Xs/021PdCB9mYyz5Q3dvGD904EfVFX0vmrEyI5BT0p1P
yyitrtjOKc9CXxv8dtKEByqnuc9qpxm8hpBUafYWflAIqzPp1htpyHawN5KKrPxUqU/HjBGLNoXT
KzCfl9VdORq4kuq+t+ElybZxIJ5mh8673+J419qZ3Mh1iN4dwXOSvZsBWHf1hCklnJiF1lqFlt0s
s3rGTVo0QvcEiRUdRJIAjrd8aFIcU+Oc/wRBfUvKf3znVFiUUIT2NiucfPzKe7plg2UukMUsng5a
3R+bzUdf+jC3Eqmx4MdUd2nmnNkJs4+aRTMNYmwHAWMLAwhG8eudPkH5wl9+OwTXiBQjL1yeTd6S
9WBe25wIhbYIpgHcykCXT5rgLCNRs9aD9GCCjsElIlw6tDWab8tpQueqoxppCHYSZWGp7QS9VeNS
oK7qyRLIiOzVH9Lf23tHgNXrpI9DLoMmXDF1q51E1xtFaGZo2qYf7oPg6Jzyv1TKtyYQjC8k7S+Y
XtbaAjrlJZ3G+NEqxrKJQ9a3q0f2zq0iZq4J5VTMNSD3OvYq7BTgLuhtsIE6s9U5+jOlL4h0XPXp
8o9FG3rXtL7Xa0Q5HD3OoOqhLf+U6iCdMgDYwTky3SAXNGJnmajU9KsDDu0ejLHOPqkwGytr7l10
eEj8scU/0CVfBqOx45KF/du7M/e4HJDQbXz+Qrv2t31V7TTp9QWKe2ZrrkW//1A7Gha3kY70i3kV
z6JBCvepP92FiuPDtAoHPrbj+9bo/BhLkRjQLWP0Cadbc/5T6sYPS7DKC8Hch2HNO0Ln23y9w+Uw
O93UGnL+mrg7e5zHwewyaQDN1GHIgxurpBNcTtwjPDP0DVcKSmPcegz1NSPg+LUGYul/OFu0t/9H
hCep66hoZDUGIdCCTJcBUWu2QyGr33fBxqVz6RSj40OYyvqCI8/aldOGEjw8lqfVfm+yb1QDLJe+
nLwG8CIhtSzeiNz6ifGOiDBDY9bNbjRW+arEyqdCbKKYnbaoCGPq3w3aJRkUGZ4cK1JvrOasQcFa
y6KRJu2cpxCh3/ZuC1CaYxTkmJfjydRomTwusLRInorUY2wUl9mqPFqfb3BcWRVSyWZD2BK+yDk+
4wYivDUfkKWXUzUD3NCHqArULKHmzyt3nK+LV2Zs3Rm8Cht+rXuCpgrwjZ9JHFyhxISIJR7EWywb
Zl3aiJtw1BRG/B0HAC8UWAViTp7NMa+y30COx5lG56Ky/nzk5ju/k2N/ZlWGtlK7BTyiQbvw1fJs
2v/vdSTRzs6nOcWOhQa4QozXIAOSe7CRy+JKIMN1XZBsNmwGuxoKcfVX3/e7Z1xskeesLyv8bsuZ
G2H5gDVGfjgCXGs2fay5AedNmlW5fQgz1OAtfp+u7bxN/nwAX//BhXxlzlZYKPRI8V5AFF1KUXoR
+bvfDGNZAoqg6E22K0p/TW02ozz24Wu73O+dsWQB0IxLaL/Iv3MrZMWoGdxHrgiQ1ZcBVPIv3Mza
9hEgVQNMy8DREsoqQed1UwIEwPGoq4tj2pSLSiEtdEE5wDKG3LN8V0TM2qfqJcVcGgP6RYymWKsi
I/41q40i3RTNOXrGkNZ0gUvKVMbyx+96hIPhZLDTJC/NO4GqyShvdzfeuFN91lN/iHBl4E1N6sBn
f8wKndrLIdJ0q20Kb4HDpwNIaUso4R9Y8/pFdrevvMarRHqO6NybZHSgW3aTPveNboc9WAC/tZ3r
gzTLlt1IY+OvgaDpXSjddURqxPS62xiQqaAszs+SCTlCPAEuDoIZzXTOKvqiDBAPtsPh1UIjwH2J
zhZGcT5IesxJ/UAqjzT+Pj40HujYIWL5QFzz3UKe2L7d3n23u5maL5A3wAK1yTEyzy1xEIDEDKpw
aOjoMhQR2kv0/ysTIoalLQpGwFEGip4H+9EoUK/L+K14shznVowiIE6vnL3cp5105BS41cHSvw02
Zn9Pdh8y24/0FRF+nO6CoREIgXitonBVmSuCjuUrUNKG10zi3/YdIBW1OuyC8o58mZDHmz9pF1U8
+AjelApuPVT1fl/eJh2DPqMpwwShPaYVOOBa5pNBGtO3Qnebesx0kTn2MyabDr6+PZ9+Whzj354D
hO0W7yUV/qE5aoUA5s2KAOGu9A2DiRkPPAbDA6n42EEyRT/Xg5fOjtUAXVcluoaVblrfqiEZZ6gF
SMQ5CKhZ/87mdn1BE7POZgHyGb0KI4T5/h5VE4lyE6NMbQNHRhGVrst7wfmEKEPqk7wPyydlvvo+
/+oz4MJri4fwx/CA3+amK7cIUhhSayG0p95k2qYGbgLzHhaSBiITLyXxWlyfNpFVE58JT3pz0tAl
HNm5A/9bMwM5RX+yL2ug3wHaZDx1knzbRy34aSqvQRQfITySBlDkDV9bYPVIGmM+tQsxq+0oVcKf
+457K8qXSDa02/m1OlWQ8rQOH0/m+MUh6/D+0VVB7/0sdyRVoVJa/V5YaH1Ws7tlLzhCzxFcUU3B
vo2chMqGXLzB9W+HaPs9vpUTXmuIujmW3nbvGzM09xt8wl+8UU9JGtdK7fNlNTX9ROTSt6n2i35z
8L9B3hBECPtJX4Z4I8b3H1nYrmb4h39tsOOVIAaGgaRVKoL0D5wXlkv/v4gBtEGeYgdcz3knjKXw
8VU84kT1s7jTjVsHvUUykm0+7JeIiaeO3fDqGHz+7l3tVshj0NsiiZLEGpe4XCAjWjza3+F6LH1W
l4edV4Gz5eH/rIMkVc/Oij9zqpFLfWsfEI6b7g9mf4BwThNLVPXIL4zPP8tBiGrS1uXNBVVnnEpE
olkM5jsYbiGjgUvT11TpHAWGs9RnNPfWRRcdMjGIT/G1CVtM8bzO4cOraP7RBR4Go/25Sptmx8zz
VSIr8xyr9TXlPLi5dhLGhSEYySYnLSSyPfzJ6ro0UM+8B7MVJFzRPxTCVvNf9qFpEtMuu2HIvVEG
JO9sgttFQpLavjDyYWQ9L6cXyDuHA5gYk3T1Xt+Xhq2vta2J/n9yo0/7AV8LD944qLPDcL5DAmj+
hBK/YwFZ79yUmEI6Op+EiluGKlOJP8VTv97/YyXl6T1h7UUjIDT1ImfwinRJLIMF79waId7/5wXG
1LKGxBPQ/DA6bqhKIWCzC1V71XDNqbymuaWh365OuYjjFYzS5XIlGJ+nOUUbqOtWLFLRgKHRubmH
4MuBflbZUSEkBj1Xh1y4QBvB3O9TgBtxHwVvW7eL6fVgN0wtVljAFExBGWucFyq2Sr6sZAEY/eQH
aicFpW3JNBMzUnGs7cl8hYbKnN9CwUl57Yge7/qBEXZCvRay1VxWTegIfcLI3N54WnpIW/uuhrNS
XHncbrLYKTwdT/7A+8DwW61MhkN1/ABtj55CpTE5eWvxsxniJ+E9yK3625CRMNPgiW025ybCn88R
eyOUW0TrtDTF/1aevayju9mB2MHmT/lvh31zsGPGJ7D2ebjsumjmbHGq7kf2oqq2PVw9M96F0Gd5
piF8Goy5VGaWosI5/MKuC54fZtcroWkWlx8w98RfmTS3WECWAE3UIUU2Y1g87IZOXCN0A0Jwzg+H
598W0NzHTChXCdJ0DeCsf9+LHdAckm7wZ+iJn3gLpgWinSmquRtSiI1AVuVE0m4ejcIh8TWs8jwX
chnGAX93QzOTiPEzQbshLpkKbGHFaHBJdrpvpFXBIAIz1nclzebwWw2YNxfHL8LjpJpllxx+oK5V
TaNEZggMexdLEhiqGK+9n0jopUDeGeDFBtNd97xRgu6aaCGpGwgrY9ZrD3lxAtK+4EEaJwKMYuVT
AybY62Jhi6LqDYKL6UIxxsSp7zqy/eVtwCfx7Mvc8CByn/NLBcaW8+nm83yIz2Q8ezqWg5gXlEVS
R8oMsOR3DQGKXIeI7iqhsWcTjAQGlH5bwwKupsQeS7XakAoFuLJ/6G47pCJcUR5iclYZ1lgl15jI
M3gLSUNP2qzCwZKkCDHzSMvO/Be7QRwNhyaULdm17Q9z4uwj8BFi9tMZElqQxCBA0NKouJ3F8YtF
lCqs7S2AZw98mRrWuydNt5mrajfRjbS2o7NJ7f4/k6VyLYiSTkxYZiczxEFFloku+avZoZFr+b81
FtG7Uyih1lUlA0FJjz8tIc5AKtkF9DTZKKR2sdo2ACkj1z2laXHGymCvuXOb6oKKMChKaOgPM9i2
9sMldj3lv03m8jEuImncUCzEctDNZC1RvjEITQrVmAYrUsNWWQNR1HrxDdBAP3F6mKdayedErOiO
CY3VxG6tPK14JtyFEYK8XWJC8XL6keXosa9GHY8zqJjB7eO5vlHf+G3H43Cplrk/L4MSG9JlkEyZ
xbWalmpaJ3sDeRyJNhmuvR9g0IgNdy0DvtcXiZFToAPGdJOfrCdPvVpQloOUMHXpdElLjOoQtMnf
Ad3ddyTyH6u7SEblFclahSbwGtVCrjvdQO5OcBM6yzj4iEPWoASr+35Jo/eavFyAZeHuaKsZEDVj
3FS3WhKGUZljImr0lB0z5LVo/U/FqaR3StvE65KaMQeFlMKf5+Ff7u0XBHF33Fmn3aoM602D38LA
B6nAN9/fbF8UgVBBrhhoJJNYCNg5YlkRL7Nq33WTsQraIXvV2pN0ap+zz7eTTpJa28Qtna4d0zeu
qInNtxCGrlfRGhm5c7Vc/EyzFMvHUcZIttNuToE+Mw8Laf9MICsz31Uv+18zv+GfnoS8oihBN/57
HVHrj+tNmiNYWW4d6AjgSaTXQCcLxB5VOZMDAKC0aj940lgF8debLEei4GPRN1IhprAOZ7ML8O1w
H8p+PF+Q48WvmpHzADmN52NECM4lhyHZJQwEuJU+WWrVf3NXiIwmxhFaKxl/E5Ld9WLW/1RAprzQ
RCAUPAahLg2QqIv1JUQHXAuTPBSKJQePjMjT9XIXBwnkImdptEMaLXV2fe4ADlio78cplT3znvZq
WLBzOAEQyLI/cVxyxfrPjxT3xN/MHFB938Qx4EzYdTwMVuhuQojRm0zkon4ZCal4aEiKGYpWcsq2
rqstP5TQI927o3MuaosXiJnvQS4FdzpVQ1oXAZbqGjjDWVHMem3QbVhgk/bc2aEYSlR2j64UDoiU
BpDPOqzTKla7RqOcn4egDsPG/eGdyGWtDMQYw91443D0HuHcYAGwCJhFjLPQISFxADNtQDYhKPzV
c7iYPhybeVpgQ2MLwHRomduBHagQxMm68FY80PAWZzmgLUJlRLMPP4Cqz4qDEN3PXrrqCFRykDk4
K6f+b93NyebXBUqkXKH+J9ii/D74Y8Dmtq4/Iddl3XYpWWXJQwdqXQcV0KiUtVkMlIEROWO/a2Bj
ry1kvdtsYEU2kS5QYapLa+OlDV5/A+pcIDqEwFf777a0XsA/kb71d4/L6eF7wBEzE2P1lotrFUPo
EgHsd3WSwcALXEaVQmcbMWKKd8BrEqOY/8KaN8nk+mw3nWr288JiZ/pJfxJQDv0jIppAMF4oYk8M
qbBwc+Iz4jr1qyzAqqymufYvVnjxLzlK+VacQVBvgQ4A5F+4TAk4lkqThejgRngZPfL4Ls7rYLEF
FyMo99xikH0sIEZYYsFusWrpiy0LLZ2oWHadnSZ1SKZ+7KJFcLILRSHDVDoOMqB5fsVRLgdZPPNW
lnnevJbY3d8qmy5OpI9L0GlPEnfvbKvObnuYBaSMejCOS09GyYuPv/YamFscnxgLVGGVmIuNiQG2
02SbMyDlqZoLHB7BSbbsKovLUj5uVzqOQC4Yaz5j5DBpF3Z8MTkRel6KEGvIT1oZtOKacRx5e9vn
bzWibl5pe7nY++kzN2vFpYnABSHbxwTm/215wb20XnlPVZVSYb1k4xqOY2+bGA5Aqm7fk2llUAne
UtCMBlV+lL8ptgyWPlj3RIk0vVlPFzzSb36+C1YMbNCVXoVWS5epyWzthrgC1QDZAMJEjLUc1pws
ZRbkkZYpnjSPMcJWg356sL2+Z394wA7qWBzqs8JPQ0aLst/Sb2qjiUeh8HlDWDal7Z+/3xl1uoZP
CkaKResoqP/GTuDl7jpJUSdpwFmFzCWHZrkqMPmB5L+0fv9xN7bL/zXWkKly/zuXh7P1bIFfgttU
ancyiLhz+AERfXy6dXj3TWo1Ar1mc5OLgvV5pA8J58PoOVB81RXHp9k2Y0oZ+nJVBaiKQOSAIx4c
/xSZ6FtQEe0ZSbtvwLLNEKX5r6F6VLP8ueZaLeqBnEF75L6CVOecOzOmrZlGp2BhmSLtB8WzzHwz
nvyRP6DTe0JWoYXiUnXfR+Xaf1zQHWNnJLFY0FWbHrrefG0u8g8wA5DjtdmmR1da0ow/93SAFuCc
0n6WXzOl3SSyc6p2ORdLkcIa5ZItUoGuToB8Zn9aW2UeqNhO0cHzKbLOjdxPm5owKb5GdMabB8Y0
+zyh/v7fss3pX/JNZ00yhYmoySxNaLQv5PfalgsEDCWVgdtQwCWH76xA4lsmT+PiJe+J4BxdsHcj
QJjPzQgkMNb2jpphpnocawU+tbEJcGol+W5g8nihmud4UN+j6iPsvqh2SgNc1Om6QVcBHzgfYvaV
/jWPVHln+wIw9dptPc6Po7bpx/DjkhtTW+qkBLp1DaR/ssIc+u733LvAst9SfS0OYiVn6LhcafKd
iR7SXrIys8Wa4GMyEi70Ty2j0tDI+v5b3XHS7Be4ogGEZRrOcuz1/abXyl45vBkWeaKNMXSQJ9fw
+gMrFsHSuS8i0J7X6m858G0YzyN4VKVP4UyFjY1/vz46Fa1i9nZPwpjSgYS2Cob85aVvXleGM2V7
IRWpW0ZCDcstkI51jAa/olnWnUseX54zn5vzAmDWwylxqSDNEFGt7i8sb+9arnxeIR3+8fYtPNcg
L4v7G/C/M42Ii/tPFK0wWY93Z6G8gV04p6+mgWPsqemK/TBefObkC+EKze3CHcCj4KweFQeNmBpf
hyFvuw8LVFPiOu0XsOw2QsE8qhkrfavNXajmhgVchcMUrW5gLjblsBGwqBgeQZZgTK1B6VVnkha4
Tu9QmkxNH35bgVzq+Fp0dnDFQCuKaq8me7QNOl4hRP136qX1fduPwbYv9AZTB79EFzLjWjwVean3
XZX7vzyJQr+Dmo3Z+xhS4A5oC9T1EDORkMLeekB55Q9cH+9lOSsduKS7RL9BV7Cw2HRhOunm/Ccq
l5PEckovDlBCW634kDWhniDzeWSWId3TU2pswR+9Cz2Y1IUqy02GMkPSUsFc4lvhUIOPGg/LUmUy
AthvbeXkTEMTJv9dDQtXNdTGuWzY7o1aY6rgA5vnglUKnJIidPN6ArS6Z1xxUtOJ2GHRxFl8G2Ex
H+c+gOHQzcILK8yy8TbZMcMmnoXw4cWE2IqD1bCugsQPmiqdxkWy9LPcjgOT7770o3n/IzdODmW1
HGnuslZllVkij0yKbplC2g6STOKp5EDgRyt9IRr4xnmtw43pNCAGKzKYj8uQGPd0U58TXJHEeEpl
RmkG49agUnzaJU7UQMXsdKdDhb7sVuP5S/H91kRI/9wTFTKgrZedOMk4snyIcNZRngkY69ewXpzd
FMpI/Etr5H9uRliyF+ly74E1PsuBEcZ5zzANhKFzs9jFUptMdcrF9LUB30oImS6hLJVggeR78Jlq
W/sl/9cdHRw/3OI+BN0q91JId5kUm40OBximN9D2PyZJEY3r1gbg9OxLXjfeGPxvhBbfotKrtZEq
oCAIlFxq1blkEwk2T57gzJGju22eefqRacaz9KLEGUuYebHp80FeiKtyQSlWH1dgDTdiEvLau0pU
YRYM0cnwU2Ak03k4v80H9NrioBEqJOpyPdkECV/ArSyi+lOzRISNABhNc3+JXtlZxTY28z20P8og
jr3JAwoE6OOPD6RG4SuloL/iz/TF3yB14OQOc2gdR2EjDqPp1QgSWERmyqVVtbMil4h0r+KBzq9r
jdGcPU1zWiUZgjx/nFGsdKFYcr32qQ+L5zs42Hp/Kny/e9ZC+q8a+E20UbttKU69fjLI7gdwotTh
eLonYIC1/d/vEqENNfYrZliKsyjUiEuD3V2drVElbyY8FhthSO/TLBJynGAdzZ6OrXt5pAFUxhor
plM9AJ/eEHJcsKCmYDfbcyAQrjVd84FR2B1xQVm8VKH8aXjANyW9JqR1whHwoxJUoacCOClUYZQs
YWSYaudynSUBLFi8NsWsu+bIHqIC3hBHngo7Cww0ruDJ3brXt72E7b5OMwHTWmP9hwg9bhT18h8v
DaRnDS5p4uuFg+aFX6R1AQ9GITze9b4s/gXyM5qIORCnKYqFEhuAy4B4l5PXkGvekswx46qcjtYz
VLnaVwNQp2El3d+Z7Ol7RutPhukFLE0mPg7cWvIjBGsT3/By7vAm90GRqzLxKOMULhBEwNljeh6q
4xQNz1k4CXJWTzbqbC76lEjYXt12/NmmZ7wyGXA4FGdynGIFS794NCmYoQ8kC/IqSw+HMVSAFV4s
spKFI/cnitdN0N1SfeCoDFns+VwyHcCD7dFdShRYZZzHdnN7fkTdB/LGntjsTIbAu95SWeB79hyb
Rbppw3OZcatbd8hs+Yu6nGO5DLP9Yyu6LXXkrZSyH0VsSM7c8UZ1RI6NwIqYcbDiUyQPMUF0gsba
VN8QoyFqMvzZSsPmbw75dKVqhezoFWA6y4n6hlG6t2OKpBHWV/+ESDH0EBWW0kl9fE4j5faxUwr2
7cylMYuByjhvzuQIjB+3WKiOezw3Tym6LDyamk9pRxhEqPb2bQYwYULbNCDunxeClydWpSu9J9H/
fe8FQN0Lwv+qm6IyE4ki7jARa0zbgEPXmrzc2ssn785K620ZDdc1JdIKYRU6g8FnqMgcRVDw4UTx
HtIuxUNocG/GSFj/RLPmxtHMG55HzPOdNW4lgk7B9gr3+jRDjczrWeKdWmpmIPEgoA4wV6H2Cs+p
VWyKrQfxXT/Esan9pJ5qTTrgDLVUpz9FI+2XTvLahpsY/Ruet2+41q57mviL0UCgKiCZ89RgK57O
I8jE+Tb5s4XkaYYfivXUa0TuNkWXxnqY9ZUbjbvQFvIa7V1fV8ZC9fuHOGVI1l2kdOKMw+A2BnDx
yE+/F6p/77GbcfCvQRkeXu3a/fZNboWpS957F61OhQ0NsWqYK6qTzHulE2VW8l9YuVQhAP+iqZ08
w9xxw+7cqhT6/chIYs0YwMJBbXg9EoGSwdrwTumEmIrC3h2VWfMwHuIbMxKZVlaV1MyWw9DWhskr
nLx18KHSYgDrFCD8CSvaV+BcJUEDeiVBvgnbErKfvtm0+foZHSzi2ypjPIW8xyvmIdz3RQuL4+CS
/fA2wKZCJS1S5EeDeMFvhc6mcH38p/eDPwtVLUb2jySBixGY6COow/tHu2dzYD6W9l+v1CRCXLPd
jVZWt3kFAoLeWC/7iIS4DhK+TlW0+boLEyyl2Mr8X8V/BOIWRvmZ3iSP4memxYHAq151cMYqUXMP
xvbENAABNWeEBSscZTiRNNiZFdAsfBiHhQd2IYpuUmd79z+EVeMbEuWO/zeU3ZtfSTafA3du24mE
lMyIhf+Eh8zoj7N/cu7uQvdTIAiuxPJDRJQH72vmeCuBjH2Tb0xSGF1iqRVl7k/mtl81ZPQJqmyJ
aq1DPgjzaFUYSPB/eC6uSQ3K5VtWun7adTUJdOFnzjHd+icnHo+03eeDJ4/yicy6+n0LyiX44Mok
uBNz3Kb/cGddN6zY+GNjtus77U5AmRZ4m758Adijl4mlxrSMUQaiQtKX0HNnvIUmy2aRCNI0Fiq/
3ZaYuKuCSr56fRD+k7bzzATee8ouuqpaBwVdt6hthTFZHuiTE7AOQUhUNBSDAAsDg6z9ZABZZNDO
dCv5H162gHd8xoAXsBD5qbYqCbsiU4j7t/hjLI3q3pPhxGxkySdZ4xnlUGrvGchFotuCqHLyBZFn
rEnALUP+2sRV76tu0SHHiXvvKnNLiSd5PzeVW86qy6yQgudFCYf3aegllTS/bkUL3ekB6U9OZohf
wg5rHnUZ1SHiivk+FS33/tc2vN8xt46T+5UHID1fUveoDzzHphTkcZVZXNZuDjH/zgRMsmCeMwWC
/UmgPu0+pIemUYkz3qv73KL8f3uIew5v9rs6/Kj38zIUW2YlE9qWdVvKiqb+oOGQi0HxlXz4WKYu
bQD7MrGu59uH6i7vfNpjJo+MmJfhWlMvvCwuDKqr0GCECkzRO0iBLNT5sotqXOUdecM6CLWrx9W4
gqKpL7ECgGXtcN0PG2hObQc0jGTIMVf2dcoYDheb8wpaI5v9AwDzmgDrUE87VNvE6RdcV2hWsSfj
6sqg9nX/Y2iBeggmqJqaNuJBFHuElHh4XSEWNNEFi+Bp5h+ye//xzg3KSVmg5UT5wecaPY4Zd1j/
aOs3MD3L68TfJre6kSzQ6DT2QPb2e2rdeSASY62Hz8RPgcjeGY5R0aI94GG1HK+7CAeaevADQ0lh
za2Ntf4c9n9PiN1uD5IkSk8CBr1OCbkx3h25OQRAPyyJ4t2xWziyuv+8dvk6YpJJDNd6rj5suIR6
/24N3csTi2dp/HmIvEcqf5hehA9DKFGP2ykvuFMx3zxAiukb0HMrhmTqvN+0iyWI1TRH1smO3GW4
UtTa5eW42sDnpshDeVUl/quFrWU673se1G16MluGaeG6oIvPLE53kVWZDxK5j7Q54njaZNaeFo3k
3KxJErHpCLW+LAgP01ggZksB07MiQ8nUfdDHxROkSpyHoxymvrvEX+6HmCxDafeW6cRohJdmPW4u
7lFJYGHOC/yp/YIhfvV8ss4S53WzoY2NMqjmWJefbMhg7JZfAaoJvrafbCLtO3XollPUW7ysRex7
V/BTjZ/zTZ4v+hWdFMBncgq2Cf4H3kUVmQjpdraIBu9VA1ZTrUz643ee5IHTczij80LY2j5i/f4C
ikL6dyGyYVkVY5oHsKEwDNd8DYfyzonQCDdyKVUcrlk/mCbnn0cmGxTScPR560tW4BlRm4ycUeRt
QDfcYPnktkVPSX9B+t3sFW4vtzbMBlJw9XBPDSOcgET4Xjdn2v+G4ewsKEBTlO4I5UhjQm7Uhygp
Snen8PmQoQzfMhjS/5C3UU7jN7CAEEMg9KJa6I4G9HTXCstQ3Fzny/SGMKPrkGMDa1iz62S5bC2g
ecwilm+Lrll0hjDWdbAvl3Po8CVvs9I9d+C8IiFA2eJFJkhj/aAF/P84Hv1VlYclpPQBNeMleNpf
Jp7sHAKEQspYx1INzzZR94xzbrs/2BKXXYG7dJhT1vwQzwLpM7J7B9WaZkLkEu6EPen2FKfQoLep
3C/h43EiOu/s1qhw2OSaxeRuebK1agXrlWhmVQbefR2tEUwVzRzW4rnhrO1j9BX3t3JDtK59gSyq
V5iBkk0k2bmL+KEe6NB39LbzPetMI7fA9Uwj3508KtSLmmbSIf0SHnWKkGLFAxniD/dVlosAwGjh
96sLFZ0V24/8PpT9wZDUdjm6UbH+ZPY5qDRE/SbpXekUeiZ8+ec7mGJHnWJ5yO5xvyzGtdRe6k51
lTwLlef6u/+TYmSZm6XjXm5yljXpae98kzxkCx7PRB1ECfHBSXEXvnmVjmMZnPBkoY9NYE42aIi1
faCn7Ouoba5GyUJxVw4ub2YLoh3h9xIIW0vUdmjP8F/CIUYFWYyVS4xw5PjR9uu6SVYKLk+iQR17
RCViq3Y8wvqhixAnSpugFVCiGgSACSxu7BqaJJ58oIAZeTzeFhhooVE6kuzflZEQ8q31vwWacGzL
3cI7QTjj+kEUeey0IYMSmS7FuWwHKZs6ty1N0m2Z9H0qGozwkXmVcNN2k9BKxECUdTimWNCaJ7p5
BWF3/PDSxNQ74oMHj/HhX/6fGhiDj9FpzFdjR2TUDSQ08n23LhNyTNFOh8Rti+4ERCBtpwW6/C42
7MqsL2EKyG8F+nn6c1vv+DdLyALQbmFhcNhRNWlEzo4i7V6tx3sGk3ssb3Csf8PTPvr6Np94HSxj
r6p5rFhqQI/SE4NlXXl6xSXREc638HGAD2Uz6UYKlEPl9YImbwzW6EDEwg/1w3rW0vKt6W+XvZRP
Pbk5pig3WSnxWIeKRYnOBGzdCcWX446mb9SGFfZljwH1LLuVk7WMr6POvu5Pivj+5GpQ9W9uvhGv
JYxsHbViU055BbG+kLqEK8ztDGWQ2WdUKmn9FqRdpKvp4821gigP7zwrwRgSer/2OS/WnxgXwH4W
ZF3vyZP8KoKXhW243e3Lxht5ubSgtEsmQos7yqo82UYkMLUMMVcpHJyALay0xYMi/XeoHHMgLy+V
oda3mJs8eGCgS1TeTFrDvVPtjbpz1YK1YhXtxNunAQpASgu8FKZ1ezx8AgBGhpMKT4JaT/JIz2kq
FGIiuc19u8+TXat8ZG7OuarSPiYiTKZtNASpSxVP47y5DjxMkMDJ/4ulJRMtFSS/ECU7vmpHUpBN
bCTtwP3bMC7M55S7WxlazBF3Vp1gKXh7WK7JcSmmIGhqAKpPmvdvcVkcvLhCeTmzt2rGzcw32Wqw
lC6DetHeLg8mtLKxwyE4qYwY39uEsK7VP/nsV82TkpMNoPHZHdwC1yXSWoUJHEUTrwbUaFN/xsji
g1HxvyLYjsLhNyI00dsrR32fc2+JjI3D5FMpmm3dqyMeJALwCg7dj+NWYEqB8JsVdvdlX0op5p/h
sdi9df14n2ndLPhrHfEkAkQHFsjB4A/WYak1HlPhVfOFVvcR43YFiOIKeHI3rKB4r5frCvpQ7/Eb
JR6lHr+nYv7JsHfUoFy/kpuYiBGLWlriCHPQSn79o+HuVCuxbMXXjrZ0jzjT4JPUnkNqtQzD3JA7
M8GokzG9F+AqNHeTGzie+Ec91h7Pm++8Z62+N3WjvANIqbYjH3/wrTT7StLoD7OIFLhf3q4BSIfP
pjeS8WtXHjgH9DQQsUb/K8/YLqExs93DlARPZWZha0AM6A/iD9MP0EOkcizZIeCWPWqytWrUAOzF
HFNzaYHDkIm2goN/Jxzzuf8rt4Ag/yP3W13J2eH2LYOxoXUH650WTHtQY928PwBX5gwe1yd9bXS0
G+mAIOAK1HdxJJa9mnrROnc/cIbgzceKUrj9F3PQVo9Zvfb5Y/AiDBgDTS4RK1f5fjaVygOwNmsf
3E4moG7uO36G7Rfjv0SWsqXtmizZFetUkC29NYjJIlU9upJXt76XuHN7tlO9CjuERaQ/GpLEHF1x
krWJODSDWzZTWYfHSPx/DNPLitjpjERUuMZBWMmTajnCEHZg0lnDPRl5nTmKr6jMIXeyS/DdXn9x
VgHHW/zBcJxreSGnsV0dv6Pw/szgI48yreUvyWE1hrLJRZaBesWAOjHrK2ifwlqwG/V+qk6ToJE1
t4+m8WDfiEYQ0tHcZHUKuraO+78306qrJKqn0M/Of5RG0zCUfd6YTnUYHxUXeFGPoYepTMMpduA9
KjGcCwcfzS2GTLtz9ALjTwl4J3X9OhrL2slTYGacq3jSj7/7N5jucc2OzkFmOM6k1oGR8UCM+qag
N8t6AXPb5MiHewplkdeOHA4N50iXE0xOE1XJmekND5lediaAn0O8LRXG+XwAvTr8MDaqqCbdkGH5
Z/2P5DSTBknyh/lKe+CTALeAujz9PlwgFw2G3upwgURRvOYnR9GEIKpsMhb7eFYg75auq7sLcdLm
K5Y/KT0PDJ0o8pTEudf9Tq80gUkgexkc7gXMpLmK2H0xZxU3t8arIOIGhBoWB790dCofw+RH02wY
yF9Cfn8HG9tjgndXOUiFVcAsP1Wj+j9Hcs1ZuraH/XWVQYLzzVus25hzCDL8B1C5XXN77YUaq6aV
3JMRfBvMOQQ3DpVW2NBOXmPfJfpi15gQbFkn7binDSqfFLKtqYc36zFmctn/sXGKsXGj6zcwNPeQ
mxHSO2K9LQSNfrQStmcXOuxisCBdZnhUnm6CdkBAys/RvWjmh7M552qFwe6sej1ODjIIiNVlyAm9
PLoD2gmwAUC5lyiULpELNwGzy4hGTlHFlf4/0neIRLAWIcJZi2OKad4BUSXtKGT8P4FkKYiCWcmi
fLwhAbZLGk3YQ1/VHSteJARjQf8eZEkkfvilO9Y2ufnlso1Hv3ZTb4GqS0srNg17FZfkgHsMS656
/n0I9aqF4YCPQgC9OsK7fAiYeWGpIrn/9L/90+SQXZyEiB5JDeQm71CgpbmLB6c4w/YinQftCAV5
JaQIWFl91VERK0YZNFv8leJEKUjtCCwd/3/4yaCBJuWbX9C3ZwlaDsQAZKlFtSbVMldukh6R7KRG
7g052JqngM11vBNxQFtmce0lqbkANlaL0qRsNVhipe8VE5dAPCSCX1zOgUBGF1CIn8OzWcGxVUg9
91XnYMeoo7rQhDA/6RF3f5GS46pS6rY/hS/g9jyvXs7aKNYmXyAiiDLQR5GuLFDorXCVsy3t+9Vr
aCaGXPGyewUBantgfY+iS4AZl1WmJICuS9leJrMzj6XsQ9NEF9r+sNiGCLjk1CgZhpUFKgufYQUh
G4ROBXg1VSem0fnbDW/bQ/jlxhbXSiBfDdj/VzbxbeZogE9dPD2HaM/7QgKA18aE/Cbf6/Wdnhyo
nDUsptd3zSbesVc/kKqIHMo7IskRDz+7KsBvzmy0xWND7YJ875D2brYTGvXiFNI27BxTtdvEeSe+
yKgC1rYTioHZ0Vnq9nQixObsPzCxFxcydkkcqEmJQWcRB5JpuXCmDd334saQMXwi70JiFcKtm0Vd
YYPK6LqfeZMZ/KnkTedrQ8osuS5N6jFJjVO5Nyo0oTyKsHw46E0hzXCsTLLj3YIG/kiGXzr8WIbi
qY9kqfEDdcGpNyRxgVT1tSaBe3aXYTEdU2rZ1vQaj4kUnEUOLcDDvDs+3QXOryaWBGjfwamSSRC7
TcVCAVctxRoPU0rdBNBfE9CqkLWHde9MSQcCOmBXBOn1PfGBvyaC/+yx9UKWl+DxPTEbPWwTAMp+
Q76YPh0ygN4tZ2iSdXYvjXsOfi89nYYRQ1QQ1nJnXkJGTM+rpqB1nfnW+1pcG6Ca2nGCwZtIsCDc
Da8O2hr7y7Jr7aKIcZvUtpfXr+/NW7rqJj6HyyHWyu/2eLk+JCpUVis9swyiy825QGDsoB9r9r2p
tP9tguA+7E6gzT7Emd06RMHAuy0Jwa6G2jv476o4H/k1FZaaVMecBfBeYvCkzDF3PId0WI5lgbOR
IPM+EJqTJhCdl30bopHm5tRG8N7Sc/MfdjOPIMexabBENFJpiU2s5RbdWwAvrC13YGiOOK5ALq/1
+NCsWRNeHsCkHrrfrevZeTXzipP6Ow02Uwf57lyNKPBMjGbTMoxgtTo1h8kK0fMYioAneG2NIPE7
PwdhqddNwNtaKHTp8VZGOH60n7y2gsfu6qHl+M0+5CvUcu0wureAat6auhlumVvkEAuzmqDd8bdM
UxqI27LNvZFziVHqZUK7lSJE2XeTFPBH7tB/ODqwW5Ju2VPWGW26UaCeShWalHRmvv0e/gfoR+cq
jwmsIhGCkATZUNUdeHcn9cNuGl0EFycAYHliFRcY3lEWBcQ+KfdkJSp3p7UGAPUgSnTEe9gmH/18
h3Ichqn9JZI8KtpzVs0Rmo8bP6rwB1oi4GOlIuAxzhrV25vUfEF+/oY6nxn6wPbIMWOSVEZnvE8S
2cxOCpwADBk0xLQsfKiH6QZeqB9mCGUb6oEFnaXgqFXniNd0Z/YKcSSpRew7SWHI5hA3airny8Eg
8x53Mdfy8Qy1pNiWINOYIhK3H2RaNOnp+CUw8WlmGidisAqaz34E5s88tGv2D7jPpLqvIr1nVCiD
PlSYoIUls70dt/lq9ECkEIoMQj2Lj1Mc8mZGjybzBheHS2I3IPidosi8qjnLfVP7+qcK+6Gm3hVt
3vQTxCtab1YYRj5R5yhw/V7ux0/1PL4Zp0mUQWoiQXIpgm7Xch/92DVy/YkXlU+0YTiRvZ/BdNhu
xixrE2vVPvFygMGfWpp3uLj7/PhRvWOo3yEF0dCzg1vPpxiUZUv46ecLAdBxQwPM2CxJfDgP7d1Z
o7Hth8imTj7uAO+jGYEcWARWpayeV/eKF+bJ6WinjBvCe0P+yFJNXrmundDqbtSZeZVnJFVAOxYF
WshkhBo3/Ijd3YFlxpM08n5yf+ll8DR3MPaCI9Nh+yO/sYnEJUAx3pJPdI/6IJVD/x2HWaYU+I13
lwjmIUl3x1mpRTyxPjk5BNe4a1feuoB3BA4a9ibiKRNu0jWw8q2lZ45ubga1BZIXck+tDZcQbm9I
Ea+glWvbZocjimITTg5Gg4hL90/MD+wWGiwLQEZgGamiLRciqEj+djcTV1r+8i2siWZXFi023YKO
MviorMqeQMXnk54Q1DrtlrO9Rep/K6FEU3vDtZb8woi/evd2X9/nIfNqHA46a2URHVCg3v+/pRGa
Fk6fegwxd9/k31l7aursOtsKi9MHRuNJKYcB3qpWdhFEZIM5V8JCsIGnQaepBJG0MCb6RbT0D/OI
lDNP2BMSM2890EijPYDDd0Kw7nuRLjoa4Hkp9kbEG68Gcw7TeEwRV7XJyi6fL6BxnN07a+Aeb+eC
vJK+N5J3xNQiL6IpoNxZO4F7vXfrpnVc29CByOfMzwKicuq00O5YJvWrxcitowh4IrYC9UFytMxk
RRSKxhSvFs0DslegRxsvP4DJRTOMwhzPF919HCfZGv4z2nOYvrqzE0+1OaapKI1QkxnIv1gk0ynT
ONEcVXZwF47o+4TN6isPPVfs38MbI0J6lSxk466LsD7UTRpCIX/zvVP8ec0ZOa5Ddy1FUFv+/hzT
FBbIwSVpXNLz6XR14XYypf894voIUHDDgsw/WSzTMf/qIcAKYZxo8UbZGPQoN5rpmpB/lzPfp4ps
DW1L/At9dfnVG5euK6zWL0UJaZthRomLfvKRzaRFcvmQF6c1uK/spJBMC+Nzy1baOzVJg2iCXY9g
I9y2Qyb0g+55VNtf+EE85KESYt4iBgAN+N6iqqa4IwWYYzlej/zUSVCQLv9MHe0b5DvVVUUI5EVz
AdBPyxNH+4q9v5iaBkhJG1dQcg9l4Kly95ZP21g84+mY6045F4glUl/aIh9gi5yyGWhwrtnXaVcx
uu5/Jc+AfM690aGlrmf7yPSmR/Ms7eCs4psS8jf1IDKwfPc63eKr3spUm0fMGGTYuQ54Y2sfBBE/
QlC5wJCCohL9njvHfnwP5KAKUKHMPIls4dGYHVaKqgGjjbSSGptMzW+IUZl6CHT8TqF7mTDW87He
ebsPU3AtR+Sk4iVGZ9dcitJ1sMZ6dBMHdDiZ41KxEh8dtrfYnaibj9sgKKk5yvWvVxnPTiin1T0p
ZHFGSaFlTcA3aH0n6r6KLudKqEPk9XOYOkVIeYmCcOdBXHwTRk5O0tUanxG3hGoerNsemi1Ph7vr
rw0kwTScBE9+B6lKzne0a3tmSmzwNiUQEC2VrmVE1d9LjFBcGxwAjamjIgJqZbG26rNue4McDRDj
7lrCu8PDVe/Q3ViM8DNNORjeSDS7Az/RQ6tRK7dyHHTEqjFKr6tW99aYxA3zFX+bLcHUHM6ZolML
9dMJKgeMWSHu5NbZEMWwtSXA7Rkk9OrQ/NqT6nYmoYeOFyWRnWM2lT4xrstOPIcW1lypN5c3YL5N
5NF+l84JdalsOyzTi92fLASj9KpMFFP9eHc//LK1HPBdDDAoeYkZ4H2aJepLCVX9uhLHvrjdIIwe
vAdAIvgu6zAoL2pi7VbiUiLwAvngxS6Xe/H8lKXYXnVEpYMxKWrHL0alnIVgeiOWeSlHfI1KUmug
9fGyxbePRNVYRE5q9EkpQNH1SPEEmkmZL0Vud7mL2wg1j5+sz74zgANvxsds5guGDY22yQJwLU03
vOgrx5LJ0V02vOvG7HmOUqkDERQXDDNT1cZp0EStAA0XcOuy7zWbTjtJ+Qa28CUuMiBmXLfcIxes
icxOMUY6QvTu0gC7Wl/lmYMg1BcV6DZDZaKTw4M6fjBSlsYb9Ay7cKl2AAe1LfRRMlK7rDhlj/Xg
dMeC91WnH0IpK9fjnQhKESNLBQT8UMrwZYwrC9nUuzGaOsCAeqO6rXd8yowcug6o5WW+mNphfo/R
ddMIBzhghnhGqDqkQ1pDcLL9AKO2Y3AzES/TAbZssvck8IaX1MxBa3I6rCG2Z6Dw3aXtMNflyrj5
Hv+oW64UIA95vUvb/AQ4hPHkw7PX6q2qM/eQfNmiV6D0WKSfwsuCfef/jwATv2A17mvt2uC5xiuE
mF8HQZW+dLlu79xg0dwwyEHeZ3Od5gseJssRqy0pAnSXLrfM9QoQsyXndUCor9ordyjBNl4dRho9
vC7JHxnsOXt/s7B1m3UdGoLZm0CFOeLJ6A0TIy8gbq8gUhghGyi6605ZUJoiamgvmkrKAgG1/CEb
tzIVGcrddNsgQEQzKKTv0b3qJUK3jhFder8oVi058miwSKl+BzdcT3jIzKN5zYl1kRCZ5rrkcnCJ
nqHe0Xi9if0YRK+kTnJsHikPTuvR5sb9JSHXC3gIf7E3NUS9vDzOj70yAlZ2vAVJtdCx6xMwp9mJ
h8EPGWgvq6RCZFseVTVXtWLPxHmL9DoogFatC05bxDpFC7g059Ks5KXZYtder1dlxQgR1aFRLB2M
OZumCrha8uwVEQd9BPHMtL2gB23nUnWVoTNTU26ulOQuyyZywTqV9dDr/3xELgN7hxqneSJajdn+
j6jFE+iEE3/4JzhFhWX1W57a8jrQchGqlICzq3M3uIfPt/KJuXTy8mU83sW6nGmWP0ecxOiYHaV0
9XBxUHE3Wzv/qn9cRS4GSSa7qB/8zZFJ3v386JPE9uNuL5Y96LlyrfWAEy0bVpteDsaR0Kaoh9GT
eMrhAxJGgU9fDVJlyiOHmgZaZdqr/j0GdM8eZi4aY0gK8KijLbotydp6TyAREQQTjVsCM/s1kzZL
zocq44GgExzrXi3VL+eFH/J/ncXJhzJd8buoThrvRjwRmiFgsilVNGJlSw1mf8ZLFVtWc0voEGrT
Phm9hL2YH+5pva3hRvSEXpDxP9lOOmkB3LZLVnk5brD9w2bvBDl0MizEAl4YQMS5VD56VAOXySYb
+DHWN3yg+Tiy4BOve0Ix4NQqymunQEE8UrKERvgYT/mYFhZqahpp3ZTy2tQtedZg0gvJurpJrzFo
doqMa/ZHvutEk+Zhc33VCJJYbdhKqbc4lo0JjViess8lKH7oFaVqj2LiNCGY6S1vO1RGyvxcZVXN
u5gqD52437fwOX1pMAz5dgI9TjL4KDmd894sp7LegoEhGncOnFy/CmZj2kCO58UGXiUvaLbakcbg
VfojaXVk/geWPmC2MyRNvlTE4HX6Vkj1nckqylZVw3n0kOZ86/9XdQ5LM5hNTuZdrR1PC2S1h73T
z9NCRvie/x1R+y+GRNXwe9zeiqwjOPzmUVxVoSA+ZooMXa+UeaKpIjWMVfFHQSNQykO4LR9ABenP
iNtz3QRIMyaOhGZAZ4Kn7d+HXHyman5APe4wr9Zdhc9KMQrLqcZ+0TGI+vypIAD+kElgW4WOD9M7
BXNwcK7HYWp3bAueJQ/sdTB78bHzcGfflNfA/tpqiLIEIKZb7C5LIg47FeRYZqkUp7R/UBtFzByV
tmc5XSnzLiOQZKMr//KGs52pCvKbRp904tUgEjUuPbDxjfofndLQQ309YAJ8yrRoFPd8Hn4r1Xgp
9wNvu1YxmOBxn9T9caGzyqNB9ucYz0ZXYbNEKj1d2ZH0hFkqYHEdCmQzaOVl3ER9/L0qGBlnqxHY
fx5aISWYDAkg0T8nLCO2Sf741BRfFsyfXTMBW3Wy6ARzFpVHGeQEfI5OrxHVRkffhl8kad5mMhVN
WX9y2+u4ndUibm8EkDRllhm9b3mY1AG/fTqMiwReydFRUj7JsPw+w1Cv5y/vMoVqj4bgcKRYuwP+
DBsaU1eDGOqboItW6P0ew8y8dLDTn0Y/EjWRLSNExTigcF+EeIr8oHEklE7/e7lwAgKkSeI23OEZ
1rE3ppeeRdeej8xDeMDB6Oost2TrdejTdSpj8QuAorn/zLjeJ0Gk2NzOoMZ2OLvzzfxfkQfoclsL
F2e2hT37iz2V8Jh9Ci+7POPd6yjdArDQjVhTPDTlxCNN1yjgiQ7S9Glgkc4y65oDx6QtWblG9VbE
0J+yecQN89TYZsnm1HUAk67xuarFE/OVIFdNSuSQUWIQYmgpFZ6lyG9AtCTeGPZooeovJtezyjJH
0FmcTa2SBIs88tL8n3dn0BCAukfCGpr3EjBS2EZg58QaP2uJ/c0HsmcBDWJ80qFvil/2gqk/FH8Z
EuYhFNt9Y6k6OMq7/Gt2SnJE3DmapIpedc7usgpZaMQ5UExDuAuqkL+ltcgzLCV/N6PuKv3y5m3s
0U6bWm30+/UQiKTw6W/xAJ+RnEtoyspMvMll/i9gMXUpdykLiaxDLzYTUWXKTsDXj2f8CC3QuTkv
l075ZGrAQHKlMxOEQm1GSsLTUG11Ciwjx1uhy7laGYeNujtrvcjh5QDRnCREWxBiOKE0qggysP16
o++gVvvQZlFNzUY8KqzlEMgsR7mQI76o9qelZMlBSzzmaajRE3WTiGyXM6NMyK9AJ/tPldqQ/LmR
oYG5W7TYW7f4R3MRCCKayPjjqA0p4r6UVpvjbqWKBV0rM0ZvzmS4+KRI9u8L2+uNRt9qf5zMqv2I
wtTcNE8eLC9n0iU9lL0Cr7OVeEN1YOHD0KVM/wt1YZo7RnHr4Nh2XTe3r5UW9GE4Oj2cfVWnk3vi
trS1yKVVAlmqUYb7N4mezJYSdiIJ6YKKMmeA8LVQDMCfPmgCA9Dw/cktQ1aN7zDSj/EoIpK7wufM
GZTGCiM3zeyGYmSw1cF4tBDUMueiG4nf1nZZSarTvXMAfgBmWCItvIY5vOHbZrWAJKN+8C63e6HI
e6pvt/YX+m5tbM5G7c0neUm5mMXjuWKp5Sn0vUvGGDrmWnhXQEEd7v0KNM1xtWoCAk/a23WNdRia
5KONk8VilpmuGz90zy8J68quSeP4G+2m2NHnMueBf4BKVy1RDrf5u7Pyf5UZssLKnW/uXvl+MVY+
2FlquphA+SCsOnY6F4jRFv6j6eWEvQR95HMtDPaEHY1kmK8GhDwCe2NHH5GTjNUFPxKSZspnxZZn
np2/6ofUH2PylWlRIng6Hy3m3z7vw8Zv+ZPwS54qPSxGOeXdfqxnRNPUlEg3SI9ElvwJAJvMwIgT
2kZP3vQyIWyEaucf9l1EZPc9fNGyz0hl69UrKX6YJ83TPf/ufjxoceRySCRDPgfNQOFNhT12YZ7R
J9f6Vo822k/oSeRAbT3NWnq3DNQZN0HWeIw1hOeVGzldr9ldlTAwvxmkk7Y8onvPiH5AHxcRbCKH
qjrG0w11CR7Ksugxxb2obDyazIA0R8Hz/U2ZM6atqecPKF6ezUXzE//w8o/ZWdX1eRakZ86sggjm
rKHWNICKrw+rzYv8Oza5ln47QCGATEMB08K3l970A7mbZjb5J0zwL4/3mqjtqyzINeWn9EUBZJGh
ZMDPMTY2BKD0/YVIbzNM3bV5rHgMcuSpT/dml69PpAfH16+5UcjvvvaI/uXfPy6K12XCIpUH0Bvd
ujkVOTk7Ch9OgE87lTXCqQjJEAzqWEDpjh6spfPENXaqgsQkjGuxt9kKuDJbnTRKhVvSXwQQbU6t
gePxA/kLIDWRVeMa0nSWwSgaaBwynyLsJccw9FAESTTDBinNET8pTFOB1qyp5vHgN15aZELEeJ1Q
93o+cbkzVs3ZOWoKnKEOG0R6IrbX4kf1GLba8z6wcIli4IGUuvXX5GRlygRiPx3t5zLdJfiG9UeV
7/r9g5DDj1vIiXdsiNOeC12SToIxseMJVo0TbD5xmw+BYcEMcu79tz1WBc5ffiR7QAs32ivrL9ng
8datZWezGG7j6VGugNjHi3t3yX6IXPrg/P4jaejU5ArrMkbtAXI92QVVhAQGQCMi4QwUg+IVvkDM
ES542z/hGQQTTEnWfzM27kWMHwi86YitVW/Gv3/X6cMd/X9Ca7pGiC/Iw5jNC7VEFMtkrAlfj0+Y
DIdR7QsTxDt9EaEmSTodmOd9hXoLl3VboTLzBAe1DQFMMSFkO99GXgQjb1usi1Yjc1oiD+5MCcpq
arhCITlG1eUq0nRQC5Yv9sFhk2sA7CG6UIpHaewqxtpCt+vJRcFa2Ztmihc6AmiFapfRYL8ZdJL6
BBvWeKr58hIGub10bQkBdhz2aJGtRXKmWrs/l1uIniguJ6PYR384lx7fTZU1OSMZFSj6XI2c+SjL
Uz+MUrRzV08OVyTqUy+0VlEIJIFBGSQZuJ7GMPJqTxxJzuoKoYnD6JkTGPLgdSr4fVhnyxsRLKqb
2ne0jDmtz5l28X9+1LyC6jE2M+kghgxpovGVt/UMRjrqgvfb3mbAkuXP16h+qwf+vdZof3OO6Y+C
JGM8S2ofkxKN71nQ5ZeMT7vqEkVX+aonH/tHVVpSSSbCMzV69RB77n4q8dH4MeJwa6qHo3LkPfe/
TMuInTv5rm/2Fydk4lA+KdNGnkhs/VJzdzipCSahTjcbzyiA+c6ecrBhjpcRORkgrqm3R0WJtPgJ
Ol3DhS4APEufg0yWbyB09mdlDlsQ+i43dw4xrh/l7S0dB9FYjeT0Y3yUHze068GR3Xbc5BDFBC9Y
6fbtoe2MM33aa+N3gob4elV2196QTeRu0xysEBM/ko/8ZvXa44WdMEVDSIGxy1pIVK9eXyqBCgRG
oK80WU9pEMlN0bDCAHcTp5wLsdTdZhn3M2X19En2kM5HYd/k4bA8lsx+7BzKd5g886mLn/48cwAf
IDOWSPx7wZK45e7DrSQ9zVqkWH9x0hwSoTs7xOXxUM8C0aSKtj/4doxzDQJFYpeFl8BQUgbsj8zm
n1NyhV6nD52O7mtzZcAx0bSn7UstBiibkw3taWLyytQqmolJxC0/Q/NUuJCLHNql8IzYDmLGAFjq
xZO4WfHbRDzHCZtGzzsmucrCAD0AwNUCMcpsOY1kzx6IsTjxoO9Q21VxII6DDWS1LE4WeYd/Sug0
AnaOIVSoThFi5JRlL+CZVCnTsI0MnRuQ0Xs9+LuXQviNNEpEn+V+CAMqEZtkAprDmAgMP6v0FHb4
/Dmbs5yYEwYqIKHHnEEx0OpUo4lATBifZ3urnHgAa681JkrYdK6aOJKP6674cr0b73myM4LKuy67
TYRrfCbQv4m6m8ZUAw5v6Je5m+vmUoyYJrfaSjf2CNcikOnIobf+r7CeSRphf6kleAn/Q9nU7qHI
AFsjG0Zg5EPcN6xXUNc7v3j/4+VW41w6/zm3/yba8KpcDtdd3y1EdbJnUAeqSqirCdoME69tRKM6
v+2pQ3J5YusTfpjyFscbkeiWI9qPwZ67ER4Ujs94z3pbFmn0F+/QH0RU8sNcek7A3B2lRxZmuqPO
a+t+FlBNEPsLkiYEtH0kTeCn50wcR2mYFyhW435S85lpRGchAGDV+HJ4lVawlmimXe6IImCFPYOD
SstpnLFLiX3fgO5D9jIFcgBycoDg7th1m/AnLFE97skvJ0SSAIQ9ggWBlg0sIFCuo61gQ46lafjw
Ims5bibWlG31LH6ty3lEVJOyr2Mr//oWwCZDEOXRn5ey/PykbhPFt8j8x9URJOvcvduhUFrrCTwL
2C2acPZJOtn3kyefaBd2Z83wvd2tz9yu4VpePYegnGiNhK7kzWfOeoVuRIfpDKe2kHncBv+rUwOI
G+JMCWtE9HU6qfwcIWbbi8+wV1G/REYh+C8ZzxerRtjfcKKThxn2p12W5O7VZY4qy/VjbfFGOJX9
W5PS6u2JjsM9rX26mY6dtovxS8EfSmRoyqXkQNJwVAZkPA5QO73/m5RnPv3zKJy5BOYC6VHE7wcg
D5BB8jEX2denBj/Orbf1nZeTVtUD7fUor7QGK3xJGab6mufPlSgbrm4SVRX/2OjrO/lJQL9KHrQZ
ylpBIp4dMAzaTVTWcaDG1X0Cx/CmbkjBsvaSyLXKFhTSlNf12ZXMP3gYSy3r5FpbEXNF0mWUaZPq
s7sobjrwlHQjceqCaNAoiEzMD4H4Ovm12ZV6jWpbxG2syHYbbFJrw8lzz8JNgC6aZlhvYTt4Keq3
u2fcYwmg8ZJSxitOZOFFoLJ3/r96QBQXdZsy5Xk4zXrf5UhaR/QFJlg1VSgpKBMmvsPRn7OSvytJ
zv8ZUjy+Oo0QHtB0xAqicSakud3lgt1TE5z7kyHAaFFmuS1QvAYXwr/r6xsQAW5MGjKbRIkQivgH
M75xGN+xEDqL1VFHFyqKZlZpkoNV1mp6EsmSO8ZFCatznBNrFX7e6ySz67p8xoedJfGRdnP2iJZf
SSBslhkxXR6MLpRHvlFrJvTdYCx0jIJv0V6xmgaTTvXCrQWOYBrtQV8p95dZ1g/tZqFyqouASaDQ
HI7/3QLFG9zZUMTPzkV6QpuTbdkKeHjR2I43skDkBCMntcT71EIYbsap6tl4kYt/IIp4/iQfxHHt
q37EoBHEOfmWDXCykKIgtDZWB3+QKDJwXJzScquWhGEjeU+3IeQPyik0S+X3I1eCOV2i2WEYDyLf
c93N7dke4W0dYQ3/VfnejXeSEdfH6bZP6GvZGjoz5TD8zADRMrxznA3mxumUDK8YWkz8ua+B4AwA
O4sUP5T8aWn0ADH2jF3jGJxSmOkgL9NSYoHAN07PHJ/kQovkhltkoxWGBvUwj7atXkDx4lmAkbav
/T870ypDSKzDfTX9qjthYgAPfbdk4BLYA8UBCWy1hkV4UlaGlnycBwrhbQBpqw6PZEsQIRNJP3X4
v8xudLnMII1XoUH1O/uYYbZiP+ey1o7qDjjJQ460/05RCKLo8vrKYh6V2Ziq7f6g4K2kGtQYG9LY
pCrCOpDpuqTI2YP2n8yiWwLItosuOi3BERBrnznqKlk8r7pEMX7f2C4I2GLAOWW1qIUNiHCErLVM
M5O2IjXH/YIO6eP/VG3L7AF4PlZOvvQu8QKBNx4ZPcieM30IK/ilf6epkSl3J5XQZriv3P67sB6f
0MCADPLcK/GqJzJ6WVc53OqD0I4+ay4A4biA/YkpZZGJ8J76i0Kp6e1VQ6jwpzmCVYvBSYT/4Yuw
owRcv4c8E6nDIhW9siXtcqnYeFiu56+13cfmz39a8L+WYuckNNZq1W1AfOfaWmZXH8xYGK0pNJ7R
wezxFFWsAiw/WeYeaL1r2Cbb/buqXZVp30DK0buBYqbcYKNgtmLWbn8npo/qEQl7ljFhAYr1oI1I
hA3Kwy/my61sjIkP6XbdEnzKy5w/Apg64EakjWFts+nDoJerma2QhhU0j8Rsz+l9yzFNrJ/TwL6/
Ui8bhhGi5rgCu0k+Hga8Fo27F43zBHMwck7w8qfKNTVWP8y28CWx8RPX8SWqlKCmIsepN+ZLC24q
NwEtqOvf8rD61vsqftBkSoW4PWtPN9wJ7OpRGa12NMOO3qmQCE2NtuYFUgdP8CoUn0OaDgOtIgFy
EkRAOclnz6hrMXP1veYvblgLDxJCecQYcdhqvhLvG0YLA7HFAGam8kLNtIH0jZef3zjWGnqQ7AfT
s6ne8mW6WU+mpVaOFAP4fu/QBH7Szja6PpEGmJ56gdaLGN1BnLJukx0Mkbe/6vu74ijKXAOAfBkk
k3nroZjIn9atfUqG3bVzw44cUQg8UQ/cT2HBtnwwi0/dRhDgIa3S5VwXpiDNivXz+gQBtGc0H0ye
iuWPwBYJ0K/GgdofcccfVPG/W5mEt9CiynT99NLzXaumquDw5rT+0CVBIg2ttDa9Q0JPId7CIXF4
b9t1tyaQvY4CGL2HBPJFWP9T9tMOcVen7kvjxpUzHXncRXvRVpA3CF5qfpBf7Fff0Fmuilb/8KF1
Ube/3SlY7A6LfOHftCPgy1aCX5D1IvT8kYkO8KyX1PzU7GyAe+Vc0t0qQz94fmTa9eCEZBOT5qJZ
cIfPYfcu+IwzH4YwA7qts3aLD/UNC2zAaRzbhHKesdgzPVGT6sRnG4oApY3UqbJoIGkJvzgTuJqf
wS5QHxul4KVIrg+B06cNW4hxl7WZfRdiVRdY0emjAvI2eG0wxX3TmM8caidDYnjewHQcTuUaPfCq
wXUob+oCYBVHlmXPhM2dvv9GSLF7LBMVbw4IrQhTG+nX3njRcqDeCTHYEbnyBT5ruvHhokmiRekH
BWf8TOwVCuhcRkpvJ5GxK2Neg7m05UvwKJoi7APy0eV2tizdiHSU1MgrluTgCm4OzPu5mtZZt0HO
zXWlNxBWekMbp2qux3GFCm5ulOJCa4xGcXPS55mdVFKYzOfneA4JaDIJzTn1vgOYpZBrEftd42oF
nKLmdpua+qJsv6p1dMHOQP7DaiNvqKrzEBauOJlX0OopLeUTIUV7gdfmOHzVRtnTpBye5RJ0N3ec
M/RMEN4iepgk8UgtQZkevE8u1r0gHyJDIWuOzKhwqxl7Or9a21DgN5TWJh3Hdt/u+E3IFGvnp2L+
5nkNXwrP7NNJ8CBSjjSPpr4TDCoeNSZOk2qSqogg8+uX7l512UMZYStJRbj3BeWpCcVNAkRUAse1
YYsv2HEa4u8eh0AwTgOzFuWkmoMeEUmLFmCwgLLPsdM+7bhgiZ/vd3p66vtb63m+seNM1BB32z7T
BaeVXb3qwCFl4P9v4cRHhAV+VWnZ0O9j6OjdVqJLTSnzHkt6fvJpA/zibbHXSNNAmOTgH210p8IG
ufyTOHv428iGxcYKGL63nzvoz6StzODUc1tA/Jxqev8zgfwJQh5rEGek2v+D4RQsrdncVEVxDOlc
yqPrruZGUFM3mmovc8T72DCqCxdP3Jimc57Qr5H1N6+6MUq+IKEYmrkYrsjZmsiOIrdjRPZdZstD
leJgKU64K5vASNk7hgoiF4NSx2WKAwoak78Mmw4UB8b19wSoMoCaQwsJTwofcUw0NAqAZ/9sWAws
98Xxtw/+LxDiUMkU1iCvtfxbn6LCFEdaBiSTb6rNsasAMP2+QggzuXfwIK6psrK/7DtiKUfOhw0O
2rFWc+FNybR27a7umVTtIQr32I9OZdEuPn6OJHMh6MZ85JLRjbD3rQC2yBAEyLGZQExwpm/Kmc1A
vTspOv4O0/OQF11qtfRPjLMZzH4H22sAoShCdI5+3uFK66SgrivjRb9gh3QdT4s5R8JFdxihGy0Q
pBLeKX2l8RNTE9c8sjMwnt/pdlJvI1OGgG5QLM3ICGeBF6KdBIoo0cXYr4ThylXi8P7yxmruju1s
m+lmQP79VM+6uXk7FfXNCd59M3sE30Mo1RSRIhbhjEsi4L8TxD1CVESumjoTtxoVjWAIF+9GSLUx
AYxDq5kf9UOdWPfAufMhIb8wEdhZvpB4Eg0TgeWqUnhPY4rdEwrQqyqt4XMG+turk1+kkBLEc+Mw
u/9zkBzPrknnHZHcluuvEmPdpZ+e/5rjFt32SZAL2lFjJIbi1P5YzADKUdUCTiYzKXuIYm+4LHet
79b1PDoQqn4cdUy3jhBDuhhMFAXy9ly4TlywzoAtHqmzgRz+zyaQ8Yz7BQKW3IloFIYcovly/vn4
kFRmHABvtvTnoUEiDJKXaFLdXOpSKswHhjGjue2Hbc8jHQxr7MqttX/bB3e9QhEi46wSoxAgSGjO
4MvI7KJ0xncdaA0vzw0J2+r0ANfM1wWVCf98ilL3zwu3vqVdKVloQZ3p8cRQ51ymWqT4MTEje7Ta
keRhcYiwlC0Ak+7BlXcCEtb29HyFuhvWPNsJl3g2XPEKzEiTUa0mEsx+zV+pAFHQ4C4tt4w/DcOD
sciRy3cG7JAL+p2TmJBeDuStYCy3tuCT6XoA8cJv4UG4uNg/s9BQMYm11NdPD7OtjnS5dvE8arM7
yUBb3xFnNSRqWTCR2A==
`protect end_protected
