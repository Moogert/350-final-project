-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zTm+EOAv31JHoZYQ4wQ8kyPImk+qTt0/F7/fv3K/HQhZXu3Jak67SqiukynW7m2vFwHII/HIyKp1
h2YRXaX8JpxcUvVrU6nYnQCvD3diCkFHvh5iqiVG/LuZP07dcN84vxuec4RHaNVzSmmE/XJ57FC7
Xnk1FTE4wz3lheUS+hL/YxuUz3JyRwBwUC/nzTrDpyl4b+FWTkZ093we3/FPqiG7jPjPLRV06m10
7TRWgADn3WNLretfsQbtoQCyh3FtHX36sRfBIWnFXr39gXXlqTrpDPJHFve8XXdbanao8b/Qbr8L
J8wU0s3H1xV8Dv26rqK3F5j99f25jtCfUOTMNw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
hfavRTd7WvmTidu5r8ZbsSGsZL1E5DXXf0sXN6VWfg4pDagVQvhC+Am2hHxkltl/lOLXVF7ERhM0
+LTHcjP5La8k/qmVuH5IQ63BvEVKRvuk8aMJUOrhKqUupAJxAkkUjmbD8kdsFXmXf8GS5iDz0l0v
06+PohkSBrj4bu63x0ju988knNFWI536l7I0x1kRGyg1UrBHpv1fD/4/A30BcSkBKcH/T8Rre2xI
aS4f9kci+AcaRU+lWy7rEuvaTZJj6xu+PwZCWS3QF2sLI/BQOrRnI3VkVg3rcNBquKKfOTf3gbv2
Ok4XEXawNJBZCzMxIkwyEb2OKWqXsZk2QQ7KQy2V3UB3ordww8iK6Z1Th3RVv81fWA7LYJbOwEcR
tokYi1YOnjphBxykFCwTb7zyqcw9K2IY3HJuiczS/FpKovPuXCX9BxMVfv/ptRQR/gP8OLt1nvmA
LP7UBQ3BH4tm+hK89F5kjt7NNXYvedx7s7KezNBY+ILSo5NJuX6jElo4eSrsXZdDQuS0QxbtOygL
uVqhIyr4c3BzxZUug+eGnll7pkYSj27VXPm9plkzj2mB03C2+j8rUxIkknwAa4XV6r4c24wtGiD6
hqn9zOQZQl1rnlvSMHwMN658Ogcp4BGpfQEsMjjX0bW+u89Xj/k6f6bbskhUPvG+hZgfMUjeMhIL
FjU5z40UBLd8SRTcqoIxZqRzHYqBahAUC8O73eN9cPwizEGwdkKVkKHGk8o/lE9eg7Uz2fXpfis3
Ygmk+r4bvxZfO73wyWop1X24AnwpIpDxpz9e+6N+xnc9Kcnyn60JGRYacccXWlCsvR+yzD9Tlr3C
sQ2/aVHiNfCL/HX274e/YS2HUM9nwi24rJ3CFnk9QI6HArsFYEytT90TRHaUzuXjxS6+e8mXUp7t
zNWt/BV1Latk1Z4tFoR+O+bdgrF02v3EF3j2UYtoAvT5Dv+UIcuGh8zbwBBkPgrmjaZ7IWMn9Uvc
41o9WRG562YYO9CFOdFVL3imnPTm0rsvBxaFz1wbdr1MvmjSfQ8So1Kf9n/oZ4V/sn0OlofxPnhi
6ABvMtZug0JTEzKUrevj3c113hUoLr+z/+jqmhsQcwsbhCZ/VHbVtdGR2YGlDvbW1sREy34/Shqu
8HyDp/9jxtvXcSDfV4B5TwVn6EJ14oGtDSH6MplEhYr6VqPgjTlJh3kdiDLwGjHhCl6GAhyp+5Sz
Hi/zIMT1MqMHKmxf9h9T+2KPNIt+BnTiuA/Lu4CubJAko+T4CZxZ5WZWIwiNTWsm8vMU4YMKVAuO
RUGqa8ni+UQR6pAyPyXL9RfDspWDcfMIbM8cu3woMsBLf21hlfLMMs0J5zx6L5YBZw8Ilq+vPUKf
qaB9Exk9GMpuJTI5KJq3s61WMXIxppBXwpFKrZbGTNro3qg2wd2JGisniuKC9kXymPDVzSp8vsxe
KszaW8gyStKxJfKs/S1U9XmJpB7UC2ZvNJ9ikwb5AULYOjPCWe09XMiZxwe8yPNxsu5QVBHCZTxb
MmKYoTbTPbDQb+pzIvpQe7+OQTfnfCmxzkj0vssedpApuuik0JA9zcrOx2KJh5M4fLC02VU0pTf4
C792sadNg2kbRLuORIC55xgzYbLGLXtXO7eJUIIIRp+iWsdvqrSaMdmbGDb70vTzoQHAvCXxMdC1
+KKOm7enIPuU2/al6pqz08X16ifbmPtt+CIzOpyEVNysCOfdgsNBUyuaggeIUNggiJ7S8hVDCth0
7pQ48nPEM4tL6YEA6zmK5EKNUQaIVEAK46YIUxGvIvZfKoJ7ZapIyjXcd5nwScn2/b4gk0trHV4O
Ry8KW6gb6kB6bEfcNtYfQzq6unms5zbSy2bop28qv2ZMYDMkRzjQChB3FNfs/dXbhc6g42/cY+jv
tDSIIAySJh7YrQk86byNStNn2nD6D5/z2ZuTTXosIPICBqbaGj6PouApO4Q1UKmgYgeJG/ZHn+Fc
8JWIkLq9yTD15ZxIisDYixjFOStL2iGh1BwH0R8vlriQ9d+6aD04wVa78J7xEFdJlDXx9nItxfcq
rxkZF/voVah60QuQKeDk5jr53bXzkazWaOJuIAejwGn3KMJ+kdb0U0ZEMWrF+xFTxDuB3aZat738
iiK3NhALVBhjbxZgovaQFuWPNSqdhH8vekn5BBhYx4tJgT2ot0fWe9cTKxv+iv0odHfVHj+Ogi8q
5F3rNhWg7d0tLLi4KTTJ62bwTj1XyjOohAGT6RBnZSMZfoxipoXkubK/IJP0+YVWgYip4PrHHWOU
CBDQFLxT22v8HbgiMYyMRTNr+0vUoqlShOd7UZ95GNaaXDRzu4Fx1143WF8QJRW8rk4n5U9GEC9x
fqtC2ZdxuAD4mPk8PznCQOahVnhzUxkbY3MF63KQKCgQJwWYzx4DOtCc3FO+Ljen1FmivLktpa7B
r0YtvMVaS1ZXxNfqpB8Ym6JCkymndm3D2s9b3+48fK7vnXa7CwJPAhBOj1d4kdr3Nic2gf9r6jcz
FxeNtYw5jUTabbLLYElylMhcyfytTp2aakOBD+cgjaCW06GyZ10Ys9pdn7rPTew+00VKCtQ3JIDj
GMJLf55XEMslDVd3MmK4naALDPaxqDIFf6cHlnGrq9/QDuuOZ8/hhTQw8FjfIdseBg++k9EcAdR7
TwKga4fFrTXKMkEjW4rMOne73tr832w29uDEmjEmLeWNje5G76iQF/nNArku5VvgSIihcCCacnYk
Gm1ebqKN9xL6Qt7pWzBQIZkkQnDNuqX5xWQH/NdXQzgOE0L/ji9EIVEqoxyhyDbEmywhnyTa7Pwp
YfYH9LlNudeokjeGs+55cc+/pEV3jWJw88fuE/USDq7fEJ1lXMXwL4TFntCcYIui5IDktHW1XthE
zMBLVx0BfUZ8asdpot0oENupbWBimXgJij6rKqKO4GJ2pD1YRK0FeIjBXHN4MZIoxDGKMvtqFmYZ
zY7IpwH1KvdEcj/VPez6LktwK2MErLd2nSb/HrolXXxui03R1Eb9bSJWWTY3GiE4vMjdZB0C2Gqu
/Yn85mRhoPKK5G8KugrsZfjBHo9D/c55+S5KANeUu6QBewCfseuxmnvzzy3eVBwIeWQKyziIPm/o
h1cU9u7yel/1NioRMRKvr8GHnXFLP+kb/CBtMEp3geWin/Bh8E574s6tCehzSnbqDu1fIKx/JNMC
Z6r3JdzhqeOo8GVtzIuz4xqgXQbe80ntYFnrI2cD8NnEdNetd8ESkHlzBMQ33eQlXCND6zokfSug
RsYATEAkqlA8wyn9myJHf+11OUuXHDi9/ZY8wW/h6OnG5dhVwJptffKMhnyQ7v30Zh/Q9r9MLIhm
zTsOgOTr0Iv+73i2NuTJOJbx+9sPMoWBb2zWzxuaAblT0r4sacVcjqISlLEsnfT7YKlRwzRzWAQ7
/KCHWRaVJcfMByuNddpFFXPF4Xp4UjLJRbQvXyHpGU2ROjgH8rz3ECfCG35DOjTuor7pF9smEOal
RDhd/KjUskoiCthixJY0owlkYU7kMSe4E8fCRLhJ42dbSHeaO7mxnvuU9xfxOH04K2g46LR8v2Pq
LmqUpUcBYeOFNI/4B2dhUHY0V9gGuNwKwScZkAlu8J4GDFPQyu6R5CowEtH4RGMjZZ1Q7t025ucu
y/AfUxzBQu3NfhyO6qgPTRVjhm85JMCFrsfJE+khmXI1B8XHs3tAIdiwfUqiqe1aDrBFnxUGd2KQ
X1C2gNjt1wB8/vNxgj8Av21JzsqQh52fXkwtTohJ/UAJ1vuN/unLq0ae8j70EAjGR2w0SP5oJnvs
cgOAuk2C7G4IgXBuoKXUbzgv5M52sPW36UAX+JRh6sSMzHIR741i8LrXa6tabIClhmdmnCW5uVLi
aZFIuOPvbAnZurdREPssOsF88b3KHvgG/FaLkL+fU6zIuRaeB4gyLcKr9qd1WVtqeH8oo/WesIPL
DnnCQUHIWI87aT4rcxD1WboXjZULqO6/s4MGmqjwC6R7CCt5rORpgIPjy0wbN/0uiArnce55VOQb
MIHFbkEf5yJwPNrWrtZVkGqRFv6L2AQDj/b9IqheMtbcBZIyk2nYhTgJxzH4aiELRHnFGdT0+4J8
sdAduCbMjeFBj9bGhtELnBRIXpt8C1jrcPKk6D3NHZro36Fn3sRoltFqETBBXL0qxIVVOG5+nCqz
XudkcnCObp1PK/lfFLZzRUuFSRsfVJi1VmXIQGXA95AU6EHoSXYTsoKHkzMOeZqVQkB9HzFzREfI
hRu6CAgG5mZUiRnbTkrJFKYnHj50YB6+kR18KQpAND9yrUqcaWxOUY2vAsPopn9tb+f0Xall4V4I
fQOdL3cKAdlCsTkjCxK5USixVLfmBWT9NBxj6vOr2oDXrZpfIVEbFcqIIXlxA2cs2vIQov/Khr/z
7qr2qD3ssQh/cZ84c4g+u5iY7O0av+plvGw34eAnWYldpLWA/3T8vaqd1qRQEpo71yHBMKOUDrNx
hrpins/+bTTqnUFupOvYa0dO0b0uanQgxmD2CDmpEpFuHeLzMd6WKdufIiP4ZWsFlyZBs1BRhuaA
q9pYW5QiKfEiFKdMKWiupQ+ZTFzxMnXS3oyJHa6WV9ulsaxyfm9MQaOV/5xbRX06B0X8IRfcQSBK
lfqiJuz8zr/h5qbppLvzXGNysEX2+i20HZk4X7uX9yX6CcHLSmeD70gAlkv4JWG+EyjhqQ2ncn+z
+7g4oNlV1iJRRo4dGKhpOng0f1SD+dS176f8RIfOjR0l0/HdPZLEYFHnLpmzolUUIiu3EyoGJL1k
VTbt52d8KqRNrGTJ18OxXMhY8/7KwBu2KpEEiOSYermROwDxZoHNYvQJqSwzMYXYk+RTSSdaVAaV
nrwopqPYUIQ7/QHO/5J8jRHCr5IwzFH7h1I6GCkKeXeP7AXFyCFsDXWYL1MIPmVIwoeSjVHXGnqF
BTObTJrHUY/IsGsOqTvqt18JcE1VT1D5ukeqAWS5pKwHpuqxbCl0W20ssaQtS90JGndl5p6ih3wK
WVs8N9VvCJ+wVgvFhaV6aBdHQODaEhlEWJR/ICBZNfzQoEeNvYYHL+j/E6uKBX3ZUJt3sZ18sPPs
LF0jxf/RYEkMtbX21PVIFRXV27jfxSSXio94/5xlBQtxoUhVKhGlgCigTh1zHm8roVg+7uazHiF/
5LTBpmkjJIy05jMVYsacVPz58KUTeQjnsd9J6mcrwgZf61Ac+5Jr37BGPJGtU+GrLM8WYei88AGg
Fp8JfFnnXtSdQFR3Jn4P+jzG/5dOeJc02CeMOI3eTVYpKO3oPMdHGX2s70nrSMk82NLCsf8hl2JR
RLb2uIljyzHa8DOqyFYEwvIPWI3U+e/oH4wk+szxLTTpI7cyGNsXGPnxoANGOwT5cv5Xp3mycB+f
jwpt0Q64oE0fV2CaCXV3GaVZ+dUnv3vXVOaLazq+4IuPeIvSFEcaTVOWwjgfGJnVkwPzj8g8X5Fx
xaf6bt6nmtFK1gCf29T08SNnCdQ5iUXkVvjO5NCekYoLLHexdwAJN3Ykb6Ns53NuLT41WMlhLMgZ
NcLWpBgMY+PpsRDAObOLnAEMC6uAfcZx9Zr9ubWo7jNUWM9GCNIW10Oc+leTRJIkzhA3YSGQ8WdF
CwbDphdNEs3VU4CfWl4PMa6EQTkTeauzjQ3GVyr6zoer1eRCYgH6OxcgylTDZYvWUVsD/bzs6aT0
hBV5NfHd0p9s5Ob87bi6P5m3AaKkYkzwvoI8+c0l5JXQrPh7XtpuBfWWhMlfIqyG0CzqwgMe0yGU
7OpEHWV1wN+MGjBhD9kHA4ccO3Ajklr4wg0XZSu5t11f6xxZdFDsvXcJf/FjjCsSy+M9l6WnQZoQ
reIyeHiP3Cawru1L6MCm0VLL9T8grRQvrSMDBrINw3X8XW2qtqB30Dv7hG/vNBkIEPRrGMjMnOBr
vs5D30GUDRKIQ5ur8T7LA5ckvGB6qqDAp/EcxiZpQKB/A9hX61xhY1yTxJmACXvGfyf/8qynraTY
yfOMrwkpltJAt84iQijrFInn9XLrOucYtj1DWAVt00muLe70kP3A4styfO4eFc4tXC8HbtuUaXTg
cOONeGBf6CtjreQlVbZMdc4ci1+bFUOn8D/avk50Kx7uyYpw9+TqM0cSr4s5TuHcrDwUwZJUlK+9
z1qKzLigdcGGXCgjU6LPvJ4NzMA9y4Z4m923QfO0ajPDIxoKQ2RkBKu0F4h+hDuVltkD9SjgG2h3
YnLuxnnGkU0FEcbPivq/VypHr2wTdE+tRMR4XSqM74Ya1Epe/2AE05uvAC516gFyka7ihWD57OBW
7uWfYDGDhY4lLu8RZi/V0yspsg/Pnsg2pB83TrNRVmB8fCU5uUiQ4Fn3tbeso6s+D6id5hZ1w5Ik
CEGlX+oEajRgRVTV0ArcwCSNOe5LZ4byx19bqaTv7GriEP2GDXraBZEYw5fukBPunQHvmw1+1cvh
l80b9tFGFhVemxMvKzQI8QuDGJSq4VEgRLLXyLH+NvZPAnAQ36OvSv+PTG0tmE/3OVOkF3qk5aEm
kBh8PYGGa2e4SXJOwMmzc12Az3+fNF0rr+V7iopIV+m/2QQVvcFgMKC7R4Sx4JZWtbi1VdnjOqhT
yzgEQ28iIdTSF0KY+Qr2EbnWqLHZLC+OgH4nO7vZB9ueVJYrnp9hGM0jlHVMryDpCdu/LgZgrD14
SnctFKZFIgw18zDlK6Z/zFKnHTg4BF/71Gvh4onC7HWNsH3/dH8Ey6bboccQ5aWuuCewLux3f+P1
vQ0jX6c4ondEs7BzjsmNmO0mNqNFMOP8yZ9F/GHhOBj8FXO5vKG+FOqCJmfVdEI7rjGXG1Ob5bel
8HxZU6UVtMq8Opa6ZWMbCa+zf3fxz+tKDfy2xaXIfBC3DtLBuUrdOa256RS9vM7fmuDa1samlB/w
HwcsJ4PLsSNmOa02De6CcnysUR5Xrfd/bzxTgnQrXpdslG0LqAufEWtH5Vqw9SQRDREEpGayziVE
pm2hdt6Uxw1t+tWIAAdMgNaoCBVT9JFInCIh74Kh0FlAp0UpUYI4Js6uauAVxtoaeG59lVQCkvIL
xg5s75/3D81JYmM6wFS6L2zQY1sRqUBX1zrea8O47uUrK3sbX5xbxyPjCk4KuJQljPp/9blRw68r
Kj/XChmw0uKMwxcxUGGufL3R4l/SrGYwVQQIWVPd+0TMms4Nd8W3urj1WJtXV6qnq9pMi4UbthYp
whcbzghIz4WyTfdCw1BRrIOBrF1COfU2cEaAiN+wOgUMmZRbhHAiLVGxPFqNavkWo22dGeY9VKEe
fqSL3MIxVi/scHllcNhkhnD0MqNTBoeDNTPJoMLjobN8VWWhq6sM0aXnKEPSoUMqBnK8MliIWUe+
TfdmYUolKAdYEZydQReA7eas2ip+xquKYK1zrOFng5suDecooqkZJTcPbitxfrM8RExZzDUHTkoZ
z6EGSqYB86zgV9bVGzBVcDI4iGroc7Gz2C7Pq8jhZHbCz7XrrK2s7eYme6k1xBMc0xMGOoQZ5Y7a
+KMtthhevbM3/mpAAa45DD7a94YHywjFXwYNSPyQb5jzbriCnIGeHjbKo/CHdSwun05fL5VPHwX1
M1VRq/9fRhMrWqrDr0mVo5aS2N8WUJ0bqcmI0rJ5jmUMhTPqioW1y1Ap53lNvcl64VrNE3IhC/Ju
+dWbBycZf+pCB9LXHU+G23GOm9o1DptmUKC1vLm01kVQhiJwA/GFqIeVTCreMMgUhrEng2T3bzkN
OyL92bKYDFXIRWB+MRTRlu6R0RtqokEhBMrC0waJKOG1dC9tHl0qgN6IZSFwHO3mfQsAHR2OW1hC
AAXLr8BsyGHUv8hqLjy5G+/Wz7pCs1tbk8UUHrbNdOFIArYHsSbDc5IJNIgpaQMZhUmfXKmbtmRH
fgTe/D+5ExCwozmpAMOqbOtlICM4Pbea5H2GAwd1uhW51Wx/x0OUP8D37uYJs5y6FDeWsGFp7+Vj
xmaGXnI05KMXTgbmdbRpF5/FYcCm171VMD85hdpkm7jk/banmRlPoDyAlOa36H1/Djs0hvfZga5z
ui5mUZ01IH55FpM49ltgh9XnImMcU/K0p1W44oCHQK57DDHfB2SjeewspuvA+JBJMA4RpaK2AEl2
3xLvG/Q7yB4uC+J8Hcl0sbRdJJ9JV8Tfin4EPHBMis64tCBSQ8pTbWNgNOSlP2zuDZKTs3nNSAD2
uunFrGNB1BFwDe3MXT9Z+yqHcyTH6/DefUip0caso7i3UPkFHlLi2z7UDShhMhIN3xXq+s7xiYq1
JMzWh8QqhkOA93jFRARQR94mNW+jwIz+kj4wcVNQQFcnBxsKL3Ty7PM7x+fXKFVUjYfLxK+gUxsK
sWeJotAsXyZvzVTNPuEfzBdsMrthH8/fS3S4zfVvtgmduh3RcaHu72A7ZDGr3kq0GEIbpO27EXvA
lCjEYToyhHLwBBuETuiZcwOKgK43aGMQvwB6ig2j/gu9v3gYtmZLetJLQPeR4hebg9+40Hp73+Ov
9zyXauR5mbPtvqEUNJyQ2UJHH9hmNXZT7JZWLdQQeonyXOpjtqSuPLqpXkZriteJpgX6pZY2wKzi
AZGCGBDRCGuGI+fYde0LKO5D/brWvG30d7/7JlAdvcYb9Uj72NTB3QCva6FxzklilpjZeEW+iqTd
insyGg2VCmGZzxeVln4PhS46k0tz+7Wp8DymgZfr5cRF3CX8p5bqoKudthnxdxem1UnGzFwXyNRT
5aY8VdzfiDJ2Jl6gIM3zytFkX4UDnt/1xZUZ7usp/U3WXogd7nWsh+ZW03T8j4nlUmXSMvzgTZdH
9ir9WKkhMkz85VMp6BpTBxw9T9sT7ZEp6ePtSn4Q6M+MjpvIaMDBGyE6VixizUQ7qyrlm1O+SxQq
ysz6wF7+g5PWbBCwUz6mIOFI+N2j5LXSRF4KUBygrgr6sdajdTJVq89gCbL7/yEEq3kZgr7f2h5j
O0jUznVDzxynm2p8oQBvsXoP+DpZ88OIm5mTNIezyxdHqFaBSsVyBm+HOF31qekKBxOIWWXydkpP
oCmrr1hBNN6I1mWg/NgEjsyfe6xX2Uw2Nzmix98YMLJumUmIElj7woHHUygyx60DUBd0NyYs5h42
1dJ2MXOTAsli79aPEovlNYD8JhLytelsQgLYAkop2tXxDGJEkSnljTUlqhVQUS1mdyoCnRmgUxhW
qS20inFIDPfzhhFBf/D+pm5vuUuddJr4T9BA8o+xBL2MyGUFxJa+AOOPoPu+iihVJOtlgOFIKYom
MecYh9C/I7/OF4DIcG59w3/Oie3CK+HjTBae7PT7ptWMLzVq2+RwsDHzooJvX58SQbbBOmRHhBjL
vRbRQiVIf3nMsgyYbga9YJYp9LWV3lR0jPfmTezzqGL/0DT2wZdCA+laJYPBlOW7YpZHpMs9MDt6
PAk0M+NbAOUYX5Nc5qMTGfpQsDQRaBUckBzWavKBCDzSUk/wrDclcwS/f0tZAQ+o8+7qTUWuevRl
5pOxqOjFMzZkCgKk6CTxONnsh74yj8yURpbX+gSbgx/o8wsiOfX6sW2bD4STX6DsgyN2OkPLp9Kt
Z/y7JrNCswL8G9aG3LA3kcVMiWospeXbGLhEVnA2t6FXIO5Wt1JcAnzP4lEW4wQSVGnlHu+rbRd7
aaJnN47nXJ2PgA8ldAvtkO5K0ldN9s1/A1R2H9qLSbbyoqAAM4dKmdWoK2JVe0eTS2DBOvreOqQS
ZKKv87A90GbKACOkfPv05XEvTwTjfpb/fYLVKWY86XD+OtvJWdwXSMRMjjrBFTKqamYO4BaBPqtd
z5XeafH03GgA9RYILerGlL4aHb50JnwQL4kuYfIoa4eLIxBB/2HrtJ3ZMLxChZOJZV/4VddaCR97
+wnx8wcwaAVHTtQ76Z0LGOxUQGmBOiX8k5XxfqaAthGJkdOTNLJDPAVrIy9b1TpDoJk1zdbDXlCS
Xn1r7pHnPsp3LRftPrHU6/8D6o2NHayudpik+5rVXl4mxZC5FiVva3DPXQf6IzoplcY9E/BEZc68
A2tXaCpDZRf0LUVc6oNaOxBwWPQKdL77LRenLvF102AnsDkSJIgskHh2gchQZKWo7fJkEArRXJ31
3WNmbB/zvmG10uz4t/msRjyR+OBdo0AKhadblK16oQQcI+eqjWlh+8LWzSC2ZEwiLc+YeJ8DYKhv
yKb0tjv3mSUcppbpe+44Zp6tL/udYPvR7uDif/+dcw+k/MgDRZAABQmF4DLJjWVYGsoBjAMSrEyT
9FIEpqmO3zDC/w1uY/SG51r3WIWw+31L21AaXpAwcWWJOyIyQLYgUtZruPGQEUTh2dojTde56y8K
Z2BBGrLEuJXq119/5OEirME8/LhLhVU4C8IlLqvbe8S4M8erzTL7YOrOBmZMIjya5w/S5H/h9zVZ
HMtxY5EY9eEQw5dM8LfSmLkIdmLRPY5jCObs4wHrgYrYyY9BNqpKqkugPUAZb8YigXHFaLfbQhrK
xWmh8HW2GR7mRuHt7lly7DvKh1ZLnTYNyAIcAWubz2cihJPo3RgtUWbguXSTSTpdxeHrVFfWvzEr
6E2ADKxNsww/URWVVHqn/SGw6qrI72TxTlZWS+Kpp0nQe+JBi6xsWBPdXLruR9EbREPQA4swmVtt
m2V997WIsgqm5aMn3WjB91Qpwoy02jrOEn/BlsAdVh8gpQcwYcWKPcRf1HKOBeNq3I3hUnO8DIb3
xzuynAUg+EInOYuLVdAC1wgv2EIDDgCTBq9apzbsoVV+DyP39PL5CWsiwQNK50/brWfhKFcKw8nQ
f7Z9QGnu3nRnu3Td6Ad1NyL5dw3E1Ginw79cwEzvHNamohE/D9sTLXKkKH2GK3s+mr1X0X2qaUYf
FfinGgJgGIY/qCcMzpOOiuJ3Pw6S2RZVMhjFqMm7X2ORqJ3jdKb5aLdA4B9vH4TFKjHnhU01sk7h
5taMatM94rCpqlr9z7sTTqflRwjfNUuOejJzSh9bP4LzGAC8Axpov/34JQDmRw1f49CVDc9fFyi2
cZFS3+J2+r2Q9X9ZMbc98pxUci7uiJkTfu0neP7NMyRxiEyig2NHPvreqL8xRtLW6znfizH5Z5Hh
WhvpgfpWf1rterb6Qe/4TnfZfS/skEYARBbEEyASTgGq8mqHluIZ5ngNhkWtSL1bkARBTHUbC0hV
4jlsR71Kj4DIoRYm73YBGuVbWjJhCCTc9LZoArBheAy9Rmwz3NnGb5SJu7rAuVhVH9ticTlDFds9
sCtHEUlX1+q19usJgAMLFKTAGEPFbEtvnKllWssR7y71oBgOroV5o1fqfmPS+rY9Z7jaApF9cOqO
xie6ThAq427a+MKDBNv8lnZ68YZdn30K66WdPPaeXfFabo1N8KAkOIlP8JXB1eDdfj5QUf6XYgPe
9RhqGZa1Op1w1C4HnGNpQJguduy2SnxQRaVRIoGZCKK7vzTc9n+Tj0w+h3CvHvhyH2B6WImT5MS8
denzEcLjWR9hmTmtN10Coa2UXPR0pR9m3yMFds8Ja8+A0InBtimdCmQPMw57lNYktcn2sMtbCdlv
korZBdBcx/CLHRAIlLDTYhxfYRBm4PvAypQsXfDcAUwNCLNV9isx69pPoMAU4qsBOCQp7eqRBrlT
H3Y2lqSlAW0gt3Ntjz65ba4+ksGleAariSxbR6g6HdSgFh5k7aWT9c+XHBeyg5a7MPHmmnzH30DH
60LTTOApg0ZWmdSAdC8eVvUu4dgs4rMMAnQ76YP/wSrirVOFo03FpW7sW6m7K8yth1cyjk11r/9d
yDFTF+1DDRwXO5bTwpT+ks9/vnn1qN9z62LRaMMhvznkxVr57zFjozedWeA4G0uOb81koJgho+4/
9S872sER7WGAeMKOPdO22bPHZHYBHUjgpP27UZqgVSr2d4NjuLAFEM7FjpTsYilxt3KLlsoGDrvy
RqqJPdb5abVVmXgRj1Vf7XuV3SOHIM4kKaTMou5q9qsc4m6MHCaMANLIhyqU104c8Qgc6P2ourA1
S0Zk7Eap7yx82VUaCHllP6faP2A0u9wRueMDtcQQr3oOHaudiYFQcNQNtIjEXfZH0ycNZ7u61S2v
FqPQzFRzd2tdljdAgtBwwbq6Mv0RknSupieSePl+0UHsSOfGmHZjw5hSsY1T4EFAnyIJGoAf2mCO
cqRi/mgVBBhYH9+si/ARjdqKtTMipm62xOqVgrEhH0eIrEdp+uVJhTga/Swv+nxpofGiOYozrmJ9
yzH2whmr/DnkMpvahikxpxAVPbLppUlxnv/9E1UVWb11+s7BzY3m2rtQj60j9UMAY4o4Q8f6BcW6
eBB0l7k8Fxduv3UYCA3cOtTfJuMMmT3aI0wwglCxLCzWLjDlj6pBDpWsUgSHJS3pY4tQHU1OTSxC
cSjST8ppBM/hhZSDmAO4cS8CPBx3xaCqjT6kBFlTMrl6WPj61WZ9VV6K8r743hotHPeDZaqu0/C3
kCpyse5fEqYCAq65doEbY71LV5+7hM6ZAvN2Q1l1Q0KMvS2rb69h4GpJZVM9EcYzGQP1P6i6fvIA
seeuAOAEeOcULyGpvFZXK1kPJGNkz5pcOQOPSoANERuJLhWznKvDTPsXyMTkk2c69/+S+C0MPwPZ
JB1GZ982L9m0C9ABrCIYrvHPz+GqouebVtFY+KFRntktIzeJ3PX1A1ZcThLhcCXdh4Eu0GnWa9mA
ISN2DQurrbdciHTlScOixiRo4u5RiyTcokd7HVJWppsVaa74Cwggwaf8mGWk+3tnuh6im2y/yZ41
Imzswg4dx9tRqbcuFO/S6d++xzdzK+CKe0kd+ho7P2GDRPMwJxWa6VHpi+hF11Gnt0XefTesyJvW
a2m48/pMWTl1osgKmc4jukQCXhy03ky/JRq1EeoJqTUHFQBbj0YK6cyl+HI6hWUS1FzFlUAt1AGh
yzWcg2Fszhb742XLActbO8ONKg/UJikpkZYswgU/sroNoAEl814GJM6CHBLCbRSvzDVVgT4402ub
tYCh9g09xgXDXO222OxoOAgbc9MAHLSOcyuboteB8g/dAq3udNZxGxXSDiHMj3vB94RtsAwk7MB5
IipP/KcbX9eaWBG9ChFUqbxr9+rVaNW21IieEwIMO7ugFYR6gcjRQV7It/ubByCzzkttMuityk0U
Bebt4fUDkzzqDFg89Xvv/G30ATTjFzf1ijWIZFgcbwY/V4Cd3IQNnR8kfHzdjO3slvobaiV532qc
N/ZNcA8GcOrYYB+XcK7ktI9m0/XXeje2sNoAAmWDxrzOTzDEYrbtRzMHruL4up02zXWEn57WVOAV
DfVpPBnXgkvX2wzTo+DADf+Yk0IofXAOGHjQFeAJcVl+adUbFGlY41W39+EaWLQlUcyDKBi7x9LY
IZonPPMLiOvVbQf+W7vyHMR2fdogQhkutNbXV5/aSaUv7ny1nVNXztiWbRlTaGEqUusXLJWMeWvp
uS8dwp8Ic5ws40kerBaNe+zEraBLVu1hbw5GNk5ZvrQ09Zz1+DifBeIZhfDOnwHp/tmzrM/dg3wm
Y+sqxSJ4NhmbH2eFMB70kigsPWDFlNzr/tmNstEg7BBYWds9Gf8KctjMOEHu7R1mcjKQ2DrPQPPr
l4oftZl/OBmE1BJ69+ysd0ZLNi8jVYc+208GCsBfTHEI6CZI2rhuqcR4mamIsT6ldpUaO9g9ZB5v
McqBA5PhnewlQjA7D2eXnnh1Q0KFal7dvZwVyArnaSCC8YaOzK7qV3mv54M9VFImOn+lYA0iMLah
N2PPmJdg9i8mnic4LIsEjL9sN0v/P6RtFEz5s1E5EuFpizju00ZypY9WH1nUTS0jrEOwfalhiha1
O3SeW38TTvegMpqpI/L7aviEoMhIRx/z7ITM2h0eAm2Zj3JDgNliIP8NlFmWCxVc10KZ+3q2x6aN
umRASdTCTkeGNHCoxxndeHrUbcnhMdNMR06bkJGr4ZTaxhIAzSyk8o/eM1R2Nx2taGsoG5SIu8SP
/0euTJj6taI6hD29z5Fb2Ej8ouXHdgpTqhE2IlmUad1XCYg2ovcbW0UcIah/bF/oT9KFb2FdaGmk
XvCkQ+JXGkAekcIqvg/fpqtbW9Hz8Z23I2cbFbv64gb5iWdAKDa2b4K22chUYeqaBYoCe0fH7Gym
YaZfWKLPposQRkvM5fWTjwk74HUwB65w18PZBMTWBqjHuP2+pkjbVv2/1C1eXy3e7QblIRCpTuMS
lHKBhA/oLJx1SZedEXXcw/QnsOIEQzr26YgMZJshdP7D9OOJY19HVE6p7CKlTbGOKFMfcQ8PBL+K
s7+V1DiO0CvozjEpLTTbGz2fBFXh3P/uCOVJ5chC0GRw8qFNwxmwVgAJq2UnaYMd566tIsCKY+4l
yb4pZF72IFlxQbp7QMLKzObno1uXIQvJqVL/HTKHzgIIQDYlDTNY+PCNERt5/mvtpA0OtYXbI2Fn
pWjleh83qJSLu622U7sJk4bELAlTtFfa4DM+cv7s/nwGfT7EcHLRhZQI3cQOV+RgjxUf+iPShRFY
yyz+ZoznqhVqikKsECH3rvqFTWxtWht6CnBZIqHxZAlBPpUX0iskBWPeYF4ki4LTfvWhMWQOp6fG
jRyJUDre0XDMf5lkDsgLSAbEpTQcxxv8xTrt/yZvrpTuMJnT1zxvtE6TqtctmmjSCs8oSfglORTz
yd54OPeFFXJ5McN8h/4Bvc65SWzVcicudsrhl4H73UjKvuuvk3RZnwTBd5DkDsEYl2bN7GHRpelv
qc3a/8cqYZFgAObBmJvg6GIZ/gFlW8RJxbpUnGV6kWdmb1n2B/TUu6lc2aGHzPpzz8YV4ZRcH1vA
speUGfqbyvtEU3lw/lngBP4KucBANThbZFXBuwRYBwKirBmL+SBuJU+/ex5sQwXc6RpEP+NElSJN
uAwJeM4MLrWPsrFs4g0scCa7Yr1eAcP1jd+lh0xIGHvLefjTSYujf6G6dDZttBHZaaoSWTHRFlEs
IA3yDbYL88QNVChVgKCcTi7O6sf2vl0llyE7dxrEHmnmgcKVY0xRPWgbuyXW3MStSOgahjJFygPT
3w9Ne3vEmFzV7iKLmuhTfAJS5l+ZAUaoV1KT7D/jzYJWZwNysGPXD1OfD2I7yUJIW02p1sLlAP15
rmIt2si9WiS5De8rqi75EJC0EbFrN8kNjTqw/WCJJFMV5ar0EgE9DxL9pbIiEsjsX/+CZM6Jnybv
qLt5NjaHxtA7spJQfrdEh3yzc3znLkQzBA4tupLp151Y2Yzd4OmiQPnRncO5K7RBY+1XlbtwRj6o
iclPeQknPxBMepMQ7OrXvaMIbvvRWF38mZNzusreWsfotv2yxbKRWYiaQ06DS717cZvkkp/QqW9u
mRZ07sdRvsRmyaw19czzNncFOPDyXWKMRSML9B0aOzFjymvVloenIyhhp44t168wf2RoI71OuL9q
XuO0on92QwH9TZeLLRuU0s1x3fhRTxpa3Wv0mrk7ITV0D/lWOhVpPVs4B1auV3ngKBO1093j4mtS
8dcy03evNWWHfxlNSHL9v0+SmhLowgpOhdwE3EpcSVNxU792DCMUWvCpzZqlymuvJPVty8Cm8ubJ
mC1hGkbQpM2HeN1ul4ciT6e9KQgwQ6CBpEkgkjyEMg9ywcMvBO0R85RC/P+oGsiOBVHJFYUnLZqc
YjcVQTfySk5PktKfCDjZNTC3v/x79tu0f1dK2RVNfzD9GzLe9Z21WS4A53aLRRwx+P7z+zi1oCa0
pOxaJgu289ACikx4smUpD4HnJz/LWrT+uN/NQM+7R8r1bD8yA6cu/NPs7js4pRLmoXE8K+9RbNrv
cDbuZnKAubjg5DqE6z/KmqdXSUdidOT85Hgz2yrpsok8U06sSubO/TJ/jsk7xK4tA0TMgaDJpata
jvWKEnKlxXvC0bSTjQOcqzonTSRNvesYJ6K6AQh1ll3spgTMap40DIE8OKb2YLjnPtgK7zJAmB00
zwfgjVdrBUV5/kOs8fr1GXwj3cr6n0EUWnGFrgzDRYdYcZ0FOHQAbIpjsqtQxxQ31ya9b/CY0h76
kvAeeAsqQuytq8vmxQKCqSVoF3LuAfDa2uH8NNTP48Y9GwJPWDXW/HhFzfbeaUJM74RcExlS0kvk
g9bsUWaSmahK9spc2/nCqs6GYRgbgPsn1kDD5uWVdmjSAIDL9SP89v72iNf7RADe1qpf+z3jfVdf
U1jRd8D9f61g+g3dK2tAFkbaywVewOgjRSUXR3wSx2I/S9zjviVYMulem7u7X+vRl2rqhqNAKj5G
8IyQTBCu3MHwMomerthisU/16WROSXO32Hh7oALcf03jRS4brgCs2P6pNRRHVJV43Go7kdVIQdzI
j0y+6Y3gd1dRcrQ54pZgDO7+FW/mxlcfHrTRaINQcD6BpkgzK+Hl56XteRHEkGs/k7k9SjxWsS/E
ANgexouyeDkQ/LmsoLt2nyakhd8bo6P7wknf0orE+S95Xy6gWw1qnQayOk1QjNtWWq3EqsE0LOAT
vXFdP1i2kHS0HmJgividTCqogyirJiw53wPHs4zAYNqxHk64YlmO7y43hP3ejMeFih0bBGdFfixi
JsVn7l0nAlwvgescKfuYYdMvp+gxgJ/EDFCZd5nVkgUBhteI5Xd/rpB77xLbBCGdrhxrdoZ8iKj3
ZFKhMBFZOYSifcPT/J1sXRTP1tAGq0K875Wx52ZKWf7NC5ejwsCr7f638GxBz5hO+7TetKDycuKw
Hkri0cskIRdSWTZb01M/13feILhdJb1nSQ6GM4ioMeyyCj577EB/o2g4UwPJ2Ipu+Qs24wxpUaSI
rHl/mx9Qwp932hMryb9L0VVIX+LTnDmtHsWbYPQBkxlqHg8AvaBFf8rJiCSheR1LSqGGa1tgyZc1
rFnqe+Z61BtzZHnrj3iQ2EwN0VXn08FCGoeEahQ2u9e78Vgsq39O8u88cUMc60QBsRyc6CgYzTM9
bRArUVi7cg3cJ9AObF0f2MNJ31SmVG5pKa7cYooxu2slivhAfKPBVye6uXrKHDtI2ytoLXo8Yr3L
FG6zvhBplmawr4V/0NFdyiNyCWhiAqP7QUpOMboSioAdgGHyjXhFAuGVeQ0CDQIgkEUrE+9FO2Pd
od4a4imc0EuuJtq7jYTVO3gb894wxxcCV36iW6p4W+bOSSxVMLJOWdtkh4mluvPGKAQeNROD3YwV
9kFwRNgae52orDPI8rsC2fPZ8lgMgObBCAo+ykU24o6aZX4627VSQGtRiHqx036IgIoMD51VB/1f
EkZ/+KU6pP6rZ+aPHTVotB41uO0WaAK4rrwybr+1elgUnx6/7eERA4sfZ8QkVXrVUInViCfr3khC
Sbbj+HamjGhu8ATguMPwt45OoLyVi+J//WUtiGB8F4zyUjwNL+PKPP/U/0LnEmXHu5/rxqOPZDYk
im7nTQTjaoVY/JrjwP4piP/iiVbdxHaPDVOa+mD3U5vAmhNR8WbUGltlM8POOuNIamfBQp7G+Md1
9E8IAAYBLmWrDqV4aUxpr9qkRNp7bkZk9KAytOc7QnvANb/Uoan17z/T5yif2+KSLxrAyl23wkKx
VINK0O5SmDyQuD4Tmv8FXtfOsfKJx7ZpZNTOAx3ZS2c9AcisNPr22Vc62AJrIds7royJhkl3fS96
CIYtTLqfvoNfv6T3HmYx2KetzPwlG7YNlpiGrtGcjjTjjx800+uFkwluJiUjzbRau4W9P4cE2Y2Q
fvJT8TgG+8lOVC9j+fzDKDnCJKHz2amlZHzLsZgG5EQOO8jtgVxSaZm/wprRva0GFmI4n7fX0Gcu
rp+JUb1kVbZZ5R0wo4xcvH6vKIc+pwRjx/frdDuRHbdN5gKL58CGe83oLfgCjygR0HBIYCJss1yd
EcGtWfIwuD5dsCX37xVCDDSuHEW9YIAJ1HLsBtXD8NVYxpjg/5sEqzKg/1Ra1mJv0lPwg8U3igjZ
tg9pZJvsP+7m3w+wfg+tA5U6O70xO5kTYcyXg4wZIvikc/KAcJ4hp2MLKQWyyImqrIrAiJBZaOeS
9ecu/fF0JQfL8eKEa629l9sfdgGtnYZpe40kKOcA1n6KbOAxn0vB3x28KMJkDFklpxYflX0u+ZGK
9SYKgnTsasJYHazOEaUKD6vNz0Eo3GpdJe2Sx/xhLzhZGxX9+FPj4av4OstU5HgUW4p5imqk9CQe
kXz27je+hYPqyk/lnqOish5xU16SlgyVBYgK40fsM8wMUEoQL+XQbTkEq1iL0Ii0hx1xsa3jgzIa
hOywza4kN6D/TyUDRp4r01IFjDa9BB1Ab99sqKLbgKASVpE024WQffXjq+fgEr00P5/cvjfz21DD
h+i3NrZZF8QTJXTeJIplhySoC1dgtvIru/dD/RL9egPKo1R8i9dl4DRObCszcgjwrC5fZYY4PvE4
NEnbDWNCV+xIk5acKVjPzz7weF/KTSEXVBpTHqKuElGegIiwqmSHOas4EpAFoK/cx3pF3BR9/zxh
RNKzkYyawAVzPkEFZDEnnIf3tzngIgUAxJ/VFzoEOeq6V613gokPx7tHkugMYwTMi6vjDvg2S487
OPsskh82D+giJDuGC8GUgoHWHfeTyViMUXJzZXVhCsWOUlWGWFolBUnwp0fPunXxZEK93GS2Nbhq
TrTn/U+3YlZXMFbIqZ/GParP9zSql+no2t37aQPeIkfj+l5uP90ZL0EKK0/xCsD0fg6WjyNe6b9/
ccyAMVOXSM5E06SEDGlxytuHQvXXEdujpESlxZwykpjnOrjCsEBDK9dv+X93Q5QJph7aLa4FH0tg
mK3e9RO6AzgJ314gNZyePF3q+PxV86w/jisMVS+0KIHXHup/SaNJnzKaWX6gcm1YnqQ/4SOc+ysC
VV609SsFBzpFPdjnzyJEkEfjzItJ3Ex56nvdyTMJb4VYUexpfMbfTvh13RZ4GBM3eBPjqhjo/HEo
D7fPsVp5pwj/JLmBR+wOzRA28SI8metdNoOeSZAUEEjIQJ9J0VNYbSz+Yhkn5N0mkIT/k771s8wd
bA/AMsCaDQwtxG3ixjPQA+dQ2gaKdZAUA65M7h0P+7LiDpBAMkFiDX1ql9PQtQUNy5ghj6xt3KSi
paf1ItI+bLlyuOQ8NQVQ/Zdgq4DllW1iUj91RVYncVVPeNvLKJ56hklclR9aN9WhFCurktasfCuD
Jk6kFxIIuvoxIakIjFlZWKeDyBrp/mG6Zxj5o+FJ8CE7FdDZU3Ss5WBN4iEMu1o/Rn74IHMSYUXC
uA0U6srxNrw1bulLzVEnSSLTWJoDFg03IO1mIokRU1bbPS0M2k9El8qWfTNH5/hhfVO+z3/xZLlQ
XkNEhYOxql0PItSLBV/jFv/WEuIMUHooKGKoxdcJL9ocjw33UJSji0p906gjVIr8H49gViXVF/KL
JpTpa/2AUikhsrtaLtLM9lH+UulLQX6GPK3Re8N5IxkT63YnLwVjCG3U5b7xB8+3L3aJ6UOkheKi
+1/T3aWI7jIQZOxJI+WaRZ+k03MbFveei7ob+DuspQ5hgfgsyZn0usgfv4feCcRkv4ty/e3w6WlL
/AAoG23c0UY9d6r1lOl2Kwc6bYkUm659s0csMVW5LJC1h4qbgdNf1dsAPB3oZGdg+Bl2tgc76Kpp
m6EmoqCc71fp+8QDjWXzaCSx/tx/qMzm6Ua17UqWexhsGmbCvo4I9X2PSE/R0Su3MP74w2UxgJ2k
W2PGqisC7L6md5FrzD6pVB3LwoUC+7JcF8G16SlQ6D2UBEAsFo9e0v0WimscWxHdIBGLTs+otDP0
5fJBll+rEHuGZgLCFIsuopCBq/4qn3RgBbe6RACwfVxXjzI3KgDx/Qm/X3oc6rtCLtufTQSeZNk0
rUlcO70tw1exxoBv7iJet5qJirzl/Szte09YZb9NgeAOqMIyMMaZD4nz1zSYKrpUlEqnoqKYUSVw
jMQsUxgscfvlojtymZpRRyqjI0Ej0/Vwv6EIQ1ZlUBns7DSXKLKfARdz0dR2ekdeaLSE5GrpzudH
K1xwvxdiA1HKfa+W9U8SFjg7wLTfvgzzMhogmFRWs9CuPkGwU7m+UpyJ+KK6mKbezp/UpYlTkF85
rYjfXRCIXB+jApB7NGVGUdCAh5r/wbmAOAGUFhL7H9dpDv4mV8nIVsqKtGT8SEFdAhwnuFuPcCYk
kHSOO2pXF/sH/f39uhnvnICCEtx+/iZGeP+rqLUVlH6YT/casUGBTS3dOZBlTlveabKyhj7GCdct
7H/ccct6fkZrUzGhAhSJ8z2LNq4bXDQG3GsOuAnG8N1SCyz8Fg48LZGqQabjJ7bK70r4/77h94Dr
b6YJoToGPfRFanb+Led2V9R+ssstMl/JS59LZN1v/CyJguF7+aAyVqzRRpLkhCTLaRU6DVgKW1Oo
Dc+krYgN6tuycdyFd/4FdRQlnXt4OGGmeShiHxk3LlydRKj17oaJ7ZHjZajAYgjEMBpF7MFO9l9F
FdDO0Y4r4JkLK9+dKgWao7F+J/qVx6Kg8FO5UAc31a0mTBz3FK3UWUUAHrhNrGMAGZMWHAfDxEkX
feWdlQIL0HzgG0DDNItK7ZcryeiQLMdqIeEI/azaja6lcKCENVVEdm1hKYdzoYpqcC7kvVT5LuaT
mE4DOXGVm2yFxxLwqRUKZuD3uwvnZ3hhu8VwwDivy8OYcm4F+K3sZg5DmUHzY4s0Nn2UHSN9UzMj
CQfOwNeFcJHBIg8Sqo0KUgwaGo4/e+6ug+nu15Xe46Lj+bHzWta7MeRsEp+E4SFvXi+fkqvw84yj
hIQDLS3H5sW0k/NnGBHb+Fqp8ZGqsR9NZAK+N3hzdRCE3+QDSud7HIeA1sxfNS7ZL9JiO/mVyxk8
gP+iXiLbpglMCnYovwTGjJZaBEF9cTp7EY5/6bNM5vefGfj8A/ugQb11BK9uHuT2vnqaIGugWS2L
yI/h5a+80YAnzrCsUFnMob9xhdFpKt1ZNgFKpV1FoAnsmHZGQwdL6/T2d35wRGXUdNRPoqnDT7MO
k1g04Q/CZWK/R3kBBg6VLJt1iTtpZ62DgCbMjs/OeRCWPrw/tdKM/BTbeXVk9aaEFvHiVK6inaTM
l7jUBj+c0goU+GcBUdRwzQB3SaXmMeQsQu9iJwLWhaGjXBDjMrLPyCAPEox517V+QpzkY5G87pyH
JMd7hlPB9ov+JPh32Iyogt5XiHabcrQXAE4x/syWcdROTAxqGXCuupJz020kRpqy9N65jwbYLtBC
xDzVtCJyEb/3p+JYPHHPZ4wT/QWuymvMwVo53XBIJkOPlOrnb5fGMAfl1052ZFIp8mGqNzBP3P7a
q5kB+t8c9TZfZsbmVb5G33k1enIYCHI30u7jj7ocTNUya5Mjh/W0kLylR8SLd2akTIjDisGFZcrj
2wYk247TDngWkgeHJR4VoYaK4xYZya/httz6AnIX8YDfGassBRGxMGfjtRJM7sXVvrQyAxi1wIMl
g2mr9P5ryWk+cgv0Lb95zWUT4Mxb3TZscb7f9+89FgGcebPMbjIeghqFFyYhP3AGombnHxzBLCq1
xsxPEloUJZvT2g8RuhGybgp85gHB4Id25/Q+mo7ewOxKe+K1N03ej8kbMBofSmAsk8TiI0AoydrG
Lrw3rHkko+eplsp4+WcBvo/Y9ScIoIRi6ctuYj5SHGfYVeBVFbT7yXnNCNwsIyv0T21iiXzVA8bg
bazGpA7mCgnaH6bV5pRIDDJSzFQTopt26X4e3o/nZG7TntDbAG2apIDhhO8Kr1VMujOTSI9gv4Gp
U/Oc7nNANXRWuPbUJRx4L1PWt6n9hZrmhM7y1V47+DE4PUb9V5aLT7e9ZcVbUN7lYH2nPThMQN8E
1JvfiXfYwKf1RtJbWp7fQitqwXTnQvfpl/X5U+va11AK/TR0GmcTNaGyMxX7I+idFSJTmAB2/kJj
ikK50tuFhGDANbTaCb3uiiqDQtI5MqwU0T2wIVV3Ib7obz5yen+gGrGTwEuoXu8279wzSLZLuwX/
i17fWiSjEoXvuBHzj3Nz7ocxfLHCuu+ei8OzYtYfA3akHfJYFiB4S4POUXvy89wuCFiGzJQ0wk6P
uSjm7IlVKiFzarcbTRdufnf3qeN0IcnmK6CixWsnXMNH7iZYqNIOG7gJ96F5h3CkKU5DkeFJgfz+
4lovpHkuGqaZ1ewsg4X3Df3G9x0ceGIo4GSiw47UWmCRoajR0gKXYeHttqpTi+Gpzvkt1ExMKhXJ
oMuJ9eYvXcYopJXL+CccVAFGgnxZX2exDvUBcMV29dgAqKo106b0ftGdpHLqu4SHLnA4UzylUx3v
eP1Ai4Z2QYfylcY+RpbWVktDeskYy+hfOpH/gdk4NXQcGEdtrUvKUTZsTo3G4Kqh137wxr+0p7yv
oLXWcQJM/GU8F1e1jh4Ryy93exJB6ldS9LI8T9jiJa2397WOJ9vQvadv6HvE+Govpzy5eak6SbOr
i/ZvpH5KeDrhsqH99+De+fnIipKvTh5GmJGjs1U7LiGHwtmzcjPWHO99O4SWZEFfVGGL1gr1FOwe
yIEZybUlpocjhOt8Gf9J4dbREkexyNbBh+aWJlekBa4WL99+3ADMNdwAxPZx/YwIFYgfRJ/moivU
FvsSo10j7cWCS1izvuf0KMC7ZODu2izYtALBu1ReDOQUjaqFUHMrSBnK4vyJ1M+xWa4cP9v3kU9R
FTs5ym4wuelw4/YK/dGTF8zwwqMRrf6DVD/ilV/mhTRzPu56XZesVwYo2AHEoWkdaNIJuBh+XSX9
iLDXwIv+dPXGuJmrHsnI3JkT2eRToRiF/tWNZuQBDz0ZWmvUt7Yot6StlnJ0CZ0JO5TizPLCapj+
0+7NptG/jQwhMpiDdvdJ3MyHKB1QBWogUp+TY0n7DPf9FhZqXQ4EDe7zUMcL+Lo1OKGnN44yIXkR
ipNJRcsRcYuDFWHOIMY6KVyqiOy+DJk2aAjjO54tBNR6H1WrHbnjQCRjJK64PNpcWWqa81JT689Y
8LWsa6vqEXrm7bqc3EghRrc4t7CPPX6cc0/+JC62RtlyBWEkZ7ooqNLzmw0xc8RrVewGKITlGMn+
935W+bAHPqpWxHuzN5VaXQG5kVX8C2Niu4rsb31LpYViDVvV/OWQWq2TujJo3lP7gtJo0Pax6Ljv
aw04UNcrLRmcOFbvEHSu7+zGHeRtJ0YeP5ti0mb+mbniFHs6/rRATor3ToV2YODiLBSS8RkSXqZi
E3n01J1RvDaY9RM6vs6wVHLex3Lc6sAifK+Ve/c7eRrsuNbBu3sXMOdC5SbuN/Lb03BOyObD3aHv
O+HpcoPMhwm63v3kv+5hLVEoK0GQuFxNWJp2ehN5US9fJv9e95M+iHaEybXLEYg5byWlz4vXUJUU
3Bm3UOpupKOsWjlOmuHL3QeLKiQwSR4iIGKdZ+XbRAfmjzRAyYLPVx278MbaT7qCvC6fhsTYmsgK
mCXf2bFCY2QEkuLOtF9ZBUOT63Ku+bqmCjIms1WUDiyxEIaRf1YJgEjM7mHqp8e0ZWGewIfXjfQZ
p6P9tuFYNaLTa/A8oyWjuu24Te7eFFRGUrPdKAyVD9uAXgi5qSQms83bYtaPwPb0lW3wzjAnYgRS
GwEuTvEMOuEY6JaIBlshwQRvHRiWtGRxPbrEqp2aeMCcRt48PKnak2yGtMW8A2xU6vICUDWKEwqa
8th0FZz3dqrYOZBZwkad+tfIK/JrSYjuZxYN6vt2xU+K5vOWAg/xr5Q6X9kZm+XoVqC5BfL9Eic2
2+UHb785FuNcQzqDxo2jhHpF+dZ9CBZoEip3PiJ3u/IkeY+oWUsmvYBGlY1yfVYfUFLNMoB6tcs2
xq14BxDvl1Dk91XGgMiGMjoQbUrokMSr0bo84kp7fsKeE9FzgnFNLhxFgan+NHkbl1s/aaUk26vG
Andq8ZObBnnvF7Mfhvdq4JE0ddW33MHNziPgPdz/apwIfcq8j60N3azASaI984s02WHT67Ejxv++
aCSBUckRPN+JlUNH0DTxZWf3hf7JI9JmJ0SHRt7csmNJAnlVwCG5i8Y+ETwrRQR4f9PAjFCP4v+v
mAwvbZo+VeuByKc+0OmgEcAoDJpTdjj/9gn1/ZRUlIa1Kmsb8XZ+bU9psGx+lPaSI0Hldv9IOyoe
L287rnfc1Rea51T1aOmc4LPi1WT549BV25r31LZv2eUsJdV/QVFHP3zg/LqRgKoG8oW9OSCoh86l
VzXd30PmC6zN2q6dbY0gOSOKLxzmhbcapiAPREvdCciZIcelvse8hF3FBdwoNaF71hzhLNOppqBs
K+Ho12mG367huruU2jupc1vLKpDAkUc1LcmLtxScUflSlEE+29xIB9vr6GvllOpMhES9M2GzYhJn
gQfT1Ne1M2SsCtrxZnfkilQFINt11bSl8dkKd/iOExB1cCYVPl+MYJEeKLUZ094jgfE2B9abCT2W
apYFsU0AP5g1QtBe0Ls17+9QERNVfOxTY5dinal6v4dwaDQtG4jKsFxtdM8IUmq2me2PavQO0hf9
aWTLWZmfiwGJoL+7KOLePyxMo9TJJVpKT2vICtyloPFQ/3NexLdanMt7FMLZvjwnaEdpUwssxQ2N
xNUyVyiOq4gumENaW3PhTL4iZIF7Q2N0edBBur62+USvoUpTflebGOROr9f/GhoAksZU5tLgWx1W
aAJ2CSpm20wvkh+13zALlJl1dNOy4+pj+CJ9oyZwXyN2nZgrH148Su0ZrhNPgRtNZa17q7JNX7Qy
XP75bOkj44fAIZcbmspxKQac+PbK2mEBRiCzsWx6J7T6yvGjU1ELINfwbNpLKMW4QJONx/o5Vkhr
gTjMKkU6Rs2Xc3Ybhd2kDTFirFFi7kUr6z0s0KkDqv4NX0f9orCxAH37E4GMXd1ySvg/U+t4OFxm
G/zg6NEGP/CC27/jHkuRuXYwQLiuFhK5owsb6Z7+s8hDrGtJ8VoTDEkI6j4R/Pb+ugeKIa9g32NP
DsEwaVJKpHrgQ91B61v5KDEbfQb2MpiJlDVW0bNl8TBPgROlzyv6+4AWBeBo86rRonwe05OcE49c
TiaZtpbpnKa0mK3vETt8wre0HkYLIvdyPfjEOEbzzOMJEs00MJrR11eiSrazFef5m05ci1Xl0Wol
/OM4QnTmgC26a6appj++W89SuaM3KpmQuT904CcGu/ULqL3kx/ygyy0UKqtYbxDtdhhdqc3ZUmAi
/dKtGrwvqEpmU59U0AaCdRVHsvWQfEOzZtde8j4RZEJybRTncYvuDGZ2ecYzdXEvia15SczX9AHs
eYeiKuTIjQ//5nkUiyAFSX0JvM0ym5JQJa/GYhsh5MS6rNMFLhyuLXvR+Or8rLb549dFWf2cxHQx
aG3FT7YzR51wLdLCKbFAGTwDKgPsZLYqDOOwoGigLMaa+60PCZxEvrVmbZtxi8EG4f/A/32WPpFy
7DFIVAOVXmnqh9DX9I6ejN3EPNYB4xZvUguQobL4M6SJjWFzM9uyL2a2OtBrLj6EM8zWI6Z81WBR
VVmowMHm0gsTNBn/A3rU+KnWV7w5v2SLL3FFRgrdU9+F04p82gOKfpSY96wsKd2fTB5KPpBah+Uq
9O6fr694X10ED5Dyg05XIPs54NEHX3A/yiQZwdQ/DDQArb3FsZgvRpADU27TBF342NDgmi41hWLB
ogMeEvEIgws+N6iqfxpWJjJVaQQTgx05cbQL8QTVI5hZOwKp2hNK5VT5+RWWki/Ivl8FW3nd/Mxa
To+UfzoZLMWyNMpC7uFlBqL2TH1uA+JKQYnGaF0g2OsOLYUZF7mw5Gi1lB/SbGqNxbNftrQpSzhS
RUuI/z/KKKyCUUHwSlX/A150eHDCaYuHI0EcQ/4aCoxMK9vk4xe6KM/IffJKHBFj0ZFlpiTn5cF+
ENHmvvI86hoOj37XAjWnetUcBsolK9qgSQT/ivWl9ctsXdAyCV+ZOqyGs6gNeIWU+iUwAaboZ4xz
umrp58Po5mWzuSswCQ6/6rWT+3uhrUEeK8yURAf7R+UF/0k3/iK8THtwNt85iRIP6LSxMMknmkpJ
wibzk0ZlFFZYBs6yYLPowKjQaXcj4snon5HbkahYlYJVsjloGBuH6gP0Gu+8AuQZVNl68YPkTGpN
W4bQxHFCXQgbS5osJjE44ee5fgwWus+aS+Z/tE4jnE6obX2b7qAyIVwwisNJ8/NU18l3qL/xwbON
Vdv8ueFQ3aO/f/VG144QNjMNxVhvW7H9nF70HGdYb0FiP0wM3hQcz8ZahrmQRvrxKg9S1lOqc0yv
Xt/5tzeF5BUXsPp/CLOzJTCVum9WM73xGScqnUXJBCd3dAiR3UUzn7MCyaA3xR3VFFMYydKikuAr
BIHtPaNvx4Jf2cAnTOGSvoUeTyxHYGAZ/EF2CC+0BzUi/JpvkFH9wANSuJ/yJ/dJtBSVUC/llk02
v3x4M9877gpUBDDPnASAjxBtyOPTSyl/MBJ9dXG7KPwfyWyoXXHlb3M83piCLUkAlx30RbhQKvBX
35QnQLCu3q6h0RjePHnOno5h4wFIM9UuGs3rorcvhSkFz2ALrsSw+/IZSphchG1unGb1HYEFwSj7
H7qa6h00S735QNjO9u6xa9UnuuSnZK3V/oCkly1FVTbKZlmMG+W1+fvlEm2t0eXSVSBM6Zl9k2xX
WDETjrC13NQBIGrQOHVkQSSh/crIhxjPEOvDoBCO8lUxG8yZKoiemar+BjMp9jqbKCmgfJxJniWr
Yqw9jLQSg9qrnMIgiZpZ+EnGu8y1VRmK8l5d1Wf9VruLd1NgRod07je/LkB97MablnGSAFujv/Aj
QnFZ+FdM0vfbdpqHntUxZb0kQ4wQ+r25eUoauyuYSOCUTcKg/9HNKwITmIKAEW3rxCFgdQvOWsm3
em1xjf6IaAOjGWFtW1mq9s0SDPfQ8WXlLczzNtN8a0fmJLQ1qefupOv9w/r2I5Vl3+9W8wMMrgml
KYdQyuzSa12Fb/b/22k2Q/WFYwo0+wRETEiESx+PdQgcAOlYy03TY1yx9/lVZV6amaUgBgp9y0En
XybIF2m2H8QmGG+WzA9g+BMX/GdiabIbCv2oDeMbFDziWspvPWZQsohlVtlMANvcy6szWuLDLYae
glxM1GVlvcEGLs+hNy743wLZHUD8Dcf00q1711BS9qWDnGSOx1biPv5vSef02/qsd4X6XzoDTkSU
jaavxs37mKXN9pN49kGnc+dEqvteDqkNMq96dQ5QQy+6cMzmbRWoUWOG3vGUVuP2jYUdOc0Vhb8B
2pbKuoRFtN9H8u6C6ol30EA51BNIa7XnmlMfze7pTMd3n3p8j5TtoOniYvP37scd+suvR2v+Q78g
31l1xbIrimXV83EAevbsZ67GQa/3tJABSJWh3oqC06Mtqe8ZJa5WJ9T9SxKIOPalDwZGXN5AK1fs
Amn2iOC8/YyjmxtHLOUNRZ0vMcx3ZkqsVumFxPRQF91paCKj39p7+Ifh6yI/rN9T/py+r7vb33+M
+0DBYLBGOOirSlmPMiuMSljFHLHS+4QxelMwCLkYxWHNQC9y0CQuzL57zkYLnh6Qrsjn1ZvEiSiY
sV076zLnoyOMz/nR713g7oppSYo1b4LjA6eugGBS5KReIc6Hgphj4GGNmMkwfloevL2Glrap/T17
HXdRWIlZNA5QZLV8Pmba5edLSZa3Qn14DWZcN4x6ynjyf7pdG+ZcSorK+Qhonr0w2jW599RHa5TP
+xI107onS0+5wm0Eg9pz6VHaONCoOSADMICtffLwS7i8RhnhfhC3qa35GelrO2xmaHbznLFhMa7h
NOnBkupRyc9U7PIA5Ark+LMjMnfL5Ss/O8X68o9s0Q7lMlA+x8mC0muwlBxMq8IcT7lX0dXsOLyx
1+SPQ8CQqHii5AoStcjKHXb41Vo3R0M2UWvcGDwfCszDSv9RAASfCJ9mcjo4whrGHX8HSH8Lknn7
sMF9ne5HphOqFis74kXDNz5ilQ5FsJSbn5WivO0+gGjglnWMjqLWy8ySzB+EXHJ4CxGBi5SJAeUn
KFP84P9aABc+QOq/cJeUI6yZ/tL+GnpraZgPxXclfNuBXzxxD9Q6njOPT0c4tnfqrpYoZLSjGZXZ
T9JFWV8XuBzrdtPjxrcae9h/968+VAjFrsu0EYz2/EWoHGAStLdd6d5t2gcfN2d80PoBPl/BoPMC
CG/N1+ir0yKsbheY9ILsL8ZQSc/445EIVA2en4VU8gvTvbBo16n1l/jfILll5Y/BK0vebXQjv1Ag
pQH70xQr/BzWzn9+B7l2gnKEx25pfqsYylp4D8Rcykd3VhjMo4sZ4pQtAUeTtM/i0eI+E2K6GMOt
gxZGJbFvGIz0D4SkNGphLOz13JhSf6ZQVMeIzfDyYC0ubIItDTjWVn31ZVvcg4dW5YgCBA0887aL
tsjGlGFYK56F8tKMrsMx0Y6abfH/tBY8rDMOxo9HnKnZQUlGDLZzAIUmEt3z9eBDiuEOjNNxWU4h
bllQsgeNBtRDcB/IMR3Jw249+2eNjV9NmGftp81IdOjLeLZRKh3Tb4Ope2PBavk0wM2puDhtNDDA
7zRM9oU/xWTdjDE0W2mIDQeHbpE7W4rFOfBLofU1WNdyAV6C0vJYg3uSGnv9KQ6rKuLkZ3JG0S4A
hXZK+ZNvaoHF+7RuN4XjLVhP/dRcNfkDN4uvLb5mv1kDS79b5yRYZ4uTcmZ4XiNcIWkjqu2EG5dm
HrvkwGcf7nkS/Ao0uKLOnhgRxQnXlA+QvJHUVE4MVwE50/68omU4lkneOXD60QgWkV3tO4KnmkR9
tDh/Nvr+2nJLXKZInOXhew0F10Ouj7PYrFJzfYU9GRqMg+Qvh/t1yaHSPTOHL7+dOyxcAdetHvLE
JMdKj4+VL4AfSO2ynbL+wFs5mtorijPoJY4Zj63ifqHWWkT2qiKxYykVus9lFaxnTd3z2yHjqM64
AjNAnwpABtP0A5MWJW2SrEQZ4fwbJe87kTsaylmSc90IsvhWvesqS8yTxl45Qs2kuvr4iqlaiYst
P7lmYiPfpjKjkHbLf6T9XpQ9jYYtwrUD0yB0+is1IqE2tG5ePrjAkovr6pmUYiJZB4Jirlcns9+U
fnHj8mqJhDnGWs4PD5bSJH2SYVPq09DccjIr6c6L3DGTbKPUXsrQJkT1tIwmJh/4smO27hD8V3w1
rIeWaUR10mQrtPD26+FtEQfYQqB/l76e53HhJAotbx5xBvm5j7qgr/VpBsEPazQ+S11xQ8SPTeaw
aQfrCQS6N9SxpGT0PfvbXOwkcGKemz7bEalTNQyy0UJ5sY8RSrfffd3cMIEwxvwbyIPka+cOYnV1
/njh2BnEXoP3/XFnegP9aonis7i6BRgSDwPIIX2qvLsI8kT3Qv5nNfDN/ggtTjf1YVJDd/TpBp6B
s5o37FNuwxJnrs4AIE/N2qU8OJ5nsKAlxasu7i6qy9YmMrGSZ4LMT3jQby8rLHVMl6ShukMvQEMH
P8GU6az/0IR/9ejPgwPAlU+mp1gFOP7IRXf3yVIRHIVXCaDKUU6pc9sj1+g//KHf1CBzCoC/JGyw
815zcVq1Xks2REsoxR8gGAHnZ3onrHX5s9s/DVowJUqhETvbPNfRSa+StRN4VVza2/yr0kL+Wx5b
/6JDglVrmpStexS3SvtgYTEnO2j5bAuEEnXomxRN+D2+e5OQa0Iv6k/5WEejkbszL955nLAsvcwv
7m5t0cMAX7mZzHcTZJiA0jXsjT4glfe0OlKxxfltXuMli2SqJtfPHHzWYh4IvW5megmgfxMYX4Ti
q8SOpWpRvbHZKO6nM7c1WAk2/uHxZfsL8z/iwYoynRTsuRnPTV4BaN08GNGP4lAkf6fnbMfMlK1N
5g8RzZm+eqDkd4vIQoER2eLnF3lTGyRP/nR+HphOHXB7G1Wz/VnrPMyKV1hvFB5H0f8qLfIpyU5l
VbPaAqBEw11eP2MzjKZcDXIGD0bqKx7Y1REDXYkfydxHWctH2GNwwdsxqMefUhCeRcZlGkplaBFi
BQHBwcgAcc+Etvlug0PIzW+SomQ7pKoXdPfFlI/yaIv2ZhgNLhvkOrvD9/AtmAKbcGeYEVGvKGI4
jVkSu5+754ic3RkpRdAoMTfMYhzKlXI3oJTvaaBrpb0cPuCJuY1kwNFv/TiQpvTs9Geks3WFxPPM
gBvDwTfRmWi4E9vptTqMyWeoEjI4MZprfTDqvPhPKm8FYxHtkHzP3o5GjMGnVd47nUjHV51LSLvM
6nCg8zZuBuCJYnQgxU2x7oaOJxb6OfkR4dwbtkdIQi8YKw39geywzNmZNvoxiSiMbRPeDT2HR6IJ
2zZe9fjABkcWN5qY2f0z7ow7od0QAECtFmcAVY3QNqcsUxaBlKcuxAmtFfANU3cqqwnTvipw9sIg
RLc60KnkPAQ8lia6HBrShpiF6ISq3H23R7s6Tp8FqBbimEv0T3zHaIsi9qJuRtn8+FQSnQYOhNUP
ZQAPBkoQbWncQ11bVNntzXo4dewDw1S6U4rkOmQW/uRu6/iFzabzikQ2LZy6hgB/zVkY4pKwkZS2
DAKQGsej4gGGlZTN99SRW2muCuN7CCuAYC2oAcwZMXIW/AAkRs1ZSSFTpkTcN0rxOW+tf4CEL2am
muIdblNCKf1wKJ4IBa5HxW2/0TNsaYkC0a/jVyZCaHgSpnFmbWxizq6/pkyT1AiAlp/8l4dwtrnI
HuUiLcnSaSqsV0eEl7V/NjjG/1GSZAvqTHthboKeYhC7IpQAVHAFF4PuyOloU2pA1GrWTN+sRtmU
5/cWZcwT342SQ002XR/t7E96ViVQZYWRK1sqc83t15dQPB/yOuYeWzK/cQto/pCOlV15niGfXUcH
a83F51iuZmTk/R01vjz8gcTZOygJimU+mtJSG+QtSqFXkp6MxRy0ubHOZ9pqF5j9U01hIY/n32xD
y8f4uvYN415g3Xhx2rjVi4SBGcx9nCXTOsLr+7sYdZNzsW1EO+/vOV+uD0HnbfHW6Ve88QYr/X3N
DrZC+bpBwmmhvcr3FH6U2U50HfNtOsowJ3vqeklSn7HXwO0X+NhraL2xqzCyoEvgn15okEK8qILw
uA7mK59caZxrfLx6gNfl1fHQuwgQWjKL2yoDK6LbAPbKnMwoGxvZvIpwgwF06kzTwFGfJx+eSB6V
ijNw4GkSbJkvSt9dwKu7FzOTAlQi/bncHUa8zDszlXU21rKCh7SXT4eOXYKWWXP1h+8lWjyQaq76
GGRW85mET2QOi0K34U4VE75YU2QE0Voj0I2w09w+GL+EPWaUecF+49DTRfAAUNB7E1TsX8qe+nkd
gGdlPcN9pFB54vlVQk8P8LwkCrhjNptoglE7ZLuTiKoI8jTbex0Katkqu40EE75BcRFecEa5F/5y
aYinHdPgHwyoqhyrpHRTrhl1SquCLGSbO+2F9dpBzD5gpHETEpwM9qnHqng4T9C0l8mPCeEEf3RC
B78fwDUoNKtyQtWlNrehO+q/YDtnej86Zx/tgsuldIt2GvrTlej34O/v0b+HDfj2nis+4+5T0oR1
P0wmBnCNBftujqThN5XHdmUeHncwGKjDbu8PFvArlVa84gKg7fyTuXVXNryMzdKHorEHN9EXj+zA
ieU7PKeOeEkDcG/m/0m8nlxuWSgzdPnQWAuLRqLUX7CMQyf5SYYEDIU9xqO7qN+YjxGioiShAJ6I
BHFtDL3bCwGuo7ZLVpo3qjmJhx9ojf/T1Em7o8oAex+T7YBvzE6HNkkT+wrx+ZVeYFZzf4p7ljUG
H9MuKjxUKogU6l0ngSu/Qbggik0KmiwuXqybHcsBZKj3P/BXyMvGQXm8G+P6vBah9y5b75TiwJ8/
//JdRM96CJ1/1taP9QOUEL/oIHmqD37YnDtXc3rUbyhB6qRkUyNLW32rzdTZPxK68zMc0OoFpKQ+
a/xGExhd0ZUzQeZBGJHwETpVwimITOGrIxYV0mp2Y2kvHZOPyM9YG07vcRftCTuMORH87LFCD1Iq
S1OuUd+VYtuIOLxlN72IqOJ9Gt0tJNsYxoLS+WnaFROx7L46TESCHGSZl7GFbRirWyGVws7fdmQC
wCEXNgr7GlAsS+iwd3Z2iPjOxES3J9sbOJ6Mu23LUOlVFDKTGX+5B23GYUH8pvwDY/NbmiuN5GUD
Mx0yDAGdKNnGytaep6XZNaTIy792ZtFxik6wWmj9i79ESy0DQLgyuUxx+69vyXAwnpvByMnhVGsc
GdSACWWVsaF5txM4u+T9nkclFOZNiZEpQK2UZM/hgU1ztCoSc0BWpjMhyLtYWu5H1xYeAkR2JqZD
6kiCfuQvv5LtFGmJrhO1CN/kZbQsk5QQDJm+iZNUFmYdiya//XmmFE5BAL8VfdJtgzIjlsJKWg+5
LXTykORxmyfcyeRr1Xajk1lAC1bJhcdbPkvAr1auCm6xTaAmuroS2OUn1g83VmC0Bls7QbbXxODo
Ee92k/qFP/2lnyeJVymp4Em0clEWZSS8NGCDmIihVsCWZ+Img2Kqsx+QdgtVQXpgVqhyM+12mUP+
7LcId1hTGFuLMyE4lSrnmzx4K2sJ1c/oRWf0axbhXdDJuLTOOah3ygp9mPfzXCnsrw7TDhIViJ0Q
kncnaXl8IQb0Cz2DCziGMns6Cq8eozpjVgFFzxN9jvO1DUqcJ5i+98diID7pmeEqu05u8gbVYMQe
ruR9bI0kcvwL7rqgH9IBgc83nNVlaRDBk/JhM6FIdZ9I30sDCcVYN61tDe6rbFqbIgX6kw7iEATJ
GqINewOD1U6Y5oxWkJ0C2DdKEOexQDhGE+Dtqpozm3WIwi9JSFZKpB4X7+lAZ+DjgXcoDCfSxbJv
mJeZNwQv5fxIc1001rCRisQ8EOLGeuCI7Wsb/2vD1Hxf37zxtY6Syhd8oxwtH11+SXlcHq8FuEMZ
f6JwOHlxNT4/st8ry47JcE3jFGlK3XAkFmEJl1baeigAxxWBQDkBGN4XZ0HUOLNNZIA0HHBh8jVS
579g9fx1OrSdAK52Way/tomKb11tIgemBBwuzTFbMTyEX2G7ScWE+ygMFT/qH/c67xP31lLGIoUu
dDNXt3fmVD+kBG7lj0CF9sekga8iCo3HGXFppt3tJ1KlK9Ln2E/NbmVcfJTSjFGoM9XQObWlt3qh
ggUkPDvDnjvmZpmYbyxbjVERvfxpnS2XDm3sTHzKckAqDfqq8E7ML+iDbwkIvdrbP1QvQs17aCvU
iyHyeW9pwckK4xa1TOE19WUIwI6ijTZo2KYXKmZTMYVrWBwSofjDiM8mDVwpo86dM00IEep6YGtS
DiBYWsIZjbc/eCDJqN7b3mRAJL9TwzVYIVWwXtqfhVlBf0Yh6Mo0L6n8XUn76lpFlf8TjiQ2XDfM
qlpfcz4Oq8wsVKz5GNbr+z0jzrbyPm0hrL0dFF/K0ix2v/R/AEqiVCnf4gExAkdX/NhIJB1FpWLm
1QTf6/GxydwM0oPlgTfatwLZG72fvwLsGuAqry4f6iqUC/JG0nVF8JnQFJ01DnJ2oTLlPF2kIb8/
/qw0no/2yHU1F8Z0ZTBbs0bze1Q+M2/7scrjDf3B1vZS29MpsYVYtm8vd8PeK+x9lE/QPHFN/ue5
JY22zlFZUWexovRA3hMytPyr+H/RAX1A2Xxvp0noRTMZggNwIQ37L2hP9Cd6K4XfNVm6wjClIjt/
iTOYNMRCse0i7mfdZyiNerDrgA/6Xb46QhfDshrDsOcjlRMycRybjBjxQJwAFaPfX8ZnFm/6sG+R
4NQM08UmGqIhK0x45TNQeqKHGK8qo99dIAnCQKq+G8hBtKPndxTC/WP+/TGWJzLVIaAGd2RCIc4Z
i1yxH6uuVawWM077wWcaPyk4haW31THyQ6RazQO/XKmeA6sFtSpRbvKn6c/nwREwx0H/wuxl3XYn
AMh50DrRWsZjNqLMfXgkuRp7AzxIA1mVFLUxvA6aPWTclHshppXvIHDcURvLM4zf/SYWWMP8oZgE
1slF6rJfOvdImMHweXpZ/EfQDdcCbC7K+eOLM9GttukSNFus1emXZ2zRhEu88Qk1iJQox5LSRwYj
qZWt7l3wdSPEYiPYbAaEFwykm+1EtWmZMS/8DL7qF6q8j+NKNV1j5eQ6WsumvZ+hvJrHniCkXbP5
N8TXWCYrEmd+f8b6UDRjW63yoRCdR4OpGL65BenVlb7Q6731GuLWa2eZxq7N6Pd9xA/45ToopRt4
1bLRU/u6Nle4O0qbz25U/4iH4YoqkAiCZkm59JjO2qfjR7KoV2g1XB3jf54LR6DaqJGdDwEEOxgB
X4CvlUvQh3qAwBAeHVHx/hpF1WVUNeJ/KmfGtkXBWQEpZnxIe2ZJ1oJGd+ovQRYc8jkjwtcbJ+YN
8URcnxQftOMedqdjpmIYacvr+526x06n2VBuTjmWQpmtg1PMPDShvT5zfxeWIdujtcbpLfQzpmA7
luxNpmBy0iWGWQ9N6aepv4NlaI6Xi3tpQidTOFq3tlv0+4n3++L4Etw4iUNQEErQE2o9cJucYGEQ
xVWOuFH/86+Ehvk4RhvlWQRkVQM8qwhh8a35m39XX5j2/DXqBCF2oDsC6q8nNaQkRUvSxdryfUmW
3+F84M7KPtyT5Zam8gRAVZ0qF8BecMZD7IRqCI+qkeMTJqrZkSh8tsVJYEoncfAXiaViO3L6guLe
QXPYqFE6EVabj9jQj/AE4UnOldXB3Recp+05lYwWPDLEo+yvvdYXwoAZmn6fVciK6BtB0apOsBuh
V6Gpk0IElhLWZbGKZIXbASjoFhZdzNxk5XS4QI+uERvyiU0YvArbvCWy9bRZ5Z5nWI/yox/SMKx3
ej2xyuuwDyj9HXzQsDJCQXKGk0ozwakwYe7HJ5Ob1QvjjrIr6XpXSjCuC/WejaahrfQFNV1UsK1Z
tn6AQ1h1qG8Fm18a9lznh8SA+0B5jyL3phK7Gut044mHIz7O85CMX/RZhXQZ7PHdFaSnaCkIvnyF
MEkHxV6V+M4MPRIxl2TYa7UNMAQuJStbMBtrjJlgtXj4g2REfXx9aS13mnHGK+tqZJJUUVkIHjqr
CBOYgbo/yiIZyPKKRwcE/thS0AZjZdOi8Fwl4/mre6DtYxH88aKTLqVIZMFPEmt/MBo7BErISqSp
lASO0DQyurHip/MhPu7RqU/qhtf/LK8d+aeurRMdNTVui47G07mz8XpXxNeTMvNhlrf5/hmnXOXA
JWlKUkpfm0dalpA+NDcTeszYvIC/pnAZWisiCxcAp0MHZP1vtuKGtwppjaEWzdo5h9JHEKQtswZ4
g1hAj4qvZtFPoQG7BKx2FxqWTfGolQh65ZP+VgBf30o00vT+B9DOmdpLRtoOX8IVaI8mmYHmDi/y
dcxcjtOyAbDDnQmQUNUl8SqpWntI6JzJyzCy087cCBblVoxIIImQShlNK9+7O8kjqhk4aDBRTMC8
/yZymaIy0BMpS/HaJnXZqT/Ihju5fIHuVm69vrJyUHgk+0j6vTIzbUKq9nFcc+4DgGWjETWobA32
s7btPqE+JH8eK5svxMUpqWpiBgKvqu+EjPxeDADuFhvEJGO5+oBsKvG91p0/+jikkIcsRH9C77lu
DcT5CvarW6895u4Vco954Rv8VYGaXMoMsA+KWkYa4X0yASml5P9y/dyXz2mqid8hHprXAFH16poW
cQaOvthZM0LfX17Zy2ZtVmCXX0keClgdYZ0EKr+eIWmOVJUldtYaagvL6rOrwLNTvrZP7pn/1gLL
VaaMUOiJverf1RkN+5IqJM9EP2lVBVTI7LndsyI8qdAy5LI1MRgqk0dc5gZpct2iBv7JQ1DAFlLu
SZeTRX07ZfIdD6brX4FsF+8SJkZXvVsqnQhoPo3CkvE8mH65odQ2iWEGn6kiYPO0CWv5Ml0/wQLZ
cPnoeMFpkvTWvh1r62oNSsLDF+Qln8AkCcDldMXu0ulUgOi1Imf6WtQFJ7IZI5NAtzuw4PgOb3+I
w/FnMAaMUklwwHKkKUOoOy/rzi2X2xEZ0a/CUPenja/cbHKYvFp8t06Ceh/B7PDK/KaY1gMNZY99
sv1LUtTvsTRY1zWEuOpZlbTGzG47vfJaZBQILoT/bq+lsu4nhET5Q2eQd2MgUR4qPd92PxpZeRS7
ygFe6Oad6GjveQNxQIaqGHMXpWZgo3VA0HCohuwupU6OFM6Yqw5Ru1ICGKS2AQvBwwIaC+NDpMin
tkkZcXXoI5CChN3sM6YtVQA4unDymDnH7y1NL4qKdizNpOVVEFZoJnIVjGANNrC2R01kL52BN4uP
UTR8yZtomn09cceAbTJwxR3VMfS3hxUI4chXuaLtInxlNNP4DYGeoKXx8FcHXepbkUHKOJAUafdS
0F5epc5S3XaJnEldKXoGLPL0hj9LBFBC0W3AgskLwY1ZbktREhq/mIlKb6nGwldC1qtiVBkRK7WO
GSLSad2s7DFWiZWnpscjWB/eBQqFmtHpwOTsGw6l/66w8xjFN5kGAWSFExwSGPpD+aPWCHIqsvDJ
nAIN8UTmfqtUA86OMYf1hRl2f5AABAH0Nnem0kM+X/aooY3QBav+vrjYnw9zj9zlEblh8xTRmmq9
zy95LUs3bVn67vE924h57x2wsv/I3mMiaS4CIhenmDDMSTO408N2m5aQq45f8anhVVJyz1JTmpvM
XXII6Ekp9tu4/VuNWCR/O+O3lr3JbCj/B55MP+2hZAkqOdBEjxfIKhclmujKV3ZTZfY9i80ogNep
Y3doUUNKbsTZ6NsUr0HHrQF9JKEWhYBZuS2gi28zJPtnbTi7dyxwwG1hLB5NWRUCHBJyjlPyQEoI
0+GT73XoatEQNnSHWgAKORtPVJmRwDZsUUEw5hQx+5fSJZ9BxKnJ6W/yD864u+lKvAaHPmubOSze
G0cAx6C3ZkqUrn1hjFWWCG8DPkOUNSkbUu2X9X6HKAbBxjpI3yye0g3jwG95ZwCKtJq0nKE7SIwq
hTlkXmSoYzfcdK7hka5agaKrFji4qEtWKp2H2+aL3JjPGOZ0h351elgkRrf/yX8XF8s1AXNfZDQh
SRPeJS/rjOu/oHiNjQLQ0XV6y8ZvXUKVhLDC+8yBCCEMjquz4VI4LebPYyQkqTJ62skpSpm3XxCA
ZPSEjjplXsF96sguOn2fJRiUqrvNJegZUH5WVZCDFPQZHuZaaAyGmgacpNyjnFKH0ZI1lqnslNxU
uFR1mvisDKo14WAUve+pXTZZ8fSoAjExCIz8afFkqHUEvCV3JdAFAHlDp5Aj3xwfEmDgxFcWQd4C
WPx9pEbMhY/T+ynhxcOX7/niz7EnFQ9wumVNXxD2v/8taYGqucJlgkmfcHmIcBy3VmgPGg0PvGXK
gCaB84lfn5JN50fjTqVt5UdLjLwAeLmGobP/rngT397D7qNy0HHA88Fjgmijcw+xqs2G4lndKYE4
osOUdn6RCOQ5V4mJmj+jNR7IhBd1oRUPmnHJhCCp9VUZKJ4FPp6pU9fFc/kcl0j57tt3AH3C0Vgi
bluFBHKaTUNV08/miMcNxJzHnSSI9zbzoMYHe3Ra6pPk0ATz/gNtk6lUgum9jyBgW058byG7wdeU
4899W0qIJSPXFc06QNHxPlRyoKOpRkSsd16B/VPzMElxGD2n/PoyxrONV4EHgmxUgPWqRqkEtgfK
fotCHp/5wOrnhRHD3ywXGxGm8pLXzqSNPLUnSTMSA7jwVUy9WZCHJXMwuEO9GMn7MkdoKcWMaCky
uPioCqt11sL9ELvk5uhLg3RAkBLYyE2bQAqiTTnhqxp+bKLqPv7euiy7xzM+Ko1NQXhGk8v7Mg5s
2JPRiMNL73777Pl5tOYyIZf4nAE2pnQbjz6hK0kQ/8C1U8CLLwxlOQ26zxGgutTksRBXcXjZ+Kuu
6Ua/CDKa1y4GYXPkKW6flzI3GAt2X/1jLgyhP2qJ6EgGpLcrwjZaYFpLdeN6YIdDnnMOdm2kq+Kc
y7XoPktiGy4Uh9uFdPs+sp7ounFmbB2H6uXbNk5b0pToUT5+zJese6GNnhX4QwDHysh89iZhMy9V
FilGeQZpRsKxJ5e44F1wH5443joku3kiW233IWhZGl9L9Ly3cXGoynp0Ip+50q5urxV8T0D6o+i+
Tz92AB5jWT954BMw2Nxu84uQWf5XkDhXl/ZtljntLX7BVROBezP3V5EtKtpLdEGqZPxRj3+M6uFi
2ylqfkycz4UKvYxpAQMs177kA9a8gsAWrcGCf1QaHbMWeAK0gObPUpFNXHL7mx7MsBR5vvQpNuZi
OqpEORpzXLTzEHOID0zlAMceYt9X0D5TcOAnoNUyxQCqmUvMxoEwu6xPdFLeE3H52sAfB099FzN3
ev85G5g5XZzJuRq+eXgmSbw+LFtMtciTSMDqZ2Saw2J1fCTaNbKWzKjVcY3m2N7KWhHpL2/9oDZo
TEIzrpRm7SRAn4bT9ZGHBYexRUnahm5Deeinf8W+jJ8ZpXsNv/EZbyRsy0qb1Y+sE3s+w9smty+M
vUc7nrspfZbehtW9yy9ybrt7dSxEP9t8QZQciY9kuCGSfLe5rh4UsY3rMTTi+F589pvGWwMKam0b
7kwwgCi/AuR4szWZzl7RSyAVnldIGNXC5aIYthy4oq+cYdRWRN09fzrpAFPY0QXs6EjUEmSNM2rK
l8BadXTWSOxxj98goiJfyquTDFaqk4DB6V7PLUqhYr8ZaCVVPvB/0T98r+tHfsmhbwK2o/ZqWpqN
Y81tiw4SilVcW3pu64FfzPHUQjIwUwGfOkpwQPgfvwI2qTpaISnQtlVxpgciRGo1EMDjtx/x6hV4
OoXm/cKvuj9/jDrOyS9EL0WhxI/Vbac6aIBSfqwEWqbqIrvTuFE/DSqNy7EroQbxa/iECBzQ/Zg4
cxzsQ+1K+fiJk9TkPQZ3zoT9NklIoNEytyBlq0s0UnDF1tICb3ZLcRvSYGsag7ImQtF9EsyzhJdF
zNMl+YkvVrFAHLzEJKE8qsQF968If4lpXbidxjgAFx683OI5TX/n2FUclFhs1I0RVd79AvvmQQ2z
o4xC7GonMWu6KjWaJSVmIvVfSjfnuC+8nXnGMgHFrUKHqVXCQ6W5bmTD4lqSK97bPHlZgsXYvbic
Kkqqa3YBURhlUlQkf4KjJLg/AAB12viVKtaZSMxTrZ8ABx1VRfDW7FQK/27Qe2scvXPkk5wDC8Fn
cKJI+GPQqEjUKe/likN42W2QDQkDnF7BUb3R990dwPVWXOpBU6oKHsddAL0j9UQHOVvQVblSc7Qg
u9+/YhE5faSzS9F//P6n7H1VbOwRdPq4ShRtBTlt7vAQfJrZL64YCaCRSxoc4IaF0ChqHQabpLz/
ZRUIfgnthAh+oERXIOg5mkHEeto8qfnDNh3Tf8bBdMJdyyN3Ces4GfHQU9C99eM/wyoU4HyK+vxa
CZdv/ysjQjU9pFedP0RN1KMim/Zk7+WF+aW0UKQyjeP1RV+c6NBtbCMHm8xHNc7hGtvdrg/w7r4c
LCAeAiqf3GFb70QkhDAuWWT3bsN1znGOoF3zlP3FvK+PEObimfJxq6SfO3HqbBkkZQ62NejwntV8
7RnmBdaRVK3B6rG03XA49ebZYNBwwvlhrXecftRjUmEitFY/dOj/en39ejVteXUAMllundY657rc
rna9/7T/3g81IW030UYvtgtUcJhPG8IEYbg/rCLOq6NWxxMOmKcuLW/x08QuV9qtIkBSi8e0QpqT
6IJ2i0xVUibOcxPcfy0gylEl+fUYeelpYPzKqUYv+rj4qSZOTJxarTeOX8QoV9ATCVC6Tf1CZ3/+
QNlreewBUpai5tPH5U7aOu8j/Cd7f5G0173gYy08COoHJRecDeb3hqBsT7n0ssNVixXM8kAW64Su
S9hpCD9qTmuUUDe/503WyOGxfsSHKcgofenx8Ztn3dGyzMzmUhrlS7snkBKsPI1z8JUGZva0S38w
eGCF5pWMCXeZrlqkxRIkd/228zN4TdIK4txbFnCySsFBspykwvMuaca/0TL1q8CjJ6lJx2+T1GMb
DZl6webwLAausUAMR1yTa0aYiFUK/eg0DK4Ez2qaAj8JjLnuB7BvyMpOedoLzjgby2rQu5OWZaGo
vaWBVvdhAc5xkm+SaAGKbZ2tOQkHyXNrvyi/TTxL6b8SJ7nacu7ub1aA49SCMtW44lhcRqUf6ueo
76AU3xX+qkMXeMArDeZ0dP7Pw/kJQMXSg9Gq13rBz58M+REq+s+ew2SZG5Q1BcuwsHQS8XuPbLMu
U52sReAktNzrG+pXcQvoEHImTxV4yiOkKd1jivngKk0iK+Vzp9bctU08rHcRPh3b/cEKPKYuExoe
51HNDkmK2VcUjhKkA2TtEvan2SBPbrkRMsalZpee8KkYrkKcgM6x5KmpzHN1maRxrUJf77/GvpMu
/gljx7+9o+ratv/n8vbO390lWXgROycd1NLS+uQKvZByxRcJtYSyEyGI+gMt9TO0lW2N5bjNG0Jj
LcNqH2cbIdIe4XQPOoOAfWGKXyygqDnMXEDdZFdETawLaIBFju/EaJryJ8PjFfVVyDYoG/rib+B3
jjuZalVWMYfWvAMbLLWOn1zomZHFmwC1XoKHCZKie62/LY2IP235hJzVzwMu9OaSuW0CkpxATEa+
VNcPo9SB+14wAk9s1kMVAbdfvR5cPfneZUimG/X5vJ8bxlNfy0yZnYyekrnXwDvxfLD1TH0GUjdm
gC2lmPF98Cr+ZYMH2MVPvz3jKAa40JV0ThGzjcmNZ65qBvC5XKdcpOjzcK9nFtcEVDvv1CA70PdA
RC49TBSwEl/ewK51IFMGes4OlntrkID9hcoVMTm5u/z+MlbI4764XZayjmJSML0azfi73s0lQ8b/
fKMq/u/NuEpdw3VnMsovBk+RJKgXuqso618V7d++iF0CGLfhPf31Y+nKkDX06I37mp4lt90wjS/R
kNDv48rubW4IgoJtdOBGvZ9Z2vG31QwL03arEcup+BEylxpKeTD80ubDUGrwTtFEYPHiTMa08giX
G+gwSyrm7tJrVUoWupecoO8tsySECG23sYnVqAD7Uirp4GfVRHuJPSoX8MwKYoLT9A5QuWmQQXVO
H6hP+aGa8h1dN7fWoDQw2VTIYZU1UYkUXA9M/zEid3THUh801cYF039SAnYj2m2f3oDyWPtU37Lm
LyIl3M7Zba8f11Kivyvcy4eI1inqaJFi/ArIcaNIWYUfCuDuzT0JHQ0YAK4CqFOV063m0mZcG63I
Rv6usNXXKuaWrRj/vZNdMdGGNG9iu/852cchS4Ft70ZmSsow/JFtxixhe28kZow0a30DCuLZ3wq0
x0poLucmoaAppzyh2SocNmf3BypsJUpHPHaDNSwmxGzsGXge8o61fMzyn49A8vlck+Q9td6YJpUG
Sr0wxBnKZRJiKdc/5jSOM3InwixkjsL9cbsvuf+iSoldX+OwxQfSSZPGJaWdobrWVoktzdqFiAjF
mbhUum3xrvKC6uj+34D2ynn4gIn4qBDsuGt5QuXJJK8zqnaUDnpztGs+Qi6gGbkpPng6c0cevoOF
UgJXEU64QNPL3ncuWwtvWONmPxizeW5IGB/UQ8QqLPJkZ0RKepBMVoJcazAN3aNIK9/hCvBfUhpc
4s6R4eYS5o5Ap8uGtp1WPIbSrCDWK14/F3AQutlp3PGO4eDpZXZ2/7ekDdNJp1aMlKmc4VHeBoqc
y6l+Cqsm6RN5X7OQ3v+DGuJlRJ5wozxWIUcAvluCC0h2B5U6ltTlLQb8V4tzIgjbP27fn4qaictX
jI51P/ee4YwMcm+WZPVdBJtqIJ0QAukqzXVSrWFxnmQWX40f/GjzY7xKYTOXiczsKLKSlhpkQRPL
MjMtWaWLxd1ecfcN2KXNgQ+PsdWUaeM4Evopo3Yo4pKy3BttXn6T7AE3LMcmf7/4UYZ3mdl3xdtw
cfgJXts7PYn49DGCTgCijMan79kVdlaV2u/d9tYli/5enbWyFHx305dgQUK/LmlQbbrp5r828E16
bmbv1Y882Rav76ICCPLRt43a+XF1rJTo8vZgHL4wdmO9tuRgbXLwWnojkQTwQtpyiqirApaFRd4b
Kkz7Lk7IoGmOP6AGeDi1iGJ1SaKD1y0d4IwhkijFuD8SpzTqlB5F3kcNd1RLEtQu8BBtrKzYGoE4
YS/0FbLQlr05MuAzWoR258gC4DF2/XpKvahKOZ7u5EKdEYM2u7AWki+z3MIBw7rdgKCUIdW0g4CU
iTc+ibhkTTSqOF/FdBBPTjo5gFgDG7wzPBsUVDczQE2jQVg3JmJPjKy/5w6CfIRWsoUyX7GnjJWH
bT+HiwlAxGaG//ONaHvEAPWwFgi1H/dgdEnHLieXkAQH9Q5kYIX02WBeKuloWmYfbJcraFtt1Wn8
DtpRjOh6dweg5wuUGmXNJtlpWGa9EF0HPN6b06HQdVyJSz7rfg2muSEabSzjaQXDAmkHz7F3mpyu
DJZ8WnUnxtATIXgFityKxCHKMDUkT+MjIpY/dG5w9a25J5q+62Bc9lreqw5fhjxeiXQia5X9JkK4
dQMO7G1T//w7ugOBhiSsffsvijQBvAQoSCTnH3d4/6Zc816c/ZT56iMuVUSwgnkDHEDS0hc/zFxb
J55Yk3mQOBrGV02/4/knRQzdnzyK4y6JEskkKt+pEaFNkmkenIXCv8OoGlyzfX0NxXdFRbiiFSak
K5WSMktmmbEgeFEWlpBaAxfeUGIBTQAhxEhO4CLhefz+4YLZC07EVfT1boUkbdluM+A5+KOHiDzw
lgDleApYc+kJeSjpdsU95icl0smyKuywI13/+/59twGOPANc2Df5H9uPv73kD/j+IvC9ZcdEiNuA
w2/2fk7wgs/n6Bu2swyiWYGibij3m14kfrFhaDvlPWH2aqNaTMkDn+HBS7h0TdWv7PzYfkCib6jh
0dW3PfkSuXHvrd3tEvYJf6S7ZudPBrdEHTEmu5NKr2FIyN+oqq/d5m0uWpZtWK3ot84FjVcFcDUL
XgdTnlbOFMp2QTciaZ+NwNVlTkQq0C6Df6G75jyTCU1Ze54cTYGGxvVxy1eXHnCUX60ca1cqB+Cm
c9cThCe+pedgifcATA1/n0mOc22v3mFU1vUCZu8k6sUEWVOM8dhbXcKXfaXDsFUX9FEDju+JAAbU
JUb8Nf4MB1WmlRqZBOz/6+DzgRIttXwR3JUkXzQr3neDmcdBgPGgS5+Lo8teNlXE0/ImSEGuSafO
lH6XltDKCzWBwGXm05tli8JpvXHXc1nHv1xhVvOD2O8gmTxFl19iZ3k1n2LWbezsoSER/6PyuWQl
xhKzg0SGFl/yFdhStRg/XetWtrmGzCbKqUJngYTEhiisywW/pKsRF+ACHfa46k6uqB2aJwV0avpS
nOBoJ2Kp1cWEA+wXkmMKQJbqidkNJ4oRi5AszvU6+dbuoT8Cix5EbXEgt89Qyi7bkq/RMXKlI4FU
yJm3WqGAZ/T28ugP3ta8QctE5tAnxu4GEDonjh+CSFSXIittKVDD7rrYq8LQQup2b3/nmWtngo1S
6Fb96ujn57ANtkxAoO/RZLK3tMcxYM1aVAUmN0a53ZzaOiU0+VdK0B7O+h/y7dNKr1YxNILkn5HL
uZfkYc02H4m1+mMQMyE0RATjtATTQEyxMokJ4+sg8CkD2C+HpuYy0A8/tRiVSfSf3omKMOuDVt5q
IcHlqilDzQ9iPQMC5r4zUun5D+yzLYQccUxX5NpKxsjK2q2IwNrMzhkedzkd82TZCfT4HlqkWiqj
54wA3H4yTrD0ZesB1J3q3nzNi+akV5tvsHHNKIoQpqwyx3772U8yI1gs3Lc55gNPnSoKXuLJltCE
NasCOfEaWkOqJFYjk8WTDXyVCnNmibKaokYkkjnvcR8DigZNynrpm+CpNdpeSI3xT6rFIR9EQGyf
pvLWBdf1hpc4rZ1WZB6YY6X10IZDOoGNuJ3Xy5oVFZUKoL+e9TyN9OQ89GwwNzwm9Ei/dg1Tv77L
VMkdkUZuGBjEmI79zaFL1YiDH0/W355sY2Q5j7UgQUFaio92npZ/dTNLJHpCtGfgCEAlzMm7hKUj
4kb9ood5Af7h0d1IZftS3NEyHF4G6OrJuaoq3duRjY31E+Oevpi9fVjevp2xsXkw3FnD4MIf1Z08
jRzHb5vlRBbI2hWBxgTa2yxASwL7RQf33BZWVDHU0cLt7Hlp/DXubkhJDMshtcZtuLUBvlxFpvWR
bZY/cvMy9E8D7f0SgnQYKKIlrA2MZFu3Lo7sE/rMNp29Fs2OAU0WNu34Cia8GeOGkbuBO3igPFI7
QuI3OYWL2RVBgQ3xH/urnReGUOYQidue24niqLsJrjBU6gbELVbXZ4RuAZEDhOQZ06LNAfKX6jEu
dkXdmUAuG2uX3oJ4bqgYOPQao+MWEJbjtguW6PpkegBb7AAY8yxvaJ7TpLzQp6gX2RJC3iZMGhcI
g3fCMwtq5Bwxb4QGLoo5CNVq7jE5B6Pi6cD6XP7aWrMDDf69bOVWpSXYNj9OjcmzsfvYyxyciDR4
1tUDNVUv0G9QT5fAacxH6oo43QLWteUo4YM6cjrKwsjz/MN2XPcUUIvSFsQnONAbT8EsFE58Ylsr
CIHeSGlLbou6bmy/DnM2uS9xLvEYlvtLVTUWPtk/BajvNNXMlcO+1UZxf/2+UImGKLhPcTewgecR
H2XZzeR1pj0v14wcHV84q47Z3Qgid8QAMg+A2zA48kQkEtcDbyzYsW7nFvpQh0FrfHLBXyoiaKvT
a6ajgSOC8zpgmc1aA2rqQ3AvAlkYNsu/s0wxte6HOL7G7soOXXYbwOew6UW/X+b49GpibsTM714V
g1w5nAUR9+2QENUjMm6b5xXnfwXJALWnknxO7NKNzMS8FCxL4huf7WfSmzbmLnXo7DQ0b2192adg
lQB81a7/BVhlsFODsIQnLUOs5QTKbH/89hdthU+VS931KUMoolX8RI9TyErrmEVvxUiAkPYQfj01
2f9Q1BAlSMw7XPsv0MoSGuM/Vix7/2IZmPc671U1WFJ51jJK2lh7pAc6xHMIhyftv/5rvkTVyTiF
bQoG6JPyRYOQ2WW9coNJsBTsKXvROhWYuWTQarUj/eUtXgELgmsS8fY/lGyWbryrdsFAraGEpUkt
0QlLLMaXJ3EFjUmjmqg1pQSnYLmbWR3Rz7NznD1ShwSljxNOFRoFmgYX2JIyVh2Q2yUygDG/+a/g
LnC222qyTbEUnLyKIQeFHGKEnaC9Ib7TRGOz1KnxkHjsQckz3fOr9EzhbDn/hAX+id6UwxWfDJ2A
FlvYfRO0Eqz2jx74538wD6zrfn/xPaQu50hDOO1IwDdID8BAyKpr0LfzjLE7pVpBZGIDAOjabBrM
BcrDvZ3K41l2SnqzlEzZGvTh3rLlvYVNEt1XLPg2dbGFKLmHZ4/2jGRG/JoYGaHPCqRoUEtC4SYB
LaCiGYMQFdibjMvPyUBqfnzTEk1CjEb4diExdjzrfu8Su2Fg06BwmL8LRkrPXRuXiGgCh/1zNdRc
cw/AHYGhxTVqkLlakTCCbL7StoThj9AssbYbleS/YXvLMon3ramDthdq7xAZh9XRj0zvtC9RN1hv
aPZ4A/fSox16y9SHRpUZfosnOICZrh8LhYv5oY1nNz7onUBv3IjqYqtG5dTrXYFQee0i7r/wnBMV
lBpwFSDsZbPpqIR2FjTTlojAif3QBUrCB4wmEfs2m71KVSToiFw6w0B3j+tUoA8TECGoUYYL7LmJ
+xqcubEGOL79toWKsZRL1tET3IiiC06xmKfTSWE06yV1HxIZb9JRuYNAc2lUoY3eEPCxnHy/T4KE
u/5fKZlpB5tNubsgPidAxR3xY3XDGqbwbOZ+gjmnfxeUlS/Hcc/ohgg3GjzfaoGzPhkoIIp4GYDe
IU1w2LYCkSivqWp0r31uO5xXMPheyeLiV9VIpelzqd6Tijj/uyxCtwIIAlUBdBn3D8fPfULm79h1
Vckj5YNITcURbgBBz0KoBvGLi/cdkLwk5rFQUBdgdyocOKnWHtFCK8i7Ep8HNyDG7+lNvmbSiaD8
3/nKYEli5mvKvu7LG83QlAzBIT2w7E9elgUdtmb0DfXQMCG8Waovy1c+9sXl0urq3Wqpi+5OWabN
6sun6iWoSSRoOsoDguoATxneWO70+XHtUOqnHdblh3HAUUwBCSAd7BRZmvTIpHYA1LJh40UxgbuG
YDovFAlc7Xy7CoJlt0qW+LUy+c+Xwk9hbfLgiuCHQUQ30y6tH/U6flffUczKFkqVNUcow847O4D3
m6d2pLk476iQnPrMogVtIZMG0PoEtoLgfIe7BmfLFYrAr1l0yHza/E5o4xnMBvQmIHhduuXAxysR
92kHZ2wSdncap+Pyr8Ut4fXVJCcNVMUoqgQ5qKTRU7C+SkWizzistgzglGOt5bm15gnU4RIkEbMH
WQ3m5QoxuHRZ46FmVTqldN5EHdV68BesyBPJxumvfiQBbGp/cCvP07/iKCviLabGIYqEuoBIHGIu
mIC/zo3hs2ruONoWZnXPLglgEUhBbJh2jJDNIz2fzlFnrTTR7DeHrAZGFyd7ts3tTMqG0LMG6lGp
E9qXr1R3uoHjo2bC3zSnJNLnCpDQCupTf3raJl/hbvSPSTvU8/Xdm6xpR09tKwoKhhTvDzm78t96
XR8NFzcri53S8IR5caWdGoPpoQLm38iKAl7us2X9dE+hmPWzSNqWLgWx8Hx2me3l/6IxcurXWI4g
6PHRieayeP0W8i+0D68J61Aze2/KI0uIqmZLHSfL0stvJHsrVZeMt5NaluED/H0Og4MmO/chchsD
cfkHII1NElJhPbAwD1G6rOMppOXifGXt0ixngaTG/BFwmJcLG+Yl7rqDajUbA7QSFxqEgk51e1Tj
lJwoT49D4WYtaZ86UhjRsOpa2szida2AoZQ07V9K7VANtbL4Oo9LLrCovtvfoQGzWDEIsSQtDphO
B3oy4Sns0GYsj9l8dZB+UwT4PJWAXTBgw4pSgaADbhsyXwxGfuiPRQx7V685W4/aI42vPXZWSl5N
DAFGQAgxxFDJwJ6cHv5lCUX4SO9JzdsjhSO6YVxtHWLPOxMxSWDUXKVL2wyjbFk4UJB5RftPy3NM
6qd+94MWGUG5YEAn2j1DBwLgvoNGjcpBqn9OpdPx7BcsTt3dTJqqqYAcFJZAYM2t+hyNmWZ8kBV4
UNlIGZLo/o8my4VyYsU561spKvv1LCojV0/XcxGZXYNlFZytfMXYgltBZuC2lD+MUUY1qRZHEb+G
/r7aAPkNaRisSRefwpqWIGPCEJyt4lSSHISmUm5jyVdhVh2GaClu5JfQPO3YXBWU0pJdv+IP2se+
8k+RVdr4+YDV4sT7iMTGe4C8e7vFZXklg1Ycf5rvQH/QRjT8/S4xHzANORYZbyOvsZQti1u9bLfJ
ZvfqAG+4dBmSsra4uWVl+E13RnSo/zHUtP8mvfuErliTseQbPIUhsnpquMxt7VrGXIi875SH+XrW
KLusNaYtsvkfyLzRqiakKAJ8FOZSzR0uHLcW0phMBADLZprn5AuzuZhoKASGfIAyNWd+yPehaTm9
aUEYV5WR7la3zAykOXa7puqujl8v8QOjsbPk32JmYzQTZGGblvg3iXNpEHCZWSyJNPSZcQqBbKvk
zQLaW8IG4PhkK3RkhLxkR83bjiytAdm2ONHlIFq2YwWYyySzXXMWEJuxe7/+i2WMIS2CRR6DJVTR
yCNANUhDZdlWqjam6AUfnbWVx3Ql55ktgdHpdw8Boq6BP+qReJ5W2XqFa/n+5eQ5XbG5y8hgRdmV
gtw+pNI3Czocd0ppEuTt+lLX96D+hizF09OX3OtZW/K9YcArWatX45D8VRoEs1VX2Wj+AwbCXYns
OU3gvqTX3Utu5xQ4stnUh++2Th/1jdYBNcwkeVDZp5BWGvDfcoBLwCuCm1qflm9C9CZ9l70CyZ9+
CvmjhTdjdXAhWxPsX6+Jz4ZiW3Y3DLtr7QVPXyZXDPCtQLeOik+mbk74fQ77TyEzExT33M3gR4r4
JXov26EkEqnT6h4mA5mE6+iCuj1LfeFvwLY5uMI+C+BZHelCTH8EQketII8uZTeCwKT3OqV/8VqE
SH/YjvxZJNZmfMtUr3QqwGkb7VVbTLdK8Yj/5H4HtkZkEKX/ziWPU6pRrAgoMc3muZUY1T3PBN8j
1XQ4nBX24qyEy0bmWSUgPm/5UHnE7vJRCRbBpMmPWDkRU+6zJUuH/qb14l4yRKzcpo5geBKxSAey
ZxUot3fOz/Z6ZMol6YevAA+UKx+tEVRD7YXg6/7nAbUedw0axDcGB7Ya6WxHmekRHXozLbP5J+gP
BysMT2p1RSWVrIp3R9t1wfIlKxuHEIO9SsECvMpFe2RC5qCIRX7QyUefB4WvL+UCpqidkruk4/X0
5fDtOue6Y1cVpzo3l0tWulSdAAhQmXtGubsOgs93iTnVzsnkOQxd0EBZMnNpiUC9d50zCIQsoUwF
UdDLgrAzt4hbR513JtzHTBCg0TWPODgyCL7FriqQzjNVh+oFudYcXS3Ua1wpLXo7vhNlcf/YRFK8
R/qLfLWMtADadPLOxwQOOg0eYWsdAmdV0TJM61UMs/YZQkmoMy9gBAbHkRZyvC9aMtEv4UirRuk7
VFaDMT8UzkWeblqd+LSkGsRvTUrU7BE3Lk76/B2D8+JmoS+J74Fv/OSIeR2N+LSljcuraTVnR0zt
M5mwJW7Mg+fY4DE5QwSJPvo4uvINYsL3w66tRTxA43AXQHzJVRKZXgjhMtlaZiAUL2zExnX4avGv
iq1pNR/2Qzb08TQZMlGilc3ic8HCbjPhNhSyb8MQMkH1Wieplbb9omMHDR1rAIre1T15iu5+/3bp
Jn7KNLm/XElw/ep/vYnsYIQ9CdVZaLYkHZeuJh+E5PqR3SGLUG+NwWqz70dvw3siB/Z92F1YA31Y
cDpe9QC2hHEF8iaRVzmSa83Cc27uxUpAzLeY4KmIygvV6iLIs7fViLxVsH/gUiW+E4GzayB1vVrX
Oxx3N66eQ6tA/7HyzymiBbqTVZagGBvKvn6A5SqSPtl9eVYZlp6X3pp4LUAKSgQBve/XDYz50P0D
VXlPjpRkjUn2VdmRA3YepmzW59bS2eLj+FTVwoxkifl0dbVOjEqx7iXRqNHARce+m77/GBcqYFPN
eQM6JCfHEA+nzEI7ShMPEyX0870sUzD+wBPN6OYFCqJfX11KXFe1HlE9zz7imJ3GbYZBDp+sjeeL
YoXoyL5xHUD25h0pH3r3rTOEcw135RMZJfhjlZhlDRrl+YFk5wHbAGLzxjAduoU9luDNgjmquHyU
QRzp0XY2TJqdga7w6Mg7AVSW6Z2G0PfAhXmgBRe9d2CBO/m3n54DkOOnqj/yOjwqwYTQeiGGRAvY
r6Dth8BSrMtWBlGTRT6TjH93wurf4y3B4PwpGAEGG0prwaDNYOOetkwCFUHn8xuYTvsqYwp0RqSW
O7uu3oia79S2XzjO11cHPaQIhRmpvguXezwnizH1MKYubFZH/t10jAEikRqWYTRibQqEzHJAhpwz
qbe0MxGT2SGMDvnyP+1VpXU1acyLZJgOVUGU7vcU8gYXgcwlXjZcjKWgvx04OH3txj2SiqhHlKhu
PMf1p9pmelE3pW1DnoTmC8s0BlMUWPDfovgbIeGcyixr7EbFEXVePmx2Bwioa8Kfx9SHK6K+fW5x
f3nJm4JfTEVnHy+2JhBr4gWXQzAwW/ioUm7RNMWRtL2Dwtk0q1ZU/96ePv9x6lF3d36aH22MUjIi
ADrk+AFjgZvtzYx3vysQqpLMALsWjuo6Bj+qNWnl9RnGN/f7gY6pe4w+2t0SmCf7l5dVxIR5JDsS
14LgsjpI7YMovQQ24c77QuG/d0Jbju46UBhLkJhUhGYd8VvALGkbL0zBRaNtfw+Im4EqNz9G5vlX
hVyEzCqfqU6ueMWEQMwCTocmt9UaB0CSNx79qm6ZjUWUfXlX9espGcoO66/7ghUdy7bI9J79htBA
jImENxtHi9kJ3oP5NeeRYhZdCh+CjyUTiABPMI/qtGZoF8qG0rYDm17uEaPs+qdXXL3twqJM7W95
+XIO90fGRAtHonY+neB4AcFmrgp3/qKkk13plEsIESGg3BAsX+PaS4jr6T2lJGw1zI/a/oSH49I2
L6dr+nZSsvhSX2YMEw20/8LUt5unWgiZ0qXAYd0+LVZXdTryIS7lzZeYje6mu4B6WKRXtXqERVl6
CezrlhkK+kkM6BEmE/5Mkr78RLImzj3FUsTPN9zeqiLIWKZISQ5e70tXgHz24kVt2vtTsyMrJMM0
I06DZU+p15JCYvCG6L7+7El0ldxLO+aKlpDVC5PnlVxDF2PoB/ZMAJNmiqZyuS0p81HeFEa8mHXT
5gypM5LwqKmYkx3eeHdtJJxPpCXwv1AUboO54OSAu9YS7TnepNqwVf1BmqOanqWmHzXgXZTYXbox
R2F2BWMCHcW7+y7Tl1jCcuFMeSUKcjsqiiro9Wxl3nOzF7vkYzt4WtGVcqhffp+6/1g3lHYR/S3/
i9d9xlDUG0kYEx7QfzO1mEy0b+E10L26w67GhOsWm+MwMlCr8lfMK1tkUhlG4EcFWQ440dmPYsvd
uolZojbwg4g+TIhO3uoVgZsIuCDPyJatDLCDAi/vPq+bFxV4wiEGFSoDuqPByJFzmxM5yZcVJ01W
GIyb2uqurYxRsVd8T+O8TOi9us+3d4MAE2LwgpLWpMSOSc3J2KEQ1Lgs+G7vo8HLj1rZlanKetyd
yDhnLpdGmzd3JzcqS7ZtTRfOA4H++uEj1sQs0FAW8X6HaOs/iNYoQjg8NPi/JVxVGAwQC8pBsdtT
xddlTcQW7lUVJdEmw4wMo2zXd2pz4QeBLg/zVJrqsyao3niLHy4CM38GZvS4jj8VWn9tSjRPsg5v
lNwQYA8G43ffRZR5mqweatXh15KOEZwHE1JKzIdwEqDPoUmN6/jcWdVizESSXKR6iBR4g205P1BC
ROjXMW8j8yp8XhVd2nzE8ip9yA9K3vgsEVQg2CAIlrWq1VaLzviJKtDkKDfOrrvruW+/xitOEi3F
tdSRpau/kJgQuLlRm9G1vnt7lBQCoDW0OZcgToqJIi/NqPHZi5Zx3R71OLNkx9cFF1FVq0+0zNPm
Kdd9/JUINQLYTLaNhqOB/+ZggBB8vqdzDzlFxQ6puaSsClvGiF9W/KY8o9W907TH+bIGkLaPQHnj
FXv6MuzJP4UXBekpeAb3q9H942DpBQc78vtC3jigElU5960kO5Nfkpwtfl/p+5HiRvdah7nLWRtO
wIlkkrorPPdLDEprljlXMknITe4GqfoikcOjSoFCBUjZikWjf6hxCDVkh72HcrW30UrP0cqCYImY
9on4cmrB/n5rm4mDBtES2L9LdNSxcf86W/ZVXJj48t7nqSfF+5ZelC9jIoaoM9mFo70gzy+G4sqD
JCVR1e7aTU77PgZBlbpbsuVy+fUbJV7qy6mkKRakHk65gxhvWaVUGYvqokTiwK4WVV4Z+u0j+FVb
/3/2s8G09qnd8f2xFCeSMGHSl1ghPj0uJOz3QAvs9zkupK6116Qe4DoaU77fGpQRQWjuHxCql807
0lttW2Y1ZyiKzDC2fkq12mJn/L7PA8E4HuAfL/p9rEcI4nDJKyqIkYtL8RzRYIXla9w5W6Ui/6Z3
BpqbRPy0wX12XM4n9Q8gusRoT/aYf9EAGDcyXAAIOLvccHkw/bFDA2pmEydcTXIXvoQZ4454PIYs
J/moj8r7FgRA1es30dq1MnBJ6wQroZUW5fPBNufeSMCYGOItmoxCbk5PGARBK3YEynBm36Cm2ooO
bHLjBCNayoAJN3e1GNUmQRTm+HkboVfx4rzzIReR7LiShLgmposRnEthykQxLmxhVDIEY7z+/ypa
9UMkfnkkhA1we/JpgNZMg+5fVb+yz12jLAgMioU7abd9CqkbaJGeezzbe4cdZ49rvci2YSha2hr3
9FEGkWOYM3H+uW3vex2SXpMumXbRjKGAwRoSbGi1gNZx9eQZn/ccPdyHAv847l1NF5LNhL1+7n7+
2VqAHsQSQXSDFbDtjnzAvU0ys/UHcRN2vhAvXQ6gJKJELhh25KFf24EOnFxXFFPYDLU9jmD91QP2
b7xujauTHokMkf/TnEV/kUiIUS+1+CgX1lL1BTDvyEvTuHUkxaXOGhw0bWrir/0ueuXNiQgZ9ddG
/tcW+hUm2h+/GgskBKJjfeunjujaMA86bkR3SWTMnd6kEb1+R9EtihqZa/IavdBrjsv1qVwcG/E0
pIwHVX6LLvWlX8OtRSAHal/4Y+fZZWV3Ud0bHiEy57Ok0GkYDucMwmlEe4exIQLiSPMYRJYg8ExK
rxTIETk7EwKmo/D3Ano7IhClsIYw0VWBnKJvx0LljqcQKINjsDazAWpwczmCRBO03jRfux0sEG0d
0/RxjchC+/Wm6MbO+3RqWOop21aoYMr6jY9DyUGvy3ct9I/hL9eF3MnBpUtuTCZ5+meJ4dudNcXW
26Ct2Fh1/QPuqJ6MQ6A9P6GnRuS7s87pzuoYY0UMwGEKeRaqhyksNbv6YStzfEt5Z2dxgZ0y6s0h
SNHDxoGT6ULsHasvVHIBqkVK6VeaRGEXBc6BKvkG32rtUEJpaFKFQX56UdOfGWmx1K9fe36LmwQb
V3XlsM6oG5LE5hLp7G0vnmDJ7LYJFyrBeQraEKuQe58e5gQzXfRLgHw3iSDU3BT0xenZwa0zQAfq
qj/yakeJKoXsIce3fCfkRf4bFvINDbQzw79GHlnn08cGCdr4L28S+pleZaGbqdML8ODQJ8lUTjPe
yp8RiznMzUtWQZSZPCwT+dpE3ZbsoJeJR69CYloQldrHY7BOujEO2Gi29NZUvCS78l9wslhIzikw
uMqcFct3PUSlWND+1AwTRBDSb0GfEykFfAFhQFCRCEJayEuU/qOLCpjEr0pHE3KFJAmDmTQz8/l8
JrIPh1msNfEhpa9zX1/pTIYEoFl8ZIWxcxh0my3s4ZcXXUi8JZW9eoUceBVALqSumdjpdt0JdjFw
LIkVZnDLKFX76lhHuyyim/HdjjZwezRkbVfYWBH8OtdLW4i6qrCAQertnDd+VLzZfcmD9wnADyBW
3QyCkc//ps9hvyuIK+U/KcSNI9buw/X/CmJgqQd9QnjPlH+M8fLmpUYSj3vQlHXChsqsFi2dXvhg
wmGx1ZrAJ3HLFxhDvXjhLDQkMlOuG5c4+nQ8CEt0/mFsVTDA9df9Po8yTC77salFS5W/GHDuY/Nc
319bDNdLXY9tIaHlbdhLinkLXyFAdPllGRqtjKcHtaXjUNA6uCFr82L7LqXwcoe31mat0rp5PjEd
BcrFaeWpkF0Vcr0Sfx1upc4rJtligxU1G02V9B8EldHaCwpFVHUKws3KJAboHCPzj/OBRLSITHyZ
ZIctgDBACo3URhDJ7hTD0lPDprTIaZAqopYNrHeTpIp9QHd3aB4E5bAHlbK4QeFG7GXPWDsS4N8u
defYyd06k9mxxGsKmSh8bk4fgUramO6IFKmI72fXRGES5ugPpgZFT2OATOkNuz0AtA0Z0+cZJNBj
D44h3PuFS4DppjKIB/0M4s324023TPZcUkmQysopJM3lUbCrRe8aM5qb/f6MmePCYGyJK8UbiDsj
b6vQ1Rgl56zzgxslBfnt1foJxKzItuhPaI6UthSDRKlI2kIT8hLlxIs9KxtzZ5vC/xESnA9GLWEt
4NkPy/ujDmS0dqJ6JueH07lzRA1n9UkpREHwBsmND/HQBOnCsaLuYEMj7fbOT9mlOV/6nNJRyPdU
UeCoe24ENFmbjIRDPE6IvyPYlg57s983Mp9Wmb4BLOWhoHrykS/NJ2bJnZor+hFdd8OQKn4ToMJG
SUfMNEvvZ/WDn5ioKcLVfM9ZvzbnYyl1HK15m+yRkSVeX0NwEsi6wj8fU+dqMcoTWLG2EuKijXaJ
tu//ZzPwKkr8srRza4F6vcpgogBThOLMszTdehx8tVjw/xJEcqVNNJ3/TEd+T9iZxtWfSZr7HNNF
73U2LL3VkqUt+DahCXKjxQHpkUTHUZajCc64ParDMaBcl34SWpbeWhIOatJktwv9VBXFELYnS2Ee
8o36zk6dLy+WejgyFIq2eE3AaIrlotMK39jjDYmar0rMUhCZXiHv+/BRMT/PD3sCKtiAgvIQpiPm
oo/3nXYX2Z7tlHqX3jLfvUxN9qI0yJsNQZV4uDj5yY+U7KSHyJt3jGFB55VBPLDHkFPYUL9OnsWU
T8jH1xLfqREtNQ84NdsrUrrTm2y+hCSELsh+9gHpPKY4ITYKJGbwMCOG/qUej2E6ZSWNvc70j8TU
NUIhuRqjh/dh2PTp/t3hetEMWMxegjn/4I1wdDRiYURZopA6nL42ozLrQPcwK2d4YtsxhXA7Kbcp
drGxdyisV+xWutaBPxddhz/y0dyCyqG8SrnXevJ4kKXqJTgwoTUXp5e0KUz0optGgayQEl+FMJql
cvA4e3hc12P1Pd7y/dMYJ9NRn83vtHxEWWb0FZ1V2FG494q/pXI5D/mdF/6/Wj7zTseqjIZeEZZd
nUT7uaWmVdPPNBd40+QNgk+iZAn/p/pWXgom+xnnXo+wiK24MZ3f2VE0ACrd86AYKaaTPVibcdMj
u1N+cy9OB6rsuNReo8f2Zg3spWfqCfdAAbKF9BzGfmC41/8NkoS2tBIW34wyPHQQP7Ap2JfKxMau
pIZZTf9dn3YRvJmXR5gI2JZ8KhLPHk/AB2yZVb1nW+/qSYw5QeBlIqlwJ/AWbooPsuF6Hyrieiyn
JT6kLt1qtbB8OScMG5IhJAoE39ZVyiH7zSgXes24+njjETU+JPqvMLytDrJzFxiLKfy6ULL/GOIJ
+FkFBGaMVzLOGHgVhhTkqsdUe7nGSsVqo415fZwAf6XtLIWAJcipxe/t6W6b+pGNIr62BFtSQLYo
rSxF3aGCNxpnSxx+GkyJgZckz+MlMEzMBynC9lA2Wz6JJmjw+ZWDWglYBQaJDd4GZwz0arBEASWk
gDOjReHO1gMD1ISVvtP2+sDr7NGtp9jmttZMqjqLpPbKyXkMbbTWh8llvHaHDieWG7erfds6eEUm
uCLnI5uMqAO2VQNRa032HT7q8rJTWUDflHmE53kRoLzIYtWnNmU0dtiPeBDRY21ETIHM5w5Q60Bh
uPMli5OD34Oybxpuq7M6tzpso7XzTbpCWstTEWs+LhadVb9R33oZCKbSeHBMcq3+I+9gXt9tmWyt
lpyYx5Ca/KPUIwGCXKaBI3uA47rkPlVf3lcrhsU0JWHtHtPtXiJV+MczKj7gG/13JFJoTnysmQM/
zVqxbUgeiqiO1BiPXhy/QOnpCbvg3FXnzsr0Il4t/iIzGm23UR+Ncd45l5oPq7nvD8ukpB2VLqL4
8RnXQnJyL2v7zMYY1Bj5+uG0cQAgoBxlML69cOSvVMVqoOhwNr3HlOvoW4B02t276dfUutOhun/G
2rCdFJs4nH3xr7WhwAplL9w6iZI7CwTDdOlc7yH4l+x6k8nqOvlBzvkJbAPfJcFaWkj4Tjvbla8D
Pn73wDpFAa/17HGYNcB79P1rDaqRKrxgW2L3cQw6a4Q57cNiOUNKsLDhngWv4U4iACrVpoHya5T7
wba1mmnfriKnnPBGZs4MC8gp/tQbqb4GtLBLrAyJ6DkCK7/pE3sBe9G2OmS1m65Fm0dsjlM/KfwZ
f6mnm5AVA9I0PHEZ+ZCbTaRvS1QrgQjD+XDnBoJYmjIAxwe+/N/AQuAkqisf5Ioh/LYOINDJLiPS
V0NGQnOSn5RK6ZtGjlnckHzxjxqyjbALNgR3ghHtchHJio7xAm3b1XLAiCj9yCQjl5HWzg+gDYIU
WCYvRRW4vHmi7Qzvh6y/N6PivhyWdObI/SWnC6n43U/8f1m6tRr4Fb1XwBpBTrijjLM7mBsEYeA8
xG4eTLQfxDgAPKbbm7tmS5XSW4a9MX42wet3b8ViSYvjbMXXTaGNIQ75jiNWZ5TnqyR4Agn4kR/I
PWjqg0K6cZ6ajR1W3dXPPH3/n8zou2mNh/hd8ehFJr9PetDNMJHSSFLJ0LnmF/N+4Hu58YokmgXx
MXaY1wZ4Bv1SqfF5xp1k3RIWbu1qKTrHDa5JcBfWx7OI1Q9z71271eCtJKEWHXfU/qARP/6UoGge
Cbb9O/S8QoWoLoHOgTfmCnyt3baonRnctCA4+J6gEZDkvkRj/L21JkvmuI/ssfmTHoF8bLMqKoAe
VH9DJidbIAy2gpu9ZMHAxbtx7u6GcNj2NY9wReHD9RWnkP4dDw8kX1i2dj+lPJVmJ5p+k0JuHqNS
sHBQvnVpu7oK5mAlyGCFjjF+8DPqZ2/JqCl342lGYz7TDof7X7ZKXVSugk4TaEIgwnue/D5/Uhwb
sNWUtILU3ZF9qejpfYcCmq7gNCnJ0K+eh+GEnfUOfSlfxpLzhN9bRrSe0u174eL0ixnlyK8ZeGed
R8dLcNzn9l2HRxmNRrHxNwvM7WMmBkcxgUTeBJmTw0W2u//RtngZdAHqTyJD49egpPyizIt09Prh
e1wP5cShcmWJpSmbL7C3aFv1265BxOAbiprq4f6MyzTt2/cHukYEryL+FKrxsTPxiFnyQcsXs75U
ov6iHKdl0tlUlVZTe02IBY4buoTtM4t1CL7fM17evq7kOhIKqGQT8JIda6lEndUGdVsjSPuHAIqM
VzaHAK7AL+d22SFnjE/urhAfPOMtnYGIuWdi39KF1rJsVNwtC6q9Wgr+0qintdpKHwCjQRxpX/39
mJNJySqQgu7VKTBzz/AYTSCade64Tl81gMY+Q+X1F1lWciKh8uzW5fnNjPvJ1v8TnCgeQmk91l1n
80kbFzYASFPG373WUHZgYAZHxD5ebHRXEi8B33P+DlKYd3lV2ry6huPHosQ9E0ikBjIKc3ksavjW
f0F3S+IoKZBIas+W1M4uZH7u7FMNgH7jzgFMW6nrlwFreKYFQ++cJsMXB+WeDweoVB1q8e9cHwX4
FCruXrurWWwiocydiwwQ5FSEqdONjT9YRPQBoXrBJb0gU0VFAO8yAAivw09L9vUBMCb0QYfKtUxj
hXludFJlKKsoIgoYXMPq0EEqlfQJ3bNTCICYOhdx3xJy1vHPJQ94SqCHcq75hC1AhYVPcY+rvH8Z
aVDufDMcDJwPcfYEd08Fofqk+OZNzaIKygygPLtcbBYYqCq76X48+vGMT5EaNj60zSADlmvl3xKh
7ockqmTOsvKJQc9UJmd9D8o3+xnhnziWSqwWhfBlQI96+I3Ec2kI3hq6TnMouoFnNkEXo+H43kVT
dsZdmuW5SRjLnv/1kph5RFxcgdEWVZ+lP30vxk+xidHftiAdh07WLN4vmOOF6xV2y1IOBK1tyG2L
auZ1k9A+vRNJsDOqLBbBH8AokKq4RpPBRPWxtXp5HSpDisnKFUaFZ1uhOjvp/HtGoneYVFEdoKnx
pEoY9Cjl1zhCg0KlETyuBj/Ybfhjat2A6XOrarubS6Ld9JLbonjCdJq1bobOmDiG7g0cRfMpf6Ow
4VoLIG++jKu7DQynYm8m1BM5XVvHat5RDuMsxki9LB6jriP8IT8PFBWEWZmYhrCVWsrrJzoip4aP
mU+a7/isvD24wwqprSzv0ayJp79SnFZ+EQmLQWBLqwwBTEy7s+1yHr9qj2hL8b7FZ/BGVFQIhYyM
T51hikiKaq6YkMCkmOUFdSMyYp1kImS1DuqjaECJpstpX0YE0tP/OF9BUXUjT5++f9tAmmB0tYeG
/AoPewW6VN38L3toS1ZJSpIfydH87+I7z1WgX7K5BwVh+xbhfU8xWRZCTQHa1i4keVQQ27R6lL91
cTknWrd8Z9xPl4QLQeSZpnkC+CknVen+xWyqh+/pCA6dzUvkwPfeNq7BnWXmLO9d2UVR2VhObP2R
Krg+C68NaKZM1VZcULK6WLSisUAjORDIwtSL9xHtuKtxfuO/7LNbT0owNgYDfYmTgC9RjF5+j5Hb
X4z77TA6/vwx0uWhNnxDm7rnYL3gZU3vGr28H7eKMdygWI7Y21vmAdcNrzqmm8P1R6vnvGNEG9EQ
L2RhDhpermfntfGyPbMBENVD2Ot8BcirexRZi3IzcaPrfAxmyhITt7MhyERIOSpo6qtj6tbnMjZ3
KuRAaKTyIyz4lDdbNnIAhvzI/SVF0uiTgmKUeANK2En2/c6A/0PcJxnamEKSJ0Pi77t+9kX9xxxc
za6BBIRsyqX3q8sclIOUHHrT/WnGjSR6WwDn6Dvd5ix3rHEq9GtdyvPKM+Y0TZIM8YqxRtEawjb8
qjT0TDdoj0YR28AiLfa7DFXrOpH1mVCrXRe8Z3XcAy5u28/0Otufxmfz9cWcWmUTe1fXKsZRPp7m
Gnq11Af9S4urEa852HsXMp0S4qpYwMMe+WJ7A576VwoPGVXNROh7V72MmWeIWeYlF7AoDakjMgR3
4IhPuNi6eengF3+u6wyaAFBN4RLGqfVRnNdz7E2oFgEvLSCq9QVzQiWoRNxjPJQlxQ7nDqB+tWwV
e4qszbntddn2fUPXmnsO7Fveksf2TgPjhHU6smQ13wb0xMNt/5wKPTPnqcvDPf/Q4cj8b55o+cuz
E6r+7OC4Jj2VlQ6b8s92Xh7mzuuEQACuG/TI0ZkfmCDw02oCWYwzDUrwJbXiEudiT+App4PvRwpt
xUjBAmfy9LL+3Gj3ll8j+LqLqTYMV+lvV70MSVHJjbgFMqP7LbLD1NJoPBstMYA7ju3NMre+uNx1
3ZFfx93r2annEzSYyA8k+J9aU00uUhyP2uT8OrV8NGG+EPmkMiskv+rtHofVU59bF89cRSr5g0B6
GtYhi0XwTE46LrTQR9g4DnN0nsQqxY10lEaXizdW/lAZJYn2rlPZAxXPSZTNS8sdATjLqBxgcC2F
s33r+Zu/XIU1XLr66n8+osN2bRT9ANcqUe4VaL82EgtUGiGNkfUd2wD/BIRX8I1evHSEqj2ruhcp
taTSTfq2UVW+Ixly+RzTquLEg7nf9C56YXqSwx4q5mvEd8v3CVZ3ttI9HbKpMXNLJ1F71E1jdLxK
zkKEIgJ1et4w6RUGqHPoCa84qsHNhD216SXhlhC5/kK8kcID2YRwhNRcqTLOFLs+GKRrtZVw1D98
mB96gDmK04zarEFz8ISHWfmwxk7bcgPHKXiHkSHpTDCn6S0vo79bJmWH+htgqDf4B8P6fGJlJdJS
VvVEn9zZAJIyZQ3/YbaAO8BMdcFvQx7hFDF7k+izxxz5dRPKD5GHWsj2tMR2OwU3cRs6sRcXmao9
qkVhf68lhk1DwDowh+WRliUyK6rj493EmENasAd3nEAlZ0EF2Jig0NaOuVBqiAy/+K3YM+KTpeOg
I7d3wQpCuXsYq/r+s2pIY3JtX/Z6yvLYnCajq2C8Bi7ByscaAAFhC8bKOJuR35M5lUKmNnT++qrw
1B6FSF+StbkYAa2cBaBFctd1l7I1DlC9W+Qt0lWGTwMx6Jsw07vyplbmE1y1az3ByXYCto7t92G+
VPI8G3nhWY6NkpUW+SSRgQovjtq9BHXW9zt3I4zUN7t/RoTdi18BpkjqAbUuG5hOWjYd3jcfKeGo
soOrmZ4OsRf+CmvNsHf+PwaKmlqX59pVn1DUJH2z49KjGJ5znqIZoo0V+2UCAe1ym9NGEOb8EoyP
zE8ky1FKMSrVhYOtby4UhCdQvXgXdpV+CGQhF2CAUn13psmSetfvnxiLFScLc52P8w4DUdaIJb34
qI23dMhIOWmKnJ5mF07ZNgVhEOwMSU9/YZMDu32k0blRBRexxNBeV9p5wDr4rGu86zqwHE/fawfZ
rqk2vpkY/kV23HWeA49hGTQEVTv5K/0k6uQN3okt/W9+3bSpJM+BNF8ZYTcnqrAfd5uJNApv8kFR
3HX71vbU/9QuL9KSNoYemOcnZ/PF6gcxUImeAzGZdt8WYg1Qptkdqg+rJnG5WbCaPYiDcaZmesyQ
z+Npd3t8cbuhir21RrOGUQlHzcmWS96BJjVOnQtOwS1KnTJl1alJJbP9llBgJIiFDrjAglvfna8F
kzviFpO1sx+U40Qu3PkEn24nlugFyUX8/OAgE1O+FswgGpqAh0Srxw9t0BcLEo2SWFiBIv3PumEu
QfIOrSCMKJVeVBNXLqYa4gITp3VI1BUhgGn9xyy2saTbzKgJuWLlbNaqguLBDbQ0jee2Lwk0ysBw
CW5esaiZ3VbFFGe8JvT0inl23JPGJW/Jic6oTeCQGghQ0lOAmXFmrEPvYz24+8EQHTVFy1wve+Aq
trgDmgMMxDlma6cdPn1g4gzRKjlvcX60nrfN2Yd1sIlsHSUNhgB9fnOWNxJMavkdwY91R4tA4e7V
jVmb8exVRPEqOs2EHHGxWoJQO99Mhwi6GcT827C1rcJDYXugMPz9vAujP1yxNoHM9nXIEMOgQSGY
CT8FPAT7GeC1Z5Y2E/PoZExRzoWjl2oxtsqDnsRIZayfoFXsRuU3AnoanCpArU3Yr7eMwZMPgWkG
2QkMC6N1cm7x9yPUf80gdWOSbf8TYy3d7dlvoAHWYjSZy8EW0WgzoUM6i5K1jZO6BuPcUnmySxSu
1uiCrS6ZCGNePpgNDiQGbApElSWu8J0d+oG9T1pLWXuFeLzIJDjzwlJZizXVHfKe+ZwlBOjG6ZPr
l3wAW3TYDAUARJ+UVwpbEgRJ8jQL8PjOUQr6JHn8xNKjr29ayWeLDpuI84KBWGvWqG9iwkCtFgj5
h1ECyTUuZRcdfxV95HwWWo4edDGkmbNV+eXrZbEjjYi+wVzvy7L1QsgTJ70Wf3JohZp2QAAJzjII
tSodIDTEu+CILQqeaOWcguSgU/PG028kh9dLqDAx1534zoAhpG67ZU9bS37Ujpqxoq0+AgDuDRmk
Wn6rZZn0X2SOZixeMh+Rl1kQ+i9acWtNioqFx23vcjK/eZAz08zU62iwRH/Jl69BFNCOe2I3Y+Tl
XepntDBW7Swj8RTARMnvm1UrzmKC4f+IImnZdV46fQMfc/c/Pu1lHO/YU0whPMj4bpFsWcij877e
ZGM7dmckL+ic0nTdqVsj91wOhQN2TQlA9mdhHWuo7RuRovhoKmU1WfCjcXMaIfST5uJAFErWw6x2
2p6eU1cRPeW1hY6qXT7QeSjxlPL/joLtl/FGsIAKm4ogyNxuhH/IP3IoKUnTU2h4Zv4n0GJgNw9H
OOtu4VRCXqSP+DC0/eXOel6Bj2qSBqL1Wkt3YBJtbrT3Ja7yJPjlyfRlYPpNEkNZVeS9u3AMsOGQ
oJFY9+EBdsigQ2RzhJ39j//H/g6IQszZrW407SCO2n+aUw0GUIq56z28K0IRH3xxjSLVM/8n466/
xKfO8wjaTU0xmBZO6XHVRvYwug7aTMWs5QkP6FQMvfNZVhhW9NGgeuwhCN2qXv71mn+98iEQXenn
r+Sba9Gh74H6tPq0sevRZ84XKD9e9Slcn7/yg2Ki1IH+6DvkWMCi6TvLsWIn8LsK/TJq3AgR9uEP
bCDxjB85tRkjVOdduMY7RTe9Jo5iqTyV1Q1OeHSO1wI35NYA5ASAs/I2qFLcukNmnwnZ5YaPfaT/
9OcmsB68ReiIzbOgiFBlfVB5lUjdFLrtUy42lHDSJJW8Nj6808SYqfimZZT3E7x63YgwHhUxt4uF
EKkLiTbOLF240fY+GTV5tNewCb82jJEHksf5DjRauBY1OLCwkWzS2xswfE7JA3tlCi+y43uT09eV
T/OpACX4gamLc42tbPUw9ZchZG3wCAWJEUjkouc2sSSw+uxPaHqfp8A7LT4Bg6uh/fxYJMxtAwR8
Wyru0qHKRhQrDjUGcWn+fNBdd3YuK72UB/BILgRtTOM/i0s2JYgWcmoyRmb55BPxNzrHOB2CYLEW
Jxm/jsY9PVjfx3Z2V9TlqywdIk7hEdbgZgkTXSsEcbNf9Kn39AQExswJgfuU6KVVueR10tyKtNCg
8cEEAPmjqC0dCh1nMYQQIdokXv0EUvgw8Ks1uDvUHSchDMlLJNxdjB772pWYf+4i4/pYphrNj0u/
d1eHreYMxdS1TPNtY8Sr9aLYdt297AhGEnSnixYPC0WuCoPVsyA5+nVK1X2w1OJcSfxtG+JYZuXu
eYzZ2dz/dJ/GjQ/CI5d5EdtGmMvnlYMHBAg5pRmQFEo+SiyPPWrJ+OwG9IIsc20MW/N8Dh2BJE/K
Lo3sKAq0jv2+FUKKoXERM6ctKIynK+0cK300HegKqilwOIj6bXt0pwSKzS9bpj3sL8twUEX2QnBR
/kMlufR3hwoqetMGf5DbEVtW4HJuBpVbNJq6/g1rprtDdntPfM8wHIM21ITBoBkk3cVPh2Tg6v9+
0ulhPc1Lw9jvYfKpaROLTjiyHrREaJxhEPG17sYU+m5891Tb+U7TosE+VkuwVU55iTN4y0gIgpIx
Hv9zk2jDpPKhAcx6BGCQF6VQtlT2/0kOFch+8Wb4M6d6+xsa2ipGkAWvg3uufV7dpXui6dTDVVMj
uUBYXkPfPf4mIGFcm86u8cZRf8NkdMiGvSpXoaxByobzWWAW72v6hrSTmgjL+xWe9Jw0nekFXfaO
XpJ2LjvdWhwhomFHBZjMzYzxiKDfCT7/4K1ctzYAUAtQv77WswrYxH8rfgdFQNJsaZ/AG9JqlCnI
A/FoklkHE9BY4ffRPRu8WfDGeeYSRZi4vpulrF6EmEdvfj3I9GZsDserTuYbhgftHNlBYZ+sTHgd
rsycJ6u50Qe4C9zcttrx4nO48wGlI2ScO0tX3l/v5V4o+y+hW2CHNZ/Js0ofjcd1pHrd/5YrQjp6
hoCo4Ip+kMQ6kE2wlpvCYNp8UWv7WcKJpQwsfunJ5tTsxw0qm8aRa7MARPstusXvVdXtniaB18uR
YL0HkVxguGhi7BynW9n0cAJf1Z2j6M6K/jakvYzeK46OPLFZWE9qDt2gki3AwvjBjAUW8ABjld5D
3OrF04FOjP1TTByp4rru108DcOcwJKoZNWnRMx6mQEpdne1ERMdQbzdxMScLlkY6jwlf2MJyPL/j
KigvGj5gAzXtqoTj0EnC7CJQ4errg+T8UAHsHlHs6MRosLq4IaK+I07lzhIKDNkBG5nvkor/xfHV
VRIChZ0GY3050mTdrPZslII2l2prLYNS6x/mgfyvq/6G7z+tSOPXGLMuiayE+ddn9PTD/MDCHWI4
wiNGpe8cb0CDZoIEULup4tQa8pptKgUmq9OYZJs4SHYlgZcpQ2pTugl7F+dRKgnhW37v1H6pMCpx
x3ixP5PHun/qmqK0XxWWA4+a3S7sa6FQI9jwDaO4u2K5cRNCjmsD0H3hActKHDMI6DBiMsECpETZ
byiI8AWkGkSXSATXq0EjgX0Q611JyJGvoU0mFIh0cp3suRp1T0WZA4mxKqTE4KfOexeGMampqS/8
jsE1vHpGDIk9p3DGroEcxpzVp8kpyNwNVYiT7TFckQ5X/z4s2N6qU8AmHnjRFJCFJFEF2FjfocjQ
K1OsHCo9UHRLoipiFiI4A4UZTGtKxs72ONFfoaV11e+2TifONo3ztZnrxB7jcmuB5PRYkuKCP8gw
6SJQAjcZTwiz+MCuokqhRwdyz9vLU3Br4KGVP6Q3uMjmeq5/1Vw1mCscnkaBnSzhcYRZY9OPwFkW
5LejwWf3pslqXmWbpqYkGEa4agEke4+yx9bc8Pm/dYp64oEA0aO79udLvUghFPDIF7u1Wsh6+Ink
JzElGjDML6SVj/JhLF7r7Zrnky0eyuWHCN5PVTivkRWzqmL02K7z/ncFd5MBynIkPJ+jk5LPKaSP
PwCGAEvRR33Q95XkHoJGIOxYLmrdeb2cmZZqsHr41UXtJitE7ZayU2o9LefjJA4Kt8f8eLRpweAH
xqxaV7WXfcD+k145+0SVDSi68nT/ziuvPvty9OCE06GIXkb2DzrJgHsv6mfNtwIC0mL2PDLkxz6M
H1jyXypHAyE1GFkybxCKFTWNuksiTGS+YO8FlnWBmOHrYn3/svq3CxgmP34Qi0ZpuoO44hO1/946
oN34t5ANvNHTVGU0VWr1b4UzeQwnr9DokNR1lrUBIC+SKCFEmupM9DNkvBROXS3rl4Ial9J7JE5S
v9sZc7NGeJHk+wJxKZaDTXFmKzcfZUQ8YlrPews5wZi8ocrFOHWbyY2YwxptMGYig6wAgTnDRc50
ECXesccWUrlMFDcOXS6p1MtM9T0Wu/xeR/dgRTypzWAIcIqdXgaJdVbtSxpYu0a7xDFDQk1I0NYa
PuNu9nSxfg8pqDiffNiPWsNqbYte9H9QVP2k6XQxCrZVpjZ86VBERTkMfFIehZPKopL4JEOkmlU5
J9uPR8RqzznXJ5fyeNaKYkK0OvPFfXvCz+UznH3ymPOa+sxahy6vlFT+qKKM2yq99cFbG2blPae2
Ok0O02jKtOxkYjK4ucnxjI+j5zlBgYEl5/NyrxgNAEjSeN64Si+XmbOTqadPjhpFSoQTZLIW7W+S
bTTOvKZDEot0p1hyAuwPugYIjHoghs3Nozc0FvZSMlZx/S1YcbdAA1Wqgjs4Z2lE5wwoVYJoApqj
TIP9/GpimjXpybsugP2DIqge89s8mMLq8Or44n3NGYrja0rdVMEpE7KiL62BA40nyo1TvBnQx/tS
c44sCFFSSeI+CIT6kehRG8Pjb4zeCbdSUY7TMAFirSVn2m8kMKQCTIZ90SEOodx+slaq/OU7ogpG
zNKNvq39clZogAhkW7Fzi+Bqq9oAI0g1eSlj1MxcqsK3h4/FoFuGANIMjJ2NmGwOWzd3KzsJBRFU
KEYh/9OUAVa/Sik+qtJuiGZY0WRyUvDbg4vttuM5eDCtjhFfg+WrfGZslGWWidoVB1olouP/7kMS
fo4+Zz+wZSv38R3krWUewAiZF8AM63E9NjlGCWLYBRrnztHdWUIkdf1/cpuPO54GO7J3I2kbmV10
51ZVAXAD4XJWjVAlnBqtZs4KktTdVuI+oyrPIJ7Y6OS+BPa5sNpb/WNPQb2jOqniQzOe0+NPn1Z2
KcrMkspgWK1jmNJUDVypwmcE32IPhbs+TGGnGXmWBB9jRqKSeU8f5vgID22G4qD0Ct6m1JfbgJnM
R7JpBZFUdiPkovDiCxpJgoHYPNsSNPbaZ4fbEDWOIQr7i2JHFig307AeHzVn7j6mw4l4Haebe5qD
GSdqi7bjAxTHxdJOlABnIyJHC4BkzYzUl4AagFckN74UO6uAVhsiWSKYbVcu1mH+h0aMrcwDTaXG
CaNQNiU5XIK1EgPcerrk47frQpIxDpJkckdrObt30D0s0EAtiOIRGAJdyCo7Pd7EKU0feIciF810
tE4bTSGnd0kWxvv0FHN3H/dWSpQ9OmUHo/lS45Z37zJZoNDvw6ik9f69+VKc+sySUDeKo23lj5aI
qPQNDF5i/qu0HB+xKzey5I22h5KSt9TYWQL+dzuejLKyUUwDucFdErvEX7E6zA9xsntQ2dAkJZlw
rFNbKbQIToyUBURdT6cia7z/22QVLExXphiuEfCfaNz1YN2TYG+kv6smRou8rAE2a4cs11Ccld6/
BrEBOHtfLEU8w89P9nxMXvUu6zhrKM4OGIbQgoUJbXSodd1chGE8coawpplNmKqH08J0HPpSB2BY
pkfkeGzSwEv0gk8AHtk+gOKxBTFaZmIX5xK1IRhy8X4UuFtu/nAEfTxHC0hbtpk7MP7SPKc9zSHB
zNUsLMchSYjKbnDQi2RozgeAOqdkwWfL8pwdtON9Z3Gf/egH701hVeSc9OarAeKSvjnj2Ze+XrgR
xDxnN6s3RyG3EURwUwrcf+cWM3vmwMzo59fZI6d6Mv595MaUDyfp87Bt+Xdg+WNSyso5I54O99KL
XjHd3VQYQiFZPP/EQUUbRPDOxUHJ1hd4oeTSKH1PL7GA9+ek664gGvcZQbIMWiVOenwbuyFS5Lsn
aGAqtpYHDD+b8IeyVbCehh16sazHSFWaFUVsNidhNey0byL1TFmijbyYr+rrf1BNcDxNqmvVrUzH
CoDS9XW3Sl4DsbrYApjPpuU6X5OV0vWE7nduRNGBJ4nHLLmtF0k5y90A/eyF2dIC9KFZ1fo4hazU
lbRhBXL2B85/CFrdzvpOEFOH5Bnp1iXlJzc6fa7jRkO56UL2ZzPkeFRZ4OQT776daaP9qTsmOczM
wLr4dyEYFpnWDEDKyC7S+ewuETJqwEktKgbhQ3P/tkaWfNWr9D1Nekbsha2snD6a6emgLJZ2KpEH
2Ya/jShWJKoWncVmRiN8WWgeIyTr6G2lJxKuR/X+OJtPqF9a6iM6M+8R76/G9/aenz0Otg7O4ToL
PTdsE8vLhrTzU4Mz/1c1nEMg9OlrydG2hbeNNqn/sjQFzq/skDdQcnZ1S6pwppRkOcb4y8e7DPHS
3TOXpb2zlVZHF9mcf8QVLAXKxCAJ0V4jH1gkULJmFnAaJ5IYloybmVjwZ2PH6/oyjVGhJ9YNZLqi
IByQkru55IcomVPhYNt7heS+p4F8KCb0nzbiOJYQSJPFRiKcbvj9FUXCd5oRoG2GZ49OA8uh5XGB
QZZit8iPHM2JA/BDNrdp8b3Y2aRL3WQhUe07s1MoV3D7dmE/L7K/gY00Yi+l0pJ1mo4NDoML6YB8
j5jAANe1YtEsynGUpDq+0NO9grB/WcBV7PClaHHCVBTUFwUkh4y0xN767MzVTHeklCrwV3WKMd34
pc4FAfrUEvwnQbo/mroeuqV0LOAYazvHEwhIwVUBTcHP5wbw+fyYpdD9JK6U64gUmPODtUW+ly7t
jmADnZSB8CZsHaAwhEdXkOxmu2DkvppiB3ZNjnJSmOLPvJwnGKFh7CBqHKaFkHB73Xf+Zi9YyWRf
1XX4kElIJcZY0RisRPDAPbVf4dnOumcWXTCSCnAK2dumAAI/Phy6mPLUD8Apem9GzXiQcplzfc/7
p6DtcHNvJeK0sJrMVYEe88eOS+X6cU9sls+Sktm/1MV3ub1/j7J2ZfnXS36LHSWpSiLuMhXIDP43
1H0pziH120HrMn7wU3jmpHiYZq+HPrx/tJ4jzXO8Ei1s550RcPfhghP/h+B4iWRVKpSdi3GZ4orq
Hgo5jcQR9o5UgXK4BaKzQs6hWVCMz2eJjBq4wr+qGw+dkmCt3+/fwZlyiq7+Okf6NyDZgkF4RqoU
vvo4WAumS1LgPrkTnO82a/kXtqC633B8loqWFFaW9qN5+2xX3bh4sX7VytPyfMKHWeogwOqsax2z
jQEWXhspQCO0tfWUBGwF/c0mdHtkPf75CFszkBQs9/JEKLBOC/mNHelCBL/zlF5s/FSKJQ2bhBAS
idxrDh63+I9RdnLdFf0CUw+Npo9+iwNFPx2gi7OZKIMj86QspHRKWhwvJhTkm2HVI1EwUxbPx6id
1BIlCpp6YVg//He9Cq7IaIr/To0qj9G0TD/xJKtt14wXcGm+kkKCQR+K+eC16nQyrMjOkBnUhvac
xtv2tMeXRzIpvvWOsQB1vxkIPvU10qPbFSCeqj2AapREp4Akm9q6qm3+cFTzda+67fB5mhRietD7
keICzPHrSMCmIM3qYRMW8SNlbeaQrCcnA/bcwmrdVmz7poWLqEARp7P9nZxgCwduwD3+2yAS70lx
+WJVq3pvy4Kp14IAEJPVOdr0wWx87fz9wIbEZ/gU0sNBkFGEP625Vb/UUI2zI5hy4/7ZTrJSMh/G
yiKGwQuovIT1OH33qrexHBY8OfPZd3emHKadAA4I2eauoWtkhkxUbcbXt3JZI3c6pQOpSVqysd2X
xwNf76Wmf2sj2mhiMy/yQ7phsWskRjdf12be6tf0QPZgt+SoEZukSBPpUsLkLk1WBD1HTWpbvBXi
46NV2TKJl/qpXt0acRSk7FcYDRfuAgJN+vYs2ALBWTMVpWARfToLiSXvI5gB+XXOFkXO+ig4eHAf
UuDnEYSJ7pNuP1kitVlZokUt2oH4y0rHxX1sovMslN6XZhBLUJmzvVcBjV0eV/f80SyljO9YY7kI
XWMP4YAZoS2I7szHnxDWxeFH3roRm4LzeCJ4d3WNYSMnAxHM7cuypMbs3oU3XFsjmUn8tlvUkhAb
2q/CZbyBMp/mYrK1gNX30HNJTLwuajMeZ5C4nNhrZksBn4pMocH/HLezIn52RfLmyrMu2O9sKfZi
hIH/bfzJIPA83jdkvk5HotzWwDHqLfG5vcTUFqeV/YE/WwV4J+HKs6N1fDqnEa1WD9fNmAkSgwVh
Z2Q/jrCKSf/seaVVlqDAMPfW9bIpvcmEyxYHrOLT8AQNe8xOu/kK+MZUJwoKFbZNu6rPe34vB6R8
L8uewdavBt17DuQbW0hSFvAS7oHaLePlz1hEFRQJh5xhQPxlBW7h6iq7aSx3nRa2dCtiJcQCvNWv
VpYDrydyoruubGJlQYPWjPApURgfwv1ibq1iSzb/ds2vnZ/7ng7mA2tEaw3N1qISOJiOOxwmXesV
hj0ywlZ6d631uo7et+gbk24I3o5go4a+1n8s8HgAo4VEy/a7JWJWwRAdL3d6h4tEZ+1fdk21qW+S
YYLbjaErUUz5Xr2+fQHKwyvDadT/zYE2JjkFXS0ySLuDQ8QYBuEIu5+PPMgaNoXgqQ7qtKgz+QML
HYpSzQQBgZs+tyyjpnpUzkPPGdf/wrvZcpH/vOF2ob+pJF7YqhpvCgMsuRb410z8k74HFzhuufjX
IBBse/1LczmrFye0ZXWXiANMSvP3rKoWNbWIz9zb6SYOrZR/+Lt3YEIGQnUW8yL+EfzYVaKV9ZvL
RsPHl2NwPD2ku+4T3wgol3jpU13MdNyWHKaVd2sdsP+Dz0KA26X037oKrOEzjqPEbmZlV/VEoYpu
d+lQAjvLPVQzDYPP3veSrFJ2Ql59Niu1b2ZxrevaNNJmHE0I1Z0hxqB59d53i3PaQcZx/FkB3hVv
ZvD0CYpPYcrMuE2952/n/LVSdMmeJEjml7nS/lxZ5o8thXJGeefu0CQzFty6TSp/5c9qj62RwsJX
lkO7wNF4iv0ul0hw4Ntw2i+kuUpBq/QT6veYnx/NW/BqZIOZVuYIWq1DjkJ5dDdjZpS0nSX9w+bj
b3dlhiEeKG08CxV6yVF+TcDoxJgrEluKtH80xELsG/AcQidIsK54c+bEp5azqXelfD9IxKHwueI5
tZJcs9W0Rt0QvZ+qqARJ0hmur7mN5RJgQsPJNqozYOVN2T3lUYH1+Xat3Hkd3Ra0PFREKubV5JhC
gaftfljqcZ4WyXSlNeqR7bTNKq8U3JhFNTdpAxwOoYAkKLKglTMWAA5lonKIwcLZmBUhMUamQylA
gboQ3Z9WUJtYd/4UBvQmV84pgDch0myawMoD9rbxXw4LK3I0hQAhi93uwILahXQKwGGyw5u5516L
h4nehAujG6bFfnY1BC1G6m9Chg+RnV0iQXevlrURn/NRbCOKEbfFSWD0gd+BuHDZjcU3r2Mh2/BR
eqQ/EZXloW2dg4J9xIpKzM2kQLebm7E2w/C4ffx3PBPxhhOr4Ty+TEm7RtUVSEETNDfkeyRgzs9+
3T4hpd/hnd63+rCjqN96gfe6FJJ0l8E86iTxZ0CXEVJacJvV+hQ6RnYnmZS098gCnclhgUHkM4ze
e+SLsbAXB6hW3mwxD98xxSyPJW499Xmgs1eHO3OIUOkVguDfFna97MmxwtjIHHKl3mEoAjWnNKUB
+BsbputxETyxePpxli/+3WSB5raOsWV7pizcOYkZD1BQcClfbN6P1osd0QZgi2+MrhC50qVrfD3D
QeRnsnzrP62nnS7S2d6TdxmwYt7k10wUp4XgFceM9UNyzovB8ulcy64OCRkGuwjjGxp2J5/Q+coi
WFivSlcIMzgqCAw+Ul0/BOx1uY3JRp9ukeUpj3WFk0DnxjUl9NyW4gw3eD8mLBa6tFJiZCgULNb5
tDvDCVyERPneJHjDfoUneNvMhp0gar6OvD+5J0sUBJ3IYO/IZKE8GTA2e27hcwFvTYxbI0jHDtUc
pgKlQRrxJxIsBOlMkrXjnoWIWi02hR2nHG8JVcK2Aitavk5b1v0vCP2wm0vIpKJvNwgL11RwWJNl
iWt/YTQ18Et7nWwWnLigWIiJ58mlrcIS/4AdND2QF9TyMTx1yIave2BdzqZDScS14WR0GTkmEfvK
XsHQVkrbvNLp5UPNy5nj2LgqHYfjr92CcwiPZkbxYr1RZVsK9+tqAaii5TvCRx1bnzLEcpcT0PQ3
KY3s0cRDyIorIWJLCbaYnoD903wlJFjhzZcfr36Bx/fg10T3iO3CJCnQjrHJyjch7Z33zN17nte1
oXfJoYV639fJB/ocb90u+2bZOcKyp5OMVADwIkg9Qab7aBosteBAj39tzp4BFLeBOZRzD2/isCNa
vN1hS91+b82Hdr+LhueBj9vQ+gjo9PuPz53k9COJDXh+kATNrdhq2K7knKfa9C5aJZN8P0uo5oLl
l/1fDCwhir0/ttARpB8O2i/mjyLopbT1y6WQHUXfgXR98tUOoM3YgSTYJOtQVXEeqJOO3dObbQIU
zQF4Joor/L1qeQJ/V+ydmKu//SbvFsULZ60VGk4Trm7gWf+UvVqIUD8SS5sOa7cVmvbHk7BCrgj2
h6Z9WH0dVmN0gag/rGf9y9xtm0K7tbQ7lzNDBOCkbzB5+yjRUxy47tshmXCLvVsWt4Wliw42q9C0
uqjgD2d4MkpBIRJZwrm2LCk4/IxkUgkN9p32JO27AcCp5ahiFDrnPB3OEyTGlMAYEQITFi0Mjib5
HXihoIWUNt/bQvZseAy65qAiOxQuCaoFJkvHXZ3iWzBFhmyICx/JKhPjaPGhCbSfY49H7E0FzI4I
17MAyTaQGEd78P7fKuyrCmaRYA4b6DVDUEvuzSTOVG6+ExkELrUaepOIwRTYMz4Jl2b+1Kil0/ps
AzVeU5zVrbrlumAD5xuLazuKfR3GResDPkYgUI7Reh+i5/kN3mmsHn1WxRA40qR4qQFCbz/acyni
y3TbRJGBQqU5qiIBI7y570Ra2uXTWElSQd/D0ZABDaIQB0aEvdVwLBXxnexwqhGbzqn1WHfQ2t6p
MmmBVUUN4Et2iHm8db+T7gsFVy3q6k/aNyZ/gZjTofANMrFTo7g652gnYB7ZO1CuUFakJCboH38k
chTIJdgYZoTjQDqhndvHmvAAljpC3OXYHiqG1dFzXSt0m4cGq0FtVZlW6/aCc3G0e8lCNDK9DWlc
q3uSIhUVgOggUhY3016PBGsPmJgWTYIR4L+irSgvyJkIB9YcEI8zY3Xw6/3FPa/Jd5u+mSu6Or8X
G1ZP+Pmx/5irP8+IqwNkzYzD4/nqgjL0ZtVGDeSM9nKNKkFp1HsAcN6orx7xrtZYWVaxy2XsIcJ6
/bTAvcymM3stzRwu4b6lVDWyY4NgpnqK
`protect end_protected
