-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gH7q3KvE/NnQBQy4NHVna/3SjYF8wiYeMV86uepigt1ZfwbgmR3fm/owKxiS0xTKPoLy3uAaOFGr
n3Dkgo/loHDX9b/FmiNl0haU4tYGoAumjCGlpz6SmwJQXhUpSWA5bJ2AyVNHjlqeWZLqc9gkxw6P
J8fdTsjRT8mPlD7OXKNlUBRBx8gw1ACf4w4ZpBO4HuZhatLawcqqtZVpVh9FJQNN4We+u3NsrBYj
OrD3Q4CsOZ3CzBi2wl+AKwtqC8HGQLX77oG30FCR3l3xcvp2Nv9U6kqzlmmhAg1Z6x1cMZLmtFvq
YRPBUr9GM4h7S0viNMmFNntKnT9W9eV+c5iL6A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
opyXXUq3pFo49HPnnf56TwxVm0a4KZbxtaul2GsURO37uUhz4/UYLQA5sPWO77mqEAm9FMwkukfk
TUu/LA92LFjZPiYyZtCOmxArbtOVtbCCdHcUDGkpUOHpyK8zhtRTrk8RCLoKwXHWz4dE/r3RT8FC
+oAxWI41cNW7fWQWEG+kjUYhZt1DvGLswp6iJ9QICAqq4SeQUvvQq5Uz2q8KhzfoMOmuMcwg2FzR
6PVq7rXt1gpS5IUmJiN1NWz+mr9Slc4bE/q6eGx16Cc00jxURypXhjU+hHJAmZytpQ5QrKt80W0n
SVJFVV1kNP9UuOQDPoUnMvzfaCZ2MGkKPVwLctQojdsTqeSi75ipWhns7PqtjZvbwxwnUWHcsMrK
z+o/yh57butIZDzWnzenTb6FKEBbP1HaLN9u8IRBGkMM3gGIXae5nn3yqKp9oFe+ndMZcs9/Ojvq
ilxQhI+BEviZZF33xThzLmrLFnXvviEx5dZ6OChA66nVPdJoJYN4KKPbfRNbQyzPzck2iKRks7ma
lzjtH43kAagHsux9OHCEWJKxM6DoOyEswK9P8iP/Oj6M1lkdJSRhkOyJmw3LmxZtk5bjjFET4qYB
+30d6mlGN5XOF7z6ae1GH7DtwyPK6bgFfM+5p6PWOiKtB3fEaMSCnixyj5VeGcSL2p7mGajCb7BG
mFKxcHMGw0vl3fDgbaH8wW5mOyaqci9KTGiinG6onlwNJw40PnKo8MVXWy4EnLDK8JBhhQOd7+tr
CPsMp4yIxKdytJat+5EH0kjobna2BokkzeeKw+ybZX4nsp4txSdiLzxfRBhd3oEgFkvKE1lc9gmz
6IzWzz4vI9sC0KCUuVsoQYtFxzxNlB55FZpVw/kyVV1+byrXadkd3kb+tYNzuiNHJ0yO8Clj5Oix
Huc3ZqtyJcLk9C8j3nI03OG6xC+zEMPm7jLMOnjaP36TdYBmL21L4OIy4AYaBerEi7Xh9Q7FwCh6
6NNVlPxC4YM8HraMMnNGGS8Y8RF3WZXejmw8UJQdvJ7+fzIpqcr0SpjT0a9e6E178l4Oej5KuntG
lOa+TdNF3RMCWFmpjkfBjV/QPe6AmTM8ZG7UE44bz/RhHPf2MC+b6Q/Ho5CMlZGrGiiW09YF6OeC
j9+oRdBT1Jk987tsLqm6vHq5IjsrWHBP+pPhnVxb4fORqJ3f/ydjynvPjoBqTxxQbcNvLIr3W+Jn
V4Cz7KsbSUG6KKSP4msVRUGsaMbG2nuqPeM+meCOoAyryui/0k9AqXHEU+i5/AwpUledtrWLirvT
1V4mBGR5PbP9fdSgXGIOvhviax2B9IVGT1UbdKrnSGk6ejZSg7xGSk3koL/aTZvl7q1LxTmHixgb
TMV+Ow0gb2RJXwRG+vrRa4QaNerOq0iCRpTJ/V1X4dZksYSdHYqpgS5UlJ8k91GEpuklRfYu+COQ
BziLY/U8sepd39nz6wHLWlA/yfZbO4qjacWo8waJb/D56rcv3sepAUenvgDuFxhx3TJWM/JvM37O
JL0VYwUEWVbj9S1U2PcImlFnPc3PiygVF+73bbP9+SCqRpZA5LrLj4Pt4RrTrJfLe4ff9z70nTMd
Zzyn2/2yKe3asEXRErzxmbeh9FNi7DHSlePOlun+CWozJZTkQIT693mDT21lxFdHKV7YQit1WTjz
nbPhyH6bd/WIBHDI+iF3CdnU8L939qtOg4e3yIwlIaSHWUrn6QWYM19ZWr9OencfpA+pwUC89TDG
4oCGwIgSuJprpwk1UhnKimhUxNSrGmAOyDGfHFO61xK1p7dHVhLSyNsIjLzuhzgXFCDnzsVv9biK
DcAvjoEJu/iyjI9LorAX6GmvRQBj42qDXuJF4w+/8/ZAPgx3XA7OLGPjaEYGgPEN+ZPsLazzBUq+
4FNU7ke68gpZ5EriV7P/GEuqo4VjgTocTZUFUYCDCnp0ENSeKUK8lYW8W86XBAWfwlqSafc73GbV
3cig7Rm4qL18G3tTQhKTG4NTFFjJL5bwWVFBWhDaBDhcp+HesZmXJyZZue+sc3pU+uxIbVHi4GvK
mGeGLechw9ExaSV1HHIDmu9utU86kd3kJxofMZNiUN8UtxwxOsqCAopUev8h5LSFUcF9Ghi32Ufm
HC4zwJZ6suNJM/suCIM6iGllyOOaMr0uFWlMsM7Dtqsz3ilZ/MGSP1F75G7i7VK5NZ9egUx0nZZo
6PCP/BkfJnOi2IIaMcCutUqNsOsiyiEmT5DW0qWMUM1Dt18TeSYzsUfM0ksZeIBWlhnWotwl+/cL
gemc6asNpCJmeybjxM25JAYKhVPfcs5K0cmYaa6pQxw6fFvHF8nP1IDKsHXgoBAI9+uPUr/Hg3V2
SCdAqD7OrxddgkZHLm+gNVXZAH0z3ItgWthfY54sFf2Qf2qEocaErH7u/aMly7UkkoMOodTWAgIQ
OBxFIdV76i3Ajc0/2yPyd9MYg5Blmt2+SNwuN7c0CrMzsxbIHbJC1wVT9w8v4lVMJIcyoxPYjdgo
3v1zLcCxdWFUen4GCyIW+U29xEf0/zDUXGWOzYHfECOGMSDjrdZoNak5kASgoDI/SiTFVn+8ldSW
hFLQh4rvzIVdqCEXT0fJ9QqdZki+G7fXmYTjq9cen2kckfkGIDWu4gdrIgc1h55dbW+87IVCYPp2
1mUWthJbjGQ3TcgEiFQdkOsp8PXWNdI2zby0n1+p+3PybVhxf8Ttgod8Bq+p3a1RaSkmhx9psrm5
ioU1EwPw3S3IFyoYuJfJhjKWGSCxX4YrbQtsgGAGOhpJPHhExVRP7/Ijz7b/2J9T+MxVTGZ8EBjI
FJ24UJvmVCd2poBX2cynwokBKzJ3EV398/pDQe9zuqh8qiOXu/9VF5kTZbIl14Ls24CQSpAnlO5l
HA8BLdY7NcVK/Tl393reqcC5rZd+CK5pSk1GUPNw0iHRJvQfvgnnW50aCQHO0/umL32AJ51x3DIn
d2SawmFQkftmRZwnXYGovItjV3lQdYKnX7f8Mo8BEjCYVuGAIPIO68r4dE/OvLeYEk2telJozctl
UsMccCFXYb0ZPVT7iRmHwufAWaG99c0tN9HByGUSU80s1E2EJMeFCQkUD7H8Zl+bVLF1+g1yJLzu
ei2P8zWXgQYtnGt/yoczYS1JUb6PaOOMLTZaEHDySPqnAvVQWA7v+COPSs7UcZbXH0RlbDatZS1Q
UWghUoVQa7RvPlUtk1CterOdapg26w3RFDpUgDs1FCMIN/YzLor+cjJK2sJgx9JwCnieVK8CwGur
zSP0J7wi51AtT2o/kRtTgPb21MtMOdu87F8pJw+JZsn3zqb/cjxANmmXGsIOn/XvptxHtYViV02G
3E+75kiRfHQzl4K9I8Bb8AMcZvItNWGJzCEJC50vKMSwXReonmoODheiS/Ac0cJPJn7T7o581JC2
CxrKRGwoEBTFh2mn1x6b4NSSmlI1zPBCjAmvwA4R0L4hZ/QsvxdU+99ssRrXj81QwAfHXyYX5Omi
SJzSm8pt6+E+JbwYgK54pFF/3N7liScQPieql97O5vDBXNkWjQJK/Jlq49tpKc9ovwndx0hs+SDa
h4ezzLhfhXzVd9cUCw5E7gczs8Zwochlpsxr+aQh/PoM87DTdW0rgA/HjjUi79JMf2EmAoyKIN3r
vPiqcVmA1htZI92VTtvJjplsXH6XbdUxVIr1ZndKA5hj3pIJAO2K1fOsRPhMAYd0Jp5A7drDOeZs
Q8EK9WUjHm4C3sWQxsH4u6A7fl/qlrMvhuRJRZMqQh67lgl9aKYjEM/r+lmg9gB7pKlIC1cozn+m
jVvpkvBZ5Y/cZpTTmuFKVVRlSaR9zDej/XnPMnOAaEqvc67AnDeKk06QFRKUuLpEn2MnZt797CHI
nKMPan1+hzFZfQ3BvpJY+kuC+/p/8nDSAdZwr+Rir36xdmvrkR2a6NaHXczc7IY4t8bVTWvLLO4B
RNE1kL7o8ZT6Q46I8lyKML4br5FA0i3CLx4OgV0wXOBxBU1jp3rvjP8xN7Dbg3K0irTSAx0rq/WV
F051pR4B9BK0sT8ke8JFKv1pq/5qIjHdD4oSETvlvrT0yb6NIzhoTvQll2c+DBEZTV3feRAvMTOA
Vtz4fpW1jwJsGSphaj60HYrQqNRZPe81pSsQLuBbPR9a7ZxJtBlqFFZFXNEd2am5KpKWNY1c1jVo
NMGP8sv0sBc5i0IAbI0hgDP54mCfrGk8f+FRG1R2bFq2yHzrMGHMRwAMwxnbm3ut6fUakw4kGv5I
L1qlhl/iFiFAqjjODI80zkmZWepl9H3guk3Dt2e0iYct0fj0QoDiPwNBPglodfTKxFL+RonAo+qe
M7LEVqyKjLWFTZXwBGgdy/pvrNldUfxuAKB+4n1BnEL4OIQ2SCfZ/q/i45Pfvw4vHzW63us/nvsE
vwZUzWFQfu0a62OqxKu1WJcFL97DAx0jx+BcBvpds1xGcKNQt8LvYlIrnDFXF8MHIReswCFbpTMM
bC+C11fAbJYpHAEVuCHwKH9Zotd7+y8/oewUIe2WfUrnlSp8IPZudqLHdfH3EmihtlYo+sIXArcu
oHoioFoh/QDAu69TvhrkJ1Ng12gygQzXlqWNP1b4/XSZAJpvcqaJ3eL8kcC72BR8dGnFDX6c1JKU
GZfmGnFQhuYwpvaUDl8ijcAPEtbcxeiJKR4+Uhv4RsYwIJAp6gCgr/zQcWFIR81TwgtUwPYiQk/3
YCmnV9ezZlKBRq/IPnwK7j8QqMBe3Igr4/o6Gi8n9xx96DQ2O0pdFGcR6dv0d7CcmwYanDLgggtU
y77uy0rR7SQXykfkrkSwGxi2q2qzd9aJWT64AluyUCswWvhUKn3+cUEV4goovZ+BEUE3u6/vAQT6
Zt3ZNl2pZB9fiXyWAmXF98I6/xCD0YpPwWLEVKXV0y64X99XnKw6OWLW4ooumULzONpKuR/8TQfs
ax66gIwauStMgC2fPdO6Tscqvro4U7a7q1hk7XZ3NgY4AM9wtCO6UHEn9II9muVKbvUAysSMUQhz
L+KiQNQjT+OKiAl9c7C8g5Uq8m9xTh7vL4h+CTy+XH9GG7IrRxYFJIm86P9Dlm4TwTqhEhM5Nb/F
zr2lz3WfYyV6CugcngfhigwNdsqjVGkcGpcI6vfXapuvb6wvwG5J7IRdZYl0hFdrxqFtbDdwhl04
i+b1zeK9ZpliQhvunujvLr16L4R6ORpJBRQ8YcUHQD9bL+7H7Jy9SmU333Vv2bh5Z0iQAuAuOfmb
1TrBGzrMbFQgbuDRDOucWEzrkrVOS+o9lpvQorG6ScLo82S3mj1MsGevJ+eOJnuJHAVkXGdCNuGv
+FIWn/IY/MGi0L3jG7Tu1UsmTJv4LtTypDJg0MszBXdXv8Co/Qe4qw3wBEguiBgGG0AT8Mja26jW
VdjH3fSE8SWbrFBxM8jrkDCNBm1DfYMR/Nlg2Ex06KsCSym1RJy7ulwcgQGewzTW5e5TA+hfHG9j
sFIq/siA2/GR7A85a2PmpsyzIYtqF3My/IiEAlew5zVYcZ4vgv4DLBaFJYNX3tNBR83IJKeVv2no
mikRMYf/G2bD3HD85cdekFnan+vQ2bjpUG/4+97yiNJnvwOJr7idcxGPGfK1rL/s1ZMA6AP8698t
7naQ8Si9d+FJv8fG1CYBPRr93kDjrdCxfdDf7El5tBpOV4G64I0b/iV6+9r+Uy92HisVsfau2WOx
vnstH2kguyLbuGBFbPC7eaK+kZZZW9kZRBiRPmuprQzFfPaCwi+6sWrgsR6IriTd9OMdkwQP3AW1
QW1y9ieQUdGoOAQAOfBEespFfe+L5WguyzU2ZtOC1V64KupBxLlG3v/v0pNhPRWOG62+B0XO+Z7D
G4/k7WCgDI1fTI1X5miIcyk/2C85HBtURKolVYQzfdFpV/gq6YUJp6oGbDJwfmXg7R4uR2FJjUjo
lWbybiD5vZMlvQAb3NLNk9vBT/mNMXsI1gA9M9AhYfkORIANSiB0oSA+VwZkPHpK/Q9diFmbOUSO
PeGJMJnF0V7uqNi3w94W9grHNDxxHRAlvz+Rsth43z7yR0gHrJDeG0eYqy44VUUi/z7F4lnFH5es
Xua0djWrZPuUi1rn3NKuVEU5GeDyhia5Hu7l5qQmOhDyv6RILy636dxibjSdeCnLdq0EgGiHg9Xq
uj+A8ziNExx+t+yCCCtQ8EMmLp5/hyDGuCjP1tufhwbQ3mK4kzfEurizstym7fO5yADWVeA6ScsJ
AFQy3UywxjXjCzYPfom5tesXKIZgrWIF2IW6gNM751GfvZKVBEbpwYXsVBZ3tVh29eEWfoJMlvnV
tTbqSV5HwLjHE6gkX4+F6A5wgy0r9M/i784Ggi8uKyCZniK6XZQ3fMfG2/AeBeoegLvTR/NxCPHm
j14SKnZAm9utfxPPuFjtXtfB4+OQW4DKm9R6lsGjTYVzxR8Qy3YDjELZoGkXt7StHapDVhZbUwMb
+wuRdXZm4hYqz0INpOKi1TtSaxi5vnMC29bnNwQ5tq+Qzi4laxgCNPzXG1gYRzkzWY2uy8n5ZwpZ
2UJBXa9ZqTXbehS9TxJEg/j41X3iQ3bDFjx4aePfQyOb/NSdWxwhzjRiLRoREFmsD9IYcFvFO4wf
jwE3uKYEMad3J5Mtigg/XWskE0XWk05zlDpHwYfV2LES8JO4d3e6AkECer8JxjqcS4akCJd1LFpT
Nj3Tb2eqxmTh+AWTViJCQM8iUn5o8/D2oX+WrNEVdEvMhBKJnbgA8If4ZtjPoe8+R1VE1yQPc31G
ye7V0mYpzyMjb5GOjPRXSq4D8R0cSS9dZ0Y7fuBagqkfk8Rr1QKTXtIG5yeicDisEbiHPa9N6Rie
5CGV6/qXpFnNu5XvpQQ4DOzWw2x/xI18CEJhogc0wsZ3V+lreyxZC5xkAwjbczQtWCvactYskFZN
A+x68WJlis7bpz7xRw0Pn2cdx1troNgn7AZmkm9NQ2erLEwLmFRFlQFm+bS0q2QNZnHmsQakf4DG
1v/o5uQr6h+MkOCcoc3mLHFYj6jf9JXQEFQboai1NdquVlCi9XC9YQg1QEykKZ0wlXm3fzaNlUYR
zxmyHPfDQU9qMt85/3VA7kz00xr9K/LkFKUQGgUeBY4IsMxXY7QNItuFAsoRO4NvfzaVeAzZT+SC
MFrba4EmBvSeK70zVaRqagYxDGQgTaFzJjOqaGfKEptYRXjVgf0NkiHjOVmJ+v1AU5c8PnCmPsQ7
hBZE7pjk2ZvMsHVdKgZyQNSYrDxmIOktI9AOalXq0ebw9jhKwif3iX9w4Xd6ASKtJ0OZ1p3sj6x6
vECHD+76CrL5ZsbaBdykcUtgJX3GhL/okJJcdxClTnXdG1JRNqAD/5RmVugBGJtjW+0fV/RFHV6S
CYrIWOmf189m5h8uhUZVKTJnzEjmQpmRQFrslWNuIeEYf3yyDOtiyEvo18enCDSocIZPX0+VdgZr
YBDFv+AnCeaDYiaMhoJOwt8qlxsjtZfpLJXMRfInnV+Xj2qLs+HnnqBklD0oo/FOq57ERxYDUPzD
8rmouuc+MZ7HdB9PoJjiBBZNW4KLmdd1jSfn2qw7z3QVuf5c4frhq/oUzXmH8hJZbDAZluDAcbnp
bKJLMooWiw0EiEbuvMTILlWngc67nwaLflwrFHoJoIRDjjvKjTJJHksMz+x/7iPIjsg4ErFS2mf1
svhrmvRXv5G62KSHFC1d6PLof1MF7M7a5YamnOtutXpv9TGeVix9KMwuBcX1eJ4OEdFUl777mtNe
94CPDbpDZI+vjt9o3ymDjS0HKoTICwTA3K8B4xuDo+GtLidZaIlqAnJrhmGdvyCjg+tN6VOTTSBj
dHsYxA6JIW4U+Odn5mWdaKF0R/cTwcrTeGdaxL0WUxnobbhH6RlFMmcJ5by8Akd4xeEleQ2D2tQL
8jSS0BmfAX0owBBWThf8iWFoya4t3NqKNKEf4Os3Rx8ffRIt4M7ZEeE5BjgTaHGn+pOBLLAgO+GQ
qePlReDJtjca/H2AZuHIMHaYQT+kUsewzbSl7z5thsIrD1we9UWNLtDry/Zc2l3s9x/R/IgIUjEA
wzWVH8bUfxvCsQEdAImlb/s/+9X10Yw/vQtiOsmApsU9RApxmlBwkRQDcbKlzFbLFqCfFRhSc7i2
MPwBF66SkJ3q6n5SYY0xAKHWRF7FQEM48Xa8XqdFiLcLis5f9ScaMLCx/cmBftodL9ai+URbgXww
uLKwucbXiRCoIYh3oguVDXPgknbkViLS87uWBEovdPq1TYEm+wdcPNYGCFKz2YJzRcuulUCmZnWn
fvZPaDYKNLFeFDKjhqxFe0FWUzo9S/mYLlucHcml/3XYUTCIQe96kkL8wWpP3xDappKUVigHfLHY
4/S0UNoRF1LvwvqfVdS0FmTwRzG7LZrftivjbouCNfcA0HLgXcliPVvs16rEVBl64DEsuJRTB1uh
aH5swRmZVQ0sAjDwR8oWDidcBw6XF5b5+a70Kx5CekVEC+9oeko4vWahYyh7uWZ4TdEnG1SLM1XL
OpcpnmoQZIf01ICq54in+71kOVEfLtxsUPfNmaVf0QSPyF7NJbX7kgjAgzsLQg03TK5yXXuvrt+P
lZUETOU72LA9uo8tGpv7NmIMmUF3+sOR5pDo3fEiqYc54m2EWROdd5BDdBSloBf9dLw5qJkIRA3S
nZZ+eim2vh1xfLIWMIWyl1fTE/9HykI5n/aoDE6qXE8QHhfx4jaQxU7YGLJfez+bF+paHy68qc6o
s0LiTTI3Po32lYnwm71Wp3CL4BxfDwqPnJx3aL5lMEcfhrMiE/O5pWOsikuDfUymtNZSl1jdTywf
OpbRsJIT/Ohw5mDTmLmN0USMY2HceVvs92hcPol258WRVK08gNZ6E4ozkF3tBz4rZaiWwBx9Ojne
uc4Ye5/1cOuAMEnoIV55YGZ1hPmw+KHTs2JOacByYCs+rgKMqmebbJcy/PVTb958zLmYW4kPGCz2
XcJCVO6J7YhoSTHQqAcz0KSo98/6UbCbey8y1iHZ+iCO6y2UnDNOkakRALElmgQtd9i4uX9z6ayN
RDXFWrtlEJ3jeSxzs2tZmKNKJ20x5U3C3vPow/webaTrv9FcbZnWNlFcW+XYE9eN0r9WgKJqFo+Q
QcDrZIIr3sMFzrI+MsbBnX6W9vW2qQ+QG8EvlROdcWeCkF1gkValSsU5tRiFDLpv1xPz0vTgwPTf
5ZDVFI1SozfidVVWEgUblEWakLvXRQYoSttYU1b7xijbEJOy4sLwBKQAM3emaSp/y5ThhFsdiSxS
q/ZX7NlMl+5z3OjH4gY/ZtZKRoUGF1lyWp49WTsKe2Ku8w/MmGwiqoI78RBh/CdFCOgAClSpIRRH
+1nZr0hf1tacE9ryzMG6X6XjhHuv3XLU6zKPzivcku3Q0sDFw9J8uLPsmicGnF8zCdADHPCWj1F1
p8GcPP6IEfIRdgbQ3Al62dUVlm6nJNFHAloS/ZG/Ce89qdaytODs+/VOGl12g39OZcF4pew87wkP
0f1zWNHhHWw/88/mZrJVpGyQojgft0LeoP6rp62IDs6mnw1wH+Srwzp1lCPKIwj3dq1iYKNEBLU8
d6IvSyPdzW6odHWuJ90fLczqz6yhSTYe3pm9q9gjpesuljI7EeTjK5/b3eHEtKEiwv986M088Q8K
Gm+ibus6K0JTfPyEczHDd2YP+3NZNHgnouB3cbheGQoSlG+0Bg0sVSNDMQhcXbEP9HryEuN82+uf
C9IGpEEPVy6jY+5ngAzVUEZg4qZ9rVjXhN9/e+/JhkonoqaovnHffv6Hi0cmwXORhOXemjyIPyHj
IMrVBZidLTFjbqugLLpCcK9bMEqO1LJpQNjxDeF0GBznoi8ccx3w7l1D0NDCop6HKRXCrSq19Ysf
9Ejr7w9JJaxkOWKfpEoPNdic7hBaxPPST8AIKd/5kj//vhzQD+1AygqYqSFtveo1pbbhVkkhrBVK
6pLBmYcJ6IMJnK9oGN17yVjiYi4bXJ5p/pqEvBMVPE2yXOa3iSVFkDtZDU5rXQ1DkeDpKQ5Rlfs+
bMwA+o93AUEjoKG+WrqDwxlp8Wft7JOX/XyeKucfBv6GApIlGWgkiMcRE4/dDBd5QYyjXrzEm8Pb
7dex2TdpJKWMDUW/XJZYo+UrSJFAy5Q5oZgoijQ8sfIE+drF0S34e517HqJ9iOcpEODEMGAgOi1d
+S5bVK/vetEYvkeOVbjdlX28W/zsmjW9Dkr97WdZD+f/Z/gXIvy2TCrk/qgmX7h15p58s7qs4/su
T6aW0OKRYOHK6dhULRqfIRv1/2jQeDBn0P9FKujgw35xP+fMNgwITYuEdsp+LC1KddfVdo+cnjf+
oaTfMDRMz+Nv5lWfmZ/wA3arLO1BhlxIIu1G/2wwA+ZQ/glXxPczqjkek1GevNVrGnQaj2sH+pQu
GmBcR+kybIPJNcbp3UYHjG2MmbbLh+EUTgBQwisepyocM8pNFHfLsTyJsTuCoWQKjhytkgPpAon7
RYeg6Byn3Xxox/nxhNOWStc3lchzfB55H5bT4xe4mC6ceglNNpeg1JaoKDxs2G1tJG6vibGW34GF
qgyg/2Wa5xgtk4bSPd8/lEieylfYsEZRfZtGJgD/9W+jxveyGQcGswYz/daVZcsbswnsOKKT1Nrw
vhH4pSmuMLy94CKa0JgBZ6ib6TkgXegN5gWiDTi/R5+Piff56JEvCPBf4SAlmd4CE9fO/63pF+2V
yIgdmx5RDxmBrPEbxKq/VQOqUiXhjJD5E4zH/CUBhqC86ALizoMVwCrO7KPdHEsSTWQtx3TwqB39
kv6GPnrZT5pYV5y4VPXiuETmPKk0sh3thZVqv5IzqVMHko5qfFq8/gIBsXBdNGY6dDSkHk9M7g8a
NvDgwJ0MvXEpndIR3NicQ+nKky/YcoRmeZxeK2nFloBqqsU/02MLWDzY+nFF6Rs4JsgJig56/tS3
hCgKMzhHAhTaj2mtYA8QjzazwHNV6ptkuU+sH4og+AHPC2MDXSxXUpDbavMXegdHCSz+kKCaclu2
or2FAHdmpnq/iYVtKpGrBmzhzgTyemRAs0e9/yb36ljnjdxqcMZe7shLg62KpYAMXSPik6+J5TOm
Wm6LQG4z4MS8qoLovw8M3Y8jvM0HnxkCkG58LXM9o0TarPdLh7K7tFTzQnxCKucxrxfjq1svaYcS
CDp6qG2t6YPyd8H1IZ39G+tcQdKnuYQqOw2ymrxsv/PUx1ac9EUNqiJPELWo7SSsZ8+pNzi8Vpql
kW6PR6iMd8uz1UBwk797cJmXKE993iQ9K9geX5rzdAihIguDz/YbgXbeFPuagQVTcAAEs+psYSJ7
OLxIc6Org8yXsUzVNFlieHOO8h9zYiLBI7Rnjv9MCFGaYhovXQcIxPm7Dkspz+18ABQ3ODBYyltn
w4+1yKmKr5abCi+u43h84S4ORQ1oWmydZA3yiwTQT9KT4YgW/D/KVoJmWgtHI8Jr+Iy2/Z1FNpaW
2PLquzbTpEhjNmC7gp+O4X7fqe/9kDhcroM1RmiV9T1Nl8flJwgfgSBTv0K1lHXXctlgKnfoZHaG
xnFRn42tomiQjvDhYv7BodA1WcJpLNdcctd4m1YkEoZ+3LOGr/dVLjstO34OZA3RDmfH6o2pod7t
Ou2N0he54YfDq1X86JSb1shjP3fsOdFUdhMJeIM887cF3TSa2KvDUnH+aryTdwdC5vT1o8gbZ2dA
QJm0Td0APHu3LOA8NRg5ZhmN5/2JSlZL4nJujbYYfimuQ7M2CL0jUkAu4IcKsXW539UTd/Jc270A
ZLOoPPgIpC7XnDcO25CjPbCEEj2V473kzOsg2EpO2WJ+s9yyLej4AiSh6KaoXgVJoeD9Hs8nDO7g
8B/N8GU42oYsHvjR43YhmfikE5pA2q0+byA6jHssBTVGxqODKhkcF0p/GErTs63bWhFOkYGvLADj
ROq3mYdyMKsyQIwSavC61BSi6kw+byN0k3eUFc/jC6aitMRDZJZwLNIuUfbRz0Q/xo0sXDBRCzaE
6CFACsgQ69zcy5sC+pNGoGjU2RMqw1fnZKc6LIDw09Gw7xzy/6N+TkEO09hfw4b0CtgptqCtaGXj
fS+I51FS4XjJ4NUpvrG6MIg5g2E7zaYQvT1Idj3IMmDLYbQQSRvEKkcfaFa0mgIFgM2t38xcHy/v
uyIa+Np06KKDDcJ6GtrZ/mGKW/6NQ1WLHjIn5QoMg6AIrCW8zJft4KUuIzWpLevlkw8pxAOFAGZ0
qObKEwdzqS6IcxbGxpP2YDcRoGzgfwqp1dw7VUNlUvKtGtnadLPmwa2dkQhyVzoFbwF1wQbRiPcl
0j2iSnDc5fShFEuzsnvrJ2dDHGb1rM/VGmN0Uva5V+WTBAeCBFV+7y9ZCRqPLyCObHKOCsP0YDz8
kQQsej7sS++yiB8SRqy+EK4jr//kS8yb29iUcj1GLX4z6dnVubOcId+Rt1iJiQtKXHRZabP2IJWV
r1NfvaCXetx0Jl/RddgJr2P/ruKU/3tsb8k2jR0GFOjcRrjuVaCcQY8KIZ9tIjguWFvStHLuFpnF
zxX5rk+Dbpw51L9atmSiHnFJsX3sJK4T+v1qaues+XrCIn34lbUJB1pGe1cSI0y2H7h/xuFiiWv4
lJz/dzA07yY1lyNxvcw1ZOBF8hMtiG9BPDO6iPpalLwol0mX1oDBX1lxrSVztqB96HEAegcoAEME
/oAUqZQ/ezOFK2wB85JfQRno8vIWG6ahsRZYL431d+LBs+6qGJ/S4890Hs5WjapCiD/GIjfn4TZj
WTQnFFkLZCoRAJY7daL+QZkEaXwOuCbnbZNqeHlaeuae5CFzHkJuJpiSBL4esCA/ir4QkcJ8s+v5
OYqCu3rVJEyFc6+fbMaQ7LvZmYtHuTVSKWDieMPd0OZUlTlc3F/ly5U+hX22iKf9aTSph+SFwvm6
2qz9holpe3JQsujSm2JV3jYIiIpGFpio3fVkbkDkUrppJIizQywM0boZ7cepXX4DQDq5us8+GwMP
ihltc2JZAYH6FQDKeX7Y9/5vET9QwXIl6khszTkFLBrBtEqlSYBbXhBUVQovh/SOcrKqAUEFBHx7
DdXiCzcdS6H3ZPAeeNl2WRYEyt7YFZf1knUMCkgW6CAW5axGFsBJeujyswQF6GhXcYzbzIQMfPMO
nnP1ifGKoIlOe+MtABD0Puc3jfpsXa1neu/Nn+huxzm7dAIFI/gDrX2ZAzn7KQvMw72dwVE+uUs2
z3h1bi+l8hX/ME/8sEk46Dz27JlYyzNa7rknc0iGMns8AGlXEj9fLOkmMb538WlJX7tVm54X3cOm
eNqCV9TySB0EZNgsvMeKRkeZ8t0ETRuAfyvavPTfTiCktJWmqT+a8yh1Wz/NKwi3DzqqwI8nKejN
L6P8r3+Z3MoOIpAmCg85vh8j4mXObnevWsNecLZ8N8cKC/VJupVKjJ0xheNB0gg1MF9aMs5enUNU
noKVFihJWBjUqXp5VOACAMxp59RqJOYwz6yUpMbkHxNzSDj5v662Mw/ljGgQoPLK5YWakEq0VSYO
3j0G8Y75xSXUvC71jzRYSM/tbz0G6+BmCWm0uUynQ7CAXsrxzaOric/1yZELFcGTn7pZxl664jaA
8SCNh7+vm/xkkgfiFBYVN+zceXl8dhKIO4FbVw/pUhzK8c2g3JiL9af+yH24J/YzrTl5bbjcRsIm
+BfDBY6fu0YLi57rY0JmS4bQ0T4pF0RfXASzhDBwc7Q08ErNmnPmax44X66drw4baCugHpgQn4LQ
YTINtEg7bFmelUeFo2+dGw5M/ZRbGTDlzBJb9SI9r8RuVI/GN/1Zj0R0gQA3/mVcLSTV3wcZeEas
dIQAIDOWf1NhQ5ElsF2upqOd/OomN8M1uIrlg3UmxMwS0XlwYzvWbZ4SnR2/khmzrgst0dhV4JJl
cuVBaCGCoF/AWQI1lsgi7Ha9BUtzrwLaxivAuvZ2JszJBeGPSkbNJyODTeIhjKhcexVqRwvvR4C8
WrhOjKVltMinz7nJcEcrhd57H0q+kVxQZrxwpk2TUUYxk4+dxGiuFjsa27fPi8vAR5Ua0M4dClnD
0+8ggpGfRtEJ2PBGfo4Bw/YsYsOZI9TbMvhZ5RRGOtIM/jJmyPtMDHItLdRGF0qle0QmvVS7V28i
IkZWuCdyTSYVRmA3XvNHJodbHbb46cCzuG/VsHmk9I3gHK9qqjiXg4WFxmmrvquwnMybFDhLWCb3
Bz+gf/DY7UXqr37WCgcsM5iUUYre3CooMGRzq3mZiVZo2u224hvWf85/uZMqcmUp7dEURNhBFpMg
tQdMNLxyyb1/UnBPjm88EA0lmDHfQwRgY0o7YWkMITYwLXcGyeISWzdsoao0dGalmpLS/mbUd6qk
eMtPb1SWdJGahk2dUJI1OafJViPDSABb3TqpZR75L7oI3ZQfI6D4fJjGoAmvTZUFck/beoQR5rMo
uIIs44ABx6UthBH/pcl2Mlr8nzp7E4o7NItwrLuSqz7t5Xwuvq1LQ3GPjAN62WIgcZnWA0cvFinZ
qJaRaAG3u1TN1NePvxUfncU/YkRfWSJIrEdG5y5LoD4SUqq9H+7vxpof8rmJm3G/HNoFqizmRCD+
YSuUaCFmzXVQpsO++12h3Uo80G6JAQJpfaULir9NonzKgxGABw+nhZJOtwlGprMqFPjjhu7WFDhf
Zmv4IPyb5yJOumHgz17NP3triFgolm/vUgwSJX1tgmy4/mhecOtjJeRMpMWvAx/Eff51sYTARJ77
WRdYzh/LZhkhfxnUJlLwXAaWYqlvWhaMbWw5292++OXDw7ulo5TBIbX9u+y5JkWulVYOPPHZJ3U5
Cca7B4mJuYqJPmdvewOydOtHeKzw5TRpDybik3nUqD1ph8Et9v0TZvxIAQeSaLdLSDBkYBZWvR5G
ib+POfwboLlKazQJrUFsMCgoJAcZZjijlQ8E/2tfzvHRvv4KP2bDEMaC32VQFLVkLezu86GSneWo
JuIYncZ7IsiomITXtQd7xI6d4ehggp6TULzGg0Di1AYWZP7n4aHRelx01J4AJ9x+5ZowBZbOzFvi
UIzt3ipL7zKFZVm7ZzCfmjwxlM2U/CmnO7+eotJ64+z8tSup+JyK6dJrralN77I1yZvDQm0A4zIk
nRvSRDATad9KTk0c5zidDSvF+2pfZmals7hvMLBoGNRheuwlcyMKqzVVBmrgCL2tLXZvgdMi/t9g
oAZvBC1FQNxkGxjKcYa+N/zJr45Oxcze/NAukwkP/GHxXLVevIBGDZE9FIuKe7ZdxO91r1fPo0yz
bs0AGR4bvuRt99k3pkLutGi/zP2XG+YsSHdtUK6TE03Dt+QTucX9gg/glU8r5zGo29cSQJHgoegY
T4Be9PKlQaZF1djtLTEfr1GzGlOT6M4GT+mcjJHtt4aI2ofLKisk/ItcZAFtz+d46wHZUFA2L9Ng
Awp+eh+FNI5RyzcvHMChskKsNRWcOJJMCTPgwELbyZpJ9nPpzCnRpU02pYGYk7iswCsX4+YZuBHr
eyqzpx6CAkYwsl2aHvR3wfGdDzg0yueQqu+GETr60B/IMlIFyy6MfGyWE2Q8Fl1n9zllCvhDZ97/
/TvLCD/MTP9dU9sakpd813o7rTD+By0uFoHashu/UJxTlb/po1mfD58oz3pAdnjKotNl77Z+CgsU
kPXZnYjmgl3lJ32uCUdJshtvm0U4kGptbR4Pn+Ham+Rah+blaTKFEFB6Wj8kILjdVjpz3iuhFZ0M
TomLIprSuBCcyjC0GSBgYTOsRbAU3DbUoBQ0z0jQVByDTsLIjRvyTusmgQVBp+UBagowS2ycWnSD
M3KN5Bo51mv0ZSvRy51aqcWGmkKO5c38/ekgBYzu1ahQVXnESvroS9/ln6cjssl31cpRvBwyrk0X
3Jq16rMEdHSiqtAmwO20TIu/RAasDadZRjFgIARmGtSC0l87dkSKwf2ujSSrWU+uScruEID6JgIi
kDdU9s2BwyrTecWPtK1iJmZsEIpaTLQa+r7xmj3b6RfBRf21z1L4Wdnr5MbVBo+mFfn8IErk07jj
+8MGVTGmZMMYiAbTf1Z1cn+A5SdGSNCcUsGxFbSJBEGopjjmu8Al0s80Xocqkp0IMCjJ0IIaAt75
N4to0jO60WmqwhTj+piErCuw1VpyWOHNXG6OE9vPLjG9c5mA7Q5oYgtkNCc8I798WsxdjPPCzDt3
i4ruSO9jXyJvlzokDpaMKcoq/ciMS+ZhYF19VgCrhzGfuJQff1g5mbJS0KGi34CN90XfKQ+Vx9xH
PfaEGpmZ8zrge2JgJ4uuV32BJfHCbpkeuoYq/Gn3VA+g8Y5AHAjv7OcDsolUSyQnCP6iuDpT8/qZ
3F+KlcP6vZnNk0dWXPP0hOZFkjOvKV3jA1hD8jHLp+DBCc9anZmoSOM6gXTpnKYUb9rtfqgUPdpT
ZI0EBfVXq/pWjYmXg5g9S3buGjGd+TKwgW1Cjs0kV371WRTbRR5nl31ulGiwm6e3Vpcuv7P1lE0l
ddovKxsFpuJZjfwR2pFR9ubaLNgPa3GeaP/KI7x2J1a+6X9HPMYGLQMD8duNi8blrojBhA+Zgl9b
D/YoFLjtLVgbKN6lfeoneyrge5vP1HPbyyKWfLMky+QF1iGFdTwXozdVdjJpDYi8ZkyCxi2xhG9n
E9+UocA72o0DpJuR4pRtguIWDCH02sKczyMQYs3EWLbdx2UmpZMtIIXW7j8SAFqhVxtJWymVU0rP
CKtR2PmuApskGn2oDFjP6IPFcU/Fi95eqFy3WpJI8RqLFB5/5uRS1/2gkXKXd8w1ICZbfwczdG4c
JF/pyOGjZd78/E6vs/8L3f1TrEBVsqNvLhQZgwd9Oi4Z52VIAAMsFDAwUJ5e2td57bencKWH0mYA
MZnpsf07vohKDGd7eF5d4bI/5ya7kX/04EAHS5z4jpUem3+ozi/fWOhUEqX/8diW7ljWmBu7wQpM
7kN3c6b1mDFsTVzCgOmHsD1RO6xrF2nA5wbDQ5ScIphJguHp6iz4rv+G41cceCZvIOeo5dxcBu0L
Iitugp0NXWfP3PAxBu+pNtDheL7YTybywqnXunrlGeFATelcPvM3BdgSiMmAnGXE79Tf9C6ezrkD
6Fz/2zvoNtWcXihW2zNxi03+6dQoaFcWUt7BSzArlj8fTLJKT8WHLXDtusV9wAk3msrPj9r6s3fy
3duMVhIa5d3qBKyZzdoS/ssxikzJ5MTbSxWw7N0954x0sAvX2o41I+Q/Ghc4W9WCvytnqwLW1hCz
sIfSkt3TuHF+OrYgO/qsi2nqTsBQsizMS3ysma/LDUeUE8354P72/iaHOfV4ennu00fW6hdn2ycw
Qn3No7KAzUUep4OAMLqX9WSXrT6FWp3htMKrUJTwbfM7VsjkLaKeSmVXI44uNjqn/Ish8U+DXGTw
R7JQu/KsjAkdIa6uOYgDWQXfaA7aRRCjW5s9fKPC2pRZtInkRC8xAy2nLmxG5ume2tSSJolCbRM+
buP2WhliC7RLXa8eV4huC+9k2sDZ0XDY73b+YaB7y6RivIcbqukvsoNJWCVRgpJuiD66c8poXs+u
lHJJHFOBcajsCoIuNUHlVhC7UPQC/92ys0WZ6W/FAtgXxpmHKQLSwzORv0EoDMz3FHVhOMrrGrJ0
9tHuppJRdJx6MPG9fCB5g1PwTJSnaYg098s2Gw8V74sqThI0JEyIB7UvJwNKYrIYfUwWp0VwidRV
iHkEiNgCLA78eYTsLZgOjqJp7XPVZmtqtlPp1LNcRpuG/lWse2uz0FBU5rmZO/8zzoQZnYGpcwua
GMrilj5wSlU8sx3EqoWQByafKfMX7HZzKltQLLaoo8XSH6UZ2db9Zkqpng1Fdv75aKdrrlN3XBoV
RUNUBN92mNsL029Mwi0A8LiGawjAt0NB2MCzpQN/Qw87r2Y1j9c3SdY1/4+gYQeL/AxCfweKeNy3
6IDn5l7r7jidqxVSv0kPeyq+Lw0bO8TCr3cLecgnqR1BadRzH17S/jX21iDFYbttXE7fUWeXAmK0
L57+rg/KBtA0t4WiunAVn0R/RqB0R967XYtjQwtbOM1+JNguS+oqwq221ZuIjnm8gpnkTjqrFjuk
QFD/2Kl6mmKfPUswnqpftbZ9SDypnwdcJZhjta+O1ZOOn+eh9xK7O9P4lHP1Nr0D2QfzPb+k6Jwj
aE7TgUx31I4P/xeEgjV6McoYURLMXEskm8p7LqK0yk/Z5n7dzWKjJvSiCmYVI7QejNZTXe4y6DOF
sl3yl+TUzBnaiZXK+h7/NWnrwK5w3N7C/FslOltMK3c7prVxF6r1Tc9WomTdIREq5H4U+LJV0EBm
qPr0Ci5OTLQomsshinOAPzDkqsZ8Xn/H9Q35Wf7c4/gNl5mvX2O1Z56AOPOSmEDwBhpxPgiRpPKJ
zkI95VEr4O2w+6KUYAdUPOfgr9d7rsLra7MhUW+W/+THmNqyPDp717QmPjvS4s5yWDF1jTYXDBKw
IIJwLwlAM3tm/tZjXf8R4HIzKlZrSk/Be/KxRW6T+FgnfXSjsgatlvf5hWmbwQy081/0gBi0wCOo
Ss50M2bd38PwJMqro1mPYtustzCSPPIWHHosNMRsNhiLQige9r5yLzrlAInW3lFnZ9HJ8aC4xPk+
teVA6cn1fjk4oZT8L00az5lJbxZDZH1yaUx869lvQg5CLbFuC8AoYKKyQ2FeFmz24uAxnUhzHAH1
UajS3j70c0nNwX82zhQQ6fZpa4B5SbV3h2yJjA+rlBq9WF4SQXGR7gKJLIPPqKajgE8NNvSWDD2r
wT4UZw7XxtVuu3b3yYxBoWApU0A30sq3Eiqqh7ZGiJNXq6TnJJNAZYKjxxIXyBlZ+uxIeref8RcG
2I8b/t8QsQYKOxoJjYywTVnSwcUxkbk8V+NuoCBVrAWhDDB8Kq4CdMLZ6I0Seu3Ac1ck28RJ2wl+
7sox6hwu7GaCLvpawKE1GqWyI6SVKAV/Z1apRvooFrTq7rSH48BOkyiPF6etovXvhLLLmNG7JpKa
VmYypXFUA8NkPIqzf3g/yz6rlNtpYmHvXLBNKkySv3mZXTR3r+cOYJ185cJvtfjLsZzcsJHm7DFI
itD57Z8O0bk1d3JlTfN7mlGiadrcgFiBNbNO5RGKAI+EBPUmFxxa74pMNvumk+sx8k/+Nez9DjYE
ZlEjb5hIx3o17XK4d1Sbsw6ZAJK7loW0qmr3rLzsBsV0A9VMMziDiBeX/rjbHfqzqymmoQQZ5/ak
5R2WfHGNep0So5okZqg0qa5JdKKQY83eQxCi+Q632oY0+dXbCDK4aZ+TN5wfBZ4PaxTXzxniBxHK
WMgNvx+YLa4ruZ4PT8xDvA9u+Vt2kp2lMrA1gYXBBft6rjjDJhNKyL0duK4GbFGqTqZUVSNz+Mg5
HIF2v+U47lYMlgvWQJpyIF2SusCVnWS3I9WIkSjVxsjQBNclYiPYSq959eG1eCQDGwTYHBjC/NyC
7SlHdxN/Utbhys90O3WTEVYq0Pbx69hX8FKbdIYl2K2W7Ucoh90FQllqIiNBoIcssATzAHYc0Fdf
B9f1a+Bsl6ZOrHvs309q9BtvY2dTEYVLKN7CUckyg6m8minYeVfF8xGDwPrIMWwdN68tgXcBq+hC
EUCUer4WnkIUH7vOuvCm6DYkSYTvRTCsIHrlixTbC6x/ekztjmx4ckT+b5/qMUg14MtmIOPHF+dE
JyE0ONpMcz/363UquWhaad3xXStm4DN3Y504yEkwEc3y+Hj1Uu/e1z1SL4C6pnW0HXXvPbGC0Ngc
yYliP14Cv6nFW6VU/2rSyfKyAROvQZwWxubE9Cg+ldl4i3Q2gi1rOm9g8o2iY2h/lUUK/XeDp+Rb
SI94uS+AM5MVcFY93gCtXMWxE5yZCN8X2whLLwYXjYb7j7nvD7wn466rbOgI74eeyADL7Zj1zbeB
5i6H50Ysy5G7cYB0SPeeER0n351DAh3AxQ/tA7kMVhxpPHi4joR1lxPo/curWinb40LKYOMSmPXp
/KaBvEc9lOKThS8wGDekSo5vcJgKDk1VeSNdgI+6bJZV1tP6XXJjeQszeFSq/PHgO7onuWQzT+PJ
5rWtNXTZr9A6fWZ4p+tqFG0KthBv56VTVPf8bx5lzCShXX7eUXNTI87ENMNv733pJxQLVC9Gqc+2
6Kk4EKGF5VyBgXgvutMtp1WaDKRogNNm3BXJ8KgJjqmzs0/bYFUnjc+bQvjJsKuFu5Va/qH2RkEn
b7+6e/XpBfWYDinAxQe3KioZax8dVEWpw5idSldt9iI+DcDamTA7Sjyrxmr8VoDG4v3DkKIucptX
Sxr8Ly1bPvpYluOg2RHkvxuYQ+a9PF6EyKFiobVv/aQAKSFatros4XZgTpU8Z3EIM0knf0zBmjIe
Y6sQDVj1Npf6v+Nj+7s6Jq7PzjvXtF/ttffhy7jor11xLJgsj7Q2oq5rocDz0GDRygxcD3Eq1DCM
bGolQDeacDJP+2uggdu2VzXfiYtPFu4ApH6Ls3orgqNCBhh36y6ODwglWZ/G3WXLqf3Fc4eUpBU3
mv1g4oDTAH3jZUINc9badtaDGyJsBLQsoOqWQbQRwlvsFp2g/5QyTO114hrcCtTDiW7GhVtmW4FD
5X3+nw3l4u3w/FY4nku4sEEqXmN/dSSEYTXM3L3kO5mD2BgSNejadAWnJAivqBBRJk/rcPLiFqda
UYMl5uo+auK6FPFyPC0Iu9v+InNDlkptLPxot8CisL87myOQRhhXiUd8dRrIVAiSnD6DoP1h/B2Z
+HGsPyzoRihGDIwOG74DO2jVcgnvJ0hOAhgnyCPITiv3IsSlAVDhH8m/0AflmIsj+QDygfWsqmyc
SeHKRLl6xtIhSXKixnb9vkS7icM+Z6FHD/ziOo7RGEIVoNHXslML3SZ72GFTjkC5zIC0iZ78BG6B
g7Kdd85FiAkjGDLK6W/DBmUwnYImZMnOTvLSLC7XU4wM/xQS2EOAs7q+9h4FqWhapA97Tos6Qn7y
CMPLStRlaDI22sOqaFAoMF37QD4JOoysHZKkILrIxDfnEHqLMwlICvQQXxZZi30uL+C7rGNdu4mE
McXsBPOFowiRI5T+hYRzeRR0GaOx4ntRWtspirZP/VhiNK5SixnL4UJTNApuIpawEwhIB5mmfX1p
tvQsxvqj8wjTps8s9Pqg3FtIsZmnNtu6+xTxcQqtKdHUVyTQDTuLEOli2+fVaB4CUfYNeu6zscvy
jcsUDnJa74qg/8x9Spl09rsRXxLu4WCYiUtQ0+pRo1Ssragz70GKl/XNzj6IdNE+wywfyemhHzT+
H+9MfJH8nIYLMkOrxcheNX8RBq3hNi3FsloL6UCEzm3dV0XC8pnwuLzwitlTbixUhRByBhgqBDpq
L8x3nDr7wHkUih8c2eSdJ6KHlx8s2qy10Xw2jffQh36wFTd4m9HKiIjIG2i9TvR5BzETFDyKzosT
IUaFF4seWTy1rueSkCylpa7eiU7topIcG5/mcpQksvVy6vmCQRvyKYAWmJKBxnjVXqrjBkAz7w0B
wInD/AkYa0QLEf3wBEwZTy8zqtLkJYSxeT4VfBsI9Vmlrk+8pbXyUs7O1tJyoSn4VvP/8J6Y75AW
TfiP2zogsof5coJ3ogc5HeqznpBYdJZ6VuxTjnZ9I27rkiONVB955O5EZXU/mWT+e8i3LH+1uHKe
ex4Tqd7lhNAZt76XNIaNt1NOXLWQQAKsx8JyH3/qXEwiRvk+jFYtu0nNyP1Ky5sf4ibTZIuLNwup
MT0BdR8+euJQ6iaOfJv8FEs6b8JGn0OL59FTbXQVCbpLJqTfQP8SCbx/zWeblQwMRbc1W6tAHQ6G
HfJ9K9m7KfV8Moeik9+hnNEuexRXcRpMcarkJV/jJfxis2PiOL3TXlQfrDc1BD5R1ejDapWSO593
7eFYmm8IYQgWt/jP+UC09htTlu84rhthCcCc+H8jenTE6Pg2WLqajOwBOzq19nyatEoAcFnS2aJH
bNjvryYctUNNYNp4dzi/Yok9hxVs74l2fcMF3RhBBG4GZc35tD11yiqhbpCy2y22XTHIQIqzXoaN
p+RMzasnTyoovz7r0wL9e6OGECSucZf/dOlv8tj+KwtEk+AUZBUIrK7Tax95MJl1IReA3y7NGB8D
6kpqV7MI6RwPzFyAkY8obfLkSQK5IRSuZmPOoTGmWmfxeGwtT5fOAN8UEUM58qbl/KwPzqqrHFld
j8nfHwFQGIi4Szra86CtRm0heN7HtVomlw0R4Td7PM/DyX0SAFpeJ5y4luSz+ESwiUPrSKwkcVDs
gI2gdPwdGeKepx3W3u/mTR5ca4GDMooR0vGl1M32GZ4Hq4yydq0J9RqBRz2IUSd5R9fZrFClPCpI
FwPKlf+lK4+x/K4YdVLMrFqyIV4ynHrmTxZoK9PtP2VgeZUk4IFQVCXVL5dWvGR9s1urjhkHTOb+
/09rJUioEN0ZW6pZhHfZdt0CZt+TrGGM2eboDkIB63K7V5IpP2Rv63yGGeJyfKcRoAGm0cmsqqiq
DsY6/PTyRSkhdbqrvdW0ToTPR7dBspEMwcaIXen1Va+o60TKo1uoWV5WCi9XCseKZ5Dz92G+zJhF
zV6MhYy4UrVcpI0Z/B/i/N2w05DWWpM1DUUMW/ZFSITNyT0iklWUi3nH/R9GT5s1DdfX8+W8kNhN
almW/By+JYYDjDBg7G7maH2cE/Nb/BgGtbrFlN8Vp+iZqzCOkuV+vFDi67eyGdzomJbTZgxYG9Sn
1mb4KzHZ9k4BK4NmTv70KOKOkMVvHcyGEo+2Wb+5n2jKks3VryrCZKKRKxuEa+WJ27eic7ZD4Koz
lG7drEOJ9RAPX+wOWl0durjgXS0uN8IFfCQrUUf31/Iqazo/ggwv3XFN/qkg62hqjE/N/+OiCDEW
WpTBq1TxvDMfL8SGn2R2lsZYZ0ndb7NzchJFSGUfApXijLENvyNZw2HhhQKGhuRTOLm3yf8vwe+O
xibryDAs2t9JaoO1RzTjBsGGux63LYb3djGzBjyJJYANFivvH+kb9jBsaRRpLuhIUo9zsg09KLlb
IdLGSnKC7fPIaqb47hVpdRR+enwQAhzB/3qGediwLFZu4va0emdO6Pp+ypFAqHJebUM+qtoXbWc8
1+ijb4fYeU0mLB8ok7eO6dnb/oP3lxEj54SmLhnnN60y+z+KuA517P7glZcnqG114X6jpHqu5sAJ
CMRyo0tIzPwqvByzyO3xFU/xdZHbvnxBtP7iUAkcmwsrsq2hbyJnNnhF+fCcXHP47r8JlvC8GUJH
93CZsgr6zaT1aOmEkYbpPJV0m7QOp6vjYscSrCj02KQO1Vw1NUru+sI8gcWk+KJj47Q97aou0Ncs
Huwjyl3S7i+64DqpCG8knecva+/xCjwqJqdtd0P+RuAmgvaDaItML/AkMJDC2sdmcfJ1Bc8vgnzR
uwDvT3hXa8I6k1Chza51FG1wK0JT5tGY8FwsNlsZjmJxzL8x0Kf4XnC5J0D5bNgQpEvvglgZ0tJd
CeMavap2TcXOphVLXNx3mpxNUR5bZfV1fhH99VL0DgesXHzImLocozUhfWCp2z9X/vYzmJlT477N
bhaF8QBONZehcjhgdGaf1oupFP0EzcNdudSwt/14AnKioss0Mlydj3LT39U/e917zxiImW/PvYZB
KQRNgTFnSW9s5QCJn8PgQDGA6PJ63+nbdu9w8edymlp5HKAqndsNnThJS3OIpEwIaImB04guWaQz
izbIDsqGUhIlSU2mES0VoYYLPujdrzydcA0ZV2F/+1D1X8/97lTQOMXfnmAXimkw1hbrmY0PK75K
sj5/kj6smEj+3mFJ8uJvwrTxcoOuPiL59V0N4X5dDe5r6YUQcQwwGcgVkzLjpq3/E/4c8dDOy7/u
dNlmpZAhANUf+1bVbgUHbgI0V/w8q2mGDfRYtSx3jrJDyxtqIwjFyOKvU18KJXz+bwsJFxj8/09z
pSCDHOgPL0VAs+FUy9rRBI4hbADh03ESWfKpox2qnQhDz4X2E+8hbc1khT6cXyhJj98jjP2AVFH1
iYV/QDCBX7eDZOfbqoWitfP5JKTXz7o2jI3ubNmhAr9KNQjs9MCLUp23gK39PeMTXAKcHWDp/Giv
k8ZVc0vUcQ2tDnM9/QR2pKmCdxZqAKqMYckD+uwP4YEA7qY05ZaLzd74bc+HYdvP3DVahY4GPr9H
QV/d3peLNKelYYXeXvnJqUrjoz8Chr3zaqOW+WwqQ69wJNLArzExWD0SQrtNKzWt2ji0lNzKFsve
ra501Kb7QRI7G7yCGyZc0t4KnamDzQhFokn/wGfCor7Y1P2lHZKFSjBtdYN1y6afxorizaaO/nlc
qvU0nnCgVbrUWW1uceNUI2sAjvAytqnEzeDr7oHIjAeEer23ORysuVy1ZQTINQ7VegXN4uQ+V2Z2
VsbDPNSd7Znn99Sd+h1TkZEi84r6HRgiJHnVDIKkHmbaG2CIEHVfv+a3gRCPSPe/HgmssO4x1sCq
m2s3v4Uy6/2sWcCq3RRQrk9wKF+XBC4BqWU/h1yt3tAxa9OGNUKxcIe1zmQSDe2eJGac4UvYVNgT
JQfjUjO2xoNmFYhhsQFH2+Ar052v3S9Eu3sX+EzvArZdKYEFY9d0BOuUwa3wTGvJ/dO2li9Fqo9+
vLY+x0YJtapiYS9NQF9JiM+Xw4/t9ehEcBWh4IV0rRXFyFb3sRJdraT1UGHGIrmMc2Ragzduet7A
ScegzZYesJAQPPk+QnDKQyW6ln/PxxbEMhyQFGj6S9j3wfSpmAJiX+2MzdaYeYF/Qda+iLB0rC3t
HKNSWlVaWrAMVtgDqkjvijkmd0YBEPF63hMvI3RXmvzghlSMqPR3dTB4552d9ncqG8G6TKm1zIRa
SNjWrUHNrmMk9+I3630pxJ1z3v8k9aSU/59SBZoKZGRSRybol/YGg84SEH5902FatLorsAtsNa1Q
Fux/Hjna6kU/Zo+YiSW6X7sSD1GWtxV60CDT9p8HtlW9yfYJKeuIthl45DycG0Jza6Ninvy6Qns3
Jt/eFPrNrBtbO9Nt3lrdaqwmgHy645mgZZMbFc3QHJVugH+UFLFXMUG5oX9gjXD1OejIZZnVSlRk
oW/OIYXG0QVnAtNSUkOw1b/8HuaoM8+2WIeLZC+MnDySP5uVZtGKFRdYwp6XwxB7ndKHrK04MVaB
QqjsNCwgCIvoGt8WQDg57erQ07pqSvs1yy9I6hnYBH7hOV/PqoWIvWZ8gdQcMdmb/99XDsaoHUAl
6h+/azUl2lrl2lkSY/0+nlT306x28EYm8rv5HRQEA0lNMANEBgpZnM0JfHCKZlZVi0qD8HipiR6v
GtY7CIDP0Nxjc8NlRdPSqKR+rb475pIwRMwusGCqzJKkUFHNVbbTl/As7za5LOvHB3RQQMkc1dqQ
MjxTnPG4pO+Kw/DEnqMU4zIgbllcIr8SP+0OkJhGJf4KQDmr9AukD+kYBhg5j8QBQCnzyLlPQGSs
xU75eQ+hlqMGrBmxiRLbZLQspa2kylHJ72CSUV+oN7fhXRrdOLRPKaPBGJNoQyNNA26LyxlAX3fe
nHudGuFDDHGEFCDrLOmchVPfCqQKfPQ4OUmYnGPpe+vK6c1Y0OcZ6fArD/1SVpUW5kJcDuacsEEG
ZSfPA3ygFl4HVHlTxiwHP1M/RvGv9O43YvcoUvENTBg8kfzoyszaBem7/U6ez3MzV2xZtsDniN5N
i+v8PtXNfvLgEpRnRW+ax6tAWzA5P2K2gxevEkpWdHgG0Ed3fdXxLfBQUbqXEPW30xG2LRyxtXHX
ifWu/jNDlVVO26RiU2szvS6JX2EYXTw02nxtB72eV/aoUhPDjj/V9DHwzwNUgSeExcePIANQnCX7
cFa+1bVvX19Wh0/qFnGJY+Ww1R0nyS/+njGmqPiLj1uyWqRtPFELaOY0oRkRxZdzmJRx1nvPCX7Z
3M5ea3ObFQyuxutHuLZPhcEa9u4OHhLnjcvXjuJEuSzL84vx5V/2YuR6PGxXOvipEJ3Omk0O7Pn2
Bodd04zPx6lGc6TXKGAgPGfgsfJNdr9mGnEcuIRWgwd1k92mcSTPJvH6h7IZlOZFvFHhhVh101LS
q5E0zt1t/X6RzPog2LBXhE9v9YxvUhgpNzZCVUV/+rcCTh0Ks/uImKP/gXfIQL27Tgd/qBae2CPJ
QHikAVI8ha/0OY6SmFkc39sfgmnwFfAzF7wQ1WlIssYrU7YSfezbIRnC+7d4PGjxblYflItfw3ZH
EPOu3/PBv+AaNWD7ZeNUUijlmdBQoRCZJrJz+1pEHhx9pcQWjCUZT7VaMiMVl18AqZ56uKIPhHUF
LC9220OMoOS6k0sPhGwsRoxAutUR0gkpo3dVw17DyYyPNbuhQZGCB7F/kXAu6JWZ0NKqsd+/H/x7
gslttbzicboihSLeWVtf7wc+CNjm0uYsbaBRkBZ6G2DCBRB8RbEzUzs6RbcuNlsoMohtOANHC149
WN7gFSj/fzI+xGoQt4nygvgvJIDsBAQGfADw46GZc18WnuFIjvy3Wt0AG8P7gmgcZZfvbRXgJsTi
7MpoSubz/pbu73/7fA9hmB3kNJAdVIkzoDI6UfOE3OSCSc9dTPITHFH/rSk3vau1y8BxBooaI2Ip
khOPswZRp1xuaQFFlXEzts5hSi3ZDmDiQFQzncKF3HDem7nZkTlvrR+F6ZE9+52tf03vWciqmIR8
rwEpXrXQtrhalUBkZ5pVDoD02vVRWmnmdxQz1ZkVik/LYqSqhgJtQ0aPmx+tfdSVNtGLqhLzS4Bl
c64rtbq6yzTsjGplsLmwlUvpZQHmzVycV7EB8n0WSgvwRDDyIneeIV2Ptidiy+7eQUyfX74nTDKs
srMkpc1SNTgv0vmfo1Yw/A3ikTvIltQHh9+I8g9tRd8lAF4RFPF7oP6E3qnV3oFb9ovrTTTAx39E
yckKmT0Jp98hvoRRaI+g8bLbttTS8aFehiyTTQN8jrfng9A+2Tu19P2xDBZEdr8csJpBK+thwOoH
jpTGt203jKuiUhCCfvanoQQ+oxOzJ9WcvFLFCpKoGYs/MjvQOjUiGmY8mAoTSpy4g4r8dDX1ULaS
1qq397SSf/BUuZYMTjphq0Bky4HizEvcB/iO25tN+Bz66+F3h4gOFqq+RPsMES7jJAnrHDhJPdOa
dNMZCgBxrBub6XYmkXlQs83vA3k06m30/ZHaEJ8BstcEXYjiHCRg1BXt35BYUZ4sndfcpj2xt6eC
Duw2LJTIvfn+kCsep1NPhIhOaGVeC+vxD/0Odvc3x8xdS+0qZzEUYuQ/aSCvA+FU7jSrBeR+Amar
krusDUWEf8MLwHMF4vqVNDk28PXR6xg+L6pMKdZL3ohJn/neH54sOhpWY9Ino0Hw45SZIfOONikr
rCFWL2OytCjMpOIdcpjYdmh7p1RwndCt9SIaeSIbREARcQbJ07R+Y2a2RK5W7+YPEQa6dDzNtF2C
kqLYFhB9AQVc13CcM23S3r28tttubOJ9WqcGPdg/9paoVbn4lvYxIrUJhyZT97MeoqAgEHEShSkP
sylthpEwuY5V3wM+sg26wF/Z6/WbL3Sq1V4Hyy6zGjZhVIWtEHTIeJWuZ4zVOWRtCVbvDBkIaINV
BINaDbdyv7FFoDrn2w4/mDSyBdz21F5mgg5j7NtQPT9GJISWatQI66Mj5Gcn5IGGyRQbvJAe2xip
cH/WmDY7ighC8MTxw8PX6QVSz1osY0S87nNQsHzK036Ud+KnLiAt651lQSLeGJqrfvQmYIMi7tIy
O6cksMPQE8o2ofqSxmywcQSm/LvL4CUi724BjAT4S8KJWK0Mqd7+1uA2pNyZ7/GorDLun2FBlSkY
pLeVZDuRRB+f8lFtV1464NvYtos+6bqiKgHEmb854URJHrTG+yPr6yXQ3tsrl1oG+dSpsRJy0ddQ
xwAEzHqEod+Tw4izYFbpdJmGx2hAAl9U5w3Ik345dq/q5obVNECoKqglchFCbBe1yb+Mp6cxioLv
Xu/WRIpUdbpGHkdcobpnFKRWWwo2TI1RKO408szIGqFxfX5xDleIo3JdHR7i7kqpAEmRaZph28QU
UKenUQcz9+qpoPKrG6IBhNHrFQyYZ58SxYTGoNggwgz2cH6w4eeJaNjN3YQcHK1WtzNLnDD8/lSv
AfED4Igp1Gk7Cye7tPuKDyZveC9iqB6bEGQzO2qVVPSOMZl0gVR1c604/DYM+gtf9v/Hkm1UXOVf
YHnFYSC7HWVI8d3XZsVtdE/oqBbaOiJxTMjFtD1vusqUemkXHdLR96C7noMmWmBrZ3wjye9h57vX
7Kn6D4H5BzcV2NQ7ytSdKb8ATwykL7M8EBJThSsNUT3POXgf6D80g27olU2k+TTGbtSq0EQDbiF1
OphM4jPPQdZmDLYaikKAg1ziKkaq5+QFfKWAmWJZ2OW/xxJ8uvz952cKFtK8KSP9HGQ2ttXK6VQ8
rNQy+C9WIwDFvXZl/VfvuAYpTAWOAkPtiXX7jSxI0jaTn6ot931F+2K+AZIUJPPKCGVDWFNORT1p
OumocS5rgi0H20Qo1y8gGfQl5CUBPDwQsf9xpz+TU0ny27RTCvi/ulrPpn2VnwS9QF9XtQcOmMB+
ZtjgT8cSCx0J4Z1BLuHRm9fvVeoL3Arz1sjIdXV1RoKrDIRkH16B7Kcpj+VLgftFWShv9NpgYbC+
3ZHZHmmCmqChUt/U56DX+5H02RlHaf0ypxVYgBoZfsqhdTNL/t36+1ghFgpiyXhb4ujzqH0XLJSL
JlDlQ1W3P3RXPoITALzoQm+X1tBjep6qVOMhcM7Zb7URrO5nM/IGOjY3i0GxZmYxTE7iZ/9kCr3F
1ofhTtngIpFpLEvn8vPNAei86OGsON1iGUm8+V63zUFfjSrMebJ8WILvyGpvi2GlkdBMLMLNgjeZ
0sz3P/j5lHc6Gp2GOrxuyEjVixN5q78A6M8Hr3mw+YW9R/lcaXruo6FZRHs7nOy6Xvcoc7CJqPhw
yArZccuXOgVr6BLp+iWnNsX9YAnNx5HZ110HizSnyf+/X75hMaEAfKRo9fKIYJB8k0yhAOvyrQGB
ZmiLNVD7AsESXMYMOnzWpIOfkwSvv5HhaygyKavwoN8IPHUE3r10wrgVo2x+cK7SXw/qrxxkObCM
cqzu3d/BKID0hAYdhp5HthR70wILTsYnzCj1VE76ifMXvUpEeU51IBu05ZN0Fxy9S6lt5UIXtweN
is/Gr7P+hhLVml5BM75jtQqfk8eC8SZjzvu7uZ0Qy73gwIROFQX+Eqkl6dsZEv4tdn6/fKkL6bkV
zL6W45oWD6Oqrh5UI9KcFlpz1AD8E85Rn9ZKRi23slBhl/IwJZ9tCNeacV/0fkJbdLhYeUxs/7tj
S8/en9zr7ycrOiKQPrZlRIr+V+2/i1hOVJw//zcC37MuBgNnn767m8Vhj//rnEYAIXTA9/cdH58n
cwFCwqg0gs/JqL8g/8IRAh9jtALU6e4akurjCKPjQq7oVv2nw80ipIOydlT5vm0R264NeVzjubcQ
DCel/glfqZRgHM3G3P26QTq9gYQSbfxA4SicGXbQ8EknH/D3jvbuxxlhmarrJprarXDmbwhHgof5
8+S6Znqgsiv45QFK5PCfWfCWHWmQNI7mEvNVQH/2r21CeJShM/xJgj7cYXv137fAEWU9DwUdtl1a
tnGvGPSElqgJf8VpQMOfCekJildfScc0Lnk8pF8NPgBG7DIZt3Wb+jKTUTP2XTPzgq2f6SLZS2MS
SNcBR1f9hZFVooraZ0hhoBUSQlG7BMivIQFnpC1sEKIeGIo2x0W+9UfjG1RulCDU+aL55iwFv7Dk
Fh73wGtQSZNNxPz0TkdU7Rdzi3Zk0DCVxnAeWbzRYi2wT00CvWDWKpYst5BPvs6g56KKr7WvvdA1
kCdvlVe99A3pYandeFJPAVr2Eb9d9xKFt4bUREPHj15e2WLabO+nrELdnuoFMGKPMhdjF5GeLfkb
J6mP9yzZTWIDjDXDyMhjwhDsN+evjflnadwe+d6OZOv51p6toc5Hkv8oTOqRaLgemIfrbDCVSG6S
93pE3xqgVWDafDu7kALzYAk3KWUB72O52Qv/PZzfsEIJ3udnt+8RqaZK+nrwy28Jrlcg9Y8ShD05
at/JWuh++WjyhXeLDVnSuPY8dCUGfQGtQAPjefOENraB80LbnEFxoro5YtT/VGRn3fXPltLY02z1
SJpZ3Ij+B5c/acz32JM6JDeUZ9hdkK0boWRmQhFniH7VDckXwMv4W0mDgwnmiHwL6MZxxrdr9gkX
P63C3+l3ON9KGvRJH92/VAiVWZYLzh15lFwCKWZbsQnTWEBgKB1VnGbso3zlzLmu4BVAQbdrSP9e
RDRBtEdWhjLdDRsEw76LUrgNJJ9GOmi1b1mMqtqB7hH3k6bN0Ejy0cR3hUY7Iizrf/UFDm2Fkr3E
NONL+fX9vfMGBoFSbGBvqUwWzb7xBiME57Gr1o1xS9DyqyDf3qFIk72Tla8jyN/K3J+AwNP1wnP+
fHBCw3C8+OFwLX4FiUwOXNC42cGS8ydwDw6zxCUbHbsfcjH9Zo7p5iKakcbD/DN7WayEPHFu7XOI
soZ5UwJ3CcFw2dKPShxbUMHzAbkmaoOHZ5Uxx24tydi6c2wYxpwdqn9MSj9WR6Gq4QNJ3tzqgLmR
gQVHPhS2m19+SqSP1371syNcdx/zQIMrur61YeLj0NJr290nsV5OqpzL6q7PtV9O2G57ScraZCmf
YggSib7osG9B5zMzklv6786ov35I8USNy5aZvHykZBq5+sDjSSmC0h77uGkviU7tTjBPFwMM391A
O2BBsqiqvjtiMqHLJ6s25/tgxhsUo7oPrf0c6gUCb/O+M6mb2O5ATYRSCoRwBl8oIg+Nv8qCYuYS
eHw3Aj7IgV/rkg0iX3+d++Rzk8k0Y8eDNqqFERKgKLzOS9T1Ql7xXntc3UV9qu4bXY9B0onfyU5t
UbRGQFuA0+T/aPdeaVsPc0OIUptF0GiEC0el5o+djidTudySnOoaA8s/X1s1bJ5vSz35cT6d0eev
fkEK9a14lxGvBVDOYAfwNKpoH+dJkyzF9l0pAZY7j64rEl0Zkm5xZv5a9tZpckRNak8WO0hX2VdT
UcQ82cBy7bESU3mAN8to/FvGZRUjTO9oyZql9Z0x8YPbXrrFn5tP4JbeqJX1oi/WrhAPjJtMn6TN
pmVr33scMgsLvlWyxP/6eW4J5ijuabKSkfs/Gh+7SiNbVzlSS3stppJWeXd3OeLrBCAj2EXeZPmw
IoAjbbdecuzu/I67N5dwJTxzfd5IyrD6NLEmDDSRfwQN1khB/1J55UXQbacXgGcdCWMbLQTklq+1
6nbeKRLoztDLaOKx6D6lYBsmgBVWacg0mMDyQ/i5c/qiHV460wQ7ss6Kd62qAyuCrenvuVeanOti
U/eV1YJH7O2RKt4K23drcNkN2WM0ETG85PYanyyk/5AHASgwneEBADYGWq/WwKMNAfPhkRYJj9S+
mSLSYmfaXHynaSq3ODiDHqPAEJsDsKZV67bfZZ5APRRADVwc0bEyOdMjcWOWsbdAmknBFMeGOF0f
9Wb5FRC1XNDhi8z3vCUNpQ4ZSszywAlJVG8/E2czFn4yB298S4lartZTLzjISHTY6OOVExsGAxli
jAhqF0Pc0TF797FntrFODSEQBvcP3cfAOwDac3nrOQHsKfHfMH7OwsoX26Afz7iYRa7e8pSDMQ/t
Mi1Lj45OFk7a1nvkivyz9BXMaZRABoIVI9WrKRhp8UZGWEVWWggkUdUc9JJGe5/JIQWIoieaK/1v
+YSlZ2wJx7uM531yOf3rqMYqxDWXbuBEjlU8F27ax7zmTdQ7Vmakd0y7MYZOlPD1iK4Tefnwz3oI
LT6IdAFHzBOLHTdqJr4L3rR9inuhDCEA+iUBBYGNLnh5n5DQia11B+0RqD1cetDj15g/JXUSkvuW
bLYL851QGtQn7zf4lxdfmaaB3Xj3RhxKOtgC9/MaM51np/ljzW06rU++fnjjVGuGB9e0ldqry6m0
a2wz3yuWE849nA0Q7nGWInun1I/evwKhc6IM7jPXg2f0aaTPN890yT5sZlcwO+ymPFFy+xDKHQdF
DmtWCSem0mTvnvXpMSwACF0JFqpq/RsaRgs3aWGdb5munvlvXZLufQJJg7TkUSQUQud7LFzycu7F
+HBsL9KZ6VXMAXtp6acooo18inX9t8VjO3HNraRQGjIC6W9aps6gvqalC9EKyl66uqtqgW1xT2sz
Vjxv/yQek/j+YD/gFXDVXP/t182LpciyKkMhwc+/Bz4PS7/9a5TnNqOst/KR93slrw+oZOXtBnl9
aibSNq3l6dFPRYhRAS08tL91xceyYNi+NOohbYtgCWYvtAXnsaL8jPQFVskLyLcJJVx0/kEae4uB
33tlRkB14LFZxp9UnvxE49pmvlqTtQ/kEFlymQKY2QVc5yP9m1hV84SmX15j0IR5fkQA30kGru6A
vurZX3qVY+ovljDcvlIcA8IPRybOw8oYf6vbMvZIDPI5i4x3gCFJh7SxfyZwyS54lIYNTN79sUPD
XAGznV6dzjCEV7gFnqSkbHOMy/1cAHl6RhZ3W19dVIoBZJ4Zsme1EthphfvwudNOxrdb5f8kTBWr
uHyg8jO1EyUjjJIcgGUy3TolDHMe4wK/87xj7JibFxddWKOPMrd5UkJ4mC8fp7hLMZ3BG9rs1N90
/jh91u5HdZbjw/2LkB6L6gNNGfn5b4MWx3+pSkCmJJ5RWz6bpm4V7k+KbhNwwIYemHL5QP8GKBrr
67zRqZmkmgu9IEhdlwbUxNmdDN30HYZxWfZP+XXFie8MpZjcl3rOqFpG28jYCB2R9/VgYCk5N8EO
K7cU1fMlrosmknvxAxz+E+ig2UJbOpWeZroOhJlrZwuhPnvrfDHM7uxJzfkhdrWyNMXdx8wEZnJg
GWNYi7g1TDHdZGbBgnlFhb2r4uXUp6wQG11LCefCIc2+x//T16bXVoLWdBa4YHTmE/FLpk1Gd2xG
MlSfpHPfCfqV18ON5EFWZO9VlB+2e0dCwsdygWOeAYIY+Va3NFa15NtHG1lBg7ECDCLZDZy1RWkm
JY2hy//XaehDWKTdFT+RNzjT8wrBAcPSYPZ/LEVTEJYLth6T/32/VGHXo8p3X9yadYdWiqNz4iwt
4Ovbl+BSg4g5AsW/1nwjZbRaMmYcfqNFNQlFyOwH0cfvQfQZIBrJeY+Q+NJjmPN3elyYq8q90qh/
iZuW7oylvFveh16COAm21sakdHqt8KB1bMW2QOfM6WVOn7ugakzW9X6VzfM13NZJ0VVLxiz4wTqo
OnzOFz+0OGnWTO/iL6ImgXi5KWT3BOILHsaiNAS7jdKVWO4i9CKdKu9LmXbxQt5TJ1gk5A70h0d9
87GIb/XzVRmo74+h4vg11KLQAhQi7Qzoj6ZQ0RtYxUN1HUM8Pg7+OSlNXTJiFR/zxU6M3wWgALYf
BGc04Yk9uH5BKH79qrYPN08NFLeQL+VrMtwuO9PYOz+/LndsQVRC/GCcyRT1jCHXxTpshAcyNdYC
N8XbLnY4k7Ra2UYE70Lc/gEwpSrqAqPztAKPOJLFfFDIuGelIXUKMLZvYLBcAg+8obRe6MN/YtYC
tOWPe5ivssGRgU1HAY3nzquHTrUKiWKq+yUxoU0zWlTaRbCtWzKeNIjf6+G1g+7cNaowpxTrPTl9
pYitbCwH2dyqYwm34isE/PLGaNx4Xhz37PV8qFeh+EOlvJYY1gLAsDHVzEHtDKqablCgs4WFImu/
9IVHTgg1lWIbTsG+zdWrZTbGHS1Ws9OqgFahU3xRu3IJ63+EMcMl/BQ/R4Qz7ixo6D46QlGl2sT9
crVOdt47q5n+7Cyv1I7ygTkdleIeKy1A75eVoyIxHkYwRsCEUcBuPtGt5odOsfst4CRMygZcNzIx
SHnhf4w9KYVTYFtfDW5cAtMeq3rAxvr9lCSLtFzL7AU+oH/KZ3kUoOk5T8PrQRpwtwlYDUxXeNwF
FvbtToXF0qCb64Wc5zDYMkziA1q4ocoKM9p3+FZ+RrmUjANc5eFrpbQ3Kvy9BMtSyKugGE0J/7mk
pXoJZZW3wm+zMw0vTLUm5GycPWfAYJ5S0wDxkQppDrxMXGVrV8eEhX1Xp99aCETCaU6T7JTOTUQL
irpMLW2BsfinWev1m/SS4YMcQLgMA+XWbmkNLnnt9hJZ7bF4K6z+sxDxBqcRbQy+6puSC+NOlbnS
u0eBMhgkjBKyoPXBwrzgzYoOft7P8v16vdPeFfjNN1IiYg0MDDHoO4e5zqeHQkIrc5xL3hiNbZvg
iiQHcA4SQFzbPuUZFVQ5XO3jVFchSIBIC+8SyGp9gZIMaqNnhj8tSpUEzqyDkafk2ebALDVOdbtG
ePHTQAfL5wa4dF14mBrI8tfH1h7B2YHLcG5rnGyrNpbk9b/sacNn9S7P7hCaT3Dj1pyDf7jLTTfQ
9E2fAhnua+RAcNrHPiS+kMYBurIct948Mtd28UBeaNDv0xKNV69dY5kas3xX4pyKHeSd84FBol2k
06MFdwG+wawz3R+gX0XJS1vMiHIQ/NGjM3qC1Myqb7r+JW73EGS2aawhsWIGkfWdbRkx32LE8uWR
ULB/0Km4zQat7IT9ZNJlyTX2bVfOVPsJ4IX+qJ0T7PXo74bFvJPy1emi1/QZZy/rd5ovgSof8Job
MAIqtHeltKa97lOjGzCR/gqY9X3J0jOTA6qsg3CvINU6RUkdH05wcJx0prYcxUQ4qf4Ccfj7XaL1
w8EgMXWxEsxL36Dyu6jGSPUuzyTG9ui9wvSgnDKcI9+nLqR1G22Pz2K17GZEZiWXxSt/qXY/ZYz3
jKblfUpqNCxV0c0YvyfZ0apX97Zowk7XRpddbUlWRHUCaQTrSkzqbfAt2RmuVhWBBXCcR+VxtEcy
SuDt/lB+GmduJCA4zkZVt7rIbnwyKP+vRfcdJo/umzXPgU1CtdHg+uWZGA84WZUFQdVkQFDWH3Vy
IdQLFFuP7UGRxBm4DYxY9pwDBAld5JK/HdzCfSN21TLmfmRYZzkQBHHF54UxCyePB6RomsqQa92/
S7x1WpSTXHw8TFB6ljfaVdkKEULlClTc8RUPpGGZk7IA97iGTN42kSoYOgv0utNUmv8kDYx0MpjC
JoFFk+aKsZQINUqsZSy0gjHs4NWcrUZMkaDsZoyCSilAQq2u+jDfe3simHNOrT4629XO6Gz5A3Bn
Q2UMDw/3LSczb0FnCEt+RM2KNNlPQiYda7budfzHOroK8QRCdGgbnNAAHZHV8cPL/5jx/C7qrM4Y
sd41nowwEPjl5qVowEh/XXcjA382+XUEV5udxNv35pWBQeZrt7xO8w8rJL6zv6EfDhP/UACOkWB/
zmBItdzczSpW1K4yNoxZbq3iMa9Kn4pcbM381EZb0Y1xegbRCy5ygcTtu6dXIPiN94ZGOyFfI4qS
GLI5LNFOXqkHdsCk+sPeniWQBCqcam/qjIeNlwdscEAA5eNl/NuHId91iyZQBfKOq4RZrHCNnCF9
rVp/fpLh2Q5/z9gCVjZwF45I3PF2/Tfv0dZPVTE3VC1emeC0hDcO6xIqd+vC52IXkBgdYl+a7WPf
2crD4SJPqSHG1aC+JiCXzJC3iLRqPQLeD3CK3cTnAzXR84/CyAQfU45+akNGPaYXS7qk3edpyo1h
UGCLhGroNZ12zrA+q7XU53edijH0OzwEXLD7PdEthUw3S3mS9J0lXjgRTbB4KVE3CcREmfJ9aWxr
H2Vzggpddf3+1V8rgZ/mpt8jDAf/S4F2MnvlH2x7K6IFuitklwFddgttjvhBBi3L5szQLmRRLPvg
Wkb31nDGukz+MaAogGJ1CQxTvCsVKqSRZKYv2X/NBazkOC/fDyuK5dVdtc0voXDqsO1WZyywj6FL
wADWYruQ8hmGS7CAELn4j3I6NXnDdOtXVPiEDeNMoeWdOePTNu8GQPIjOScPLis/7cgw5qCJ2Hs5
x7/6g/JZguGxjtPp/n5dS1Bqe5DCrv8Z0sJpbIouTkxIX2HXfSD3Sgl9IwUWeFdqIA1DKeXnoI0v
hYrpr/gc0p/ZxrolBoJT9caTEZ7PHZQ7Z+pA/4yh+NM/KofCjQVI/WWYOf3BJJYWMZJUxRes7nLx
R/dp47CD26lRRpGXZmkZNEdwqgw9uPvdRrp/MMEOTDt7kmwmA5PTFqivhEWvDLuVrtDpITQuuj6A
SGglXWI6B3O/c4aDr1y5UDaI3hzQ7coJurzgAd/DfdSIBygjCKusQPhZtCW0c0N30LflSxmD/1kA
BC/P+tbqKNqpSzqLw5Fki3eKiEG7ExdWs+85B5BuXxhLlte6J6wQpTbjnCVx+v0rP30M7XpjeNOA
RmkcdMKVUOiWVSlHAGAk2N4Z0EhjSo0qKW0DJxkaUhY00f7rmdyNHLnVHJ4TIM/y+69hffMOJeMC
WtL/pWA1Ug3hkL7rZYU1crLD2jhaT+9DkJrY5iCCHI8bwAt9ZXyQkLCITHZhSxHtFLT38GXzXTZC
MSIDyCmmhmO2O95htLVUeV2EJa8msZiTWiow11RHjsEpPj2OYKg4aj0J0Dg7RXCCSwh4z2xifQvt
BpHgfcFtU++1zcIk79w+Rew3Nl7UWfG9Rz9BUmW6laQGivegUOdvJOBnZw3uYDCdJ7Hf+QAabxh+
Gr/4+SptG0ahzkTweLVdJDvzeKOI4R0NCrRIMCeLmdmBXJ3BzFa9tbLdouOsL474tCkwK2pdkyMf
TaZUv0Q0NWN24yeTGA3DLm7jO2h2X5Bze4txqm2PpcaDeZ+Mi/7lFJUUIQBGACXLd/uPMIdTjIf4
ajH3z0XrrMsvNAzKnV7zZflUuyRknYtgAi3LW9U6+IWYCeNr07M9GL0LcEqog+jrfTtEJO00N/kU
yqsQ6+uvkK6RRAYnobQLRPIQ6vJpSp5MFh13LVDIlgGGxi4ck/Bvl/GfHBPtoyx5AnL1VmhCOzEZ
hU3XCK/7UIInq/nsi5c6jU+03XrejPR4OY84UmFFPNylRxe34hGCZgYD7+qnSC5lWtIJRpoJUNs1
Wnd2YISri8XPAkaar8fbk3rcDhOdBNIoT5NLkhCeQlKRiW1UQRn53mkq0VxbKBVCLn+n0p9L5kmC
zHVb5BqKH5NPp2ut/6R9rd69OLEvVH8DQFxg/JFi2D0g+F2xeqWpn+bKqHyX+sK59Vedg2T5giXH
p2xF3sL0Yy8biFKDCrfIKRdVdBkBL9aq0aEEB7Ih6IHj7jFbcl7IuWMz9/ZZ6ggBj4dkX1S1a9Hw
yKlz2X8AathB6KxGaD68ef+l3L9DS9eV9gvK1jej5aVtmfjxf47fLLozFrYZ06ppMiLB/pmG+4Fl
hlVeLCSKeymW2mC1k9PeVmnEP5qI69JXF4KGEQhnY86viFp89NOFR3IEhRzLvZfSTxdUYIg55vDt
I3y92Qnd4VRuRJHg/JQR4Jyrx4tAgedWwT/WrPvf9X0gYugTk9+/Oz3wJy/YeYDv1JAyzLbwOlp4
htq2/Gj7NfZ5g/16agpHMUfeAbayyY8XiEac4TovEf2lVY8goLh0tk9ynnBd3LP2mC9nuFLx9HlK
SA39uV1AEQIfsV+qyRcLlzWq+5sDIB0j6C3wZZMkcN2AadJ+15eb0ijRzF9ImmMsxzT4rcx+gKKM
48yt8SUC2Btdb1vg0mKq15nSE+CwOtRqJN8P1wk6/ksXUx714Ka6XsK9u2Q5Cs8WrYtpaUdCOoIV
pF+YOMZLhF4lZiYvzIWwZoyDrvr25SX15c0yOYxtiuEqp5ShxAKc0TrpnSuF+08YKu+EFlppqokX
xw4hnQF4Iz6FMznHzXaGu5EVCT/n6ohxpp/j3YsOkWFqVMivXz/ncxkDrXfW3xYn3KFwxduWBdNI
S1qLosM+h+bLkTW2ee6ORgtsysNeze/cXVhvvT2qz5c9VxsU+EaJAs3CnnT1WVA9ZMdGQh51McDi
FQY3E+d1sEmV1PmsJILAl3dtr0vIMrZU0+SLu5rIl+3ZkDpECr1+rNStP50rZItJI9QbeJDTprXm
iP+9+oBOdhzAxMgDdOP1cYLJ2WUZ0Z7qQEl8DHPZTfmsA7QSfWwhbnAPX5LtS1A53KN2wS8l0QkQ
45jx0KJdva8D+ctkFVKCGNFod5QlxdwI3XhxwRdYkX4VJhsLMDoj9P3SQCDZtULIy7AMpwmpVUi4
nWjk6y3eW3TuZjeiuWEDx55kV2LZMmFdoo/xKVQuI57mY1CKEKow2WsO1u9fN7KcU14GJAmCwhUZ
Qh+eQ8ZZ8a3VuO0gd5o1QscwWi8flhgdrUHa/1Lq6PLcPeC7MlzAfp1MnZb7UK4wl8Ut7Ds7zqVB
GZBqD0tzhnqTVUJ2jcf5QlQScYv6eSWD/sLeS1SPTG5u7/PxbJ6uoua0QY4m8rL8gpv4jXok96qK
ei5pivvvpbXPXhRy2lDWssTvWoKwccIdA3U2NudcuDojI8ro/lGCq1+l6Aa3juKsrn654Ol/isg6
PKRzGlXScwpPEoKmYWI3AVMPCVM8PMtInuXjOPZrCJas+XxaiiM/8VeOaQM4w5wl0k6+yGxG9gPn
PwGxFfmldD0DY8PRdQSTIvKw4dfQCGzO9WwBst6oGxUHPCmrCR+ebuoh9W6gqK0fNsdlwMtKSOPN
hnRx97wMQgX5ME/LZ5QRQheuX7DzZIB/HS7hnR2VpMX+zMbpaq+i5OtOQqNlipHfXBMecca7so7a
7uS2l/IDKv8Zq8zo6omc/UgYra+ALzgrS0ZD6R+0ol4ymFm4Cgb5hRcm4hBk9u6hGuKpvi4GKodf
R6SN+mRD0Me6bWIyEvJ0oBtMrXknapjDUNL8yP3n26bIkQVrKHzHkFDnCOk1bjJQ/BRyPBTeIidB
KBzqzdkec9bzdVRqbDQtGtoUhyWLbcUEboBPBlyMqpAfJnoY7l19uaYqeBiS2dsy4i3JRF/73gea
NX/1wyEMTske33+70cwW+MIIjKaK5f3bB9p42Cz0cyX2pWR+rrb8pLg5B1KyDpJIrTX3w3p3rGLd
6Zj2MfDn6T/omkWAraDDXerLy4tIQq3BRZB9y60Of0W7SjZ2ypZMMdz703mTr/F97lFjRx+AYEY5
dp/T/QVEFR9AYOeWqwYw2T/+middwV2hvizcSALcWgIvAj2ZzQSp4JjY8pEtbd88XlkTnYI6x2tv
ZmtzaZ/A5VqNqi3eytFoEqFygucLzhCPxaWYaVFiwo5NwcPxvEqiR5Idq3RhRx5SzqNx5m4HazZd
amibJRjIJFvHvdFHZ9aCgwBBbpHz/9cl82cFkz5y4SBw/cpLg8l1eNVlzVosz+mf6H9P0OezItF0
j7EmJ4xq8tQB7jIeqKKJu5w2LLPPrVtfN/wWYSa+ERuqyt+ypeAI49b7q9vkEeXpRPCK1a5YQ8cN
FJF7uzzWrERIgXS5NfUjAIO2UO7shuFIWXwwLTMsi99oo0sOmsA9GO1J6qzm71kJjnDSDSyuR7iQ
SrPvXC5YMd+zFVWwcOTLDIvsJL9SomIKc62U+REvIXiSso9M6gQtgD+hbmU/nYf3CgxiBhcW7IDn
kvTdPwWIz7nZR/J5W51iqJTXMnGbQanxaWMJWRcyWvyiBUwb4N9wE3gkWqijyNKF/TgfRT+XQrX2
QHxDwwxI6+Jk2MM6cW7t6KAowtEK9zZnigLvdU0MsydmzuaSZvRJXDpiZ9+ggNRRDH078L748PQ9
t29q+Vcxu1AsUBtiYCb+QHkY3Y+KIUDHRzcOTKF8q9femjFAXpkM9hEJS1/ztdZ2sN29rjnxQU2Q
YrATL9GHgeldU7U2sd1icieCR0xfTsG0ydISsuWMpT8SuiDvwtS2xc2OUMvcNEqZGwgk7G/KHmbN
tVswLd/0hrIwC1NkU/nXTIYoLQxFXD6qMsVcuASo8hIQw1AaW5yNzR4T0pQ6F/PxroiZ21cjwYux
uCEq+HKvWhc9V18BhXSZYkxU6LzcFOc3YjEA3YgFirYaG/56eoFRUyjeWjJNSg7jMcIL+/63FeAS
O0A7V6itH5oQGSy9xTOrN3WEi+F6U9AtlE8pbei7Bnfo4SKyaCeFmTtEy0GfPa4ONW6CQgFSiqzX
5QVkg46/djIxfo/z/YOT2HsXQ4rPqT90PmgGv5G5+0PMzXyhQQ0w5HaGflOlfaGhEVuDyG8P/beg
HKOM+g0pexB4UOSYXtVLqDPqr0WkXyNyHuUAPZB1erUYP3m8Rq+Nt+GOAl40wZ1XfO8fFbiJ6PzI
RjORD6ZalXpLMT23DxIUnEYAT6FwO6tZlwTT59EFRv2JiBtopjDML/lSku0R2zjyBy3TV1R7/tCB
cEcQ4h2x8XJ8TMEJB2Wgos1WoN7gAkyKf1pnTqYlDnGu69gvI5+Fnfp2D1QKQhb/e+6zPQ/GE2O4
2fseLB6yzspUs86lkYpc20lvOv2sxcJxvjDnXNP/4E+x2jL63EEhzQN7Mp/q8cssJLTE+wRORBd3
FjW/PQ4gTVohm5KVLP693jD+hhjVGjs0teDCXsH/tJM/Qj22bTx469uyhm7YOtXxvUecade7jMIL
QVg3NTot9lcTJU+yo1Tb27UCAox+JSZuX4ufhbFoEwyr3+9wXvNzBP9gJjIOOa9ineJONMusQx42
kIVqMWSQR1qKarj9g5jO1tq4r4LIB5/0YlFFd3h9OOHN9UjBfpda6NPN9wAsQM8xYyZFzmkdKH3J
rRmdidJ/gEI15RDxksTfmzBrtPfB3bUuQjXluuHKtUBxEgWsrw63dZYBOKm1JbXB1y9HRF7RERNw
H6pbtDOEC6dSptNcqHOuqikgoeEuXq9xQ8l5tEJEfiGMeh1uxIcszPbYNKHXQum5NpBqHKCLcsWa
yqlyxljprUMVbttQM1mHoelVSNbFiKJc1Nyh9cuBPtPG4vIgwFJHyuxhSswsbD3vAv0fZurm6L75
L7AF0XBd0GaPsAOpY6pRZipxttoTzgLsMD6EI90ZMVp+7PtoVAZxPSBSqjEpkVdSlponAyPb3qCG
YdVX32Xhp19jOWB3juL1ulbhDy37wGICAk3jeQZdF3bxTbPAieGhsVEHTMO/QDWGX4Fks9RAbxud
jQN03NaSm93fpBkv4eYVgMIFH0xPGl0319tYLN1QDXGg5pF4zHYy7hWhPCHOR4sORfXGz2EmvzqF
4ZSX2T6TH2qTbJ+yNTci+jPnfFuLYRiz5YqU/fn572NDUPyRB4mchE0HBY2+iNO5KCHzV71TA++r
FrBT5CJHLEcxPpuNTmaNFk48Oq/Q2frPiSFsPVV0o3Irmre42DsudF4QkNQX5A83sQbinl4mhFDh
/tWya1os8gX5yuf3/SMO4XzdvVnuUo3T+LIrd/mMtb6IKhkxD9nSRsR0WUtp2+f6lPrLC/3dLY1v
9zwTLI9BCthg40ML4ygfxVeK+iezK0CikWtG9tMjR2dNxZuRb6iarPyQHaxSRl+yxAmNtYC1z5o9
dNC+SOYPMGs1lJ17dVL9v0dk22Lp6kmg8Ay1Oxja8K3RryunLtAqmgaM5IzNcIYPY4Q+itIKvdXD
HrvrcJEZH8OzERabMCJjXli1htuy/+s2ry0L81SemxAI0mTGu8V5SI/eevfOBFTc/VRe7OWL+HRD
Ppg1WUo9Ro3YqObvfRfoymofDSb/RJGM4HCYQ9CwYpc/ZVdISLK/ykOIx+47NVva9r9o1QnWRUZw
oc55oKTMCDhzjR6rUu+wrnQ6hHZGPIS0ZmF8WYIlPstd6ufkuI38DtKspx97iGOlQp9ZuIM+wLoY
xupY80xdadvs/E+YxM5RiRIC1fmmMdXH93+d+r8VLDXB7bld4Co61+jKApm42HSSgP8Cq5c+FLa+
KROSbTQjY9hQoAu9MoyhWgdml1Yp0OoAJ1V0ZisPHVdIrTE8sZRJb4Vw1q1uTxJnAc4s3RMwdNur
9ULhOHKaqLxBlfLg1Hl1RTGyEpD/Umb3MlgXxzDGKNKesF9L6RoEYlkVDnLyLRAdZvVj8aDnpebz
oBjOiLUW3fEN82J5CxdCZdndC3Z+9F5JcBVd5XZ9F7ihf5gB8ZdEGt7qOURMaHjRmFOYXdHvK3kf
l/sOAAQ61ksnAh3HZGfk4NSu9wRE5QkEhkXQ2fZE6vP6tpdabB31QJXRwj8tsCHwMoJn4lS3r4fD
Pcy8Er0Y08bH/B5npJvco6vgXJ1iDDDwu95Zidpp/+5jc0vjnsAFgSJ9XPW4l2I00B+0oJVEhj/M
UQheEfDET6C62RBQb1SRbkUQz78m39+vT30pCbM0IifwMeCZpf3EdEXSYRIyEzP5q36s5NfJct0i
bGxkf+hJIXZAcadC3FO53VV1raQ/N4RYlukbn7vFpNNY9WAZP8e2ja3UG5ipHWdUh6n56cpz+ZJR
E/lMFXkhvbyqrN4q7NEYzHGpJSm61rsxHEZJnuEw9Dg8wisNT+mawSKGmCRGvNoTjMXosl43amxD
j8b+gvr6ybUX430zEZGN8k5SfSU2rVOWQJNwphQsf/syOAOmGCQ6V42hdMeMbmm38ikifuNsWtae
JACDv1IWoS4twjjYkxrAOLwZpGyfFEgN2XIKwZ1za17A+3e2ogdeXaTo8fiJxk/UZA6CuWsP2UOK
7KZGrnEKYk8hOYdpp+5bKoqPRlIKhQ+25UgoikwqN6d66tl5hlQ1p4sdci6NzjqxFBOAuuSrTxEU
zJswvJdeG1t5YYUvy2D8gb5uKyNhAmUBEUp8A+6hRTlbYvdvP58VFLBDl2nwBWS9UbGgVyu+FU85
f720L4Ov8Z34re53BaJBarC3DY1iJ83ENQxnhRUvojF3eDHXXGKbUB6fVc8i96kw2ii9PE93AXjH
ETapRhNv8HC9r2DKLpyt9C3gTOByfE2q1veq3DknAx52pqxhF5gqHDBGTahyDl3V2YmIyISJB2ST
k6AlrAUeyi5fnOsJhZWnzjuUtRZwIyC1LdmrRkpTGexmmUxAn6F0heze/dJ32Jc4ZdFMhwzLAH81
zTeZcpL6raPpqtnEAg8cflh4E9YlSRFFhmVaIjWI5NFJdkbIFTwF/1XmxBl1BcRg8Ctwm6xKOD1R
ntTMnpDWbjqOxBlf99XdkSxf/yDnj2wGjgvn2xNsBJz8fr6yC2WUw72nw+qVxsVTIY6f8rIizBQw
vUiuYWMt2Ib6LL6l/ASUMnuOpg9alkrLm5b2Ta9XYKGHNuzjnbKZxkMl3LbLlYWdDRz/v73leo8G
jRwYNUtzROoZUzo8iJQUKbzIJDx9R7jZFMM/bTm0Ohb4t0WGHnDV9QCpBDrp6IxXCoZOFklxujBc
Rky/Y0FV54yl+YE7Yy6eJ0QHSDWivjG2+tLAHUtQcg2SJpmjvkpzibuMD46c5DKEogAAyKeAs3gn
pxisN6mVf3T0mvUKwJz3jPg+iUVCBkBZxd9NrKkVWEFVUbeQx+UYWoJzlFc9Ci6Jo5fso0ddPevz
XBS3r8oRjsPKOM4sOY2pezVcU1doboKC1QlnhZ0OC+o5QCAouMEZibLrpZl7NjE31TktoXflwaya
j4EWasgHOFEH+PdDFnKCWQSWp3mDN2k1ubfz/Li5Sahf6/G4vg7nnxpDMaj2RlIpgxUVMyS7G+cB
2qT8y9SZr7Vlbi3VjgZ3iZ3lo5wsyzW5z7LUkqG9PLmHzczY7PPI0xh3JSFfNRa5bAFaywD92SXx
NKStfCLC44hj5K+C1JkUWTSZYtG5ah6eS4lU5A17D0+/zS6cl/qDR4jfrpmfqis/Tp/8CbYGKgeT
Q0qVJ4GMWIBp0rEdJR8OCmUkwG0DExcz+LgjdtXs2NjDyDW/fGWe+BVApgj6KzDouBkipjwupP0O
iovIaDmtB6zDS1jTFoscfosUv9e2yk4BEwlzeX5u9ONHyG9KlO7IfojFcfrrMzRh7MYDqICtYvSr
IP3ouZxV7gpRVatkduEmM7gtk6O7FB6//ybNWo6f1tm6IBovV0JGMYa35GnJLYhsRTv2j/nGvrjH
Y7q1KaKRk7Lig7MIB8/s1MKcqr9Hr6bhtes80Gc3DlJAiaHlAdeiBrgEBwE+xjZpndLoqxdafWTy
ilunfbAzd5+7hm6r+Lw+4xfAmFHOoao/Iqo/zpoXP/WISa0VZEWXxobNRE1i4QH0UgAIK2axiigD
Q2IMzuir9vxljyMWmiFpFSY+xgVOgx13CoKBaQ4+9H8FvICew/hm8/IHgi3mrndbUc9+Ipn7hyDD
iEFK0LK0ITWjtpfJv3Lsw+jsK+yooDUXXWZcVlfjjqmaRDQJM2ydAI1Uo9Kqx8cBTmGEe+s+p641
e68wXnNAxrx+cqd7UVbvceF0yJg58RuEQfk9I4VRMnGJ/p2x9SZ7tSrRHIEriZ3JbvmQ4sQVoKbe
95f5ulAMNzkfTsMa+FhsxFG2TKMa3zb0lz9w0kiha6keanuKocAnUhCBG8S8tfuzoyOawdkA5K3o
kE5F1z8+LrKycZAWCiuLeRsUCUYkU7DeCXXDDOYoWG1/Syo8aOh4sspl2E6qQOVO4qxW4LAiPFC4
kMvypDxf+EhO5/jLLgcv3r1/qyuhC24qXFYsu9dSsJ4ieSCjrRhUFnaWn8sEn97XfUpU7w/W5EWu
s1ChMN3H3LuJEU+dZ5neZhW7BftYs99CJJeG0FehINcGzkxgmt47GMlrx+LqcuoeJHfM3zK2ojUA
0EI7/XNd5hDNW2XXC+qmo0pT0YykkYGExl6ElDKpVel5TOBeXO4l2bj4zuQY+H9/zVJpdZAy7L3n
O/snvaXNTZKvMTDi/Y1rdLZ3uWKiiy7Ibv/Qb2V5h1kMuEC4Z4J2Bwd/Mjl7y+fjJFYld/4Ophsh
HsIWF0/6QZo71QlXagSobBmPj9R3sGeSYu4ht2/FRMXfyjOio2Mf2osAjzkDt8riO/9IYJVuh7Op
MusiZOy12BK/H0fF5NemaM5O6f0YQk+AMSHhn5i8WNwXKm0r+l9h+tIPN0mOrE90vhuDzHUCvJS+
nQ2v1yHDuDxCTnRuxrvm3sD9yceAKx7cmYNvmG3CGx2yoU1rr+Idn5F20zxfoDvpGVw5ne/h1axX
IizZdvtvp5IAkZtHI5fPPu0JK7HcK0JRbUo19wePHgvQNhr5y79yLCHovqvFth345964pG4pvkaN
hBaQiPqQjUT+wR6MgAAI77SweOc/6AWeZSldLNzEPrISytBXOC8XYneelas9iB6tCsZW7JNKipJV
KNNeYTASHu7QOtBbAfTFJzd68uzTY5XZutCnPDw0Y3YF/pLMhu2+ZOR2l4FVIWF6dKHc7HnX5OaV
iJ3ar93cVRsQFqpmJEq1cI45/L3yC6xA0kwK7BWsNuJQN6MbmR4TPUJ7dKwCYvztYCqNcgyq6Foy
kVOvPZJxnbwVa/jambwlUhA6XZvkJG37UKP1KdFnVgoqJmlGsOb5dEyMMfAMhsr0fVSV4GAD6nLc
MpOE5l0261CoD1HvelpoyZaQ66PjgL2vH39U+xQvCwudAuNNW/GV7BZtTWkT91GkneAlWJ1RqgGL
6xKc44k2CIEIZhmO2Q8pEPLVLWNWH0qvWv/XmjKM/05zJp5Etz5n+WRkG1I9EUrdVIFSAJ+/d8+T
HYbpEOUvX20kouZRz3APCs8ntFV9ls430RHeJfaU15qaScT6DiVd0e3sG7Sx4tS0ZqSAxWDGbq9m
7NlJOJ/K15UcULBm8loNClEoke1gcinbxKi/r3DuDVXEuT9ZOeqoUbf+1fVwOC8n5JtmYQK1k4Rx
G8wisSgvn3bUiDE+Jkto+vwcDCC2zKkz/paj5rKE0bv0VTkmm1wtAvodli5GI00OnV3s0V/jwtbe
P/WmIy+qf/+mFPtoJyCisU2QvgoGey7unJB817x43G1F66v0X5GZ0kY/Q9WhHQnV/OWI5LExaydW
9mjCIKGg/1+JDb35S+3YDdtaIrn5Gp2LvnQvnOfWTnjVnqWVuAPKIzUdI/+0j1C1ITwhBvenrYQG
uUmrPD+tWXhMRRvbK7lNZmcJPCxLmPED99AIHfTEVJFT1xuAHf3E8+22DlCduEU2v36NMobZqf5n
V7siQve0kSK9H9yjMR+zLcOb97/uoreK112ZBW+Wfx0jpfY3qWX6cIJQWK8F/6ZmIkV9OsABj7C4
xncWzXAZvAjI4c1QPDw7xU4aF3+kdChA64GCUyNlcVnAgXOZhIcTB+2wvtrspJnrcJL4Vre+ch0L
3HujD/xPyLdCClNSIcLpHsaSo0Z0OTXVwkUOw2eO8XItMWhZ9fQOS1zrAN4GSIqxtSSVJp5Czoze
fSdUpPw/fXHDidq27PFdh3RUjNLFRnOssiVP++TNDAa12T2pAWc2MtF6gYYK2x8Ti6M35m1rRT2e
ly5Ttox0LxawhbFmSFxuCvuPBJLp0zax6SfDr9eRacjjki9EmAias+8jhFW6koDTQ0MkMa8j2WQm
scEQA0rhviUIpihYg0NPxrDTrLcB6rAYJjBnb1jNi+FNGbGoDeoyN5rIEBvlQ0PyPjTKJWJBYcdn
bmuRoP9EoR9XkwQDvxKZMqP0+vQx1HVGIxWJ55PsR6fNtmtJAxFVaKDhazfJ8ppclv4M7iyjl3/T
zV7nrAmk4YXhGg2O0lHW+axfcB824WTuDa0pGAXQdrl8A1BLG5y7r50u9dWJsZqTSmcp2zuO+BfO
J/aS8ssUEEXIw12INwNHyyVFQQiGnMZrmyfZbKwdTptgCjiVPOnAllScOUloNap3IQpE/36i8LMb
3Q9bBpGFSjEElMexJlzaCTxo+iZMw87ZzZQ7XC51hmpcgGW6ik1z8prTy3GW3oi81Epq0/GIP/B+
Rb7Hprg0YFUsUI43s3rFOusQLYPXrAwYSceeEkEplOyKx/B6EepRpMVq0y2yhLQsZoITDB/JHhej
viXNoHWD9DnLee2lWAmEWvvPPxM9IqZr69yIw/KVGSrjh7NZDrolDfMhpdHFKYjE7ntZH4YqjNo7
zbnjzVnnWF7QV8nh/bQ5rLxC8D8yXWPCxWp0XLkGf52CfsOFv9zkSACPZql8ctmW7qTBkfU1uX8n
q4u2+BsTN8e/iFXp+5DbfjCHOnBnmJ0GTgSd1bk6N4MGoOYgQ2OClFIItajwQ+SChcPU88fDsxE7
zq0/Hnr2q529em2efABj/9MgvbLFCEQBZtSw7a35Iyia2HfIc7BHSdmSWbqpDiw4mYeb7UGC6eju
b+jY7H4xIX044PPSD0Z3kt8veQR/raDVUXyCrz0xGUxdZozuRunqwGFsaTj/GeVlgHqgrl7VP7te
8rFyAoqd77NG4n6VWmOTA40HyPAZ1gv+p7lMTBo9YalYyTZ1TzYtMP5Kp5PhaS8Vx84DRfFTuoMW
2tE296dX/bXhpw0UDufNM8MpX7Tpr/5LhzGgX13crZF7Hpf65LppEsMVSOpaws8EY0CMHKC82cnn
ky/IXIFit9fvOQtxCF8o9333fbhtpiS08YS/yzegbpAI78Jv3+JyyKjAAb1QBnF2/yO/q0Ht4q27
sa4CYMrmPkY83RiFwwdDAeXDzM7D7ORLWx5JgTpkfjYW+bbJ2ykN8qeynvOXO4BwOmi/3i6RkKTD
HfKPR+Cda8eZTt2Xwddfe0ZZyVcWPfDej4ZfBD/Uh64yoDNrB/0Z1Ovx55UsTv/zZ3fY7+o59ydW
xjzcRphxREyKZlhqjBpoqowdzCy67kQweuxrra7y/U/j3MRq/PO8F43jxhQBX0EKDtdiyZUaIa+t
AGE6sa/jy6vJf0p8k+jDWCTEXQhnqbsC6MWTU1y3v0cvu92289X0abRv+eD/p70JbgeZWZ+xouyN
GE12DWa/zVWN2B82vXwn9R+V/YmvM21JCWW7bzNcNhtPtoj72zUZeXLDrVWQxPWUqXuGa7rXdHks
MIMkzHXQzQlBAJuqINpqMZfze1BVrF1FL2z4Ltn1EJ6USlQsYo+mCYLMCtOnU9vP4831o6DW8t9b
RFmkFalLUrYXi+QDH2MIWTe/6v7I4WsxAAyZbsnhEfuM8eLYWFnx8WugdkCQkVOySEfNVvuUlsBI
QVhv8idgH4rTfDQuhPclBfAgG9ZS3Mru4i7SyD5YBArSd7L1da9y3TDhx7BpgCFnVZIGMWVmhVAy
CgIVqoiLlYCMnp2G7MkazQVvFkCbTzMExcC+kZAoIVwIpSpwWfU0sHwfqqdS+kaHvhrJgUxjm09J
0hdt92+9diIy0dZX12uNZbvW8zU3cv3gw8shOgLR7U5FnzI77xck125MnBW2h0nt8RLM4Yf29Gcw
OsQnybUVBJQncTblfUBmyLEkf5uM6xtHg20onh2zFkHWhDxzcwKjgi/IvVhTOhdXW9haPMbdjokP
7N2B+8fdHpvtWQj3Dx/tveAXDpWmd1h6vOOA+LaiTOMpVUd+qNIFOXVQvpDqveNEpaFgG38F1o2s
5A0yP4frjyDc7WYxn3pBl36ifI0k0fzThkhJ3TxjoOdRuKqk7fLSa63NgsyaO5ztkP2x1r32RzVD
Wghme7oHe+jEfqiYUjXv8lM5ibXe+xGIYf6BvSeo3MEKcJDczz5xhMnrNnXePX157tjUlCfqBo5o
jdy7jbkhxR+1x5L34dO5ilbbhTmXY1xfADFQVvSKH7lylKNyeO4qykYJ1daYNgW91SJusLUpBkeU
XI/26QbldQ8lJsU956E5e4zmBxak+mTYyQ43w7VPvgiZOdNkGQHnHeWFUStMdN+ViAEBqHb0tbxo
e0X3EL8uGGUsFv+btJ8FGftSl8RbcD5QgmlNoAQHbuOjjJHGGhVpFQbKwV9EZVEObBga22rjr9XU
fpJiHGQe9ESBG7wkjyq/cnbpCdvYuViRUZpHFW2rzvLYgBkLkDwz+h0fzxByohr6XNYurvrRa9m3
HjnNJswEFrPFU1XC+1MURFmDBh+oZS69MHXGTWxpPdXnKEMtyKYQqbfFvs3mtfKl/YfhffY8sASq
K8NhkQ7XhHm72lIaW5j5JOP46xagz4qdu5c94Byf68c55gWlFquVPtxarw+IwiK6MsOZ4YK+JEKH
WbwkOWVTnJVINIDLeYl/PVHFyfKgkwxFgv0rRJyQhrbXgcZyro2MTA/8jcKdAHahFNPOdyvFeJUB
hn0+4ymeQEizB6pZOm0ZLSIBNVVJX+FdRfEjjiB9g/POF1ZGzv/eTpIS5XRvw0Z5UKDgrbd4PKPJ
rVV2UJ5ZDqAykFYvvQ5bA1/0/OL/6slt6pOT1ZaAM+c2pjIW+Rq7SbtbPtBhhE5zlbVnsEMSBYqA
2yk0vl1NOFpcRdtvENr1+598AEuIJnX6YECnpiW5UjzgvZBMzjdLGBOVeCPPWhuvcSutlnAVKvYt
Noql/JnrgtCMDm+Kao4B8rZdORAr8Xgl6Wjf6DbAkMvjA1IyAUiz1JmMk9UPkuSQZlbAsU/uWEC3
k9W+t62AeJNN5c7RBW3628lmT0psb9ZrCFy7A7pdRG9XXGGCer/Fjk1NzUeVddXL+90jcla4uLUJ
QU1QxqZJ+LmF9FI44z4MfspCE3bpHiBnuSpHFH1G6aCAIM4F3jCGcg2SVTxTxdA7ZXs4Fmb2kGro
dkND/AXgbYvUJBGVwwomadKcZglbUEtUnxiDlMhA/uUsRSSKT4sbCqdFZGmszyDHmvUlagDer04F
bYCuVeHHJjQ7mFswp6BIvsBvgBEaA7JA723/5458CUNMHVPwW/okkeK9GvyBA5xa2uQwzARSmrv3
0zhk8K49MHhGuGe7JI1RLoHvvo+sz/swdzSBNCkT6KAYphwPdDbmMaMj22N4wkh5WYEWYGr2iJjj
t56dWUWo02WV4gGpgwHreEwMSGfOvEROHIMo6v9wnN1eWBWmQmnHl8V65N4y+V+OngLMSVH+VPNX
8utlKJ7R8xhNZo7dmuecWab9bEUsyXE6Zn7h677p775EXdWn1A39JKpTpTCJeshjO/43OWerr0V/
mJiTuJa0CdbQGbZgsZDkF+jhaF/gTrGLy0q2KPhtJ2hZtZv3hasA6Z8r9nVKf6rRncoMEUmY+zGE
+KPxppnukKW0UaCsGbUKKU07RXvbA0frl/HFf+UOA/NcEm9Mqf/hoajSe1Dh2y3UsKHjYpFO7gMY
Kdq8Czl7MSTkPdloO+O+ylyu61d4JYPqwZ5p6Z9CSUwwZFBPQo3Dio/g1+zxMny7VHusDtkchxiL
9itAgraGXweXMTPuE+WpbFjajL6zsK8aUZ07gliUZgZgB94s6c6G7edOeI3AP35aIFgX4ftr3ovW
bRDC6QmQL/rXEh4+33+BJn37aAx/9kZRtl/+ZtJxkiTqkZQWqBd457SG/um4Pn61WqWVEP2cXJaD
3A7RGAwqLOCKW+5QqHGc1egYzpnS8SiDMM+nnr6wo38ZGWgiySjddjcrcxxLyG+NIr0zgzgPP2XZ
ib2wVPZ8AeCbMtIMFzGQnNdRuGfoLZNmAM+wOTg0tt4wcnqiFqR1gpub5qt1SROv0WHXSwUQGMG7
JKwBLTo87UXlkz9gSUREBd/H73eQJWhXEqs5ijOZmLuE5uPXiwsN84TVJy9QUxbj41Vp91q2LwF+
G0vAN0TTdZOMteoyv2Gdka2N5qeV5ZNnFMDketw41aIuUBdJ9Z77R5ytyNT8FIX0lllG2lZxSrjC
ZIJK+6K4tNFDrgj3FXVBF0EIJj+BGBsZ3BwMA7uzfy5diwZAFy51DaFw9mcqlVQwKpiutJU88kIT
OVu1mlqa1SrFcdHv/3rexXH6rlbzCMooZm1RD9opeVKiC8NzxvJlSqZp3wtvbuN6idG/EH2r9vS6
ssyu7lO7Mjh5ChopL77pd1qSXiQU8p3wEvRI3G2v3+Tvbgc1l09ocjIjZmgtriATsRTIJBRSXDoX
gvOPTBWv4hZ176LGWzaTZA2V2vE6sI2evvJu/NjZ9DeJlSDT8KpDomHBPF7M8mb8JGwUTwB/Ly63
62r1VtjNUDvwsRux3NvHzkWAXRBTl5Zkk8KYGCUMw1WLTIBt7CuvEgLepTgdqyY3CCq48QqwkgQw
kPW6s/z+3y6aCzYomJYdgXTK5QcorIAN63l5wgZGxygmyNI7UKZ/CNa0E8ZQlzjo7sX0pnApI0z4
HuEPaYfYtm2A5YAjGVPPwVP2LFbALHYMUpX/W15OXpUV6O/adVE0A6zNN7xW65uKuY0bSGgbRH2U
q4EEjsXt7BBTkC3WsM5VJjjxMYdS+lXzI/GSCGF1FHceVrEMBES22jkA2LPBybzXLMRoHiyN4bM9
YdAfQkSnTkM231L8imrMpMCwhEoULzLkfhbA/3UDpoF13iSBtl8XZ2pfavioZthhQX1Gjguc563Q
Nc/fU6c/OWxf38MK6uol2jSXR2ESl5h8Shg50tert3RmPGjsaaA+NXW/NizXcJ4AyZtxNvMta3Fi
VdS7jN81AnDeNKGyKsTNTZ/CZ6aocZ4g55XEt7UO8SaJ+TFNRgm2Kgrm/BSvZr0Cw44bHwjZe6SE
lysT+3rWX8Qk2E8Gb6xxhJQ88lyb4rGCpRTpxTNka8P2pjXaW51C89PKoJfa4wUxZfLTT5UURafR
Q0P4TaADkCRpyrXAOMai1yQUVHy0wSrX4myyw2VPO3zYPF/b4NYW1yCjv5CNvDvE8qNfDH+XDsPc
r9+sWrJmekr9MyOdS24fMpMninjwT5MthUJujlusJ8+lqlTW0k+nJTxq+OK5yX2P8kTjm671Tgnp
tGh5mLimsDO5cIF9vs6InJ67vsswmb//u3nkXoCR22qke9cu+Lu0pbWFXxNlhrYaxL7JTH4DcUJG
ncjKmHqtDJVJ4OMk6y5fEPbfX9eGRYPEOC1MLBKbd+7q6VjBivFKesVzI1hkF8vCgJa6zem38BqK
vnGEWYbS0zr0bYsjItxSXpCXbNcC8QOR5FvK+7ZFKMQFJPbWjh6Hb3cbdDKDMYNaZm5N6IMM5Ol4
bLi+5T2xle/zynFRC3CND3zAvb3Ivfrgtc7vt04OL27E1ff1N7WMGgI/iJw9xPFUYsmMP33fX8aH
NuIjKyj1YjEc219grWr5LBMovturIdGhC27CSZEt9TRT73gKoc9IDvOtMzCw4mhIKts7eITp72Wh
69d2Nf0vK757B58WBMpLr4XoLp1KBAqhNH9mULPaJ/LR2msxXHvoR2d04tJGuMzKR1vVpzwRdjM2
bcHWtvSfc6yNNKpAoRo4U8N8c4OjjN3zcUXPczIE7rlN6nxDJOd3aFEsRdizQTXZjpAnnM81sWe5
A1ovlL7q427mMxq0BrRrv6Y5CK+Ea/PPnj6N8rxXJJedBlvNElw6lgYgMVH+8GI2bbcOGHj6QM8l
BuedxTF1nMQYG8hC8IAfqMo13oCqI7Gtcai5OMDb3KZ5ZhDZ307GaVZWjhEac1Ea9/+y8KFUjjC6
fRVEJg/aDVY0RW5Enxl3NSDlOE1otqH6yx9sXBPj4raSITn+w4W8Awzt7Zgm+bz9vM1WBLwnGy2q
zPopV+vYmSXHdZTV/Xpn5NIHH+hvm2EbE5zI+V/ZJIZUCu0JrCxoveqvbxaQd0tELbqUvURwzkZu
8ovmB0+4dpou1qMIbAX0Y0HfsjxJT8gsmh29FUJ+XhNVh7+SFKbsLuGljP++lodfGCER/OCe78+D
23Fbsx8Vtm5clK1OofszJNw/7QMbN69Z85YfR1f/HgYTpBZlDQ1AhrT4Cuq//+mQmd7Px4Rhh0oT
C09RomjsgWxrNkAQ+SdoQhImP+T4iWGJRNFjZboY1Y7h1aVDUntuMl3r4VUO6dhSIspUY7L1dx0L
OgWOVlWw7g+4do69cm/cHB1ndDgfGcrs5BiQGjmNxTYdLl8MnwfqqBAIFf46heatZxh1ywRlfEmG
H5W9RSmoVfziBJ+tEu0/Klak54s0RCX9MGGCasBUcVaoViw7MpYWe7xXZHVXxOA5S2fTU4THXQJ3
yFRK0FbGFBWLC9a5RV/XQwcNTO8Cp741Skn3Gu7K2ItUzyFdbeFDIdtW+PAVxkIE3Og/jLWtOXDX
YCHXnsvpYZU59OYNalimsjBTpkfyUtgQnNy1BNHmqYTZSRHEcug8T+9VbuBhBp+TIXZ002Czt0H7
DkVEZIpKHxG9eidmIp8tCbVKEWlUcUBhZhB7glWizIT3tKgw/gXXm9KDoUanAYDvq/NCv1tp2JUy
oFlxG8VUf4pCN74PSCkw8IhYc1vI5kriFnmGIG+PjKLpqxVwX946QDBTzHI4k+lZ79xZAUXkog/H
FNYm75KDkG+Xsu29z/j594/igAECCUhdzUjVNOLW9jv0MLuPxkA/0ZBlGv6O3uNP9HdExYWxyRPN
+cwzC+o1rBR+vZQkQT22p2paHliwAykWyn1pzsGN0Rb+MyWgi70x4n4jqYm6mJt/iaP1OkOWeUxH
uW6VICWIwqQa5XR2PKc4i1JT8+CcQHzgiPzYYli75uyQyW1wPC5kovDgfkoSwC/Ej+SfI/dmuTy+
lKfSbRAIZ9MmyFnArLX5E/MptLwdLPC2x9Bs0h/WMvTI4r405IKM7k7t5tJdBhmcati//Jdo2rMU
Dqe2oLqHoHKzOPlch+5TDgYTLjdeTHZFhpXmOjn0BQGSq+HMHeK2P8UqV1ePvTwhmiCCOudcSVnH
/zFy1yh31nGzWCouH6aoQk1/a+vnmB04akufdGBCkyX2rvskO8NurHI3nxsHPPZVQUv7FrPtIKq4
vM6quXmiy9ed7N8cau28K+5pBjGYXuls/eNm87faIlNlN71NYdCGw0nWMPmYlMKHRvsXsTsPI1AQ
d8jeibZP3/e0QVtzZz9gpuH/fGILH4a+6fww8lDQ9eUv7dHf3x5GgLCHOgpppmoHzCLKSqBewXVd
PQYX7OvQtJnt68jrQlQnp0SZm5APf7g7M1Yif3yUBX4r3/a3LFNb+JtoUXRoFLK52+70j/URGTGp
955Aaq2gDTbUGBVTUmXpHqEJ4XqF4UvsJSS4V99zW98vMwChxRAde2mpGhKlWZrX3x/kXd9yEfyq
3N12QeuNhxMNBqn8D2KZJIP587T6DAhfsAFcFoi4BttoLHp1Et0qzkV3+X+o3gMuQr4UOAXvSGcc
/BOq+DzQ5ec1w7yANtE58KzYJfDGT3xY08X8wxCEqBv099ETu0FTo0RTI8pcGloinzfepXLxQ3rt
/S5msg9sCj3zBdUxSpAXW8YIXVXZqxVO2nc5Ip3ZZsWL4SQlWRUkSueLfKqZvO9klrPwJkiDQOWz
Y3YxZjEgsTHFrjhOw0tHVvH+3qtE/SQ9xy8Y/D1eWVvy03jJ/R9TVd/TfUyXO5qjJCEfwoXGOhAc
rzBLPN6ZeFwOmDgVGqGl4moaZstetLgakxa8XnP/2oSDX/66lhwRLNnKbsKjlrzCOv5OiF05TMEw
nzPc5ellz4tiK+VxVpUGm8ANphb7R0CxicgWE2nzTChyu8BEF7xhTOax/GCUYHjkkRQIXJUPwh1L
uM8Kqhlqf+YvUSR5t0mxto0RRJr7H4hklj0KYzs9Mq+7CR6Tu0lhf+G5wAn7jZXQAd2a/aIkvRKP
nSQ2ly5s/0xsDbdOYf4APfCjXpL0ut2MZqo31PM1xjNaeMHHFIv4+rVx+b6kacDr2cRtapmBQ0Md
PjHs2s0Z11em2F33W+h/jEXnD11u5wx+lLnolU3BSV+k4XBoDb1aj/Mv1iFnVn062NOsg5+UNlHm
XtzIj7ReFaE/4P79GnpJOnYivrLQ/YzMRJsVGL/zuQPhAI+K1VKAY5JBULR7U5jq1NGO34+5G+7A
jDqFwnxwAhfKJwt5QqITcfV58V4lCG4J7o6UwGB50XEOBUEOCXQmNwxnBtS+Fs/XnLpFkLZSNBTC
bT6xAJuZFzXLsxU+CoYvyde0ptm2HVWd30mESmxnlrik54Zths9A/BaJeiCIMWcO7o60wLFUl+f7
ghGMeqHWaFqNwaf7+I32jJ200OqgRaCGpcFtmJOYP2nYLLfRugeYInFIKe6to4PLIcRLyv9KH2aG
zi8g2M7EGz6hUCR5nGMNmQFaeKWaYqxP8Lv4hiPcn1uG0GUZy3T9C+faTJdG+luxCZ5otxZZ8wi5
Yax2Mgv/UZ+tuzlibcrbukebxuo06KYD6monyAgYttq0UNrvscCv7KUIlLybbVbf5f8RxdnFV1Zi
HNAa0pk+4I2YsWb2hH9LzjCIwppmJ2dqcJZdjn9ENsfhA071oagVBsuOE2hv2WpJhGAOr84DMt1Y
1c8ozTkCB6xCXNo1wTqEEnuChGV3FnvSboUu6wWih/gjbtA4gqY46C30BoY9A+1PclpaJYqDaiXx
zRRKXqUbxZaJiehbzfIG4vGAT7OyYAhtIFDz7D8jJw+bCegyz6SiuLF4bmZUdW5EVuYdATr9DMqR
vWv7WbVLzBprK7ittT9fprH85W09YVg+sdnpk3ut4jmARKLuTXfvDXt9ft+3Xd5ou1MYQhB3E831
kzYrj4xxGOE057frHDu6JoC2EgqOwphtJixnLOO1GxG0I7RTbK8kke6ys6j6r6I6TyOlKWucOg15
yzq1nnjI1icb224J2Nt5ot82X7kx8W+o3BZrILGN93YfZWPo0sNSRGIqNPXA+27yXEbx8/Tf4JQ2
mbjTUyqKxwHJLEW1wa4PA8f2M3zLG5zqoIyHiQPp273sVdqDtWATjYawJK5hOlvduzn/74jkhdX6
+hNJdxkKl9JAEeNG8su/IzyZYbD0zxTKRCDY6nZAOky+S1tfaJJKkjtwGo9G5zJAjx+aVOuOn7SL
lI3wvE4urjzZLllMk6f5pIJom06U/JZlaGr1jCX3h+dROT/pjTPikOiY/aCil0/r5CKVvOzBDRd4
ZQ55IdC4PbraplnUsm5zxNAtra1FJQtZW6RPavUQ/SHirpvaDNheB8l9wqN9IdcdZyzkxX4+0aaz
5w2HXlYkZhTm9ZX/inMz1YPY//xRg+I2WqT/e8xSh07H0DXwbCQjYMfOyt5HOyqH0OFG94rR/Vx9
Aa/hHdxY/jHB9SXwA18CCQhIbRH5xIBHJXJDFqcRlq8HTwFKt0Xy1Kju/P/iEYlHjJ02vo7rNnWi
HWoPBV2R5ZplSNU7WQoqhyiBxQY9w03+UUDfOy5/erLSDsTaDY9G0RXUZ73Zvd46bw0zyPfHNibq
bQ/B4jTUbHF/jsjEuRAcAfWV2fmi+v5AxmceifYBIeZkw22vJ87VGvcSxNdNaDArWJ2cz/Ch0xzd
HqsUh9KY863TGynPO330ItwIrts+P16FL/UUYL3DLHfC/5ad63wxar/sWLrF26lvfAgxdUlAOmSw
kNEEkMsAX3ly2lHtpSlmqoSPeRqYfHm6MtO0LdQ78neeICO9Y7OUIQYWDFQnQ0xuAqyC76uH8YAW
cwar7WxsWiTjEJHUnWYMHaJ+8ukvHVO6InnB4bnxUvEfKL5tLsGNIFtw2VCLvOFsB5GPML4NQ+3L
90sZUIhXTnrAoKtnBA53HjiqXySDpE1+qt/T0/D/ij/lujNXI+58gSPykVyoPUtq42po3195qJ1X
iHml8Gp9bYFlhTYoaV0cTI7s9zo51OBYq/Akfm4YWGTh9Mmaq9gNklpLTfW5+97MPg6+2SyB3u2u
NvjOPLIuAuq9rpE7hD/AKeDxHCDTYPB0fLFfzo3tuZSlL3ntpF/jcgcMkd0/FysQhuCZIlX/BRU/
b9tu93gIJwnL7jadWPvnXiR1vqRYLnO2nrSmMSXcFtvjgiO1mTfKEqX6tUmSeTT2SeE+6dCyNTVB
xQcwmDJulR1TuMfvxn+1jLGX6R0cz4qHn/333/nBYJnUuE8/eRtOHR5PbcOhUOrq68ZX4Vej3jWo
AVKYtDlp8FmMvOXj3tCUP0mwLt8avnOIvLbvw2yP6zQ+2k9vMimALbgczv4fs3OpCqTVTaK5UDUO
X2EMWmu5NjKbzrpc6HV+eCGeZS9qohwsOjgxtRgyeUEXC0Zdryjl/oRFXUF7oIQOJlF+YMEbY9E0
QgZbCo91MUCkVholA0czj3iQscWqhqSQaRJYF4XO8j8Eho3aPWnj9NxTITulzUmGwYzA1ZCTBVcr
VqOHv17CRuysLdF7UCk5lOsox6m5tY1QXZ9pzPq/nIREl5dvYWytUx7vI/slZeqBuCS4rN3Idk92
IRbOWgpBIeb5C/IVbt6o9tqDlLigTQ5fmzc83zSwYPvDewX21WKVy2gA9vXOkNBCoN4j7Pv/v0j5
3CL54lQVycpN8s5KtXAM0qYA9iBt6uBlMSVe5jeQLbNSQJX7qnnc16K2MVf1ZKsp9zb2dPL78wwf
364vG/FM2Chj64hvilZ1uwSm1yEOS55YoAdP7YBGRRnroVv5NwGRBt2vb0hqwoARzN1osQWUSwLt
dmC0L2jCyizifRmaEaZPuN4ClsGunguVWo2nDP6FM5RWhVs4LhoXVFtYtyXeAJWf+y2BFtPQDCKO
YwpT8Cm13vWtOTbJv0qpKGTsMZXaqD6xhKKETZPt+u2w8zbcQr29sFQG4KIIr8Zv6TFwsMXxmqcC
KFDxtoosMTMovdd6pOjLjF9vqJiI7bC4NxUBZHXXQMy6v9P0pkN3zuCBg8sje2xI7nLtqtB6exic
0aTx/qRkXgs3Sz1fC2PQvknUUnwH99uWbbdYIYYDTZxr7ajcREg/W7TuzYFw5Ojvj/7kE1QR9xc5
LXCjVr5Lk1MMKOYnZ4sTH3Lq59lOp8XWSMHdGkpdZiA6/bJJYQaPqBt8eGsPVaIgS/KNXkRtphWK
8SNTWShLgtEFY0Il9aYuqoPWHv0PSluOgktKS0ihBnOvSvXTlpOz8Y0jsPWHSuIYDPo4MTW2axoe
ouZmRmC9Q1LnhJDWfOu6VHc6Jh7tyAVmFY9HzcVySPRl58VLC1FvI5Ugyrb+fUfqP3MaI3ewO9mJ
gPXbue8db87ccpQa0tp7vzB6NEIi0nuyD7GejfisAor6p7+RRw4mh9tOVU+85qurWorOuNJHq8fj
L3ANz/4UCTQgpFCTSrko6lTGt1ru9ag76BnMeiz2WiEVLzcdfYWs+KIeS6oQ6IRtDdZ0inDT8ZBk
vxaNDGPsyJ8p7Y/uG10PYbHSJ6mlAoTbcWLTan8WUI82/Wa+BhFqjqS3hhn3+vWTug7gFBjXumDI
AFl4AoZVsi5VAccuBVw2gmGPmeioHTzrwNFLLTVc7oId5G2dGfRB7bfzYz8+9BB9hJYCupWj1Xdy
HUV5n89FIrc281zZynGAFZcJNj52XjGUJMXgciQUMgLOZYeLNc9YG2SX/vRo9/KXS8VG4faGwltx
4sHahmpurPYCYgAfx20iSar5OKsY6JqQApT34BXlPV6/afUWQPdNSvB6TXSCzt4oSR68csX94JZi
UgIFenMytlMFplEXHXXd99uXPGuwJ0eEwcEGScGbGRXhr1z7TObqw6y+HI5g9PmY4l0Qm61KlzNi
dOYH9EvVYuOqgffUH3viTAIrjaqQ8BodPIerpt+520dx5mCkbqGwThgCbisbnet5koD6QXaPm7wg
8/dOtq84iXMAHyJzu5aBveOk8nrTU+VNsKUXmHthBSDbskBcQoZ4cK1jGTXxgZbWDt0x/jYXgB7H
G5RIQGNQo7fxR5Bal6F1u74LFk6FCmgUgFsoaT7x2u+tkrE3tcZKLq4iMHc39w9sT9hX+9++SFfj
7oufWsUGT8iLIAxYlUVwc/PbGvo6dPMkPYnlDE3A0ZlKD6oFAEnn4PhzgFZ5oU1l6lo+NRv/QPEj
9LTlNpEINUbWIgbC1veKuPIc36yK1i6JlbQvX8alXcbjTCGtny0uPJEzvVbGqmYJ4fQTyWUDzkeL
n3P/CS7FGDL7Pw+Hjdab60EIW2Bl28NQ7X/9G0sZTpGvIWYOWLGuswC3OtFgculk0Vi3lDLtS4e3
hNk31Am8FRjkWF/3JHg7z3w+ZJJ//iU5EKvjpKMepRGVMkejp5cBjmSgc5+oNnkUdNdxDhZ0bmR9
QC7mLCCgNFPCpRh8PXyWL483mG7Ylf3kpowPbp1YkxCVPEPCxFcGbGdpuxkNUjhvaJx7M46S/8PD
0PzBgXhkIBvj9Z6qsrZiFmr8ce9Q7195kvt4rmJIu0Eibjd1j5vKCZ9ojeD9EZ0egdT6rfJBLRlI
KNNtM/JoIGcsjQKOhm2oqUK7T7ZQ6ClTa/1ZnjAbzf4vIiIOTUs5CPBXWmZmqaIXmlfxoRH5HYaK
GijPhM0qh9uGO748R+na6AI6G42vCCdTildGfCqfEkezldBa2W57SWyTUcgMhLsLEb3bYDvVAr/X
X0wrtokuGIiJELySa4L0vu7WAqlyRcytBqvmqnwOC3oiz/HuwcehnBsv7PJCuxmoYLnxFN61xYN2
ipgApJL6kzdCWbIz5fw33baYf1ojvKbL3I+GUSuGmLxJboEFJKdtREzEhcRf3oj7OZ4RcpgPH8eo
VoC0PYcux0r8jboDXZDFLiwbzoJW/pRmZN5ioKHTcIo+j9wnJHJklJ6ihz9msqVdEUMvdECOMymu
W4ZNX5Ztif2cGwqn7ueWFP4FD1NbOq9RC7a0LYBJzFpMHsHoPTOFYHssqq3AmU7s+SCVNbKPGP0p
xA+PmMAUE8f9w//o9Yano3j+32F/LIkWsKVeYEP7EO2atNIYW1+70F6O6iOFgcoT74B42Om561MX
SYlA3HFJ6H8se2OlTUb0mjWdxV44OmT3E5cIqQxtjT7AbaNbgbvbFru82YRtVPNtCTxNeTXxMy1W
3Semsu9VjEF6/PplSZValBI3KeabfJeDzAgsRI5Z1SboDn1YLTAnXdhQqFhcAMSiFcU8Nv8I0gjB
Zv3YoAWJVNGiDGD8Pn5n//7gIL9c0zEtbTQivU7E7+ZKtTKW+S4BntkoFIwoSblWrHIOB4DWo7UN
MEbMBsfnW8aQHdawIfSUoyO/mdbR5CZP7mgV0SpKzlBntxlIaEiC3v3uSmZ8Bf8cp3kbIgM0maOj
jJpHPVUw7g2nNytWzKQD+fwpSP1l++H4f7a+N3+8pVB7ezhp3+Xu4aiP6ez3POXkMOu09z02xwKg
3oHc3F5jiFf3BNnKExDIMuHbwgty0e1mvVzWU11PG8H6vXFAlykLFkA8H36hn3AXP8oy9ktHmMf8
5JRRBqySl/1ZuD5YsbTWHp2Zdw9S/Xhpum3tgWGLzTkxFZOF9kElYYeT+QN3bxgDnA68UXxM25U7
CjSjVUz5Gjf1s0yymOAi0gLTWeG8anAwunBXajTZAmNZksS2Ftxv3ZmPTNi3qVyZLJZTmSne7FT6
Yj+rcZOlcF7/nmSm0MSwRp7luSAC5SPypIiSRORNxjypbcy8hsGEd01Um8xi4R5j/zcvZKNtyKjI
Vi+mlUhs4N7uAM3Mb17DYi+tdGLbO4v/JJTlcOqGq1cayUoZw8sJXi7c+DDxkpEuY9c9CMO3uAMy
SDwnsUTAr8c8an8slfACJBUX2+2YJ9HGUP6tNxXRuC2J5AzLk2v3wTrqCpjyQfytIaheIaMTFOg8
H7lfwkEylLAOjDYO0PKIt+tIxjVsGTtYCob4MmpdrunJoWJPXkkSlZ0rABn3TkzqpCa+gjair2B+
0EBSsoEFUzR1iZ4I+pvsMVPKqwZwVIMkvANEiPYF95pJP29Hxn/uTR1LA/VXIx5smr9tU3LmYq7R
izV0n0F6ACIWZQ1pDvDAocrYstXfEEKAV94gB2vTBJbGGKnIYg82SGUK7E/daChtub/tVNX8VIAr
/tNPy+gnZuXXoCVSjmXwHmOh2dvMu9a4Gpwr2iQSEjaUt5+lmhje5WiEZXrhMYkpzXReLS7BUgnR
1cfBbSoINCb7fPvj/DckDNWNh0zorC88o3Q1OiA8qWeXqWIEclW4Zu7rnlLBa/7jJ94YVrLyAhDo
VnxSmGTopzrFB/5QDFAOneCjXDIjYhQWoE/bKB/bIbnq33OqTmgJyOhJyA4RYHgCn/q1GnChe06/
bG8QsBuV06a3MnoORF1VxiCJTRrZUjTuF0ge9x35sUZGw371VbosBDLSICyP9J/q101ffIE28i9y
yUUoRWzvTNkc1eGo1U+cpSJ/YcCRHk/Abokzxo+SRxqQ7Zart3qmbUC0VKy7p8/iTnWAp3GHzLaE
RWOXOtqUcyKBNnwv4DeVAWv+lDAhvVnvC0TsvkFqockcqjKauTz81pRSLXWaQs544sI11mmB2xBy
4CFJX6RYlvsunIq8GTARQ5yYZwxwiaQq+oTCj+3TsHnLQlUkUgNbIqrs/CN2WAuxPxarExO+QWko
M+/MnC2AgAQPz3b0DGLPTp8qqGFAr7BWmXE6FFUZ3RDrF7tMaGYpm2Sdb82GA7Tc0+QCnChIrCmC
4H/p/x8ao0ncdOj3khoIlQRM4lc1jabiw3Ci7ik7m/hnqEJxecAGVUVvKtfeTcHoz2l51sC0/nKk
b9dcCbPagpZKeA/IobfjFZQ4u1w9896/dy3K5uFCqJ2T1COLV4Buhpx/56vx2XIoybeteeemb1Hm
PhwS16VEBqy0iPJOlreOQVvbA14jL8E43JxAt2eiCIa7IYu9/CZCsFtL94r20SXDMpx1dc3UXAt9
Px+P0DDNwOe6ZekYfBL8Jdw6cHOiK7CUTrShgmZMRNcaYUYXsiMcQ3TNUpxXxOwHkeg5DeO0Wtl0
rhP0vLz91JuJsCCs/0Ajjx4USenKiUufbKL6HjuzIeNwjoBBFyzgvuPflmoUu/mmZ0H+34vUM78J
dAjvyGmnO5hLuzsOMQ0Ft31F8wfjkjacB+5QKKShZXku16ndccNO2N2o6RKOZUBA2OW2pVjknqTC
0AogEBa+Csketo8xlWEHpO+QH/hHPpAnSjvK6K0UVebJ59PfaJSsGuFLCTrZOfqqv0zNOqyga/4J
KCmAaVFz8o38RHBBxt0ZvDGk2yxCJhztT/H2zEUcaHCBFxUqEsF4yNOZiCXffqdqQ++AB+LRQMEJ
scMXPIcrN1hNxyQfDF4dLmvH59nEvdMTJMo3K7ExlZAbNytk8nFsB9PLM1TG90V0ZKsMr0sldRFf
QtoNrDsXBsIbDdg342471CqKLuBG5SAADQwsKAw/LBRGJfEc7wG3AvJ+TIOddrBqzZgujAClgyQv
/mxtNJUBjde5R/+5sYU9yWQuFxrMKoNU3y6M8ZO/s4oE7lfSHVaKB0sj1eXBzt0czm61Kj5uo571
Bh2QZQiuFZ9/T+WY+Vk3eeu3Iy0YN/ckRfIBAG06K3Ol2RfEKSQV+ZfuvozGHCz8mx98DsOZnzL0
oUmUKMOD3WCSZlHYSdMnpFsLWyVc59Dk7O/0WKjrH1OJdpwDjz4/hYl00lxx1NVKgOREvOtx9HBg
SxxV6OHmPxN/IGRG6ijCRhzoTTpjO7i0lUDQvE63HoYtkiIxlQWITil28oaZPFD4W+xXJQo8bcFO
2Q70H7hQNVPyfhulSdPbza5/vLufaWIL6w3rwsgnDfYyBualMCUNVnws1uvcfsxETe5Vmx4v0pjD
aobqh+As4ecaZmqGXC4jvLPeBhLIfMONNfrEUrbsZPIsPYxMGO8S+cG1ZjFk4MPzV5uzHLUkM+v2
PyD5S6G0JF+m3V+9gMCzMNLmsylKQztUQsa4IdMIdx9ISupB4wit722zQDUkuDsC8oMDUBcNJLix
JG0XamODzUx5YwGDw9uVN6NYb3UHQ4ieiFV7JNmeckOmNq9kbHURGxgPkMbj1Imh7EmT+YNC9RgC
j2n5cQQOGYmFCP+SDsnMuxLk8aFOIu36ypl5TjNagF3x0LstMt3IazJsvhhAtZM/ZkagKyWc77VW
L9Nmlyjq6bmnBQFYxDTUGuz7FSztvkXhtLq9Nwvag0zdWhtPUVDrS2Uel3WoiMaHmnmMs1/TnVmV
M4VMes6y0fLvidnu69ptuSVzmH1nXAmvwkiJk6Zql6z3g5SuM8IO7pu/7B4Az84f/xlH3hhTPnTA
tcKyL5GW5XQbxF6IRPD3KLBjoi9QbRaO9+7R9EsSTnQQWb/2kflfuQEijcefmuz50dbAcp/NFH/N
bGYVjIO/Wj7kWzJT4FmC8/JHSeEtapBsAvLD3/WYpYTy1YHowpcBPEXbgOfDCk3Vkriu9ep2E5eW
77Q1B8XkgXzotu8ybDpPd8BNJ9nJ7wpSfkEKOadtTo7VRIO8qfm8iwDr56nIPtkRyD5c/EyXQKEf
TyGtl5VKs6bN7KjgQvuClWfH+1/ON+vXU4Ouijtt/qacZBUv2O7d72MA7FGMJupsniZWvXuSZbI/
Pykk0MM9QKEn4g72YfruKbblrRwH5EMuq82EWabR8mu866FcgmmDN+jcsh87THxYRZaXKCsXgiWN
Lxky/kicGe68VLsq9Pk1Eq7bmNV8Kie9023JEd8gstPqi66LuSFciH73IOuVtnPkljHjBUks8vxJ
IxE7GVEjgRlFtne4im21JWlsjV0qGdENZdTZN+xTPKDNrPK+cPOkTCnbzLlSnFzD/Fc5xSpBlmH+
tivDflLIbPSCgajjY0tmnobomrsXukOFp06lOR6TD41orr0hpb9DXPYrXZ2DYM0MMGoFfvpV+1T6
IxXlqCBzixHGmrDdllSn5LVn1+rvkoH8LPsutBWGRLwmxqi9YHnxKhsAHz0w6OcfOadA09z8DTIx
S+sueHHLEYA3PyKdhZRaMzNwYZwP1nlvT3I0wrtFzeLFBQpiy2IbYJJF12u9Sx9MQg/2tgcAX5qc
Wyb0ud09TAel1j/Q1igTA59b5UC8skx5Kr6IVWz+JyvsoPTweB8pREBBUnoS75p6ZSNULuhZ1w7f
Di+FSGWqIQbTfSNCnpLU+Oh3REWz+S57JvBAUd/aNwrc1+HGEXR7Se/LP0cikNR1vLFwZI7ApnMX
TK2dA7PK3XgSFGdch0xR+H4lsWxpNW3qM4qKIjYzPbtm7mzFxPVKWFJY9x3gu1QsEw1u4LtjT3S/
e9uK53BCE68xv/K/9JnrCDJYjcFlsZG1tj+l6e8KO+bvymnWddnwHUG5TkR1DueP6QlM2+njWPr5
xUd8PODxxOl9mI3edA4MEYQA2JLVhlikDO+AtqLk8d4QN4EU24oVMf+uRsKUw2UykjVRvV2lw5Pu
ZR/QGQGEYjMmrwtFCZqTWRo4JfJHZhUb5JwLCpyOWCFyNjZtK7kJsS63TkPLk9fHSbtkVJ868tU6
OWsvfW0dC6lIRjiFuholL0jveG9KR9NN78fLNduvk0j4Wx4lBt9JuNmjMVi/ZZ6Mpk0JO9zhX/RI
ttemr0pxDezzU4+YL2MKVsXApUoWzJXCWPPpC1VLhkCVAbtdkqDRupT9HiN84b7nrLLc8B+Kl4ju
xLghZTWkb1X7yXBvjrFLRYzByNAkQkQvneNawoqB+3GieW2XFQZPc1JD2hNsRk9GEeDzHQJOA0Iu
5TmnHVrglQ7fdmSGOC0dah0aeQEAjAdffKH8QreNbK2G95qyIm+mZ4BlM8tt9PdwI9aprxCNZrja
1DhXXb2j3N7+bVV6H+X3vvX8QXlriww8TsajOKGGn9A2hrxxt8jhNM8F3lF5PldGAIkjK1JTC/Tb
ARitDHJdmfvZ6FwAPQPTR+vTF0HP8BMDGDlgkdxbnqYYQU2DS1mUOPEga9JIl+FnhrWeJA1kfA8o
eET6Uyl/kjczq7ZRNT3Cghyg5cLT6q03WdMZZM4kB55k/SvKclHNyKKKznGiMI6gf4/5SvF1jrJI
VIull7hUfWHRKYyKc4d4/QBZq3UwZNfn3+Eb0jM7sn4zOxU7R3nctd5peHog74hD5PTZh8rDpGWj
/Fm69AqfvqAftlGN4A6TOR8X0+ycqatgtpluk66JaBZDYDAtVnMlsmEvReNmCE+Dhx/BgcPaxoCb
9SzPuXtCKEVWBONe6Bc2ATMH5ODYrNrh6RTSIlXlCwelPVal8cgs+5Y9UjHZAvQLXKQBxcwrzViA
XC3QvWIwiXFMvybUYn3XNqZryFilqvb9K2OGqFKrtYKPJMF/9bZUlRTTPE1Mrll7UGC3Lz+0mqgp
R0N3uOGsr7dUEGIdEPHix21ZVSVz6xegLqwUI7yiESeR0GG8tqoRJ1vIQUrJTdjY4nlGil8WGeHm
viCioR6fzk++FPV55D3P3A9trSHn9n9PFUGxqC9aK7reepvE1DPOR8E7BUTxJjX1/NHNXviR9wTx
yNhOHJdLuv+FW8TPPQ3k2gLu+YX9K81UmGtBQLL8docgK+pCLKZgOBmGjKYFc3fbTRLaK/QavNHL
Ho9oeMp5D2XOdk8B3LwIhrSjHY/z8RbEIWZd40V/S63/JVBNlDpefpbHJdGNWYc4Fu1Me1iQt/JE
6JlfHPu9ZX2r15zwLm42vKcaA/iHU4cdmWMkQrZAbdUSuUijJaW5WiBYpfZb+Wt4LYrFuiHlPvzn
p5/jNIDpcDJ+FucR+qJChhjFF6YK+U251qwDfWF2DslTbXc+7Xp6tacbBktPXNx0l6wGjpI1zUfV
/e07hucgF5ov3mc9iDV1fpMeO9RHjpNdp7XSa8vIsRBfmuWWic/pFQm1lA714fms7wgETFgjdN6i
MkflBfoiv3Wot3NxVXhtLbI327D9yMuthq9bu2OnA6JUXZuJmLirvg0uojlcigRwxvLNQbTYeHW/
xuazR+p7QLs4zve0irvg4KbjNd7izuzgyPqw3xLGtf5BaOcO1XIPE31FxRyNE9DFPPYb4ey0sQY+
5a/Gv2ZoSXuipSuErPWSYxw7HmJZKsUgLknldQVQ/NJdeqQaQs4sAn9Ib1kd5fQypdhux6daS6Th
XLcOuV8KSvJcrVMHbycig5yauFF0NB/D5A4xGSrmb++6mMsfpRMmFyf61ZyCpIZOYmHlz0bsk4jW
x8qMcZrFLbBpAts8MjU+25FOIOBNfiNkKrK4qK4bfSFRVRQ+K35+xXsXKDxT4dB8m6cZsdkxIVpG
SVSYAJQdh+yiVt0yVxvYuem3FsFnhyC8IxIL6I2Q5a0ljHEVb5Gm4GudUQT/FqnPBiqO+BZ9cCfE
20OXpbY/xtkuFw6Cj3aczJN+EpruJ2SfSH1dm43ZzT+cmTC3M0C8h6AiE217BbZ/8OALq8GuEoLv
WL5Pn8yplVhNlYrzzcxHVBZmyMrrvKZsYDqq0Tl8a0KCLG01E7qky4ejHvHimvi6ukzZrETE7+v7
1l9Y9uFKGbGkd+ONryG8riADbE3zbD0Io/shpZxXYdKBXjYWBle2zBy81VaR/bgV/atktrTqbMvC
LoGov72wUL3zGSNn3bwS9c9uu6TiV4sIwCKaL1bihXNlPM0QN+bYx5YLMLfLxa6IZkuhwJ7yc3Qg
RzGeEW9cbFIVm6ld5efzuAJ7J2E0ZM92cei55642rrayMnqztZ2INisFmMzT0+zWCC4hdiU61RU6
w3qaQ7RAFWveA1hi9+qmHd9HzbFXN3JBSCzERnpSZXnmScy8+QAa6U5KBPAYVV7tTAKuDcpmWg+G
K44VfV3iBbAvk0HX+gOXgzjnlAXOENWCrhMIHJ0OLu5uSl7ZRR2xmyr61jeqBsm7llFb7SLAEwZX
hETKazMMFC+479bu8/159CpZjUZrpaFX0gOPgejMnOG3b9/R5vEkxlEVXEQbkdzQxGvECQKbJcYw
KgjVIeEEMRbqyHBdB0WInqzkXbISO/QTu6W1bj8PV1pKBFTkEXPWmzRrjFlYUb5iIq1Qcsl0KLbh
2bh+cyEPtQCt+/TWO211BeaRaitIgx2GViBe/WqHYteg6lwD1tokaRVQPkSOyI0/Fma1QdNM/Ti4
/LvcfcwINgPHdPm6H/YVAuw2LbzdXT8tjoKv4CL1xU6c4omFK2T4+iUoupQFU9E8bzJbXBLOa1bX
P8kfhJbRV2xhWN/QMeQ2A+gPS7XyvMIxG1Gmjt8eE05YQOqHF96BUQy15IaHWxX+ez3bQtO6euQ9
aLXcz7v+7xqRZDH+6qNgkTtINcKnVnSx2y4vBZwUTSlTLtR3An9YcggDVMHd3oY8P9Svp11KKgSY
jAF0+SXLVs9DlMM4bYEKDcraFHb0VsZ/gJEOH3o3boTk8FDcDpwAXM0t/brSKqtELbl7GcvQN1ew
lL6tMSm3wrnYf0WreAzVTkN5M55/NPBBMPVauehDQJOepcPRi7tziem6PXI1SgA7y0b+QTarlmO1
aUX4IVWCbo/slqzOA4ZJPTbXobLDTAPRAIx2Vuu//e1+LpawYwvp6gnlPBqi47xxYmBysfpOrqWD
9a6EuxWRv8e2QlMkZ5PESJ53GQkuCbnc8AJ+lMrn0WZsrI7/wklV4ZCXLIy2q0KF/DBp3AAVbsTI
O/FKQU7xLMdxgmuEH/RLMJJJMcP7x4DtzC+r1gkTBRpHBZElpa1kITcsNLmRagXx7lWf75HopNmO
7QSOmBHs5hy4v2S4zhTBcr8msWYMXo35hP+L45uBJX8bCWoNcvr21f5r2WaBm7KjE0vN7yPCsnGb
srrHt4MvKplK4w0GvWLKcVW/YtV6yL5IGoNt5vhq7kVTGXEJl/UMxp1FdFcQNYFazEY5t+thRedm
F5rEyoTRLUYjOIkSfuLb4UGWQSLftNhWkbQMlNhKDgs9/xszvyL8XFE5su7+rEzFoNODD6vtvfU8
BrvbmlqbsfaqE7zVbVc+6BfABhqG/9hy1/N0KqRTFqDaeWPFUX76lYkMKS2UGl+cH+G+SwoffMh8
ukdgzeh2QplHoAtBE3Cd/bkoCjLwLSFq6TLti8UpgIp4da3KO15YWpdh42xHhW/GDyJTVttidKwl
IqAm3CU3718p7/2SgaPT5XjITpZz8/gpfArFGJ5IjclqNSZIrOz6/lRPK/Cefllam4QJtNOBhDhH
kv1p5HJk8nMvOvl1iFv8mAnSs/Mz5JgX5qN9w0Ts1q5/ZIWgTQ+ubIhiigRn2t0bpA60XKZjYauS
pGLB3DPPWa6l4oIXEn8mFt6DHemvK4Zz7cTUBRxRs7QtLcsJL1RDO3QT2EoJOLY/AZ5SgAXWSESO
EybzA5VcJZzN5BktLlqQcugjHy7w1avRmBkiBXpCxzYsYNRN7qUXkoi0B5DRulFZ+ynoFk694SkU
0WCHiW/TdaAB9fMKPZUJPkxhdpLWngoTmDpjjeL3BnU4Xb11qlHjxXl2VTy6BAiobEqc/Kqpydsk
Q59TjYAZI5Mpc7uYt4jCjddmcPKRY8dVjeOCyhxeBtiR1KgL7K8NKfgXuVEQPj2RelQk385XLZIZ
SJgAPK0CyvECiaQg4LcKDtkolWl1dk7Yq0ooQamFuzddXVU68C77PE0rGSHEjbEhj7yXepAyNkuz
U83EE28rbvC53pgmf2k8Rsyf+0/W+zDQkzbLQJ7i04fXJ14M8Djhyqp6PM4A4VwXRbpehrjorwHM
Zgy0yIsSS66CiIcHqMOXwNu22MxClQhl60vK4M7CynekumnVcWMY7NMMUDLVUhbfUPCsHn3WkEv8
54Pnf5i3hbrKd7Yv3tHwY7PERkgOQsZwugl2YddZr8187To8jmCiQcrJ1OQzR2zBpHc2D+Wi3kn3
x7PdnX0NaVe8DgCDAtkjMeTeHCPBTNc9lho6ShfvQK8fxSDRQ4f7OqL0MqYIhnL4ev0xyBtapprN
wv5kYJuCEXI/STu9u9cio0gKl1BbHuFSqW7tqWcmnANeKC4f9H3Ws3l5w/nlvcr49jZzuoZ0M23n
nVD4lQCqJ3Nk9pw94HvacdfhxHe3e74NFFo5Qq3PlIb7G06LM5rHxJLGehWeiG3AII6MpjLlvpom
GjSorCIRe1b2oMcjnmbh9fdymZI/soRNo+Xk6ES7r62EVbQfH0HKFRuUSI516+3YMGA0bf0e+l+U
oaYU5U0I/DIquJQlw2RvsWxrnFKZ/GeLWDAVw3goaoKM/9n3r+DqsJACiJDi4X7Go3FAqRCSHZZw
MjmiSKoe38Dem5aFqMxXc8/rsX2Z3by/JeCMHMbSjNv5rEs/H33m3qsEG5y3XluDJr74DrC9ciEX
dSNUXFNm1zONCiJE7uHDivA4mjKxD9I07DOIzeKc3hZbZdr0+mB9a7nxl7ZYkMFwcPQmHlLWlCwX
1V+ndUsBPJZD4QyG+UgCPZ80htkB4RG+YEgsZ3KyS3eMDCHqqFqwkZSji+tM+k4Ju3HO33TJkXNo
UHi16MlwiNJlr5IOBEnaM+PZlyALg/OmGd7RcQuk0sGmkXAokOTmEtngQH/nYn17ex5L3iZatxvo
RczIy3pW0HGpHUroU2+jQ9P3THNkrgYIQeWjNXpyljuLjUzV+vENk6o6+20Gvl8ufsfe/4topU/M
E1pUN2LjNhgqt3zdTyxmc2vLbQjT40wdEqa6aP7KCFOYb7D6FQUO9KesGVX5fbWnTbRhhzjA+rtu
vr5wv7Wiko5RuRps8+OJeOmDyWSLRJfTJCcMbZhzKHpb9VK+uyq0moATu6otqLD9kisqgG1nc0zt
hMhTTvX87CAjQyCgKBbTAY6K1CBsRt4wqZZImMFe8oHKtyEpSOI5DSA1GvWokk1wxVhhhMnZHKhz
pj8IaGZV3XwH1DrIeOAxXWOGQG6pNzG1YOlNGgc+4WB4/CLO1vfsQPXriilm3RCoBgFozZHf5K/c
bgosD00XH/teJAbxo99U/HGaf4vkKo2mMf/oKtiI7Gwkxh3h/lZKa26PHjdG2ozI434HueTnEBVO
ONn2jnapftomTaWD5WJJBBe67bSK3ZDXz/dt+kdnQLygBB/tpOQlsStpv9qN+NvTzl1FTMVYmByU
zT/OzT4kTj4S0h7tCpBjN2k3bczZAhrhWBXEn4kCpEvEM1qCwPXTQvsYB36+T1YnfT9d3fyjMGl4
0Xex9b34w6xqevzlP6a3etwUlHIX5UbFhIiJ0n/stj3bv/djiaTyWHJnsiAQJtePY9mdhT29ujOx
qjYIqmCqLGZnS7NPq+MZ3ilRFJGQXM1Gym0ach7EQNgh41dg4wl6hqVti3gmWL+/YcTb0zkfXWcl
LaLKyr5IBLYWKJgsF0K3AKCzYg+oeSNij1GXTWOLzfi7f5BUTrlwOTj+fxxIKWqO+v0iUmt2ZQvE
KBPWixUNNdAS+Bg3EiQEF9bbhIV6YsAoRqts+bEFrlXrccPnWi4knS381myqFHklULzG6Y6pQJ7W
VoWs5+2uzYpDT4dqHbX+zkiJyFXZo58N/7Z/IomDII+FZSUOaB96A1HJIlQ8rZwAcHOAtGmzF3q7
Usr4TSCortS1n3t/w0sM8zur0+pyf/X+Phwcxx7dlNfzs7vxfyXxCRtiV4pjhR6ifwfo40pAGEQh
12lg2Z1x4c0lU2cVp3PYEwO70BM5/c00+aQ4ZcLgZO45BIoXERAwbnYozedliQ1uEApZMreL/s9x
GOTGZ9zjUCvDYs7Z/9LIiBIId3EfMM3QsgoSOSsmN/EF85Z0hfq0svp1tMuQhA1t9DEDaHB1sF4i
9sLoobixvakDJTx6GHHRwAEMFYbgC541pPCnYR2TMJ1rvT0gF0fF0pssVlGUGB1DblG6GWxyJvhK
VCX1jJmRZmtvVk9oB0pEQ5hwGpogYp+LE1SwxU4NvLVDrjIsqi4cCetbVOhvChcgCL6K4d5CIKD4
Gc0vZrpnRxD2QR6kHorYtpBg8G3A6ZH/ihg8HhyAu+V1VinRLp4IW7Iv4/ggVLq53MGeVvrN/dFA
xsZxxp5uD5Hc8ezQUNcf6boV3bXmRYpxxNdd66rWV/JZTVm8vXGCZMJn1Ges3tUjdWbVRaTHbMHy
NX7OuP+q1nivPk6y6+1KULR3B6HHwAIWJzPOLLVvagKG1qhyODYYpQAt2sfm6Px8TU1JTM5qEjM6
BIxzQ5qYUfq3WQIOci5qPV5mUtK9VzQa07sqcU/ViniQfrygXTYV6PcI/UCnX2BkNIbcV87DPb5Q
IBDW+7TS1F57tdq9p1F3g0at+MjFLBF3iyc+E01H1X8mQvjro0f+pVn3hZz95zWRmO1ZC92NMwK0
DsDz5cc9Fml3bM00LFQbzVQD2WiAdAI2lZUkC5G2Pwgl6WgK8pX0fGFvPxOpVt5O1SXZd1cJHYAK
SihI5PlVTUxT5qszVbCaL3vpw34VdXx9Xu8xMfwWWfjjkgyJCIHaTbbLe00CUpnrGe7621TmudbN
kuhBjG+ZGPihtX8KWIdGe8O/T7u/BjU7BX/r5lbCXDciGiiYNle2YwuJCjWHNo9Cfmq+8QAZ42Lg
9NqsIRQX5ft67x17vp1J7PLjFVKRt3OYG2OxR9rpsZ2AWmrzTN03XLjnZdW/nxHpFdpx8k/OtRf+
cDCDwNBiBxjqzPf7es+kSltTZbhxVF4+0BE7+CZQ4Fu94Yh5AyZqkciT2K7BO9O0i47GJnr+fXPa
3FHVvYrIRp5a+Q6hfBGE38yNYV3y+af2MCr30ZTqh9gkRBgqKhIqa4avAqVYZEa0hVGGDZJ5m9c4
VYCjYzXz5EvWaHDN/kDzKIQluEwP0COyF5/RtRajrhaGJWDVSQdRznfFjsRLyy6SUIg7dPJ1cjUH
Zl5MjLUiTxyng/mmCFuYdfVOav6tWAz2YIO1eysLrwt4OmyFJT/yanXJ+ZKb/8OCZh4OwnpkQo9k
1SuqpMBjkQRbh/M1RyMAtksAng7rabWAk4K31PtoVuThCtD9aNRBdhMj8t1TYDsixEObkYDsLl6j
RVbqlsrG4lJYfVh/dQRyPIK07XngyM1hrO6XwVlNX4eF19OgBWHAQM7VoUbEblNHC8IfJllInS7X
f3o4G6PTSm+evxv/sWULduYHythyz/sEN6bicuAFXgjzrISP5lmSG/A4TT36Pb2Qpu+/+RB/hKlZ
HGzWfOzNrrGMvd4ZYHMv9zL4dDN8APaWLyXMeZ4PLVVHAJCXSC7UcGVj2GPUgoA09oXjgtsNRj1L
TARB1uYoVPtZWKP66bokS6z8Zwpun8gUDs8wVyEylFSGINI8uOmcdN26GHbxjagLwnfb8AiHSj2A
eYTAip0Ij6bqcGrtYXkzZq2CYQEOKGimfJFC8s+vgCyCPApUg+rB8GuQlVz6mt903NY/q+Ly6uwb
mIUdG7gMGCvaI4IjDBqU9LgHUZ9orepl/jS4wf9YQjSGyBmLFV1B5t8GGbZhgkKN52ecrpN4atez
Qzn5FCs+OSyZPSJKjTrw2N7tv6AwTqlBpo2N0meqBU/M83xwCLmGP+Z0sg+IS6astvNHBovLgRnI
Z3Rp516+tXsv6dL8ElC7V9PcGcN+c63sXZkZHJNpNS9mZAXBWq9zjeAFouPa41wOhAH1KplxhRiM
an0QkspRNKZdnEP175z+NWREhEkXLcOTagTiShrVhZsFKYJvWuviE6Ndq/niLHKBXxSrRlcg2CWP
PB9dGEUDPsmmOHMntCejafkz8mMXPokVdzjf/uqrkmraUKKjnRdprcDCEER/Gp/TV7WzZ4bSnAGp
HHWn0tnu69xNVQ5qHoB4GPlryQgWg37/BDeW6Ovc5pnA9diwbZSyXbq6ngp+/ANnSLcZYv3+9aaB
Th2cVZ9zSwLkws0PFOqldJlXHmB+sv/CfdENQh2DiPzlj+TD/QJTzySNyG9KqhJjt7klmyTQDyd5
bcie9Vc44XaVtNJxOAZ9nLVCp6ZM7XPw30SS8vpnmYAH/QrgsqwFWLYSwoHydmHtM5ePY13alk7n
BSIwpXFk1WAEDsR7auJAJr2Q+8FPlUJlpNxwzsYI+0Tu0lbG5IFaebrM4xSwt07ftcCopb4p9kwt
Oi7J5f1/ORNAxdsBV4qk6LCxk3QJjXjAVd4mfDvlTlq786MFBm9dGig+iFq+n89JU82BQBcZ9IiI
f9yoeLopdBVngZgGucfQ2EJnkGmoqLQGW8Woo+JKVe62JPM3H9kmQ8xSCYiqHKybWG6etCq7vEdL
3kVAYUqB17JYe2p+Q8BCb+zQIfjnCMObeWQ2H3qQnaBSaCoKurzCESULR/h95kR+fMSkuflFo/Ix
BWL8dA8/vXhx3cEhb0hI72rvvZVgneTx31KJ4jN5rzcTKRaYTbsldPrSxQDujqv1QJnTMPLEiu7N
2ZZzM5RiSiggBOGk9YsvtXDaC8ie8NYrdOC8C6tuo76xltqfSG8z/oiACo0pNWGHWCYPIbKTpTxK
JATHF3YJtCDbxahga9CTHdpF8dYjZKXoSYkrLzD0d5ivsob7qerialjsj7b5moeJ3nxk8/H/M1z+
ImYOKaBP6Qqh7ZY4F7Hr7vMH8C4orzp2/9hrH4D5F9ahxUwnrN38OBSmeNlWLRvHFwZYNLRLdRD2
SmwcV/YFoicFrqthCqk6badVnaB7M4t1NZgsVNacFbMHw0Y5Fg2ev9u0nRq+lwGH86wsiX/jvMOi
ncBq9lmOnUAtGWqM3A33vCVKRb8rbDQnRxuklerzxFmG+/M4r+BWY75zNyeqcFIagBZoFMNVB4Xr
tbvAcSmOhICRI3wP7zzx68UuYVZYbYGfMQdQuQzWaM313ohFA1q0Rnlm6i4plUbsbXAkDP0y+N+U
rBIq4kzrJxkDNBpbPTwiQMMjvg1Tw8+c1QzuJokINw5JCRYXcaeC1DZkL/xxeI7g5p8lEXoPEBDU
b44lQ/InJ0x1zoOeWKe+i5Pwkm0wKF7ye14YCXsq1elPd8DRJjttm3bt67J5j0CpT297k6bio3GP
IBR7+YkUWHjnNtdbrRaaE7psf2ajMbN4dzVqpxDtnMKpEtSmDghGk3LhuVJ3v3yWqAD6psNhXBTw
yBqV/1Px7mAC7qjh5P0AspYnjiTwAiAHaOSFCDXILiQNMjLArR39EglGYy/KozCoFLzpziD5JEPl
DbMAZc7GriSc10X/2WWGlnftA7zB3VZ/3pn+71BK4cowd0AvDB7dluq8goq4FnuC+MgvTJDw44FO
p0CLg3Q7xwAUZRKZ7h4Cs9c7JlDAaDSHHkOcoY2WULI+La4dXzPbolV8LdYHgmke2D4Q4MPYsRke
Fm3gm1zsSbJHhXTISR8ucgIjdPHb2WU3ZLh1GPBjA/21+oU5uuQquUA8b+IMDKNszAGUstd7KMKv
1kxU9RQXHbnhWj2xvpsbumSjcYLxq/1Rff53MJJDhTcMrQOcd785tqdmrnUzGRlu3NboMep9m8Kq
UMid6OzXFPVOvfWC0coa2+bdMwdpUo+u+iDg1ia6iDvYv0FPN29E/6w45QE5Lr1aqyeWXfp5I0J+
MvQPjEeUBGl9it1Gd9a2Dcl9+XlWjLhs/jyhY7O6xehaIeJLJWZlhTHJP3D/cJPE7gXuq+6nf9zJ
jI0cqrKZxRL7QKFppxeLi21Cb0xkVP3B7PFp/zf+haAn+ulGa3Z7ASDG+6z90Kg7aibbpcKsv9/d
3sscbIjflrxohWx33WOwL69FaHXRQk/w9x0Sg8tpkFZ9dZfAPhaMbgraF3XyH6Wfv4XGhZtdXXWf
rowtM7OKx727QwMNzqX/fbNRzueNcOk7lp2YVfyib56T8qq00mX0T0lZVuSlCikb5EWubMVVAIhC
wIbNNXqwX7PUmwV4A0Db1GL487ZFUAa33UqrV48+qSYtTyVY1DgW2wUcbePvR/NORtocCG07uqdG
rB+6HEYI7OnfxlaUCTprr8H6dm9fuVcYCrgzwmx9Qa9q5+Ay/QtRldVBrNTef3wvig3sUrffQYGm
jy6S63vcUW9ShfShOVopzzfsfH4jYxr4m+HMQE98m+QPvRQEJQ4eCEl8N2XwGDZMYyqZUhcwyYtA
ichz53uiPkLO9kxexxsTd7DjyIvKQMVxbcW4z8lrGj3iJmxk1O3y46b3nAsAsg38cR0ils5Yg8ko
AfN4z9SfIX6Sr2FCIATeDGalc1z0dt1o5HK3WQ6BIpnlxPGAmt96wL7TH2eR7jnYsRhcg5NVXYOQ
HCP4pwggKpcigIqcHfKf/9E7JvDcuQOqnnfKft97ABUmFTomzeVMAhBEnAKXrZJTBaA86BLTVgf6
PNSqSmrvgj8/a6uqHLZnpqfPhgelLO6dHzjbBytGv0C2PbaK15T+aD4/FWKlgWNhjJ9pNh5gIaGa
Mo7RcqB/pyGdrvfCP+zKaCucws4ZtfWDET3I7RI0KoxCSOhBXFNQQK8v7l7zrb5mwTNwzW2qSVdw
AOGVcezFU86gGJ5f4BVyF+wIHo1zqUsDZm2InSms/Pzevi4Z8kztrVGzgxKMgO5vsNA8rwe5DHJv
LsbDPZ7oleeU+BFghEELL2AhbgPOO7e81/XXUYHYmhyxOb4XrvgDPij/YjABFSttP4YxaP90UstX
Zs73NSBLgAKP4Y9bIYI/T/tdQGFAsvEDGFU1OuYgkNVjGd08NA+rjoz+XgIAI0ce72vEXTYNwXwM
4NX2Pfrld618Xs4hYvti/fUmPPqCK7Z3aBqVisip60h9mxunXdyntUewgSAfCk9IXKM7z2GSoGxM
Kj7xjW1oCyVl7WKPuSxE//EDjQKJNsZUnkrW1qujq9mKV2C4GJjLcIWRU3NR+cpP6zaYSoOfIjqM
kAHGHUpuGnwJvHQYnNJ7tNMISwvjHc5TtOUy4yDPw3iXvGbcdspe1MY1ecTPtx8TyU7SOOfqF+mL
PeK3RQkdaVVJjoEQWFYKIB0hAOjRvYtDAMmADtwCQFhM1Hb5C2MXB+JXUPwWL0uqymoKnjQ6onfb
FrHw+Uqt7OsFdCWXAWFlgtqNf3OxVfXlL2RUuB2zBRb5ibrH85a9cu66uAmycRKns2zGY99/1x52
Okw5S2bXQk6jcsVerfVu+uq+G1Fc+Ws1o2aieY+b4JzH/TXMdyvl3w02qQAis+1GVzczwZQQLsTG
bZZ63r5tjQN0sLFphAjxoB4sXTM4JGYPZug6Fjf8aTuIA02D9ZAd3RFpakUv7iNwkisPsbJJeiYn
Y1izRwL4qxYrf4zzxyQb5ep8GE1uB4O5hBoZIFAxhg0bn9OGRNS7eq/7JHObWUwn37Vc5369JLvW
SCgW79z0np8BNvIUncvJgrwGCr9TvoWf9uYNWRfMNuJyJ4YH8jbkXgJxytl6hb9WMnAAGME112WF
VrCex+TS+crFpkwJJ6/tbG3tZIaaIs0FovUftyIAumv9RXikS55fzcmy05ZEW2jT0KAcLKbjjSRC
57ZnkjjEujQAPVUmRc4ytVnRNKQfV9c8yaR/iZCuMwb8ElqUSO+mgt7pij1DpHVcraF85Pz4CqIo
xOjgiAFW13QXa1+LpVvKiFfDUIPP1MvVYekORGEHE3J9wi71B+mI7EBnIzGs4OPIRhkn+XyQb1hV
Zb67hPJD0V5TQcZBPiMNyWYNbX4MN+38J/q94XhVT9yWJzjnZqemHnxwgZqGTDLUv7C7DEJPfUyk
67aFYA0ywZdzNRYa8vSpLx1lDAkWrUG2S0xJgxlqlE+EMjiaHHUDVHGolM95c8ErHsSBAgJ+T41o
+fRJVLkCU+83ZGpgWT9GkTLzli3kw4PpuXgcdqujvfbsg8EE1j1GMA+riMRZWIraVM3jXbb4lITb
D5RVHFXElbNaAneY1gd84jImNrnpTn1H13jvOClPAQ19f3b39qn3rf2Z+JUWS1nBAzWakRyV8/kz
qpY/3toVah8waexmOvK9Rb5iDgpZPHuwwbpmg0POJU03ujwdUytwFwdL8OJNdi45UUSBk6rP/2v4
TiJmwy3DwEHoN9Kwqe1oQgjreDam7mxCQ8584/eqi/djp7GWTgSGVN1Ttf4MZpSbYtp1UyMaDfyv
WdJZtN4e3koO6GNM08o9uDWgXzhTfROxqV+pCogFLFA+EiQZPxYZYZsMVdk+ANz9gnBifYarMeHv
+4EIwgy9jM8U4G3PyP0FOmIoQXCIjqi9500Rzjfh2rPgfL4cuLz1iNfsCDeqRknrZMi5Fe5sySou
Y2ex4kWBsTM/OtX6pdGJRYiZi3/iL39B2euT4Lqh9HC5DDHXbauVqg4+jPfuPyNLS5FkspGeLYqx
3GrgPyRTawQ8qFlqK4hLulNSGnuqViAthGy0XCcEn/+HoWekGoQ43DfvBH1PK4P0A74cUf61HIpS
kSdoNzB81J/hM9K/pQj79KBm5oYqZDMMobmCOMfgbuIQR4ouCEwY7gMlVLq1VMlqfQ/3jR5tpTm8
WNKai+II33pxIe9gzxRk0xEdaLh9SZklIr00MdsOahQWw2v9LqLFQSnn/yR7UiqUBnMdH6QETGkU
dkzF/4mr7fCDUpmtrjNS6AV+LR0gZoaBlX/KDq12afRuC3c/3jKpi29URugg1hiBVyVZo+KeZBTR
C78Vy06eD+Z98cfjm04n+j1bHUQAAt0cyDrqzyMmPy1PtZKeCRwVK6mEOo6E51TbrC8J+jnnzGvQ
Ky6p5kcvKLyeG5UuRU5iOtXNCOanv4ZbWyumUNRLsh8CwIv3X0x0O3ymMfGBBE8ZgD+fmkKgoLhs
PEpzyBRDJ9h0kOzO1I2Q92c3m6E1L9tug/kfdNsf6NzUq7Pnz2WOfxuBklzzHxtroX7cFlN89z8u
YpgZsMMSfrhMBw+TbRDCYagixYKqYpU7jYd3rW6hGC0pDNNuOPMfbMtX9EhasJ6deqVSkBGlmM0u
hMQUVzzl43VprToHYLGKlrV43it3ZM17ACMAMgCtI6lq3gX5+ztcwYIfDe4Fd5+Bq37Vgd4JCber
initWXUYk9yRVuG58gwe865upDooqypgd4SSyo/qRkPV2f/JwMfxjbFRhRqAyfyYyhSlRTI8jGUz
tJrnBfUUXSvFTKjqL4n/T3g2Q6jWkmJ2dBbyrRFQlGgjUxV9hgXj9Yu2QyVzZ2xgEBFfPhpwmdCe
7na+e+1uxi1B0aR1X2AIQz14c0hUdpOYUM84JZG4SzDIDuVpc0aGPSK566/L6NPbUefqebi62ZgX
wXi5sgthH9WULa/TUcp17TDF4GaX16ISKEt8oWtdMDMEytawVPEc9aU22GJ03bg/9ZOXvGqQH8qC
rKoKTSQUCndhuHo3I3F4J0j47UKN+3+xep7zwl7GtHKfBU4L+6yfBddWRjFu7QLJbE1Jb7yoUexd
zp66NlZpf1IECCVhUWfxqFzwcxbG/PYZRxrzQE7YF4bEyPW453NTmlIkEu5Axakqu0XIWEE6TWUx
jULnpxhPJrvP3NQuji1a41/S4ObRV4Win6Ctv+0QnmBAdYA80jKilrKwc0/A/SdZL2AYz9tAO9Ir
K13J4NZbs3ogNk0K4jlI30a3eceMOSo6c280bJjJvOL29o7L6iHbjVm4+wUjfcaLlG0l0WbYDsqH
zxtJNW7azWuh7uI2x8TfvAzowniEhCEco6auqpJPdhm/bhX81uuSyE6BGl5wgDrxXPDagkD6kMGE
aw03oXr31syx2d224GMelotJ3jPWkQaIXq8SbxM8yISpr5Z53+OnVk3MGFNhvi0iX2V07YHUr95e
ZTwsPZN7EzF1noy65pITSMXIf8eGRg92h4634+qvHzbOK7IaO71HVM1InepzIBsp0UKjPFGOgARG
8O6ErLWoVfXMglBj7a0i/r5zm/LYsf/Njcv+vv1RMgtT3ZSVVX6fqyloxvmFmTjebtP+WZG45WkB
ezmqWrUHjblXS5NR+sch8pWGiY1g+8czj4utpr8v0aX6cx7SzPmVyuf7HoTCs9aiLdTxYy1PiCMT
lLr7uPCHlFV6/lmQHzNeuNVoKrnYTGutUO6A6OR/aQFs/ZS7MCD8VzG3u6Zn4cPf6FeHlr75q7zE
jYhjp5wRUet0eR9JCj+RGixS1hMVpG2hsVP/FM8KkYfJWfbUl8jnQeVwkg0WsBzEdJTMkw3EmMHW
i91hV1TAESlrHJdZ0cmsLeg/M38K1cXvEa6G76feJpbiz6t5cYo5igRrglnYpyNM2zbLpCG9Ph8Z
1aA7for02g73iMQX2eJ9PVTcvR7pjcrs0k7TFb/cIo4yP3wfGcwUXRw879JjFYx/SRYlLRdJnAh5
gvNSaiIEXz13KJYwdy2oxBrZNh+14dKd2vfbdyZHyXs7QdWhPZcGxppczFIo19EhY2aA2jYQndyG
3OdRKF+E4UfQXKiHPPYGsyULJZ+FZg6qbWsA6OOeIxKcNfoTa9q6gRx6jOBNjTzXRB3/z7EWsXDs
DiGmSsEyX3Hbs5IJMCU3RtoBuuEr2XLRwKQgps1gux4JyvQ65fwlo5M76dEh123joWyQBh8XeN6X
TS35aj8zaBTFaRDcNuC/UknslRo5Cv9PQ9cDHVw+jzxGs8ghO/v9lU5nHefJIHOqPFP6CEYNyDFc
nrgK8noehvqZr36sjtI22wCE8MVbr670eVN5Tun2fPulM4DblI/FiNNc2rPUZjBIgtkkmZjTPjch
MPMl7di/5kdPoyEfFL7Zhn8rL08Q29b9dkW2YmvE87wwRY8ySCmw1U5EKj4Gd4rNosrevhSDPrRk
BC9bYWG4TzeqO4Q5IGU+tRNPmfKUcb7ntKZdvnHZWIt4uhj45DToGn44sNmeMJeYeHCvIQSIdnL6
YdnQYdn/dITOFmbQDxGSw/gjxtmsNbDeKp+stuLTsEDMSDqbBIL1P+r/mIxOqcZyyOidDvrqte13
e4Bpr4GPFqYiEFvSlM8ufpXIepYP3Tssn1Xr6bgcVl/epWYt19KyOzsq7gqTzrP4dHK/L+wxxrAB
ACEHh+7tdQ0uWhOFErYizmg9bMxF5waCfNg94SE5wg3qhoPuHohfklMeMeaeRDeUNt8rD1pIih4N
8AX7LpDL1uvuO5ajwUonc0GBniLGm0YGantSXDKU24NhBuhc5mqLZRe9s9TXt6syJskQmNc9WOct
jeE61YI37AUzzSaZJWroR9UOLyFQnaHR+PAebaa+/tGpzo3zOVsV9ZIw5JsPBBkpWGUS7ipBwT7j
rEK7GY3SlRUlHfho6ow6V5zk53dK1vLOxNNtGvrkEt/Rv81Oto/gPhti47zLe8kHUEbw276bHPIE
hfyemX+3fUut8kKwSBo/Smf+NoKTgIQ5EYuu07f4bHAu/9YqpVIlJWubz4arVea1MweGOSgOR29J
ppuCJJUo5cTb+qkzpGIVep6coy3lYbkxb4Ed+wl/A4XMg7U/Alv7r+65QSjEpjybsG6fjJ+siJeP
q7mur1fkMMX9sHAyfQawJ8KQJXJScV+Cv2mTlBr/sIdNB3yhhuk5+X5H7DLYjob5OTXceEmcpteE
OOn1RjhKErIrR63aXERo5ymfQK0JRY97m+YlNLWr2EAf/ATMnxf4wGv1D75R+npSqf5QmMZhzYHH
MpoCtt5melD+y+keskrmQKnzEUNsr94TDU2T12LR/G8vtHaU50QooG3FtKC8qepnFNQFLts6P9ns
KUAp3jlc/fhu2RdPuOSlkdrcOMbmq/+TVlku4r5Dkv2zqOpq+Yd39Exr6TVqzTuPI9m2JIPHLVxM
hu54X3SIuk62ZkCFHCVrGhjpRTFCAFE5l2pDs20zL4a0kUbKSUixWhl99FWv8eSyCYcnffFRgfhA
QowatAsLZR4dEF8nkMZy9rnUAa6px1aKdDOXXCOOngbfailj7Tt9DouCOrtvdsQgwWQfBpASZqJO
srpMc2D9MSY9ztFQJByCB0kp1Dzum/DccqxFUyOovbXsAWo0SMXTCCaVdXFyLgUDo550L9XMX4G/
YHr+re8BkMoL/eSfgGg//kn9H6i7VPMfVqqD5bX663HM0B6JlF2plDTiyMYTTC9RntyLuwX/XYIn
E5s95oUpPL4QyiZSZ7ccNP11Dl4pEj20/fcn8NcMRpvtjr/BuRwC9FPpC7vicmXC7kmb1qwbuNCz
W9qMnJRlWBj/vactp4MxflJGLmOwmE/zpeZ3mOyGROo4BjWOy2+XPfnq+wlmJgqGNbj8WoNGrD3+
8DF+HHLX/ceeCihpSOOtc1PjvwQ34qH8Y1kR0W6//LYZCdd8EJtbhx0uOOXrR4mCHAIrI3P55K6z
/D0IvRvde7FUgUslNj8/wmF85AfWQb4RPMLZTcV2Pd8n6m1EvVyrJwzCWUFGJsu1VIoECC/SjwIJ
B+YY52SdY5nymfx4pNdVM13wOdMMIqq/n/9k+bYzf2vZ2Kb1uKxznNN8D0whXA/L/mb1b59696sg
zkbvlXwrb5VifV9Hks9qhh9K1a4EZGD3vp5MXYQ0VONc5hrl06v1ilD0dRaVdW02aSr7FnAizlJK
tIKYrDVhfcRMiuHLlk6/Jx6kzLuH2w9cLI+B+hMsy5hnSWNZBH4Rk45PwX2vT4hvAZ+IntrLO7W+
UCKnkGQHiHCispkCZNljAxz9RPKI7R1dOum62m/FM+clX/wYIU8R5H+P9P6cyJ85RbHxPEZd6gww
lWMQYZsRmwilra+MuwG5ErrU+F6RDe0Dc5ttVB1V88rKdqpwZ4EsVp4W6pg5lzW67NakjaLxdUsF
t2/gBlGSohR/SyLMIkebqNPoYGQl760KXrfZBSccD0UHvLPp7Uj4xHzPlJu5I6HRF5jv7o444+mC
ZPiny+Bonc8sH7fmu6cadZe6RVZqT5dzZlm3wIbpRzH5Jx+R7QSA3deo4smZPgcfNFiLrJePDcQ1
k3PJ2cOeFTgA4IH8fMzycv8rBAEUREaPASzy1sr3EUf5QCgeqP7q7mqS6CtNZg67cHy6dYSnECsk
FNtxzijM753Q/CEc8uzVPWiyhV8qWZEfSMdMFPqmuN2aPtZuPCAT3Llh6sE8QOc3BGngQRqLqOQH
QlIbnVmUQ4os6cuFfDeKj1+/txumABOQDiHZTNFVCwGT5J5FFE0mp5/ryUjun6R6DsO0i0LLK3DF
lvNGEfawjmeaKlthBub4LPOZMUlAaTIGtWrMVNP2TRqVaqCfCmWxjyTOM24lXP2GVMY/DZy6CyEA
0RTCIPujAlrg0Xxo/LCayFnZiWm6/gaCMyir7sfeOylvDxsVbPmDL2Y1/DnhgUQnZTmNWUnuKmPE
AwJg4pLJX6TdqPDec9Q+BsNuj3f84ZAsD9BZ4T2LG6sHWZXmSeShw/c+T2jQT6xUGPRX1zbgtKyX
LNKdJPQe51AGaEg97Sw2DY7fJx8Pn87LZVWKslCBe6Nd+A/ne4bpThC00zphbAxHBdX0ucGSl5ol
UkNFqUSgM0LsOCUpaSi3eFJIMPmqQyHeBMW7aPDvVOdrAOy0dQHqiQKXUSpNegDSkT9PjiO+rKEo
e2hDP/Zuaqb6929qfu2SOVN8APQnaCtVx5dP0MZjufdyc6l38OBqYi56Z5vFf79vKmNnsCpwkDCg
7cs5CbCVhidaXw80lmgQNqsEN9xoUY6RqS4mlFGthWUBB0FjrExpAs34YuSbIr48REwX7FuoAM52
0tYBc+eN93DEfA1nIusqAGG8xeOZqbraYGA1Z9fIpz3Dqex1peUQdeVmyVX/ENwzea4A8YBe4S7G
d0P22KJoenbUWP6LVOT9tQfCQYo3vEpDEX0vHVRyfr5jhkdiFaE9YPH9Wtq/g55m/bVppSoXIIPU
qqx2IKnS+1LeB9YjfHsiBUK+giWduBYxPZtfURp/v27zslIPTll0nkGWRZTARYAcp/xoVEkJwsIp
E8gaGA3MyLMLD21JKYAcIhBPZuQwEorZG7/34GtZ8Yz19MFrCi4+UYFwz0Wa6jzWVfH1VFUE+HG2
Qh7N9Q+6jP9C8wzkQ32Tif1GywkqJtW8SCEr5KD37OhLb4YWp3mvRcIOaFONEA8LXUGcR7wU6kpC
/7FjgC9CqBwFPwRAD4velqSCVI2VUjRLpRt9MmfiUIVVJN4vvLTyqqVJVFqElP+XCUlas4/zVtex
0IlRETrA7mzFlFKVB1TPPl76l4Lzz6ji/mNmySVaytCqAYmbm/zU9R4Ocwb7FZrhSRiqZA/2naYx
oLg9TMG7VmjIJzXZFhVw8hFm00wn3AfF4sgF/cxCdy9FZHwtuqsbrT2jn4GqJFgLV+oJXTHfZC7H
7OLTTSt9hfNj/hcDxgTPMlBUWxgiSQoWVDT6xFET6yj3f1Vm02stm7KyNIH7hNK0aDYYqexAUX4D
6xlhh6TIcFx3+/m/XUoqPfauVLDM1KKIe7gJ46YHMtvP9GcpBxYPIYvb6I6DKzwPYQ5hZ+FzyUaw
10Tynz5olNQ1U+cZF7WyoUEgWlObTFqLBbfAwhrLCBRy34L3/ilAuiOJe5mmzLd1L6Jm6GblhUAH
RgUZA7Bu4sIZrtQgpKlIMQsjiY5rw6UEDylz1Lh0ysBfb3R0Z8ToGJPqrC4xXz1XBpAuSOAf4efT
+FBtGLCBl4pKTipB3+DKyB40Y4uNyUSuwNjijmjfClwQzOlIsXOeR2kazv/B0uiR+Y5LuD94hfyX
yB36ofWQgU60tbuKSFes4+8WdcuKB5dqOo+T/Gjlt/+YWB/3poXpd7l9GLIqftRoUS+I5KmHGIet
MrfMdrjcZh3sCa0oaSwaLy/J7PuWLaS1elP6OvN2cdcBui/0zjm2WUKd38X/1J5AT1nD5PisVQR/
lnuwCYfT0JqsVxpKeSPipW6Z70ifSkWFopiuh+HdgO8yUecrCWLGsz4Qk2W7ijGXIi49W2aqEJRU
p4hTVjtsZd8ZkNFop/pKahIxY8QKl4UmGZMmScFfWRmGE0cUXuqvWjAo4Vepw5Gaw+FH7ZAy1Ig2
+kghPqUhTxh5ZKkYkvnizeeis5wW8naqWQU43aaiiaH2NtaOBoivMsOwX2ZLntzzDPOGQailCyzT
4NbKkntVdY3mWixtdEfP3AYwagf4j6/N1TdszFfyfRLQmW3jpEvIXkHE6EJi9CcT9mzyn9aJNPl+
bxnXCApiGAhWAnBOaxZvi1akyMdv3PrQqspObRXs8+3+XVWr5frlngzRUZAJKoaKmByk70ADU+Ip
m25H2kIIdiKDf9RjRTOdaqkYSFNFKiUqbBlTbBi7HwVTyyLQ9b8ecNo6naD1w0qIRiid/CiBSp64
Xpa/wK+Cjd4+MQ4ZfVQ28noR8xRztP6mBsEWVtgPgskm2PqWMKdWLk1BeybRsgIODGm5LL3ChKHd
chDU+gA7lzB0I6k/JR46L/l2Bv0xO4/ioraDBOvZDvOiRX8LKKvPTfVGtGVoPcODFt61GCvjLPU3
1TSrzKx5zQ9s89UC1OirqZn3UPLGAvn5+bm5n6QcKRt8+auMK4A+5tcHLdYE2xy5GHlPy0/aiaKV
yEhiiVfAsLO4rqmFxn3e1SYYc6ckdbnLYJ4DRXfFQwKqOm2WDs67wuxqLiOZaOE10aajRvRQA86T
Q5W5lhs9n3oDYgl5Kt6YRSg3RwtYkRoaEEScPJdLADLZTlADoywiS9mxrDeCEpMCkEqQh5Me0KPk
9NvsKrcKz578BeZplTraVWF3KARIYzPb6Vfw6G+aLL55khjzm0kXY4NC4F7L22yyk1JFv1m235J7
NrfYN3Tu/ZqZa4Nixw9O8+HluypP6BlVww3sZ1QhmmeCB8lhubOOqtuoroZElEoim/SqkfiBqhFS
chYkNIF0KQHVveZQ6GTz9MUzrEHx8UiGhnl1kzykOYeFpXLBuDr3E3bW8WCJEulXKD2a7mU/f2tq
i221xmuU7P35fh4TErAvhENaOUKOAfZCIZKW2H157l/7zhGI+wcoprMqgyWPjpC9wrHq24oYZcMR
6vU02CFt7TUkJOJ8ug7BpdNuCfaFmLEt8i+L/6OCL/PWDF3tFcLkjlO0Jh9ph6ft6SrRNLAXZtPD
FD06horxE0muk1SGnrGCRCoR6/dVXf38ZgVeBUlqv9gN272o74+8N/1pvx4nDgKMpfWrX/3c6UlE
yQYzXYoIhe8vdzMgyr9cC6304FmC00FSanUHRHWLR94xNiSDtJHWaZCxODSRFsaOZW5r9MWIey3d
kmpx29n5Cf0K2hSOtevOgklYVW1PHw/WVyE9Dy4kcAxU2Iyj9GhxvRbO8MnN6rEl0GhD9aSr/j4L
AzXecrEzirjyKe099awBHTaWZcJpmH9Pd/kG0paiyhVdD9xE4cwcxgSI8uEusLNNjElhqcc0pyYE
M4r76/RLLxK7LnR+8eRBmveaptOWgN2fn8okOHjui28Ag9NWI3du/ZGSotxyfRYsopZrr53pa/BK
BtYaF8dTldpU0z5Pc4AmNMQfipcux42AQCmdbNjhbOv6MJcSj+xj92dqVKvhdi+UQovbFIe/x8tp
VjE5Yceyoh5KrNUw335Op7wLqAwAntjwH7f/rbbVsxo9SrXgTmEG1jtjl/TAj7m6o3doVOdXj3tm
881oUI4P1Jy3qu0/btfWee2j5lm/BA5bM4pqkUZ+7IP7yGudYaOio41g07e+tZyDsmScEeriEoJZ
UpGkzSQo/L6xldxCxanPHJbCBmeSP4TaSv8kpSJwaFDP9ypbKj4RT93vxef51giJ616/QcnbmVNM
4cgF1FiYOxgV+HUAgUSox5zBoJbAdnCVSNHq9qJYg+F2Gs5uK0pkTxbTpT+3zLVtoVD2hHezgS46
qSD105EjB5SwMWm/S1xR/A3GRc7X4s5CtWrd9VdSjDQ6A3nOIIIS4SU6qMNfaNWh6Ab3HShSrbCf
2c+CqSEF7oYkZzYJqC6mUnTjrJqxdJAV1tQh96w8fZYSiGYyWrQbLImtQoTwDOHkz3YLjYMViLTz
mV6tX68r1O3yOCDqIIimWYUMPpRAJTr051WDu5Mw1fvwIaTKtrlo1OBwITIeA57V2D74gKooEb0N
LXic5/9XAWrr6ZbxkkoJXzwYLwOSRXl+PTI7lJYYnrURI4KJHNw4iuK4j4uTcai8RvA/MpnrB0x0
4pGEI4hOxsW2ZKby8eXxU2IqIyL8k5fU07wKDvymuUoNs709CfczCAikk7WwoCTVR6CrVVgIu/eq
0OgLzuLx2SzOcYYPU1cucqhH3ldIoaMgqdyfBbjfFHDJDMeP3LCoi90NtJKwj2lLnp2+sqP5dbts
kMEWll87mY6sV4jxSuTYOLqANk0YsK88ju6h6HHoS63xYnTv0szEAleb7T5zOJD0MTplwnQSK7Bh
BWC+YnWy0qhfpND0xIYmy45oSipklhksDLFSC8oOgXO/6UvOvGY4F7A5sW98lzBoKyvRsiFPNKR0
PPSr9iKaVwhSkWfP4ebVh2xDxgzCCB7CoJeo/6ZbJxaOnbz98PfNLT0s0CH5TSBdhaJ4aDbDpz/q
/fjR6mjgqQTOO9M5eFYUndU8Ds1mdwpyBRtg/tzq1x5MdWJDlEV0UUoO7FuDnXmewJp8sljmlwU+
9ky+3Gc0QJ+Ml17pBoR8MY1qoINH7oyNC0QOFqqkjjgjcI120HO/cng3/UcH6EZeFGOili8K4OSj
vJXWv4ialYC2l6nfhLazcAHJv8ZYqhlJPKpvjK7/cDN2K+gkiqnqGTdHkiaQ06K3z5ET1bafq1AL
IxHtx5EgTw0VLMsHJAYVKTr2C60sS5FnhsgyoE4UnPpm1/jLimSbjXpoCooj3fAf3GaoyMHJwSAJ
mjDa7v+XPtBlAIxg6B3JT7jJtj9XM1qeYzFD04hQIp8WbTJnEuX0zDsIU1s+h3+vboK8C5pLboJi
LbLY6CLSQaAuSIzBTS3vtDLctyaUrXfVOB+5fjdCppxhDpN4Sjsbiq3W7ETHrpFqafLyuPkRCrJk
Z46Nnql2XttZWUbOqwTggvWh22L+ReQ/K/qmzpj8TVkLD/YE6IIBc/MGerzdGMm8ieODSYmdns0g
JE1sTSyufcCpto/PhF6bLD4QaynG9Isn00TnjACeX1/pyPguNF9oQ6L+7xCnflN1iAwWrvbUwEg6
eJL4O+A3oypRbE0VcTvNIa2DZBL+hJotvMeDdjSuo8iJVx+UmgZXAOog8cENYb8q4PwXX5w8tWna
S+W0DLG1E1u+CeM7x4xGpyOhdi9L2csXaATSogvoKRww212jgH3xr0k1ooyB0qFG/h5ikSEgw5am
3iybW5r2qlHmFd996XKan5C3/wKJcdzbPSBcJcJQvQsmmOaRx647cgQcQeZE6oGev5pfKJXDzsq9
18dRB6nIQFr22Yutd9a49xaT8Rq+VoDZou1eZWtXpQCxMKtmPsHjndmBtU0RznUklW0msKw098bx
lZ1y0vI1wWGTS0QS68FQiK+geN0qiXbzAWzGU+l7HPShd8FtXL5qlMuoEV/WqEW7uhD7EDAfPji5
Lx/fp4D8vjCW5Bad8nVp1jxwwdYvsjCFwWWV4lgol2wE4CCxXvxRyDK4xaJyJI/z7iCSVxCnwrCy
BCOZiQb5/k1K6li9Nw2aPhd4Q9aXiJ8Yw80IyYZ2NpXmvc41VCv//jeH+llvkG2ojhQZ9KWFHLbU
PRuWHPhaaxR/wNnuFMNoTzg9ny1XdaRIzYNNr5iv01WM4eTTOqdvNG+TLPgulC5RnKc8jE8EDvj0
RooOuafVyTP2TF5o3pOhCvf2nvYiLntiuvl9Hb7BcSEzxK53T5z1p2BDNbPEZuSIDMaYfPJH2Yp2
eicnjsaZH09PWsy/e+aZI0FI1O10r3ZyIXM4GDewXyrL6jFahTZeySD03T6Ic8q9/0515rnSjVbP
POyFqjXSBv46+AGoaM9aDqzF0MgP/ellj24let5xp0yyDRB2O6rF7nOx40YrXp55i682xd/1tyM2
qpyrX2EOQa8+z2TPGiZqz3EF8+IojTZhwIDwMa3LiDzz7hypux3f5ClJedDPrWMQaAx0B+vgGMm6
DFe57B8wXukHulh3ym0d6xNX828QMeBT+lRwFyl7bbJ0k6GnyZmv0o1Yq2mZoawDciMaY4bcnvs9
c0KaSn1qTV/3RwT/BpexYP7BwGMczYSdLcddbqH5yaJN9DA19IOtEGr8f4LngxN52DZ8ekNkbOFz
MWUx9utCn2S7RDevgy8TTmcSVY+FSjfGCN0v3QZIkNc6HH7uxHbGM1X+KwlkFfW4xnFSvQQpF0Ae
Ehy6XdTVXqd/RRiczXcobVQFGsHX6Lr4uIbQy8D7wZrqQemB2aS5TznXAFS0/OsiFo2tn7GwNTdx
Mq1nsRwnGXNiKqHWzMj5imJEvSMSAC9KwiTsDx+LxenPtKCyQAgpE9hqWNcKbAqkek0kX0s4YO0G
YBnynE3VdCSUKSna3xB3SGqFSNJRkVzJ4VccujsoVc63sefF+gE0ktHSHqEGtH/zqmLERnaDHOHR
hVfaURd4D0vcbqGw2uFB4ZXry7NdovL6llNqksayZXBFHTz3e6JuNDK3pBddtpNdgLtqZoz48FaD
30+xQmQQKZ7r/0BjMICtH34ZTSKsMSzIGQbQyTLvK+r/WwZpgCMiTVvbqH0Z4hbecWJxbqSm7pd6
amtbRyd2P4UDhsrjmDMeH8bUT/XaGj0Xmjx8gV3gA1fqynp/b2raRaxxFayP7q1qPVVwGwwFKcTL
B0yDz7orBRcXfYXhVpGYbw/eLj82YHXigYytg7DkjKpFO6z3kD8yOz+oD2fLJ1U2KmApsTZTxcgG
v/AFcqUhKfjyu/PJThAQq94jlQwsMEm8nNYodzZg4aIQp6K2zKbBiGlbFlmKID4Mof7F3pcvifli
GFCpaIVEziU/iZcNDwmRw8ychJajIWlKX2m84TNprt9MYPeLCCnQnqjvTYk/bAdSPf/M9+ce9xgQ
Aer9I0fHffoLUEBLnMsKh4hSBtd3L91jLiYUm8ffGFYvEO5cAPK1ofoJhm534y0NA70bFzEYfltN
1qbX3/Vds53DgGdsj/5KDEytjMMCccXgAsCxg06wwTkjtwiCk//m7P2J8BoJ0Gups9+EOGnPsqbI
bouaa40ChRy8gZ4+/leR8gD/LIC2w2kGH72U3s3jKNRC5kiSXl+ajwMD1bS0ZoDEJaJNIOLspmur
YEp6JVQB7TiHHeXcdD9dIHm9dJKkfO7caqj3wnM2L2OoOpbD2v8JKYc9m9nLt4RBF7860C9xP6mL
LsnMxd1XV4gITWZROeHqFv3uy8FohIRs+6T+qW7D03fIpydKkQ2fJJ7OE9uF+Ad5weVhB9BmW1P2
/4qU4+ZHSOdLC50CXFf/mq05B/E6CfaftlAK/39YxeNJMKLhns6bkwqAadlmciysCy7yL5LiogqI
IZGBNmpJUhFgR/m14FBTfodLB0WmnIUnG0JbpO3/4bBBe+vGGWNL+kATQJcv8T21ImMfPF0teuQo
8DpQWf0XlqMtKa+GIt5W3lNhr3ird3FTrVNipX1Uc+RSCsYUVJXoqcobK20Je5F8nV9gLdZHGcA3
72IBwG2G6SknxCG1zDL1o47j+xnVPYjPHVegN3Njj+W54Rrj/+z0uHatKL1ZFtLD8IAUUbQj6mIJ
EmLw2SD0UWc+dtDQk97QS5QJdiKB7bVYDrfMZIUt7fZjzPLipyL1XaM8NHzcHp6OxJTT6YXgdiir
ENcTpUHTEOYUVHVxc8Hobt0TsCH+LawvlRwD3qbZRAiboXMRMsW6rT3W2bFnfnEoOuR3+glm/Sgm
xGq45toSwlG0GeRZxOaXuVMxZKZXaYtDkiJganhqY+sIazvTc0vsM+2maieAVoxYE7NrtMXOQ7OM
bKYDAFH9Dd9+PO+K+DyavJgMysaXaKBKNPA67OTMJnds48bupSEpFWh3BQEIRpV2rzoUUczB2XvY
b0DNs4UvrD/Rz7qw6FQVaghOxvP7ycbuoDiQhjiNfp+Ux8sdjSabY0iLxW7L98993dGGwi2jR+fM
4TINoktQ2IaH8SYpERDRsqPPto9N+M3UXJhhrizth16knbpc6O5RaD7kY3syND6Gnpe276Ln4c/8
iTeQdFYze9F6hm+DYosp7yCU6QClU2CPhLM9zINyWSX0CAQ+IsdXpZlji/GKJ/Pu1ssNd88BKWo8
jvOB4/YSO+cwCWf3q3sYITnmuzRb3c+PqHWFRsenRirz7dt82Zfl3hmHg/hFkxVLEGZJESy2PWsm
hEDTjAQBVmKTFwJhJxJrx7dGkUFalyOs0b5VUxOuFJx1l1I1NLnP4N/j7GDZzEUUg89w77cKuiMS
Ebw+F8eq0tlgFIBUcxuiyjRGUvtxNqF4jFWRIzzSxZ/YfOTYAxKyRaZ41P00Difhg1LoFDVFM0sI
5PbhRM7/Z6hS31duRySuJC6pW8Hkop7mQse/qeN38guoGFeK4TOrkauhm2Td/VC4oEr3tmahB2Vq
cs8KTOXY7kiljNSIEwwVwfbLQT9QnfFM9LfmcHbtShIPfW6Tq9HbF5snxE34ta8bNpRfu2panXCh
ooI3f8CQXzOYFMJovJIhNXJRXkNtb11R0kZ6CXII6g1tfHBJuXCj7yXXgvtY9CX83hDF+mfinXS2
u7/UnSfNuAC8RjyWmpYYMCWRep1Wat1xFFoAXKf5ssLzkdczqTLEw3UyCMPMBrrxd+l3fPh+wVHd
zllPBOyKQO8B+LnwGFDQHO7NueOebWzwI19JcDWmRhptxs83NoNGgQyVHsAnmDSqHMBJDEVHsaLx
iwbOrR1xDiea0HScLOP5kxbDU61bKwT4FFX7f4ZIpOenY4FAiXzIKZ+cIs/EbHvgpav0aw8xsGbV
LezUAGLMj0AwzifV6TA5DYgFtn/01q0YPsaZcQb8KmXXRw1gteCxou2qN1es3gyvS40v73KvErnX
shln96dUFymeYmcs9yLRgAqC2T/wfUwrpPSIcHOX6ENTAtcKsGzLPU2LUoH73TgVM20SiFen3t0A
rm5SKNVp1JFfTuIrBi19Q8LBFF5uR19l1fOlG8R92QVy2WvC0v7EfiEUun/VHoF8XWdNw6qO9kWH
kFj3wsUQQogt6SGWNmvYUPchtgyFIqCfjMQno+hg9rErJRHRmgbUCCHkJYZQyjpK/m/z8py09nd4
dtDsG74JdMIAQPzocvjbUmGsvy94Mtv+DCJMT297W+Ba9YsIxkY613tZVD79yzoVuf+5v2ZJ6wa0
+T67okK4jgL2QNoyRHnHjcBVbGB0tOIDvGm2XREA1ymWm+OYNf8KLe3PhQIDZPFyLaMBy7S7NN2R
DJq/f8eLjoqMD6hen2W4RR6BDSRlOw5XOkSIB1VG/jZNRNrbYfMlUdD3nyxDut9N+87tafGf2du/
m+v7ITHaWyN6dY4yzzMwkS7YGUQBvApdkTk6dp3jgGhxUuMqLZF9pXXIBDAD55vTmSIPxFSUFSQ2
EYT0ZUDriEiNOA37i5UWdhmokBoH37xTR7cJdCqTA+M5Hw9JWKbuFa7dF4/cBxJaR0lrF3bh3N/2
PwR6eJm98bNKZqMTrbyh7SdByGkYDpJzLh+zRVqYunQ2yYZBF/p1/6DIOwCtS95/JHIYg2eRCI8V
2bH6IqblnNfCdHF6jH7i9O0MXTy7mfzpZhZoHS9F2w/KSDbt4RPi0BUrRJmd1//RmGTjb14SerjB
sK4gX9HIZfVmVg3SdSQvnwo5NlGsQTjhk20BU1vZpsJDqNXIDLsKneU6tNDccJ1wLLVODfnsRBAA
wfz/o28OTgYRECAELEO6RcTYwYFDZ3P6vZXv34qjRyzWQLvq+0GNMPboH5/HbKfBbK+V6C4xEN8T
PDj/wT+i8ozYnRcIkp8m3S92FLbYpnm6wcUAMYVHPzgMFhCkHK7nOGNqpNiJn949ecygKqoVwwlq
YlZ0GhjHHAxe/1qixZndolPFcu/IHuxWYr5mCknEL8KcjB71zCaWC1uc1/ufYbdANhQFiQ/h/gzb
FCbuq757/EyIBtC+mRP9Hk7k7Z8hKPFck6XOU5VgXkYEcWaGvjQSlU4nfZxE4cigsgQjH4OL61XY
HGeHLM35ldK5pBy9CHutQsK9rmmzX24yHliXX3yu3ZCRduoHL0N1Z+KoYTWAt5JRta3Mmod8lxzr
g2ARA5PfUBOj8gzPuO3gJz0dfiZDurErKOZxuqnO/JZ99vR2OifKliCA0ro+s93i8E8x/ixqLDqq
0lfzLm3Qp3ApuaEgeLwQX7Q1/HIaaiurHOCG+bdhdud81VvTSWOLalqGvRJKh4Vqpm4YH82g1Q/v
WyasUapcSdYRdvfGXqnwo0FozsUDMR9GEUayLeU27KCT995aoUcvSKsTkM99sOLvBTJM2ZWTZd/j
3uwznJSKCKz2vUYU+ZfwqAg5oaJJFOe8Fv+zc1AKwazs8cMyXoFA5GdZSYRyLTySEJzn2ggu/b+5
UdruTEs4FCxuLdU0fgvFWiq1t0Jl9ZeFP05W60lMcQoXHvZ9rD3WLRqv5cAwHI2kxGiPVdRVtzfQ
3mc4mZrsv+iTtgwlHIBbzETE4nW5dmQI4v2vjlvHwY+vSlTEHUCCl13BxGZ19gRrQ+wHShkDtJKV
2svcKPjP0Yr6JovTaBRB4ek7NgwoP97May+dbUqFZgIrRxVnJjmuPGq/659o/o9aTKgH/IqImlc7
M8Ad+ZCIMzweI4CoBvDphyQiFTRRqFcF5yCaBrsI7shkc4ET0+sQp0+etp93c7xatcRKcUo0dcCF
kZSQAdPs43rviIKa41+UaYARL/Gw/pH1aD8nFXat+n1Wa5v+67Gh6EQWIYZK9S9wuL2S4sVlx61L
M+1NiRHMj3tISZfGsmqFWZc2nz3qMuOOOr9Ur269ynN7O37rOPYS+9h0AnAE8A1/B1+BQKS2UHGx
3F5+EwOMRT5mntCx/RT4+OQ3avPXlDHgIsNWdKpWzGUy3uWKSWCg0E2IdLZDt1mgcRW81obYW3c1
C3fwYckpuz/rLewKQQLi09SVjmZoYN1zvtL8rv2MHvqfMZbCeOAJeK2v+Prsw3vocx7D5gqtW32g
D5Fc6b3TGH7RXzDLcyPl2i6KSQRgflOMxT2XxnWGCdkKN5KhvlRQgsDOxw9pFfnR+pSt6yGqsXHg
LXrW7szF+knJwx9uq14984mE5BOf8mW5F0pgLc2ErlrFgjeD0ybgHb5U7s0zkIkNTBCsN6gmmw1h
FQ3eworKtfqdJd7JtnKCLgD1ryPEDHAPrsz9goJFlUnZno2EXShqn3TqtZ1y2Tz69qmozeBKIi+O
supfPE3i3tvJBJ/ROe/efrmRF9oqmd3sfFItAa+vOxlThtljNRW/l3MUqkFMLIDzbtwkGcqLC7RN
79ECBCYj9x2eHDbuVTzxQPvojZpNnF++g++d0Ft9/A3dQUx6uBe5VHoeIjN7dVRiRaUgoclrE8IH
05cRMr4XUC45IexPWMwWxgqWzwekM52U+VeRQgqBI1xnD2AirKfE7IECXnQ4begQftyEW1h+6Hx0
kQK/dTyZy9jqwgmQ/Qt8nrcU/8Lg1ttFy2zomJxpqawBljXX+Dl0jGJQusQtcqjVhVi5lSxaNmBF
KyIEM6WUXolRUttmqyRpObum2DKyI7t3S/ZbSCWA86MWbyv3pbPIyjKfFHk+i1RLQSI76AYqFsa5
m+wpYYcrbbUBdKskz+g+TX1h0Y28AqOUP5zVKjwH55a/3L5zMGD/sQy8ahzlF+1FFhBf1tghmxnc
PvyjsgeBkwtvDL7SVj/Z3EQfUjDjYYPCifXEJoT9K894JyJbiTyLtvLL/lvS93DRaG2CCdTJA7Uy
Wm8QEI/qkBoZaOqeLcgAI/7rhmiOmGOr+9ku2C7Ud7Xab9cuvmjm31btkO0Diqr50AbzJMDA4vAD
w4UZRUUJkH/51WepbVAvQYwjB35clBGsIxjyhsCfLqsnRgPiyzpjfCSZo6O2AQ8fpE78I1eZDhEe
6M3hJVbHEnM/ZpHOjzHPQl5BWslJAYjBop/OG+QASanp1PlAyqt+kk1sNApLYyI8Phv/2+wNPffs
zuClMqUzl0dkzqSz/gpuGeBGDse3L4PbLLTXHt0xWdvHH2HtLeNQ3Z2ldFQFoktRcrQVkeLhKXLX
KKfQhUjgNhKd07xfKXrzhcOmc4H0PwAPb+iwWU6rS6xb2BeXFex7N2anpnal1mdLkq/bg2OxMTaX
gzYoLJXwbHU/e1asX9oAgIo1SpfJv7CFlHFfxKr7vq3JTNT+zTD+WsCpJgcGAqwF19cDnMThJXFK
k72fWdOLkZ9/SMrMq0RXoA5fme7UXjRgHmNBA+Xx1RQzdaK1UifMrnMF5IkS1tvXWhcsTwmPtoaB
2ZcOMtwFKnx0l8IA+y5FHnNWtFz3sK/FUA+I7DlKB5tjR05dD1JgZ1HmYPfBzLtK1ySqf5RlkFDJ
2+cEP0zg3Nig+TdBBgGG2nuhkZ9S05d9GIewUtcSh3SNxp/rPUOXR/RFsYsIdSfWONpRTfdW4wFl
77heFQLRC2TXWP+ZZLcb2KdewwGVO9RJJmN46vMOsZ6Xd4M06p+Yl636AV8JxR4PsgT1ctKQVgxl
HpobGpaK4gxXhgKSioZyRnhW7txJS3sPOLOqs8MAhCXjwo3u8phSvAa5dDcRHGWd/1mCy3D9ts+L
yRannQfyiZq62alFxFzYbm4/C7AvN/CldzkvGx363Sc57de5K1PEMnguMozTgIK4etfogGZLkM6e
Hk19jj6E7hXtecTVLluCM/a5HbTw4lGCR1J/DWqPR3vZnv8d2bNMXqNfOnbb7TBpWf9VLx0FIWu1
gtnGjyhA/FxmYy8e5YkQ7qufRPXG5dTqR69oO7GKBuuihp5mKAoXBuIUYIOYowgo1xQZbLKYH98W
dDP/i+VafIspUgj7jYekV/buFvZmAm6YIQQ+/YdmOlD6utGvZPL5fPAqU8rMq8M0J1wWHwDNUIOT
KOYzIR6Mm3JIAXFKhS5EACMK+5DuQoJ7IlRP8O+J77P5zDOkDvj2O85XvnmIzrZG1bxFgR42jhN9
1dhEFbOFsOkEUt9bMTC1GM/Ir/bC8Us67Zn91HwjvY/xFj+NdeSeqg4HFW8V83JVd+YLyjP3v0Ii
SOaSbjLMryGUM7KyHDh4kTD95kx5muEWgDUm5TlzsmGidTlQfqWnr2heFEjy9xb7EDqQ4JPc+brk
yl8bgZttJcIBgQGjQH0PiNYYrZrpGCsM42aCQfrSkEIiCxJPKRd2Nz1wwiWFQ3HxhFS091wuZZ11
G2M+gLircDKB8YajruxeDGX8zfoqaNLhxGnqSj/ml3yBiA3huWcvl6VjPWeAr592sL9piYUfyhsy
BnU6IryZzlD16c7PKj48SWonhQELtyGVw/3ztOVhVNQzNNn3gf/sUZzpT0Da7f6rCEJ1QZFqCKK5
fQlnGN2hY1Mk+oqqm/LOTP3mpjhM9E5XDr1RJ0/4spsu8HiTj4/wCBeb3mG0pvFs2vx+8CMFE2K8
wptBVWJNO5GTXA92enkhYGVP/QQ77TX1TMbz7pguOUSmnRXrTm3uZMGkNmuQ5wcH/bcmyYyHl3ON
5gQbLn55WqdeIFOmj33Lkb6D0T9q2wKmyIsA0kfTtEgT1DlHaZe1RPTkzhumtFpfuMOOKQw2Tw1M
44C21w+8Exr4ZqUTddfgHkh1NWCtKgN6VHeX0xFMhE4/zsVgdRNfP/VtUX/ockbpq1eRaLW+fE07
bV8KcD2qHO6Rt6LaElPxygwfAdsGlRAFPX58RK4duWUyEy8smsrNTFsxpIVtkt7XyLp6GUAEtZHi
JSenVwwdLtF7/KirrzNCU/ffMyOhwgM5FZQmPbmZQlIzGc+fWX/l7iUC64iy1eWqJ1a5x+gDUNid
3+nvrgI1D5GwYsBrOrmshRW6pc9nBcZtOs97Ui05YeZHS/hnvJab7zVXl2AQ8jOzyc+jkXizQevK
X4t/j8AQcJ5wReFuX0bullMFSNp+p6i47iIA6JZGZ5aMJd/8VEDq0JhPO4Or+lMWFbTnnSLDaXAI
RJC2hN0J7TcyW3ggwPJcnSTJQ+Ys45Fg0Vu/0YWWLrwKiXsxk2tXu4qS3eH98IdC8+lBjt6U/AHX
2jczG87C/ZBjeRWiGbCVrr+xsia1+VF0nAc++5utSai2zYS2JM+oOvgS8ZkEjdzo89AfC5Zb/DR4
lOkcrnvrJq4i4rh/9ZYo3NL9FQ1toQWX4G7/HgKcSOeL/E0wz+Q8aiMVLYxMAfU9pS9gC7KmIhe8
qLY3KUzLkKA7yyw3Ia9E0mMHIEqEqfW1q8Rm4QQTs69TctvdsLzFO172hUVnwrrGi0L499gqnbRA
t/XecSNI7KgO+/aoA4MSQk+A7FrHakeaw63G9klVdgcFirF/ZdQdeEXK6z5b3wXBzggmdwkv9uHZ
B8XiowGzhU/hhj28eYVHdB894uSJ5VIcQO8FGZjJTS4PEBKvXcOeg5xMOLmS6MJLTqelcxUtytXS
rE4Izw8FIDjx0or33ecnNwCJG1S09xjGoOf7iCGDg8LuMlxXyURR/Pc8RYmcZGAHVGK7MmJGpeKO
F5nN2CIAAR85nAc4hTzY6dWy2OW0AGhmxPGxwc43xtf1T3sJE5QzJ/aNXoR1c7BZf4nILU4K3tRM
+8FqYozyYJa8ssnsvDC1NjBd6FOLnkCg4DQxaSVNDzQdT72S66RRCDEsro7T7W/l6tDYCAF5Umsp
rOobYEXmEbVmDA8YjYp6I1DwZZTidv9nBLsfmMEDDqIBEU9c+qYnYHs+c62ZmFx1V2b4fP8Jk27b
8gVx5Uux4FQQ/+AJxpqNaaZCJzk3l06oBZYv+ke0svl+i9PDLDwjPwIe3rM4E/B3Jk/cAy+PxGgV
x8gJEkIRpNI2g8t2PBqRxGZhWBvcnSUJ95xkRmgzwIhStfeC68xIcKMIMdqx0B1sW0dMyEX6cYz4
BJZXNgZgO3w9pXAUEJR5qfmLprjvBMhzq+fvMzRWr5Qvey0LOFuCLXSLzue1pRROMzHy+xOkLReU
ZYFCcZTEZTw57KwLygqq12xj0F5GHOlmUSHjYTkKjwiwt302GQY0gMm/jMmXIR1cx4b8xUY8xLkQ
sQ7aCnI7+Sv9uZCJGzJkd7/W+TxHmTQD0Uqtby/xOJB+6mC3u2TWLkPlLaMsX4zGWhsoA1sSgvaT
btN6YGLq4dyohUn02DMPUyM32+3YOvrkHAgDQnuMRdT3OxOpONm28TTxBhmyEGN6FSygNh98zgSu
+NMFR6yLiVfPMLSDz3V1JYJwb71Qf3N+26SaSoZyBDsoe5bSWZR/6ED4dbMXRx966JsNJIS8ay8q
tcUUUwzqHOhd1tjp5W2ukbuCJoYFlpIJ7249yLybLa0T7ON2H2ByS6tTEq81t2aI4bPlyp5U4OIx
EnIX5pcbvOufosMtyC4V4HjlaU1Pxv7/SrFzJotDPlpPryv8f6ZpCLIeIbVsaC27PuNCUpXKe81j
N6ITTDNOw14kFqmGwwdP9kdQeJy7q92Flw2Z/FdFAz6DtdUWLa55QBjNlm38kzfKdObMc1B/XQcA
oqEKd02XXSK1j6rK7pqJlKtJM07qBQ24q91UC96nBjCkeaMIyH/FfQabV9buACuJH0zVdeRGzsyc
pK83gt9W2o/BaFV4KsyKF8Xl69URzaEYG2TcCt9xFiO29oIxdVOsQZvpupyW7SgmmgI2J3TxGnGL
tgG5rGU6+LtT/nj9chqLXMeSmsmVupfOuaPXDqmw4JSIAupNEzHOOjwM8Os6aiu1KsY7Pou1VJEF
6okPclXPR7BW/PQ+TK2CQ06bhvdspeS2LquP/GUE/MnLUmu70tajUtSJUOQc7G7/CosedHN9VgMj
HM+zACpCT+8Y+f9GwpB9a70wE8N2FoN0Abwo9HWrzX3+CrDCkQhts3PZ02hXBv4xeOP3V/wmzc6m
EtsHPMiE23fEviJwkN9aBzeQeEpE3dl0m7A2RZKEo9fESGFqAS2BnPoIS0Zw809WMIiSlkekEy58
yRH1OIowCr9TiYYzrq27N1Wf/Y4BeLNCbnzDIucj/cDb99SMRSFlH/qSdKSWEftXmiZVL4/CNiLb
xnW8Z7rscSBIJoP48N34V/1OMC8bWWOKTBvH5MWPHb0bKiBEsFV8lJ9LghUimKKdsVl42EJIo3a2
814yR51chiU/FnIQMHrIoKk6YisxAgksHFhB09gezHMj2bJSdKxR4RmORKmN+EGp6Dzqy4iofr05
0ejptvSDOFnXmAtwvnqNU0nRfPM4WqeCzHX+j2QIdJw8vTqJllSv21ju+bug5nWVWf6QVY81LPmn
I7idW8sGZxJ9EFZr0DNAM3hfvxdT27udnZv9okqmWsMSd2fq95cCkX0FqW2k6aeZNWCTXI63cRkM
EEeVdGnHMpXbrb5DPKuqDTKOd7N7tk7dJVh04x7tGSF9GzgED0BTUPjA1SWxl8IWYNbB0jVKDhGl
04/9j5zKQEJBHi5kzI8ppUaE52hj9+qw80fGJbeeA5tqdhZaXRXVIqDJ8DTFoj6ZpqqHZg4vfiEi
FL15AkBWmSfDtPkUmiY6gkE/PEZ/sO5+nNdSp2g91T0lbg6pEyqxZ2xHT4p1VbLRzTi9NK7prK4R
trv/rr1IrsTN5LUGG9DzB9w1iq6DVLvgGHG/2FZhVz/PIbF/uS9sYRJihjjCasxMnNRWmznuaFv5
fqZOzxN7N6LEE48O/oZMVI2rbWt/IyHyQQR5iJIFI0PD5Y6jWwqWJTpxvTQiykwHTcxwtq0uw/I6
kzuTwr93PhdvabnlkxPZmA0vtBZ06f2NUI/Vjlq5QulKWqYtxw4hkS+hBbicCq0OMBAlEmvpDNXX
ruqkkuav+v9vAX7FSu2FYH3EYgR0BjnW0o3JonGdokJTJ9DsUwKzbE4TvQUGAZ9s+rruaHsAJ5Pu
AvQXmzifqpgCGxgzUxPqXbOsz+lHysHOz0hLg37/t05E8+1rjQldRGcvz7OT7YEuaYRJw+5jZkmJ
5Gofx5kejP401UbZ2HswUVGrTA70SmS3VoniaCaK6EMqLGcZypQGUD/z+lCp6gmNBpXx43uKRHMi
mDbrBikT7/qi5wNWop+q65jyXboPEvaifvfKo1Ap+EQMAhz4S4kX+loyFc56214PhAn7k86FXwev
5wvIrGD1M9CNN0RI4XmR1SPCsFXoQ+KxJP7874sR85f7zKQwGzNwsvtcwEiWzBaboGsNBJbM1He/
i4bKemcu6nG6DBOqxwdiZzo4zi3zQTFliwHFnX4GISUY7pfG/x4HRnxZpSKPF6/0BpkR2GXu1kaq
DWa+2Xf9Psa+Wqv6B4ZmlJvPROPz1OLMt7MzCNwzPt5dfs5e+PZitYLkrYm6DhVOZGN2HOCc/pgj
E0m+vZQ94hFfMR5Bll7dhxsQpNrsYe3bISkH0mI6T34iCSlk4sSCAftiHmjdeScR6I/Q8Nc/HmvL
ZFAQENewYfPEJ2mwxuLU0Z8omE7xL2DKNJ+eXhPboYNccHNdTSbQqhGdAzguSnnF+5ahByYmPPSx
pz+aMff1TOSpQwsBd7/1kBabXxRNkUN8PJ/8XqjZWD7kqzFsvEbr5jrMYMWbY91rr1A7/+CO4ZAs
dJ4F4Fr0o+FMyfUsXwxmSjnLc6LQxbWtQBOUOUBi26PPYkaF6aB5ErlSPMj8LZG7krbemDj8tmOE
cWBVGpNyn+9bN8ANq1aq9C+FAhDPa+q+EJ361fbpTQ00A9mDmLPGI0smhlOGdYSssEwvACsXuKcD
v5g4Hfy176MbtRhThmWjUxoFvbjRmZAAOvMKz94i3Tf8atSZ4czQXRnXA3c6mfRN/K4Cf849MkMb
Oy0eBkS3KlWoIoiJDGubGtT1JrTCGBz9kzpdHD+sgEkj2n+Rk3KF0TNIcxj9iyBmWUtDFNYDJShP
eVj/bB4actQ880LGHdp9zoWxID9ZbkHTG5jIcfmZP6qoHRm3eF71/tW1ulPca/uoyIE9v3KVXf8g
ZlVCt278g6ICbM6MkpOcBZ5jjDbW/nhGZaukcLIOdENe4P/tUFsNZeCzq4edRa++zVxZb3JSaMjO
DXLZXLhmnmkU+v1vitNGhPb7jidCZQJPwyLb1V39AYTL1o3cti4fFDBftoE5R0sqhucBpuRf00i1
FVx3uBMpMHtLHDHOeCtDuaaMd67OotVC970PRTz30R6o1o6214EFTN7szAvIXokq7NdET97wOkSM
4qeHg1l2ZdFnQD5OIQAlCnb295w+/d4e4w1qy/yV58LmsYBGWPblMwFpyrc4ZNdtdgLWwUDkMe73
BzoQN43ZufDRHArxxM8fDnYn9YDsSyHG5yvWTfy/ygwJwjpznUmdEErSTrG7WTSohdf2sb4PGyiF
XvVwxntnJbNdv+9a+ehAmftdOHV2bJlXJLk8yQ1VA+FBz9i55Mvs9AX63m4ctxkAuK+lgiRAab0F
+HJLaTqLXicw2JXjIf+Y9mP7dILJcuVl4lURPoG27GnLUv0cNWV+naJhRbbuWOapk8l6eRVDaIBZ
wLQUpdVtM58CSlYaSg3cHfD9Ee+yxzqWe0VfBlMxPR1shly6EqD02fTDE+fvIcl80cDwe47RMJLk
uQUyRofpoBREjUkzToPPhIC4U1BAdFXb9RLYR/rHHZZhMiG1tSlzHRaGrEdr0jZtWcd1MA+I2/Zz
t5eO2UoDyiPzfGD89c5gGkq6LAF21xsfSSEWqHCxeZ4zwsry+7ZlnSETcYPuNBFnkpZ4y+1ZRaFo
1fV0PUy/GRUFdHn0Y0zk7dyNrk7/d9E+ugOhieqp+4odK8i8MezoDPUAlzEQoyzZNYWu7cINtElJ
JBGq1fXWaw6KZagCj/blU9INk6FwYz9tBtUYYzs9P754xclPVS+REW6nuVvjoBkHXbbaqB8FToSK
BhtpNpG1icbgRbBV39bSODRUkNPv6tKEhTYx2jfV8AGMIZQFVBqRuXl8q1z4qwI+lPSG+XoAY7sn
8OJpmoQwkS7WGZ2fp5vwaECKmvY0e+wqOxhNDLi6xqjS7zXd2lq7ouYzceZW1uJhpkBcJFJmAiOJ
YDcHOJmwbCkJXonYImDB9+bxG4HwiJebhsEtqXIvoQV1LcxiRMgHMlFDI8GehZ+AqgGY2Dh52yio
9ZQO7aZ9T4/oVOHVwOVtHcor+Ge/j/uB9b3T6NGjP5ySjwfBRLn+XaPO8nVBsdV83RRdXEQksrgF
XZzXE5cZWzSH4nsiTexBn+34M5qXTIubzg3MOLjOoDdktvPDiMqrfRLq15vWkU764c0mTLg6zrma
/ITaIOSF2qfXrFEKVgxHJDiIxVFSdTAn/BnmKYaDOy7l++qAfEkvbtMXi1Dg1AH08jGWhfVpSc9U
KhFD07mtNrhiM/ATvw+l4NUgqqshvozLklao32SADCFrppFd7ciWazsmEZRucQKJONuLiNdPcNkP
flJoSQb3v/9etaFZHXkNUPnJ+n0D/lNocqVYIL9n6Xy5nNnimv0t1KpZVTvUvvXCQ9bihcURxrl4
JU43KrKRJMqL2vj2kEc3cZeIUnCalHH1P+Wd8M4tiRxmoZ9pOSuezKexoNWen2P/u1ClRo/iqb5P
aqxW26ZJs+xJpGuPWtAELzvSiQDWU486jvS1YlE89wfNOo9XU8BQn0B58SBJ5ZTkRg1B21HGkZCA
guhSj2BXKsBHVBbZzeBwQjVNQJgqrojl5s1zZWtzeojsBpbwGenVEcIlw5DL+02J1A6XAoJl1Vok
owE+6um3wUCDdmHd0ScES3ncOoNBS79fbEQvsb4hJ4t3u3HZy9Tu3ZbKGYfHru4bdR8wkRd97wDO
0UWArQI9ZvmzdvBF202+rLDmj2muaWpiEYnJUnriAZD9/f94+awgLdO5cgq1eXK38+EXiYCX7VGc
+Q394RKV0WyiqUuFdNM9zXRSQnay9kLlfq4MsTeMKCqvn4/8s4rCpVCB+lL4eA3/nYK2dpnpxNWj
cO4A11wCfyin8xPtl876I8ED5xJAqhie6jGfUlAFZABIYo9/zj5Eadz1KiRvLHkjVZ9eKp3SRmuD
ke+Y5vT+7Zn/Ctbg58IDuwHvnCA1k8GT3YQolPRegJrWkISNX2fDI0dtVqTzg5Dwu3Nv0gSaLVmX
uP+QV/ouVBVTZfJWFXlCZXsCFAUAXACcN9s1qDJ61FRyhNKGWxFjjhWMq71mFyVjwrK11XGz7mxp
JBbNF3ukAFvl0UoOxd54HysZmqwA/9rlozzIGicMz3wI+vWN+g1+fO64iWVIqiFiNXBwr6GKrGVq
s/k7Dr8egK8rVLLn9zTYdDxR07eRQcQQbsBPhaZiPVZBhhPmqeinwDycNfH2f/G1z7Da0qxzeNxg
F6H/5sey5mzzQhnirpVcPe92eUHlsUcl47nN/9u8Hi3K8v5ywqkgGlAcgi5GSMKLCH17c5WQ4DwM
q/lVvj/OCLuQaMF57bAO+npj9D1DHjnLv3aU6C8jvKWvhgGCjLJMsYTGa8J8o1lWfT5PyfKjG9Ox
I95+1/vEC6310Ucktmi3FF4wGRC30S9I7n/Hq0ld9fTBghZQSUSE56e77uggrkFSd4vXyBwXNU81
tz/Z4Z4GnNn5vCu7FRLcG61aLDltBd2nCl5Lh01M8fQhGBJGy19tLdcAK8CSaOdfSWIZLX8tO/sR
6mCoB2p6ZgngxqASqeDtfV8oAQCNdecKtsSMl7Rwq/7Rs6GY9X7yNsRS+qxmTOWF5gIKQg8pw74x
iJS2/mhJsF1McFzn+UC0T/BRQ/Ibh8k8Xs1jxi65z320abF69ajRa0UAUGnm5wAh8KitFkrNpwXC
DAM/h+rqcxemNQ3w+RDns7i41AgLEq3DZLAfpW2e/VPwdic2wJt3Qk2ieO4WbnW5fxT0XMG9C3di
LlU5978Yc/LU6IaJko9idfDKVBLHRNgcpzlQPqukypyhoCaN0OA/GcDnuABTHxQLFhZvgiZI8yZl
Luq+MTIfAjJzDS4OQrCy25iLqRC+EmKnOPnM06o4aGH5fzB/j4Gs+4TpwlWVZKVU0r2Z23Vuura2
MYDySISJtWGXhXoX3+1aaon0aw1GLCC/SpOcQqcH6zgHkqs5QjErg6BdjuuYmANaxmWF/7HEl66i
+BDeNd2G3emi0+hNM2vHhq71hBuk6XKen7mitOiHL5VN4Tz/rChbPmq2VlzOdIQJ9zJu7FYf4GyT
o0XucAw/2nEkr7HmvN2EPwcaU/nEDomk8f3cK6XmrTvVFItFtOouxJifSBwFBdjm+7GZyuuD62wU
XrxRaslYo6N4NJ+iY/7qJbv0Zj0EArKrpM7Uzn6idGE93S/yGH/B+M50cwPIpCdUx0ihR7i7sRrD
GsWwxpmbs/umaru4OQgeFehCHyBYrIbZWRkadr84uX130+vUMtuacJsMZCkmyKiVZ9kdkc9GlW9g
fb7pcUR7D15AKq4PWO9weoVXQ+AlvWZbMflWEi9wRf3rNPQiB3F58egg204ruCMA3uxc7xiacL68
oEkqfJtUvsRw8VjFjklGyl90dFcx7YDCVP+h6mkvZ1ioveJMROZQ1GQyakFkwOObWd1b3sYHjCS1
Pc+cvxHR2hCI0HrvzO2x0zsxjzj/egS2cPusrGPvV5awbh4ZoZ0I/s3z95RKrs16dYm30Wl/7u8U
MHwMrVBS5Hjd5qL9d+Hx+94svRJ3jbNX75u4TPFgjzLCdVZXCohwoIlN7dHCficlw64rUj99ruLq
C4EVepnI/9HkJ9eQ3kU1C1xP/+BVwMnpesRVY72rxweVJJRaicCWBpseu7PPxd/x0BeOY0DK6tun
Gg3XZKQ0P9im4gL3uA0MUqaKVnhSbJXgzmDmHP9C9P85/gjK9UHr4GJVL8BKYWguf7gXyUw+Qe9d
jTWKOYCC400GaqAa2qxLGzxFiHi5gjnFb4Vnd3O7yitGr+0zHYStCcrpC4OkjFzRLNQWxcuW6zwj
S8shtiMLQJU7ukyvvYaJC7Mn3vbqFK+T8DIhNqM9fEnhNjNGHyMkkCOYPZZ4xIRcA+NIjXjSm9bG
RHqTw3IGPPhiETi6Xhp7L8jBD4I55BHSNmSqhhC89CoU31SfP53xfi03dthSn1pQg9Tc9mCE1h85
SGo9j6+wP/4txaGNP7yoedoJ8qQ18lMZUmu0FkjrP9ANyfbbxjgHxRwKNZyfig8kBDBtgER1/cET
+12zp+vqTKVaAsIWqCL1bdoO0wmRTHl4s0RlZSwutieZnGbFXjBIAaUg6h+W517niGFOLirrNMtR
/Dz+agxQMwGk779TXz4S/iwmXt/QCc2mlJgQa4sxveFps0RY4nBKXLj7Og8gnKCsvdHfH76s1/sV
pCw6A2ECMfu+AujeV7Rs6OG1RxadnGUpkLrJUuMFcyLZ0kuYBtRqcxz8ThU647Eqmr0SXxDS0nrT
ueHmJ6wvigw+18w8chOiSb72gSsXjappMHJHPmFtLK0f+d6rsvk/5ZnT6ZY4NYPXXDMpEn+lGm11
el/zPQu2VKgrtli+0szrQoS9mPc9tpcEiFdnXwPDxwfU63S5PVzwXxqswaUnKN4B9bMi2jInDVpg
JXTzbAz48HjxZz/3HamQR6XMoqT6pDNh99trG1jpbnk6uxmXc7A1MhcXIHB9/035UXplwcjK3OBu
3BrzBxDlFwN+PXhV8GD31fnwr/jQ4H8uqLK1IpI5Ru+INXpPdmlmQ1ej2ki1SAVj8MF/UZg3GpCe
i8rHBwz9PUuEnSJDouTAigYH5gc87KjEbzyjK2IlMM+fJuDI+aN+LCaxhCebCX+NJg/IuWoIi/Xu
I0cju620GxHzc93SbNMEgkuq55HqIooazjpdARRghTnN35VPBCWzgirLqcaSTzluTRM1NJ2XkC34
PjfaXE4SxaJZxYin3kn8JuLzBTL0poR55NhvfWAhv1q4QWgcwGQuovCgnWl2dyY+QwbyRrpOBSGC
yUzpqFB6JH4wyMJkdKZDIQqOxBcZIi2oiWVzEG385ESIzOS+ZBQcSBmd53jq2uMHPgTHZvFxUoRi
9jk+ybXdtsrsv5D3eP25HmA5fDLK1rLHNayRB6DrdmvATFqfsJdXtUkVorztnsmaQbccIybNOdfn
Hrsgg2dPk3kkCUjsTIWgG/FhxOlLM72jL7e5muWif1q4+l1qiLQGkovZa9ZvXLNz+rqC01Er2mQu
UEFizoMKsNl6WB0gMa99435t9691hVfGqr4TiqZyshhgE0wx6YV8UczuAZFgkrKEKAv4i3el25dc
Kn5V66Q7MpaH3YxWxHAZPJR8Tzq6h9wrjWhxAfTrxG6wEKVjaCxGsZRnIzoYF/nhvhNX9R8gQcOe
ucpHAKWKmaC6/uHd37zGBHmDdQw1SMDNMHWOSYwJ7skoOT1/V+rSpRCa9VwJiNA5nG+pYpxvanHS
iQKWeVVYVlPuQAsJij2ZZt7GvzSnLzINlKkbsD+yr6m/D6H3ReqrAn1imKtnF7mtmme65LoNzYTk
rak9C7u6cNswfXFdzEJxGzR0INZquoDG5ywr/49P1DMzaaqaCBAaykQ/RtgPGxauhFO2RQhkRbc+
X9AIE/UnkRLqTyR9UN2W3FueHCA3sM2dtspqkSw1WJw6cvNWtK55auVdZW/nX4MZkFVOIMhAJ3d7
HghrbuXSxvNqcBRWzyOnNlKyq20/w+etpuflCcotGWAz2UYLoUkVu4yJdrn41ngK7n0QDzM9Smzl
G+Enrx/bajiiPgNaZXuMwYowARUbW6ueM2hB9TdzRyfZkmaB/iCmdML+mMiorO1MGQUoDjmyOfM7
hFINObK9dsft4d8a3vwFwsAcUgRIUNgVh6pKokSWv12iQbabHYLslcCV68GM0dNd0VS1nj2ksdlb
gjiXcKuhllE8DwBSfL3FLNk4wpgHgsR5Yvcdi3c32fH6bsrTFZ+55DN3lmEPIsU4yZVVm7Ioo8za
dAqKE79MWF9dt0rB2yXQY/nSJ1WQBV/N6uGsRA9sRJO+FoEgZWGH9mH2SnCt6p9Z7Noc/0K/phHR
/OYL25O84kpDwojBWoL55+/zJq8gjEsSh/Bb4Hb8wMdeL/d48ewx9hYWL1QsEOaE8DCe6lxxjFGt
PX9UD6ZEPgLY7s9+kP8fVgMRZ1tTajAApPZr87pPPlb8XfMCrYYYO/0aL4wPQd701+hX3jOj/Pnr
nmV3VTxzVI8nA2zbgeuMizvRvfdsIQCc9xREuNuLTTzfslhPmGqtwrHSeJZKjsygkisa0OjmMgDJ
UmWHRM3UQflb8116sCQdxAght2FJ+kPtO8ibsQJjDIwDf/QWAzQb5b5w4VnbYVdGcOT1tMZNe+uP
vfqlIYubBcaJsts47ktgf0CoRb45T7HeLnXopgEvbssIs7D0xh5AQzz/zHPMPxmSSvKeOMJ/teV+
j4QoLbLW90gHPt18TrDz9hYICZk573tgpFuxjqCEOfPQxR9OLmpVFJkpCK+8B50tmpY8T2A/dAur
uM1OghPkhFh7L8eXA2D4dI/AM8Nc+NNfCUoAo2GbCSYdryG2j+2G9EyaAyZqyhHC9DiefZcLHhTP
VKpETkYN4azrxVczE2Pz1C7UcecdEmczR0Gt/2yek9QnZf02TdcA8NK+Ge5AKl+QftWz0iWJSTGe
D/ABfjZ8nDTiAvhtmcS9WfXpPggYEmmqeSqMybolL+0ZkxiD6Z4lrg12lffROlTX+US44AC6BKLu
dmv6qr3uBeP/GkO9Mzbrq4P77pv+yGqw7Y13E4ZMr1pWZw6jJZuwL80Wcz+my5s4pf+sCppk9eQC
RMgNi8nhR17Sy6Px0eB53PqChtZDi6XzHKNQ1lXshpPcllEmfXzUoBWXB5tuQVR6p5wVMmehzcBA
I/EJhJRnBkRovlGVQAlVQOHK96KPaECQEeE7IoTIo25ZyRs/uQ7LsghB0JBh7n5VSZQo//6EDYTI
FH7Y4yR1py7xBpOWRuCCyH6gUpgVxGLoUpLGKZXFa2km8sHPNhDoGPjhAza0bPsiP43oZFZ4Y4po
y0FCa+ncDsr9k0doYYf+dtX2X84fMTFIPfbNbBq1syvSW6GdiUVS1tSj8FkLuDsbR234ghlwQSVR
ldja5+4RvUA6mwfy6K+mcNtncEfSv2Ffp6dlPUYyXs4/1Rm1fW3pstY4KLYlFbWUTIMdj6v7g9Zy
PtesiXbCbdFioLC33pXx4Qi4JdAFW0BC8hZw5nuCIYYzNsiZgU7MF5NE0l+7oitYTHZXhhHuFl1I
c7vprga+QGBPdpH/ASpryG+G2n5mHx9sbP93ZnTEaBQtmfsyG4tl7ZNEMI+iubR5oHR3t4i75cnA
d6Fp+KFw1WB9c/awKKlnrW58KYDT+ia5glnNwPfIBBBk3A7Z2KgHud5p0cTFPhTBO0CdwiUKeptH
LA4JrYVD7FJ19eVk195s9YskO4Jm2Gb+BdCKJrFJcWc/cY4pnONm+M3M2FsV7dcdiH9AAut9rW/M
cPlVvh4eedrtLqKc0PrziRGgZ+g8ZPhlYT6WebvMIPY0GDLIk8lgK0agFXyebC6s/fTT612IbaSU
mynFTQnYDOAElVv3xJ+2vDtRMdHQFec6VyA6fPbknIvIPB39Cw+sQ0fmlTlMERj+FgVI+zZQvUnX
OGcKAyeG9z2ucfUCdWbiVQl3/m4qYkmS5LBi6QK+gL4xjnjT1G//QESSqVBQVRLbQFi8WTZUTwn5
YhStZv4PxhriODo/bkl3OGhZ1D41f90JnjnULAIx/JTW9h3sILjjRDUbG7+Aaq+/AmJ/hOqkUfi6
YE2aS10qnGt0cKTEiqKjfBYtGuXvBimImvZBDX7i0tntAbhx2DFpQ4MQjNq2dnqsDRgz6BMKa9HZ
i4rZoE9q/SdAOzzb6y0qnSpYF/cGc+kX0sgH2otW+A6cTkUAlD7cbw94ydsr0i+atIH2FMuQkfjR
y4siy5qSD4/fiea0yWKO5KGQLNRWKBnA+PwpF5b5YueLCBSMy3d3ArnrD1gVFj8CJSyU1KmDLqx8
TVSd1RJ6o0ooPo+Lihjs52r9fm8HezE/7VZMHnhZBw7wLqe4TSzChY7/w7kCPcrAltzIpC4o4WH4
Iw82XwWLuzJ7RI8135Qo7Xgj/cCae6j2mmZFqIjE/qRt31Xfx612RGNNeKr0QKk3JyGqcYivjy2k
Qu6JMBO16fZSeVl7CpJevW8VaHV4qvnELdc58k0Q5WHdVaLYMER+Bd6b72AZmXmZ+keuGkhflSPk
sj4QcvrP8olXvjI02P9op/yGmm2ZCHmTzuWyec+OSnPnyhMiCcNRGBPpZIrcww8kCeWc25ROjCc8
D5YHZZX7pHLiZyUbKVqmRG+xEYRUgg21oazgML7BLpQ3vb30/xpc9x2dNbCxGHbc0U8RSiUdmJlE
t5uVYLJnMHDxSdUgsCRM8Q2ngsa/e2FiFP2R9QnnGjT1ew96GScZNvyjWmIa4IWx05axMaxCa3N5
pkbUF0Q6seU+1KwZq7Ikyt8EaE7CsCD1fGBqeeThA6Xn+Ylgr0EvgGpaYKoJYLNgoERUfxcrBR23
BrcKwSeMDgfzQayH14vghgSmPN5RhN/lxyNqvr9X8I26KyAqNyIM6q52UuOY7OVcmExz+Lwzt9Tj
l1oys0M5zDde1g0K8Wyo3KiqseJ8XUzWk6tXx22ZuZ3L3wGHlc1FlM9ybdOvd6baoVT0QfElgRIj
EhCfO2u/okbXk4pqOsP24uBw45SPK3UNdBNYdjqfZ1VFgYQG2TE9lgdr+t2d2sZbOePS+NcWIeB7
DVfdrIq/PVU/OdjYEUXYPxf/uLr2eiOQ+9EoUMDpUDGuZjNyf6mnLPYHx77B9xmE7mjhqUEcESVz
/RL6Gdrnzk91g3+uYf/ZPJV6fik6HlpLRbDtKZtrzTBdPwfEVWtQ+6rAKFqk/QyVHlR2X0RDxO7P
DXu7LlfTeCRfOxczfYRrQxwwQKceNZ8yGENs0aFMPh6k/7RwCB4eodx7SBT+EX+fMqGlRop5fubX
mkoYOBa9pSY5LNiwQEwmPXOnG9mwBcYIumlcJiaTVPZyHaniNRk8zuD6voEABcA+e5UvvSzHpTFC
L1s0oXBf3cEl4ajPbtixVrf8dtOqj5IpYcnlp5vCgQuM5FZ2sAZwWjZ3zwUOnWreM/fZYtyh5rcQ
mjx5s9w1i1pT1fHgMxyPtzOegydkOW7WUK3IBYp0I4kDZQq/8MBh57l0fjl1CpXdpeD1C4NnFYOJ
Ukl6w6THB1MMhTNUN3RyW709cn+ydByMO1xCz7eUPYgFsVVw/5FvAKKUNwEUoW1ALXKzjk3GTNCy
/6mH036AL8E0AkmbmD9kdwdqLxGr5ffBewC5+Zkxe7+2hyodxahR2rrn2+ZNDXUtdvw8Km55ZjnK
fNnclmqca+SpKXWLnWSH93Ul7nVRYVZfLl26Tl00rqTRyk2nAF1pGHqy37Jxlx6JIucUat1ARTyP
3SZdxpFBXZi5fcGT31hnRZVfn8MMhLTPqVu2djKCAvcP0anXLvzzrZSpugA6Ks72AMOTnJMimzI+
p6VJmB16bZuYvHmX2m93ZrxDlwcTDQiWaGA4p8uhpBZbRRLYiSKUsn4zKT6qaZHiE/TZtBaTIx8t
2ws9uGz96mHEIy0uU1nBzx54XPlg+TAFaWQve/9mPjt+oIaLaOZ5Ns4sXv7tqBYAMPNioS4O7/TU
Vme2ClPQiRakdhohxdnibWwAfKw167ODIkVclbqgBYX+AZ2Pv13x+JwLOvMJEwb+K+Gsn9py5y1d
Vn8g/hk3Um94IjhwTnu1LFMUpdpencPFuRWf0OEqWKNAFPIgnzg8d7SSWboMMP64Y/cG4fvQltu+
pJqi3y6yxeNSdPzQ9zq4g3kHAGuqBnJIy0aBxbJEz35hBoz6Asz7XhTP3gsBxdwPlKT/yh/sBM1T
k9sin4CrYXPL31VkX8nLrCD/933dwv0bNfjMOAnlS3B7AQRuOcolTYyRIfBWbYIj3ty+lKLuNjs/
DvGpv0kiO8xdoPA/skM4i72T47Pjhd6O9dY3OVgxS0i/qTn54D+uc3ql8uw2S5b2vgL+m6SbCJtJ
MGM+77ZhCt7/fQmFqg9noVl8YxZCUfZAzINxMgtByxD1Sd8PYDj9L5SjmpbtZddxyrPhr8ly0fM3
1tYQOgt9Dl4Qas5ZwZjW4JeqDAzumhb20FuwbCs9lX6mK/Tcu8Rcc53qyHZlNLMtvr2JJBIhY/59
5DeAgC6mhshDAgLjWdE8/VupgP8Mm9dC8Or0wfH+sYnN9hI2+dCZh50rzEAEMmVW/QGdQTealK9V
0uS5vN/KVoxtp6NZZUCviY9RpQOgIv/iAgx8OR4Jc+9h7yey8KztAXWTYgSICkNX1VrILGI026pN
SKVFhd5K1Diu5l2qQeDIys2ibseWBJXKioZptx2dAA7T8EFGTYkVQjqP1KkbscILiWsJDkLNTPd3
NG2kJ5ljC20yAnRCkyvv7jA+rnZ73iNZujX5ahhaEHREd/S4ZK+Nazzp/n+6G7XPNJr/+JyX7GQW
BjUDFe1gDqvcG23Qk2+6DAer87Lo3cDO2SE9gF1lnnMQKf68/b6q0xLEOzjOc4W0GNkcAGH9l50t
pRGMw86K82i2ND76ULNk6skfaeIai9z4fkDrplk8y9Y09vNo3XACcS+tgsAvRDoKp59ZHGMSVS5x
f5TWtVTe2n7ahdkzCtpFO95p+bTL2gjQIt/tUCVlkHoZvoo6decJWNT62U1NfseXf8otmhcNSnVq
ryAb1TfhD1BoBNtQQL9v+HDyzdwYC4SQGQWTzd2xB0Zpi6AAhZfyuk7E1frwzCO0gD+HuJAPFcJQ
tUBtiRW5klti0O4L8L8Uo4x/RVb4eaNpLPuapRrmzwPANF7P4qxOrJMbT6LnYgyKZdifR4zeWKOR
wEOEnChrU6XeqgcLbkgA9S0zV+8Qd113snOofm7bDyRDDGUH44hgURrelQwe4kMVvc+YlxngXRqm
1lQJTT1Ka+PUVyyy/v4oeh5ugTPhAXiYxrLUJQCKyukno5PHYQxoZVvBWkGuWtHYDhGNLj7Ev8sQ
Zvtv2epd3dJpa7klKpZml4lD9Nk0nGg9j+AAtxtzT/olhUJ2/9KhNOFFX5bNFTikI62Blk0IffIE
KcpGsKTumQynrTmjIBMvU1D/NLCptZw9YDXMR9U983P/bOksp/bCECFRDYutHiF9oH3q5aNshKTI
c+yW9mDDw3GotZNQX5MU7i/CLBQMYGVbCmfX9qGBj89cPQwAF6vrBb/Khw4/ob8Xv3hI6T+uEo42
FPF+JUK6KSlwYENkeU99CoXXFG4k9B+7hD3Fgrc3nTn6+dogNP02phQ6Tt+O1Yn8Na4tySHJuxBj
+PkzAdIDNHjSh9EpAITUk4p8N0HJbwoY/y4SXYgZgj30+Z1JAkDLUang8sbgxMYqHPDoVwJBC85t
2SD6x28BQ05AtrLT1NB0rhj+1O6Lte6pVMpMwj8dpSLOPoGq7hMXpfuWY7gJuQSSioV1L7XxNC3b
sGzmY877jUc3aKaquKQwh9nKqEwTaDOs1gZoh+MT9mUUjP9uQobM97k4nYXrQsgG7m7U8QLagU8A
XAxO9JlXj8suJQBDtSnoA/BzAxIpBIqF4Ot6uMmNds1R7SfaBo226hb9ACTt6syr5gao0yWAjx+I
tuFQYwkDZq473s8nya3YyAEhVIHspFaFBWN5vkFiwO0BuIi1MMIk24BwwaeW3WPWDorlA88ynT0A
+1zQKuWWtsPu1FiZuFyBMkcXnfJT0ZsrHsGi3Suc1oINQElvMxEyMQLVP0G8dqvAtn9ElWsw6ehu
bURgnd6nzZ+Qii08b77W8wvAZ2Fx5hhhQvgeDcrkCFWCc4Mgenle7zzuJC+sJnS7Ndw3WbTmNTul
mgXkx/VJW6tElR3Skt95M9fs5QpUzZdXMRhii9oo9MejRqQMP5awZ6BDBh67+7QjgYpzl7JrRr4V
ZyOly6Vn5Z5WcqzbAFcg9VIxy1ofRu5NhO3XkBe38z1rJyRVdRjdruhlNYXB3f44+efFYTuVYXez
8027xB18r0vRKDx5f0QvS10TpA+7vU8t6U28/rznveehz0drSkoVlq8rBnqwT8tIXKyPj+X/JERX
000ODjShgsmgZyJC/GUDz8AHXw3nMD8WX8Xb2gwuWM/Fp4B0SAD0XC56CjdZKUxuQu3s8Lz9IMr4
aF0O/+EOt49rDS9d1MGdtjFL36bRvdXZIEtEP+ztq+8S8cKIuzH5O9IDljuxf49tq6P70zjZMG5w
ar4XkBf4YmH+Tuo1w7O9pKfsApBN9MuxvwaxWVoFMmJmbIz/ouof0kbPXNiS0ChZjkizqFc+toTP
SsEnurC7SrrzvLs6XE1Crv5g35whhGcbaEE3pL9yE6IENMAUKHWZguCuAYncPIJwnj1eVhpBd4WA
yrP2VJD7PZzTDVd+xGYdr/bnNSfEk3+L4VcSsAQkW4FgKarspyzcJlC4huWu4AGQZKYU8wiJwM/s
YLd7cieiidfDmNsUgFRjhVX9RUiZ/jBkLrRe4RHop/VrawZx7pmE/41RgvsQcQRhPSQ0R92aoGsT
EbI/4tnY1Yb7VL3t3HejpZWCXWKwdxAdR72uGqk02Eqc5xwLdR1CaPFEy3eLCfXN9ApEWquU8fgY
/dn4QPZUn4T94E6voc0Ohmr4S9+zdklPvzXnA0CbTis3d8MF8DaLwKbiNNkPHOr3TMIZzwE5l9gq
O+O5Oilrf+/tKqjqMm595Ld5wisvx3OrGXje0Mj/ws4ktiUzmH1seVxLqZD++/zePET5CW7RcSNk
ZrMptqkj4cGvDNL2zgGUleIJhNaEwNNBipESmprQ4Vqjv0dbWUDMm7zZE/gaNVEb1W6alzxWcR3/
WoX5VaLDRrJf7Z0NZaOA4jlL3UheyCsmACMrxEuTIuKjyJHTkd6pOR5/10TaAGRg3MqNAAiNOQn7
knSHr+HalQwmKnMMYBMa7RfOUXyWcemraEpPqV12HYLlQGnU04lktl1NBeeDfl0lg1IYbJPREMnb
EqXMq1ilPnTPQC/GdFvEVQinMUh8CBoBcVwoxzFsc4exweiCFf7gZr0XCUyfmWwNQkvgXR37xAyR
BhMVfJILAr9TKvrcueGzP69CGFqU6Vx6gTAW5l0/rpIFAfwfHTFUQJkvpOXnUjLcIgmSq9NL0we3
Z6EBUItx+ajl7P7LWEyXL3aaRsimVayJh3czIWpArR7kXYoJVWTZ2n8u4tRZ2L8hGqmDQoiN6a2Y
7HoY+w7Gs2eX2FNz/KFrfOea2jti+lI/e+auiVELabwhi6rmIs5GO3NJPLD3chezAYpBYhy7oOlV
CqGvjGKA/GLjGj0NPk1hmCm/5tLc0eEuD5sE62DGwEGb6YJsXAc+ZrlwDbi9Qyu3Jqz+0YFmCTuy
/fvw35qS3CzhWtpN/Yz1huT1m0zfGRccu+zDU3UOUd2s0bR37iwPMIhV6LnCLY0o7j+kCcsAJLmN
i8PlAXFwGTJYR0e/3t+Y+EaN1ykV9Lv0lGPObTLjsCXbQ+q42kjgeebMD77PBsI2vRayfyX+JUEA
xsFs3z6TndlHI2oqA6ayL7jzjx/QHGKXQxBWCHIPrxt0iwe+TL5AElJauMskthAU+Dobb0+KQRBC
hb0YciSTKzSJLcL3A1Y85hCj0r1+4tFLZmWu8h5pRgc2bsf+p4UFUAf+F0ZrkVbyDquuv93VHP3G
sDDZroAmUn+lf6El4kiebggA9rc7TA1IAU3aO2rC8hhnoM0Igh16sAnocqelq1xu3qrQJwfFoud9
IXGI5gfDPtlajlyrlWV8ilI7fMupPXsuSgPQPrLnIRd214yOIULy8TawgE1KH1+zKreEHId2EIh9
qtuqsyzR3jpr9hRW1d0yfwL03aPavmqHGzTpMIDOB8BX9/j2RY1utvE4FQqmeDyEPi3RVFUBNPeU
3YicD8joSfNmIJMoe00WnMp+uU75TB2QY2SRBUW6s757fHyaCeo8O7kdUk19Wfx8wijPz/9kG9Kl
aCefmOxH4zOx9zmyu9MKNNnm5I6BZLhAXcxdZVhKb5uvuzptIRWebm6rI3P1PYFfP8pLndVRhT6u
WVVzt9XPU+s41E3uBQwx/eIXtgyL1TtLt/flhKrC7qx4Rhmnig54VRjlTuKGpTfCtAU2N/plMeHq
Nyop/XI1a05niWau0kljN15YnJD9v+nvs6HkWkDMy69akfZCnTxahBSe3huQdrdgMzEgT9h6GXGr
vZbjoWWp8iSX/0fpX9suXHR30wgqtNOP9aCmFVvVzgpJiiTawLahgh+dg4F28VV+IQIFpjeHTgOl
H2c+jf7gJVLsGtlXc8rWytpv00lNXPHCJSgQmVvKq5CzvhpFCsPYWQ3n7w3vIgIE21vUabjhlhDr
AiflH88r3JLLcX6S/tbvxsnnANQeI5S3AiMX6+lJ8RqQLl6+hnNWzFJM8wwlXkFmr1rvmg1u4zz0
mSeX/J9rKjuvlTgo7/O7dihfRHHBvBwCG4RugdO6fmJKkuzhTTasUQo7Sp7c+ruldHuV/P+u5Ooy
WSKUHIlIj8dCizZ/L4WnbQ15QNnk9Muu7AMBYzCXEfIlnxBTF1/jABPM0w/vXgnHYU2tWkkaoSlL
3IvZ/dQ7IbqZgoR1i98NYQT3bSnB+N0NyKml0gFVAPdwqbXb07NlRMaU3EzMIcOTUxLpP53dQPtp
Ah8IROSMxfwOCVpiRTjCkOPADJRrrWOVDfwQctbFN6/D60BzNkCMJbMU0TD+tCsZ168efR1yYkXL
ltK88GRQQ/v/RW2R5V2cDcVy18Q00LWbxK/n3e9UYQA0wRnpD9DhZyViDb9B/KrplGe+SrpRX+40
LPiuvuDvsWGY4+cQGQ4l6t0MyjVt4EWthNmZZzitAuhi8BDBeCagUuO4d92MQKTPVKo/7oilH80l
B0ik8K2zF7x8tV9SOVnt88zhaWd3jnjBYErYxIm+0NL98f5XMHl+tRhpurJQSTCEXwvFbPTB2jpu
8bRe7vtxmZEtavAVopPvqBPYAcNC2MRNNpyu2Ao6GeQWeX50mz+UPXIvzAD1l22YJHZy73d/EpYZ
yEnrbMq1kv+lO03JwrP1GGn+MkgPl7qEc+SnlRs4Y4yVEW4d2bm82xvOz3afJ4UPGndIQhIo6tab
V+bRoeF/kBU5AqP/yJXf1FJXZBGWeoGYpZAPapzcz8xdi2lNtSUHCJ2GhsSg0qnbZPukH3y9sxnU
BqoRtSSJVwKsAD44qlSYnKDskEqB+wxaa+qk+YEdyEhTKItaZup/THMxIUmo7OXF9NXR6UQ5er7j
pOCCvBrzJRRTtM9ZtiDS52GkfdxoIEzMivUB1ncxncdaWkQRoYaEnNRgKIf7T3Cd7InzZSbhNpd/
hlQFA4IxZw1YONMUXfsyIWJPt2qDqbdnlFHjNPsXShDHS4olNZ2XH3tBastKSRGXzsg7jDK+fQaI
NJY6pCANdd9DR7Bu/YQCSdKErOgkGT0vehOFgj0guF+TbKHXTcMr1JSmLZHPJmTs+u/H6zJn1qs0
hsjZyp2oaBWZV1ZpcvkAhUs0A7R7IacqN9cVvbr/eYC8JzX0XaJY8Hr5ea66B4EmHb1V4LAgn/XI
RmC4XLAOanUK6SKA8XDeGKMB3uZe3RAfRWyDav1FW4SHxx1nKNfCmNAdqdK9IMuHu2bzXNTbrH+v
dX+tmrqaIIl9Sd1OaENMb71099ijiHuopiNC1UXo7zgQwMx7fzucmi+KdR3IWeX9YQuM6KkIXg4a
xrQA331h02dkSo7kLBrDKwGDfZiKjYkG+ETA7i1WdVAS9oGnngzjMLkAohhmiC9e3dtD87Z4pc8k
sjJP15JhLJydANldb/xrP1EKO5AUdF2N8jIDN6gq2br0TDhHlhVm4CfkPw7jDySDoSBTsTJkBmKi
ZgHYNoZfButLXUo8JXa5PnaVmr+beJ2ZWdgYv+JqCs4GI6WZyvPssua296H0B+iKXfD3mKnVJOAy
1G2QTMOYmsGX0rW0qMjLYIjUQUHs+Gq0zHO1slr4TM8+YoMIahAGOX3Wi/n/JBktGY7yuzeV8xMv
jedizvMq2LtwUKlP0uswsiFEhINWcpEGNLF/CiflSLNf0EC2gdTY24wYaX2yiROw4nlrhG3C3gKM
MMZXNNBkuQeo3eW+QaTPNMLpMv4ABLB0Ee5pWkVk0KY2P1wbvqfSX879AtNjcEiXkPD6uXn/HH/Y
GPVdEZnnen0HwcUm952DB9yXWMzP5KqCzQqWr8ixA+NcAbBbWBku6Iv4k5es4f/+y+PmVRI2QTCU
7XoJvtGtP2gI8WVPf05A5bcE4jUnuHKwwr1bfRvdXcbaqdzz4Myi2TqRmOF7SNLCH1biKMzV5fnK
7HFSe3DfKqb9KsB40z2H8vJW8eaMP30l+Lcmex6YNW6rqQBZTAm8TdXbmn+Di0Kh/SsVO1wNO44M
eVLQv65ntIjg1Wf+EW5kjK2sunGn4ZhPR51IyiHh/GdvPzIIASd1y6lwGNDt2uFN3KDuVI3/ON2l
onJpy0VJ4oZpQrRcNaVGc2+1Abt5dGDRVt8WvCMTvFIC/eqoFENQTYT1ucXafJ9UOdRN9dbxkQZ6
WDKC7nb5OXcx1D7bM+BaN/X8qlLgnQsUlLAxDZ/Zp/kgeCgXsr6znZtzzncTvVYMcNwLq1XXh9+Z
WhE87wS4khK/jeqi1ll1appIw15JeDBe1doWlKFH3GuM7ATzESotF9F4AvfKt7228l7hWWx62Ywr
CsNI2XUaZFm/url/oJ7b6hnuzEcqrXsNnBhvSI3BKGOAs6OBgKeulkj300O93fePd8L3UwD0nKFA
L2Qh+fy9gyS9Kkjoqhz9F7SwrqwBv2G8FIUmnnHxS/ru5qsNlK39aaUQigfY550INM3wnYi2l36l
L7HnsRzz28USCp0AHHYSjGtVGQo7gOFgKdRJvjU+qGYVgQmRolNQaP3tR7DbPXVLroNj1NOgSMIT
jMx3wnNccJiP2NwIUnr7p00slb5y4rDAUoTV3eVoph3cdkakzeoTKIau0K3prwgvOi5295TKaJVE
42gZFqi35rYU5lICtubrfoxe9uMlFo7ECi9t/erFmTpZw2lrFSzYZbQ893Z9fbEfFEemeuOckSFb
SeHXGJcxJpj4e3ecHLmM6vjNGL+G9CbEgsdu37g06WQ+s9ExfBgmKGkNZK5oKgyltZdTd2RPND0N
XOHgjjb7h4D+ltpQZphAzAP0MGJKTxgVNVjONvKVVajyo5pvnJQfp8+KEepq+8zP8tEed0f9l8nb
v9VMgT2XHW9um5Y0w9m/oo0dT3M4mXYuzRaH2jcA5H1MYhgRaO1Pjm+gIdgDHKe3rAxKFbPux8gU
oi60H9NhcuUM/CdOIf8naDtqbJStWWTn8W79LoKlHpVK8lPRFQrMUbHyzI05I33A6jTIXAnDWB5l
019UaSSWL0MoaUNcbThWkY9vi6DB/Su5+I5K9R1Q38JHaP72qm1d+0vZVbp7mD6SgPeun4qosxTk
D3efzCbY9KenjS97HJnPVxvtv8Rl0f/lTBKhGEVdhJpwvrzNc8QZo51I9KzdEriGrnTPrfJKqQCn
Mwjg1tMU4QYmvDrX7k2GuE0qpRxLMqXs0dabphFyELiuUQtcdLHvYFQqiQ4Goncs3y7rjlEFg/5P
JzOy/1qTv720FUrQOpn0W3FL2e7ckdJ6iJdWFW6MIM1fXj6v4IwbOKMlTRf1bQ+DecoBwjgNCvPd
fW3sZuCbbruGFLk32bHkpZqxyIQ9s2PlCQKOaMxAIoJVDr3WAPCW8DzaWt3pbvYSlwlQ0VH8ly0q
cL0yMyuKzOdDAzBKYWyZXFsZQeKRBHLLFc39pDSpDeFaNTeLhzzgcdfnWzfdNoA8UOSJK6y5bc1t
sOidmyhoidFlB+qsYyuWQDCHR8Jccv6HoNNt/FiANLIhOJeSY9giU7icJnWl2vJ2u+qoPMFcP9F4
LkOkpS/UI4EJbRyeCIf2JXr9DjeWeBU/tZL4stmbc3mA8WD+wAsi3SSopbv8eFt9djrFIEV/gRSw
uYKikGjKbeUxVxC/1Sbjz76WNeIImLXNuZxAM19bWKmR15cW5OoPfMNT9dC8QPc797sXIXA92azS
0qAxkglopbi3i0QG2FLocUiwdApHZWbloOv3Iqb0pGe4l23Y8ZYUob/vwJfQMtbQKsy8ciyqXFWc
vG4Hcywk+nY0uVmwIoDhBsZNMK4fK41LdaPzsUqho5+whaEj1/HBPSCjWEgCYrmNF+kk9mCB3+Fe
j9TzAt70EQmOaSr2kBhdEbDyZjvg2UDMxDOsBU7cVl3EycJ+kteIRFNdCuB2aRggz1AE+SG94Y4c
SbBhOpWT87Emm+4MuxxHZzsPa/RwFHMDHwCWWSYi9Gimlrml3l4qU2XVD6kcPkZQhCIrUMOqwwbb
hPq2frz4Wxwd+4MVi0ulhKd9x7RdXuGxsN09lAksSvv0PPywsrWF3AZjfp01PNVuQGit1pa1xFNp
XLbcOEvCImpysCyy2O4BVsHU0XoGT4KJdm6wjx6IO8K8GdgRTi33QeRUrK+r+QbafU69vkaje4xX
kY/YYbf76R59xC3yCQ+z6csgU8UzuPdxDmwrGte9dyUziwFag4vzfL9kDaH1hSQf9qxun7ndUcWt
JE9UShpJrXl0Vj2nqKv36cTbXIhToqNDfZaxG/gXbrBIGQSgHBrPejZbJJ5zZetlWO+YGZSRIUJk
jG8s78vh99TgwEShNPxEAOa2QM/ts/mYDCBHilGTZhH854cjyrnlhnyrZEbzySflcSFc+cEJjSeH
NZSzRCvZIsax7Wb7t35dwu4s4B2Vf57UgJUg4/TBAHz6jOVc+Yqs1vK1RZHffA0FfEmoNth868OK
FybPtlIEO8R5rnVHGmVJXfSzCPAHUtQKp5veij/A9Ml/d9fpXKxB8EYny7Sj6XSDergL7hhKBt2m
y60tM798cDGSJAkoR04rpcLjSMKM6lYqBPn3QTOr8Npym6TcvRh1uNshKks55ARP1pQ4/XkS0lFN
AJjzTbZDrGvNbXmTBbwQBa5xyafa88KLRhLLChZ4ISCxv9oAn0MLjobq698/ebjZD6CIdL/qCNNn
n7FhwFnjU6N8L+TPVQ64DpUQe+mbV9VYDFd/gZn8gT+XP0ztrYJmoUzXeh0eyUadqU34vHK/RZWo
ehH7ybvGE/1eF4jLNM5azre7Ol8EByGDGovf1PxvMWGBHvJAP+SA4Hzvu9gxkVc8ADQ5D7rbVtjv
1EOhMWaEFTkUxkR0MJ/FdV9BgfTMvPrB6xz59CzJjZa727vI6rMU/T6tWyY8DuGzrbYCmoHzMmc+
XBEblOtuK4aPRcQdzFC4peq1wpy7NEr51KHiGY6F6gEpEMAPIYRYVWMKM3pDJe4wT1Qzlb4lZaQE
EqAy69GgubE3QcG6LrZ6eNzL9gEYXFAtdKCVyydODZx3sT/O4Ozss1mzieBkxugGqboYyPPHSssR
oxKi06Pu9DTZ/aX5kP3G15Rz9TnNBQuA7FjDYeQ7sGGaAQH80REYMbexk+m3cs2cv2VmBKV0Hn2i
rc8m+XHoJkHFsotjTCFkSxZ+WDIabhbmgh19iHKHTWZ8fwktW0dDRk5IzzfSwU7QNxt3P0sbIZxX
ZtkEJNNACnZuxSE58XQTO2aqIxvkdV2E4S5nfYU16EWkbJ4L5MukbKcrnzj8F30lboPlMo0KuE7X
gynA45y4PCbSeUYPVimLduBmZ/tjJekVU4KHFRoRycBbixk44KyEEa0gpHYWINYUUurAG2PKZZav
s9iikLQMpk1hUiZD/vpILhF+8T+PW149VwykgSNllpfdvVFbqn85EITZMknyE5JHAUXUTgk4nBgK
YKtwgPYD/8JNJYFnC25HoxdFVXSxOY/SjnBUxadwIcHgRX3MuOZWaBuS0yo76uc6LMWik/R/HlzP
+kgKpg3p+fAXeJTFhZ/69rcGguYLmvuY0Z9p0g8UnPb1T2nsKQRfJSXgjbcZJMibgGyn3lDQk9V/
ltmRVoRuCgFeoJEZ1x1K03bwoKgZb3ecAlYEZv3sDJPSHmGi6k6lQe0nK+XbpkjWXDcNnl9pidqY
2mWbcwgvbopNx9YWTI08J/+cLT7Znz+nlH75GtsOWpkW/Nqgn3hBpVQGfIfhJzCyrkN0Q2AsEo5A
D8gpCLiFf4SJkcZ6G3avStPiw7TF5+dzLxgf6Yb+4UgKD5EzkZ9nxjusNVg7OywqoGYIT1g7jB4k
xEaMMETbeVMi7p7kyfx7DGGFtmN+meenyNtqMCOA3abRqjxiVT2A8qia0mvBqZR1odj1TKjCAzY8
GCRHmdjqflcNNDrvBSFw0ndaNrw445KSJxDVw1AkPxzF+GElCMNjafLDkul1lBaAj3/q8NJflcTv
OZb8hh2hqNWouFiWPZZ/wbtO0jkX1SAJZeLS6atzDCPWCVXsiHVe/galkWNeKmEEM/M3TWIIJvaK
hsUCdhbpngzj2fcBD3dgkZPUvzpEO9nRez3CF+vAQIgEbOfQgQ1TW/h/41K1n/dUOAYj08NLJZ/Q
5pIrAsu600MSVDCDwWvt5s2BnTIhrGE/SZBOcLRYNZ0xrFkt4rFK6SNVDpEI3Kmem/z7MwblFzBe
0lDIenKjRYSuZoDSMZDFLlmfZS3nrAfY1eTws0LrmZ+ArD5uCqzf1HCczCl+K0zRVm9+82rUwD2d
uIARPIHuoylOLjG8KuFpudlFiAMsgXjY43RQvLs0rXNfNX/wfWskGDtOt9sL0vsUMMFF/edRCfBc
+ZqO8T95XrCX9NGX8JJbJnlB4KvpR7QTxxZKNsjMaAWoH57PT/VgAu+DfNV6rt5e8DcQ9/pQSAoC
py8DcCWxdlbkb5C9h6ILWHlo4mclk6IUa3NZKpEWcTc5sKK1yF1uQdODipJXN1n4ydgh3Du065ao
2n+dTpDfLZdgKDUCBulUPLAgZCHaN+8rNPvwHotBTmIIyVqSU65gCQd6vQDoJ7tr1zl2sIZUoze3
7QWG+FpU0pNth9y/1gPYIUQfgptil680oV3zSWKh0rQwnVH2otzC8802dF8mgAiTtNBBiEPwxvU7
xuR0znemHHEwm4AcLiVvkUDsa+jfm5jQTUkuwAGA56/SGDrcjWiIGH3XRmfGZzXFlyn5paC8jH7/
GiJrWnotKQzEplmJXB4ofx0UgsMu2waEb1A4B6OyeeOtCjZMv6O6rgtmMVviB98ISR5iQuXTiW3n
0MGOqxGOjAErKnOWERyLa24+A8btUruWa/4Oz3qXHS/7F6EGtwWWlbc0GyCBInedrCtmmEU8WvoU
tVCIofg+QdSdHRvzf0YINg0p475B2xHTKB2QpBgRxa6zmoP+yMqt5uphmcnTnhs0vRAR0FpBphOH
0jXhvPuHfwXzy58FvfbnDkgXpMUIL7Y2p6weqf/9EOGqgdzcoAWGkKCse2wAQHg8dxt/nLtb8M6W
xPyry8uQEdsUV0S6ggIgWeKAtrA/NaRxsCiTJtHR0OACJkKhlImqsKBfMMvZRI0pTuLP6XRbxt+T
2dSPbnY/DFVSKzONym2Dfes3v//W3MzMZeptGuO5HiRKmmwGu4qPeCcQKDnG3m5gkv1S
`protect end_protected
