��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.hW��迏�\�U�A��t�a�!Q)?u��%��΄r:�Y_���9����5~���$u)���{d�Z�E���E9��M�B�T�f;��iU���wm�1�N�x�b2��L _)����x��MH�$�1'��)$�������.f� �P�3��C��4������}�T���3erj�9"�^F�������u�p��9I��ck�8������W�%�F�H�>gds���b���`��n��Ϝ
ո�s�L	2h-�&Bҧ;�h�g����Ml�ܓ�4A�ica_'z�i	����{�]�A8��b�U@��7�'_l]�d˵`5q���ة1��pL$�<DxhR�i?i��88����|�w����h�-aE�U`�Ks�z� �@�B�� �1�_qB�Y��5a�Y*����5~�iᯅgW�����G!���8��z�N�~Һ���Po��%��0b/S��C�P`9
z�MqQRSc;ܹ�c��=+��9'~�k��ʬ�@�Q�qR�T}L2�O`��	��E�B�
����cV�=�i�K�� �V����l,CdփҔ����o�K���7���Ew_� �aU��@�QLjt� ��ui7%f"�՜Q� �(���E���H`��t�k�VU,���{��v���EBW=�R�!�V���甆�t��)S:y�Qp�q����<
��2o����Zo��S�$�j�$�?�R@�%*������rEF�Jyqho߱�w8�QV��q�4�f�6x4,b����D�͓�7��%�m9��>�9U�� �v�OX�����#�@�M4��IU�X�� 4���%9�ʧVG��������γ�Q�7އ��4ն����{�����P��wƆ���������Fp�u�Etû���w�)=�9B8�{~3����j �+�Awu�� �5&�Z��ı���w*9��ٱ����o�׃`z��T$�-i�-U��kho�W������q/O*�
<��ց+���d���-E���0Ʉü��ۑ�2�u*�Ap>�����;	^� �*�n���������륡w��ɼ�W D�oNu��ﰯ���g�<H���<z ��5�	l�p�]���ZͻT�Z>ĭ@����6���q�����~�������K`��]���C��y�_Z5��4+��#���k`���L=T̎�	[���A45��}p��:�al�pdPV�[��BA
�e�*?�w2�*�&Ş��7)c�����B��3�Ӿ*�D��^�pD����w�<�t$�Y�����A+{{#��6"-2= '�E�}j�Lb�2j�(R���*>U�z�Z�B&޻���ę;i��0XZ������ZV�$V�2���n�� 98\�&TCq�N�_6t�EfD�6Vjw�d��\���U)�:��j�И��w}��#)M�V1��d10i��C]�kk�w빺�q� Wd�5�:���<t�YNXjU&�R��R\���w���ز� �����+�2�U��M���}p��˥K���8�;,�)�L� �/ږ����JڡJ�,�����8�uŗ��T��������2!���
�#�Q��PⷁE~��T��q�6reUh�Ծ��t�E8��-�4~Z��4S�K��Q� �z"Qyu�c�y�^��L2��?���h�Z��7����O��Rt
�]��uݷK���7�#7�����}�����k^z<��u��n!�I/G%�1��^�P�BŒ�wi{C��(�I�l?��$�aۯi�5���ֽM��W��Y�^4���Yn��:Z^��6�G��s4�}��ٗ�/�w(��-��- 7F�<X���\O��O�e�φ4B5Ӻc�]-~HN�=aFm����B�9�\L@�"�ż��Ϭr?�]�����1}4�Kİ���ldz��Ǧ�l�}}%�-Q������}�}�=n�����k��7�F�V��$�>]H�T<�t�z'u5��Np �.@��hY���]Æ��<4|��z�cv=�`��k��ҍ� A c
�xn��,l_�)��g�՘y�@I���G�1H�k)jk}T�tj�rX�� �j��y�)�_E�Z��z�}򝤼�(�Oj���vh���޳(��v�i�u��3���kƀ��&U��o%Y�?��6'jb�R,���dA6�x]��,g`�l���@���h�dOݭj$��9�׏�U����2�)�נ6��%�1��+�=���R��m3������Rb����/������~�I�lHA�m�ޒ��W�TH�ī9�T�1���L>�zƽz3�	Fj���@�΀�z�q,���,��"_��c�/W�����b���E�  Dx=55Z��`�q��#�8'ne��V9��Xې�����F ��n����2킼Q�ѹя�&B�GU�&��}��|�5����
���}���v�ɮ:��xp�Y_��L)Q%�8�e��-�B�j6/1�����y$iP��D��s��m��
�ˆ�jHbf|%����"���O��(�?]�����`*�T��r���O�t�� ^uG�;�=U{�
U$%��,ߒ�pƐ��1.]}y7��xְ����hhhaݔXi�Ҽ!w^ߞ�<q�p��^��fPsՙ<<
n����;GL���=oIT�ʖ|F�V�Ų	�%>����D *2׾��c�f���0G�\7��Iܓ�<�h���ϕJF�P9Z=����T�g�CZPk�e��Ǥ{����2��O��
%_ԝ�D39�tQU�}�M'����.p�SO@�Eh�'%�ˍ �t0ը3� ��ۍ}w�éa:x[�2��fyM��1@r���g�_�!�3_���1F�n�����G��<�g�� 6�:+���1(.��ND�s"qLjk�)b�%�ͩ_MTYΞTB�]��-��C����+r^��u����n�����O�xS�M!���,�y�P� 50lѪr���<�C�"qEY8�<1�a/?c{UCZ��~6�oK��_XH�*�����Þ��E���\L��@7��\��J\�C�-�rY�@�	z��i��L����A3&��<��I�1����\��NϠ ����������B�gm��am�T�"�EБpL֫#�w�`w�"T���OH��s�F�m�j�'�����i��E��ёS����H�DVkT�S��Za����%�_�+�����s��6��>*K�W�y9=@	�m��
P��v��X�F�k�*7Ί��Yf�p�}�)����Z�$�S�'@7-�v�V�UI،��0ὅ�ꌋ1�^bT,��=ݥ�Cf��̻H�h����@�q�'_ɻ[�̺Vl���䔟]�6uD\���X�t�<��1l��n ���uE-S������L�A-��/ðhB%�׵~n��P�����,(�S-ֆ,@R�3T�{��{y���Fp�L�c��-,R�n���8+�w�V��gכ�{�����wwXP��]��fF%&rk>�Ń/]D�ф��9�"z4`O��^���-�ȉ�ަ!r��,#���T���@�����;c�p���冩j�sy��'�JJ
��V� gb��T���j[������KD�Ri��se���zu�Շ��G��MF�A��k����I��f�B~����?�nq�Jzs*v[P��&�**�����voIf�?0�ݎ�qR���1�0rޑ=��s�o��+^k�O�\�#�A*n�7@������kY�X)F�$�2��>�i�v!�8�����4Γ�FX�W�@o�0��*T@���;�F��̃�'%�7��������l�<µפ~�v��̃˽n�Qt`�L������W�wM�?6��oB!(���F)c�Ȣ���I�%�ej���N0R`=�[a@�Nzt,PĒo��o��D�<"��&h�y��M$�焊�tb����W����6�rT��D�������xh�OE*oNx�N��M�C�*7�Ѡ�)����P��e&0E�bڝ-T�Z�ꢧ����j�'�c����o&)r�ڢ3a	�m���L�VF���2gó
D�u���߿��L�UdH�v�V
H'� ��7�*��т��U�[6��u���\8/4��c�b���ٺ��GDS� y6J,���S� !j�;���9�-
�"X۳-�� ����qG�h�k�kO�_u�0�K�o�����)6�O��'z���:�y�F���o0��B��y������(3ձ���J��+�P�����h����R���,'��	��#9�u�<skE(�=wW��&&:�$�XJ�� <Zݏ���Ev�V�i�k�zhT�o��{�n}-�ĢɬpiJl��|%�V��/TM,?���
U{��Ś󓂳������VzqdȾoO/M]}ͨy`����O=�&��?����?�υ|����=�N��Z�\V��1��<~4��'�m2����
sǛ����p�T����.��`Wr^Ȩ
��AbJ�} R�Z�f�t�$zi]�V�kW�=g�4lWiT���������t��.����&� n����1/[+��g����p�{u�g", �zb��nƼ���<���t#4UY����#G/��ڐ�0�7^+���T2�_T3��� �
9)��q�$�%ػ���c+Nv�x1��,��J�y(��M�����+u+�l@�^j�f����yᙎ��d!?�J�jNGJ�f�ʣ�l�9"1�W5��c�tw�^s@�F�p��	 v~a84�tDW߫NA�}�Zf��ܑi����م/����?
i0�P�^��6�*��yS�;DL���v1b����;0ϊ�;��1��^�h����Ē0�"=?�I��S4k���63�H�a�}�:~�er��c#�ʻxr7IN�`2f�)���B�_�ׇ�=���-��Y���eMK��7	>:�������K������ؾL�a�� ЮTb����!}��L�<Ċ'v�a���4�#9�a�?�J}�s΂C'�<s��[i�����X��r5�Ml�ʌ?iN�9�O�y��[���M!Ǉz{?�M]���6�0ܖ��|�����y����Г:�AhOo-������A��l�.��*��@�lI�o]�P�,�bd֯��WOܠz<�z�5�	�NkF	3���m8���?����u�ltW|�>�W)���)|���lZ` m�w��j3+ �s��"0O�s;��)	��a$ef��A�r=�g��h��I����2XO����:��'͕i����v�B�<?��)V�zS�ٶ�,�yf1��4@����i���9�HH����0���0��`�%�c]�����H����w]K�˲�q��B�90�9���9S\�ހ���_a�ʙ�>��Qu�&��M�dR������K�R޹U��8{�F=������?��v�`wl����a�M��!����蝶�U���^��絨ȼ6�!$���lgT����"
�.5cf,v��l)�zE��9s��o��C��p%%SbJ�(������6ÓIs�]��b�߭�7�<�r��|�����<�m=��8%�"T9)/�K{V~��	��FS�2��L/�Q�(�:x. sЫp��}���N+^�",:Z�F�CME]�!��VW߯D��߳#G8��mq�in���V5�Vt*���gM�6���g�ÓQ��?Nݏ8�����3���:@<��x��F�i�!� ��/����wU�lЄ��� s�/�="4�@��	���JW5�i��n+�"�	�.l~Ԕ��A�����ir�yܚ���}�� ��/e��6�ȏ���MDq�M�=�{Ƒ�G� &x�k�-�����76Ƽ�I�9iz�LBkQ�}h�y��q�����j���c��3�����t)ٙ��D��?b<>&s[�g�W^�B$���za�D$��R�$ALo��:sQ�T�t4f��a���!�qx�|^�!������Ny�����N$�Z����ín����0�|����ڢ�ċ�T��!XM��繒y?֑�t71��zc6����u�' �b��Ƨ��t9h��K2$��_A�ܯNX�5��7�NM��Ö�7�����-&��t���n��|��GR"b0#�����cӽ�j��m��4/����H�#?��&����G�	���u��� P�8���J�4���
���-��#:HQ�Y���P��ǝ�^���#ʭ��+L����%�Z��T_,���ҎS.������͉���yU|�{!�3 ��W'�s�ˍ��O�'�n�7u�|>䱸�hҨ�ѱ5����s0�EŽ[K���ʟ�_��.0����g|*{�Q���\��l���\,N��B�!o���ч`��iZt��^����ԭ�)P����d7�<��F���_t��h�6J����X��Հ��ϟ�e:��>�hR��-@��T�И�WQ>���[n��X|��k��"2/��:\;'�V>��O�J�f}=m����/j�R�WLw�N����+p�r��
�S�|���şO���5�[��?Ȓv'U����L���~�-���h�P�iAi$+���'k`�d9��̋�%�O��
�y�M~'����h����ǐ��zȽI+�}��$����,�2��s7n�icsA�����*�o�S.�oS�Z�,f�o4x����O��h�q:6���QOu��>;�wE�lZp�����o�:���������x�wj��Q`�2�4� u����܊�1��_��3H�FE��_�<Z����'���H����e�����5H�j)�|�:G��k�l��+�V�<�{������M�ߊSϡ\�y�Eǵ�$�f�߭��LKa�9���KM:�v�1�U�L��������ݲ�-Q&|	�F��¹�-	Hb�r��t�T1�䭔�T�C�y~<)�L�	�G����f���Hb�Gc�0�ON"����?� V��>K�(�5-�ČS�}m��BZ� jM���d`�:��p����]��������D���g�H��%1�΅�fh�Hto�T;>d1���E���?`�i+��R����T�^���0�{K�?��1uE�1����'�J�y��,_J�������DT������򗽸�i� 
� G�"�\�z[	ݗȏ�ݖ#Y�땢�|�MRBLx9bf�vе����⾝���ف9�����f��h���A�j�vEݩ�� >�� |�1A���ͷ��!as��ߍ�C3�C�Ƶ<c���n�]��uṲ���*}�̹�ك��MÓ[�L�険��=v�ߒH�k��&g��z�muA���/��Q\�(��ҬG���s�-�k]d�3>��i�|]s�	.Y�!��U��l�ȏ���"�u�G_ި	�79&�M�lqTC6"��Ō���I���L��wPW����-�}hU7�VX�(�������n��3���v[h����ҩ��o.c4��O�Qo�q<p�?�dsə
Z6%4b��ܢ^�{����qb0SB�v���3֏�h��ђ�>P>/)vg��B������s��~؏�n��)�Vu� �\+`����yԮ6�
�"�Q���2eAWb�*>�~���6XsdM�1<h�^�����2߃����?���y�����Y�!����oD��PB�/t��]T�!�d���!A׉�O ":�лUR��'F��K�:ض6ɾ
�����W+��%n�{s��� [���Y��#�-ѿ��� l��y�T2� S���ֆ���I����m���o?�穌s�T85�k��6�!�O�NPT$KlD �1�m�+�q]Ǎ����o!Y6������TOQ�2����ߒ~)@�=K��#���P�K��ଞ���ŭ�|#���&e�P��������������m����J� ����
2M�xOf-�l�N �2e�6J�U�+s��W8�"r����q/u��
!s6X��"mh�Ea��K���a����e\;D�����Ps���Y�����,���/ٜ�5Y��Q�Sj�qH�u�P���wOq�6�����D����v���j�e"�y���MQ�#J�Q�v�D^�fVF�X_�t[��b��ŝۀa�`�Șd(_����{]J���a�ig�����t��_�?�� �#q�:�SϘ*��q����Ռ�Sl` n��e�;]= 1?��ח�7`Wb��vN��db��@O+��tǺo!���"��;Hx��M��,���E�7դ�>�Z�������b+��}���{�SPjl�����81�UA�]����\W_5�:{x|�� >��q��J��*B!�u.rD���,#��L/��N5	��wr�����mE.b � 	߸6�=�$q�
D0cT�_�A���[^@�[�E������I1��AYQ�D94Tt�^���,�kZ^+{��+]P�m���2�2l��a�*��Ѵ߹��>(û��������/FLZ��|l����j��H�eo���WY9ޚ��F7��U4�&p�ˁ��o���>E��~q����;�X��@{p�̾$(� �����.J=zm5P%ha��9�2���@2�{Hl�C�ħr��wZ�4�֤
�6�y���^����x0��q!?+<ǟA�Zy�����h�������} �dR��`D�Lޘq%���/����Ij�+���ȩ*��~�&z��oz�������?��X2�ma�j���q�	>�2[$ �'3�$we74o!���M��%%yS��"�H]k�J��u�GnZ
���:AȆ�-��7G37c#AM��C�2{��:�}��#��i�恠h��.�T�p.����YX�=�D�=T���K�hm�@�*åa�ZR� �t��`��0@��t}3-�`gf	>y"ԣ�&�W��|6�V_v�iIdq�?Jȹ�Lhv2;�\�|5PP~ohQ�5��<��Y6�y��M��FF��[O�g��{F.�0ۈ�m�L�n���i�i�S����Nq4Ó �0k�TK>���7��}�[�P��e{�.L��怃r�ȯ����5%�-�禂���׬��E֮~U��N��n+ښ�J�i��W�1ޞ[H�e,p扳�1x	A�0 (B$[*8�2OVy��C�|P��D�����RW�:(g[�7���6;ĩ�^����5��دo%��Q�0�>���cZ���.#=ZI�����.n� Z��a��t�sB�.#J����	�Y#�"�<���n^m"���v�5�R%z��Lg�B�N����hZDR|Y����]q��"���Iu���' +�e��H�����#�tW�נ��C�S��"�V�?t�E+b�=W�Y}co�`��)��/��M�[�>i�lz�e6���@����?qa�-�� )��?l�O�i���a���X?31�T�O����l�O��QV[�����^�f3!�A����9�6�dUJ��A��)l��C,\�Id����Noٌpwo���)��AYe�1͑Q������!1EM���v�].��XP�~��휯��q'�5�O��HՄ��"�>d���������hx�'ɖ@:2|��n�W1Gğ���!�\���^,��d۱�b�+�YP)a|�I^x�ь�j��c�+���HݱБx
^�"J�C���8��XUG��łs'���7�H�_��j_��4p3�4j*�_?�����ύ�0G�)V�'��̬�I>֯��[�g3X�r���A�F��3��d5�|Jq�|�����QO�����c�Dhi����򡎏�(�� |���$�=�py��Ggb�=��:!��&=�kK*�뗆9jn�½�"F��Ԁ�@`�'��%wY�X�%T��R�_\�b�?v%�5���ͤaĩ@ �{���1·dBi���u�D���u�K��H@q�S�~��$y�1�Hg`���t���j���%_��˄jղB\��1#�d�[؟ ��'�~�T�s��f_Y<O۔lZ����a ��ꬓ�N1�w�x�U�GTFP���RPb�q{�nΉ�T�)���gU�|��s�N�k��nA��\:���T遃W��Z���6�ْ��T�ʢJ a~L��M5&��X��1e;P_7Lz��F�C���?3)O�; A�m�&&�?�W��m��=��0��<��'��B�}�-�����7�Jy5X��p]Ý��k,�k�_��K��9�T�i��[��E�pb�]s>�z^U��$@[��D���r��ǀ#imX�,P"�����Ѡ��WK��2i�d�7�e� �\̾y�Y5�1�*d .:�6�p�t��|bv�Y��J�oQ8��ΎPc���E������b���ޕ�,�V����l�-OL[@�!g�����9�fƀF�U.��c����E����k����S�`�RNR�C��~SR����D�����).��W�3'��<�YM��7��$.6��A'���='�|z��� ���:D�24�=a7�p~��D�X�)x��n�[�)��c���/��g؆\ȳ��S�����,�^�v.�s.�%���_���H>��k���㮛|ܸX�`)aٯk�F�7����Ĉ��c�q��]�B<S��`oM#Ń�,�:.�c���"��n�ֶRs�!��ŅcW?>��~Oor��
Y��΋�fJ���!5v��d@h�7���+����P�d�b�y^�7�.�8���s�e��'=2�$�7g�lC�W]~>�E邮bF_b �R>�P�|+���@��`�8���l��k�?MMo�҂8�l.x�?֣����8{J%;M4�g�(���!�9�>1db��"��_-�k`���1[��1�j���g��Vzo�iZ�,���� �X�=��)���iV�c���c�)!�;3�Q8w�T�#���]a,�e�r��pR�`!I���Lw:�[\p9��"o����,q#�蚖�Q��<Ԩ|��*��[��=�Fj��-�V��ݏ��<^	���L��0T�ts�D�A:]k��H�v�kA̩3G�ym5�� b�!�7�O�p���T�>�d$�e��uh��k�$͠!�XWpκ�eKh�oWՊ��#�S�
+r���r�d�&h���+v�PO�Ż�뢰0�w	��</L��"ʀ�n;iZ����Z���O0�fY�~A��Y�Q��Ow�aL0�(vp���)�e���y�c^����%J!���8�a�R���8vpw��ݶ�MRU� �K[���r4�6 ,5��m�C��s��)�Hn+�I�U�)l��'�"�;����T����8a4W����v|�@�ӯ�g�/,X�M���s��$�c2D�m���Z�yg��b5/9�
�8HWk�(R��}!i�q����\��]&\����
�2-�͘��2��'._�B�h���{�