��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��Q��`3G�tv��-��ފy�|��5�H�8X	�c�ZlO:[�Y�~L�!��7��Qh!�_���2X95h� �8��z������}�Y��Q� 쫤�Ili�7�	e�p���dв��|�F?�2zə8�U�I�ŷ��Gs��	�(O��'e���??������]ml���A[�Q�c�\3�'B3d�&�����.��AR,��`������|�L�|��Ҳi��jr0�$}��MR?ɒ$���Z�YC�
oa�����U���g,+F����K�y|�]���V�>
S#8bK�ns>�?G���з��8R�7�����Gx����]F
z/��� �4zq�tW���X] ��r&���:�}�,n�<I�(q����y��u�Y�D��qKp*���wx�N�H(qɄ��(l����w%�)��5��Ԃ�f���v8�x����y��j�����S�_�C`W��&
��N[��/��E����ɩ�K��r8���/��h��'t�(���
��Bj$7ۈ��ni%�$f��}�#��oz�F�Zԏ��%�D����a�B�q�������� ���<�]�I&�ň�+N{ -�s���*8��gD�� /\R��\B� Ėl��Gʗ��piM����I2�e�P���n��=�oj�q�D�>��^ K��Iڜ\�
�,�2��ݚ�ӿ_����ם�b��DOĉ0AYD�ujn�#ّ����@/Q".�O��Hˮ�o*n&S��$x�>��G'/���,3�����೑[l�k�5LM�C�����\q����$'�`)�H`�3�%��o{p�8�.Q8�ÅR��?��A�}��w�X�&�	�q{Y�}/{���[:a����0��6d�h(q�?��&�\֑:���<UrG,*.�9/�
�o�xw�tb��'4'R�?j)��,��o9l�"�,��kr��_�k��.��^ع{�jxH��&���+'
�k���_�M�-Ԓޅ�����Θh��:$^��o�",��49X\F?t�3��G]�7U�6��ڗ��:�6Ѓ�y���?�k|����Ѭ_��|�͌GV,w\��{�j���Dÿ����ZL
������h�wD&YB�/H�F��v�������|`>����O{>~�2	`_�~X�w���վVt����*כJ�U�ـ���V�i��H�~zB�3B���t�O�Qw�o+�Fig�� �{��=Am�g�g���<U+v�Y�����+����|��H�/{�i�h7I]ԍr�u��"�M�Fo*�B�����W��	���٦b��Y�t��s��'�E��3B[�Ey�Pߣ��N��#�'�Y(N7TS�MS���.h�8)�OP���d��aL�hl��ќ)�$�:!� ��Ì�Ke�i皾��rsk)�օ���V���gM|xuF��(c�3�k_��Y�+����3�s��0{��@�g�K�8�sOCv23�}������h�'R�0Mk�T�E;�r>���w^!"�e�r�S������g�.c��r��ViK���G��Vd0�P���S]�<՜�z8\�\%��oּ��<A���{�'�E@��V�t���Bj3��~�_⚬s�ԧ�I���)фuK�/i������5��VU_�|g�#I��t���1�w(|�8����6Q}$!L�l}��#27o�®�=2r�c�;׍�����
����>�ۺK������+�>�[%�9�[��J��E����ڣ�.�ʙ����HK���E�^A3��j�-uq�v��_b0�i/MBBJ�������Iܱy_�N�sQ��D��BA�굫"WӚ���������%�fb���_�O���f�K�^��"M�������4�J����.�#|t��[U$&o�\q.Y4e�P�ǃ[���sz��˷"�	7�j:2�*�5��{h]��0�Dؖ�4����$�$��K �<��Jg��WqΨ��N�B��;�3�7U�T�pp�K.���P=�CPo�{�Ï>O���Z(���~͔��8�e&���f8�vqK�pW�V[);^�6"��*��gfy�\  ����@q�y��`�	Y��.^{�=�9�k͛9�m���B=:�*�ƻ�������_O�2�z���~���r���G����%��X^Y���`�c��aw������C�?ANdĠ��=ޠM�q�� �������1�^�g��(O�S�VM͉�)e��\�o���@j�lp������~F" -��Ʌ��E�!^f��B�W�΁�`��φ�B��/\�J�ԆR�j�#�Φ5i/k�"�1o��9q�;YH��NrD��Wߞ)ll&{l�����~�8d�DH@������o8_� 4��?��E���`��S+���s��[E�Y�ٛ����Z���o̫��4�_'eYx{�4��^��Ĕj�[~��v�v`{$�MJ����!�VU�)��ED��+�� �q�)��B��%�OB���4��I!W�r=�؇d�B�:w����H��	���_��K�YK����c<��&6J��W�i���\��8f���!S��,�*,� ��Ɩ�ߧ#4��̲�}N����� �1M��!/���a��{ʊ1b6�mۜ��ev��`t�y��G�ʹ�~P=\�W������}��^����sq�,4k��xCޔ~�[1.�Cd_���m$o�~�ί=��ߨ�Ŧ?t�fQ��X�N��q |$,�@��Gօ�m%��/ ��:�t�@�{P���T���i���r�;�o���y��2uO �;!��iZ��:��`9�D�)da��@����C\04n�(0M;���c��2W�vL
�>5��e��Xp�;��t9D����1.��U��X����2��g��% %��2�?b��]I�͋����8;�vy��~Z[�{�Mgl��������/�7��F��n:��P&��19��}i��ʂ6�Y��q���'s�jf���H�9�(��`������Ty�;VY�x�%6"�g~>�&/�a[��s���)��%^�D(���o3�ҔH�k1~�^�ۆ��}��B^�a�u�]LUa� J|2���8m�����|�
�?ѯ4��ƛIF$�#�9�z�u�m��)�7�ߟ1@�����jN/�?4 ����, ���`����h�^�-<�k�a^"~O���w;�0��g�~_��K��LW�-Nޅu��9���v�"'���|f���E]O�U�� ��<��Y?bV~#l;X~p��Fo0��e?Pd �[��Y���{�pq���䆈d�xKl`$pL/t��-W�觌O,�Ft�~xX)�w����j�t],�S������y@�В�ܨ��vk��y�Dd��3�/���%�F́5�qް���|�y�Ut@`��I<֗��˳h�K���=�[$�g'?�Z�#$��G��(W��ã����KD�R��ܸ�%?S��,�r}��g����W'�J�^��w���{�ʳ���^�ﰤ�$����&2� g|j�O+��Vb#��a I.�Q�p;����iP�d#-j�e���E\pZ������\��8��y�;��>���<�l�i����(���6�P-��Y�y�u� 'R�\��������J����<"jj���[���أ�3�|�KMGI.�f���5sP�Mh�eN {����g'��@�r_. g�G𘃋�S�1S��;$�ފ\w"&�����m�i��,5����1��
Q��6��e�DL���ø\.1|sA�qfn��%V��f9H�i��Ұ��)��6X���SM�����W�:�\Q�(R7v�/��yJp8Z��[V�>.`u
_�c@���_⌭�B�Eʈ�`ɨ,�4�b+|�sׂ�Tqs?�i�p�9q�?Y�|͢�6���{z���4�%���07;�Pص�F>I(F�z� �F,HGJ�E40�Z)3To�v�ajo�XQ
�Re�\��'�h�z�4�Ř��nĜcG�9j�Ka��Y�5���N�pĦֺ�T��Ҹ�O�3��=^��^l��^�h���ԯ�R�L%K��Z�O��9�NY{&�.�3�A��j�p\q�_�y��c��yIs'�����[@ �hhp�껜�-�1�+9���~P� "O�ߚ�+�5�'J���aQ!�.�3_�0��p �kI�}�aI�t���$mA\��;h�(0���Kx�d�9�t9�y�,�@(yW�Α!�O攳�Z $���}U�KYz�)(M�Un��R.��{ƥ������e���<�Րv X���4P��S��v��۰�w����3!~x�Z���?�sȆ!��q$w?⹷�c��YES_��kO�����^C���+0+ҤǤ-�M��*auFU�?�����VXj.��{�賓��R�u��iǍ���-�h�<=K�p���n�v\=���R_�>U��C�;��'�X�y������^!~8c
��#���~`�d��L�mZ�K�e��eu�-��j��Rj#��|?9%�x%�@�[-� �Qz8t�"w�)}d��b�l������j�| � �g��~�oڐ����ͩj���'cdnK�̆ع��E�b|�ۣ�%7�5Y�v�a"76щo�[UE�J�<6�5�!,��d�D��4���i�����sȖ��L�^A��\�;R"��u��f����.�rH[D���������l⁅�&-.7Z��H�涜[�5n��<�e�bF᧘b������AvMji��N�W� ���K�F��F5*�]�=�mH^�vj�H�y8)b��~�`�t��߭����l��.����z������dI�*��C�Y�@�2���F^�Eh�9��:�i�AX@:8���ꂱ�jpr�"�#��Oa�,(�>$1�!R��g�)Cq0�3��9f	��C	:b�q���צ����B'9��E�lw�����΀m��P[Pf=!��h��Z�|Dc'��$��U�-g�L��41�2�b2�P?����X�G��p��I���gjO���q�z^��ȞS�@eqH��{�_�[x~W`��_o*D>�_�%8�90R1\��������ڧg5�_�89+�ٌ^)*e�7�� �L� 
��<�q����: B���}��d�	����� �H���r��O�����ݞ��W	�sH��9�n�8��O��^���,��� ��!���8W��H��tH[����""�O&R;����j�!U.���%��Z3w�}짾�Ve�z���cʞ��>_F��>,"BT*A�D���b�m*��8���B��� �׀͐�S��V����j�^��=�;;Ǘ@=���%[Z����3=?Q_7������l���NW�}�M	�f@��5��5q�Oԁ�{3������9W����(S��~���H�n�ŝ]ȄW�N�|F�g%����q��QY���Ӭ�O2� �ДE����� gy�|�(�����k�C�1=��`Mx~%^fڞ�Z��b�9�X�`�(2�j_���~g0O3���	s�ݖRIgO^86�,�k���� ��G���kU�W'?E�#��ʊ�a���bJ�@�Y��cߤ5X-6�K��?�
8��S&�4�}�I���h����`�,:0<h���j4q�R����$o�.ս�<����ൌFR�!�������N	����3g�E��נ�+
��Q�_ L����
�Ů�1�G��6^�b��B��e]
��3� �\'T�x�ѳ�2f�o8�OE�{a_\��h��%z[��/2��v� ����0�Nc�w��d��ڤ�Z$Z�WHG����Z��� ���2���8���ufk��LM���ڗn�`k���:*��gvL\:��\۠�B��qw,w	��Wm@@����z�Zu���L�D���pr��纀�sGL�[�*����3�E\�а9�6+0�������5#�m;0�䲴_��2il�%�Q������Ex���x"bey͌T[I�E��%�Tۄ��?�ws���E�P{Ӧ���b��ͣ0�WŏA�Q��n�XM�.�r,R�=���?�A/��U��<{?5��*@^(��V����',;��H��e����;�L�ɣ���E֋}�Q�WZ
�������evl��,1}�^cEdf� y��uY������b��r������@�lj��,�.�
�b��cf�ͣ��!9�z�c'S���-�P�.>��E�XGh80S��A6V�$��{똳'5<�d�P2��*;�ɰ�kp �n��)�mמ�-c�U V��֜���=9�j*����Ƽ�S���]l�Z�2S�q�o�&�k�E�yM�a�*����N��~��<!:�V6�<�'$
RĂt�Rs�~⯝������Ntl7W�]�H��[����؃p:�
I+$��E�����|y�I�獳�x�ڄ2�^��u�t�Ǥ�ٙ���o�����V!;�$/p�L��tf;���\�GޝD�\Ri�j�Y�&�ⓙ��J,�Z��~sN^��׮���T���xVԉ���I��wD��$K紋2�h5���PRB�43C��Nؚ��=���p��z�����������+A���,H��Ո������>��|g��X�fI^�b����*\�O��vm���tʆz�z�����xO�UN�B u����B��:HOΤ/�Uv�_shp6f��R�̠����Y���(Z���(Z��k�� �.��o��^_�BZ�9/[��k�W`�,�~>]�e�W���3ֱ� �]��|@o�E�y�0�2�˸�R̕a�ǣ���� ��&��&��?�"AS�6�M�� �	���d�����9#�\���� P̟^B�G���L2�]9o�0�Y]d���P�Mc�� ���[�u��z�|%�A�i�P�旄�!A����iE�ɯ*x�������}2��m~���+�y\�\]'}[�mF���%_1.�s�k�O��+�F1۩j��s��H�1e�8���?g�S��i��ǍV\!���R���̓����̃p^+�8M3�J0k��7�#����Ơdӈ9y83���k����ʋ&cw������U#sR�\v�@Ch���'�H��m���v�P�tKj�������@���tX�����*��x�&]5�)Yp�<d>��o���7z'ȼw�J����[9{������q�Xf$�T:3�ˤ����샱y��K��t���6t&_K�X�R+�کF�H��F%h��*���A��?F���Kox�� *����_�|Ǐ4�m�a���� �cb"�`m�g�|S�p}S��-�[�Vp�קyO
L�[���wm���;'��y}��c�Ĵr~��^o���/�F�b����G߉0��V�<����^[~���⢶C��c�0�c�ӭ�L�W��F�J��?!��.�H�ǔ�i�F��L��=�ӴϾ��@<&J��c��>�R�!�=�+#3��p���&U�\����ع��`���\��/�`&�(�w�shb��:�*YPMb~ـj�8���
�
VG��h7�J�0�+J,j����Н+��ǹ-�Ѯr7="my�����`:�W��8�{>3�C��s�m�*��+Id.�5�МV�*���BC���?_�_���ЂQ�����CA9m�����.��c��i`*�8��1U��nZ��Akj�jet[؉ȱ�ͺ�pT �u�m�
d���$�9ؠ�fQ=���*K�[�ʟ�Υ�rf����Ω�Ϟ�� _6i����e|�8 $R<��hzg�Ʈr��4�ޖ��|+M3;�jvGփ>7��Зc�[�rj�ì�}�8W��V�����E,.r��69�ͻ�6:�f��I?\���S�����R+���G��EP��5==�raZ9������R�u@Gi�?�\��F������`r[�l��0"���Β����[�N;���׵���m�-3nD1����3R����f/�f���p�q�B@�-�/��R�6̞C>�h�G܎���pN�� �>��@!fXҍ��MYsB�J��7��)L�(,A�ՠ	��	AJ�:&{IA��ʟk���>��`�㞡�q��8�hP伀۾&QT�wе�۳����.bǋ{���v�P��4�CN�d�}�f���A��c:,T�p���O�;c�P�C�Hg�@��A��Z� 2�#��X�QELY�;��Ae�=-��X��j��q;n6��06 t�0��?A��/�r"(�f��D�Q����bS\��vSQK3/f��3����e)\�;EV;�q�ثpzr�����%Z��;L��"��)�W���C��q�)�	{S��'�@��UMf)�_f�����i��L3J@o]	;J�Q�K�j�d��]��$����5��ٖT񁹋��2�Ћ�k{�����L 9{�Qb�3���bS�əQ�K���S�EL#�~�l*�`�9*3��W�Ԧ���m�o@�p��[���[�!�wj_¿3� ���p	*<��fȈe�H���u�#޼*׺�A��'&�J�ye����N-+�lL��� `ݨc�nP��:�qC�<����B�A*�3�4�#7��S'h�~�y�V�	�����C9>�^c��1�-�5Ϭvp桄�G��F}X�Z�E�����"77���
u��XebN�q2��Di^��}7bD[�Q��o��$ ����ѓ�����M&AQ`4n��J�x��C"��: �2�D����b�5K����|�u�h���s2�G�Mb�O�k�"�%?7-g�/�.�z 3 �8ҮifJx]yA�	�h�$�� 
�4�[�ݰI7�]HV�&�1� �D�5V6�����K�߄&���T���ɖ���@K�ar��+y�.����\yR͖��q�xo��i���HHun3dٵ�K�w+���(y�O�-UԆ����M[�U���v�Cƻ@D�?�F�v/ěU�-r�s3~�_��}�ѣ�Ʀ�Q�k�C#ѿ�P�\��Qg�)�)�pg����%D�:��ݾ����/�������&!k~�	��<��eI%��nh�J��Ma��zo�ہJ��P�jDXED�*�˟���بƱ���.�<d5W�1���Px�UYM!��H��T�j!����-�y���������`V0,.f�uM�ˍ�6��}a��aq ���y��+���n�)��p���J|F��yC�}B�V�p)G� ����� ?&v��[�+�p6w똚��L�0�gL��si�Z�c��ܮ@>n��ci����_�_@�����X$�(j��D�	�)�N۵�i�e�7ظ��@[XG�R���g|~أ��-&"GB' �,:9*qZ�ߍ���,7d�����o��Š4ƛ�3_�DY����|�A�p�{j[W!�%��ۣka���c�0�Z p;��a�f-�����C����kca8!��˦�b�C�A�u�5��a���U��	x�ǋ�0��K*��ٓ�2n>!�Z�R�����~�I�I�6��ˈ@���2�^�ꛬ�RX=��@/;S6KHl�n�A�Hgn���6J#u۲�,2�����o����ـ�o�b�v9��No�R�������]��#�gR����A�]�m�����]���H_|n'0H"r+�&R؟��>]G�4��{]�����"c�zQ�,ZD0/�#����������ap��ɭ�e'���ǝ��r�+��j�����
�(v�1�-a螠2n34͸���`K=&|���x��ɖ?��Њ��!o"���HÃ)���rƿ�4�y���e�i�|P.a��3���XrR}k�V+4���b㐣���<~y��ݟ�eJ��؎~�����X�"ƛ�,a�( H���?��4�V~�u�(��"����~/ϹWŊ����/c�6ʠ�7�K�p��$EU��;�r�3L-��K�~�����V�3�(*�������{�g��$H�1=/޺j��I�� ���X ���#Nw��Ex����(U�>q��23K����3�{���8o&��?/C��R����}�`�>Q4�B����2��L��sB��@����9zń~�m��ݜ�z�p��4�ޛ5	:�J8�a#V���mМ����lI֏�A�K���8�A*R�2m1���X�:�iv�З� ��M�	Ҫ��	�~v���+4b�|J_�z�.#xQWOل￠���¾�XzSO�ı�Y�j ���.��ӯl������e4���Y,�?v�V��V,�6xig����m���d.r�ZU�� ģ|H�������M]Fh��=A�>��)�]m�_0����)��j�zV��dԚr��ɉ��T�=Xz�ED��Pu���r���݇v鎨�`��R���ԥ�p�XoAq���N:�ϑ��{��mPǽ�"��y�6B�ۓ�2�X���w�B�--��z�<����\�J%����6�N�%��!l]�>j�C�J[�p0V@2<D�&� ���c�L5����EI"�〖���o+��bv��$TN�C�����vB*����K��������������L��Ʈ+�&�}d��=�VL���=�ry��G3�����0�*���$��f�8~v�8�U���k���h��K����c�ҡ���3?�o�<�{�����n��wB���O�D�o�5P,�57̐fܛ���)tM��v��RT�����X�č}�����&��7:٧�ic�U��������)P�f��y1�/a(@.u��{�:V9��Y�@�W�)�L?�~���F ��{9�<��42����Wړ_,G��|���m�l��
3�*�7�4&*E�/���mӂX���{#P�W8H�.�A�(��F��7m���^\7�g;�iZc�����H��%w,��bʙ-�w��]9�Ժ�k�mV@��.�+O�Y3	?����6�C�#�8�;.w��ԅ[n����'5D�56@Z�{"s�!������Ü�n�绑tD.pR\d��"�;6Ԕ�r�Q�@��8��+�e� ި��Q�w0hR����it�`"�
�Ȱ{h\y1��wb�ܹ��.��a��~`&Е�2H��b���⃒�dm���|�"��-�Ɨc+�*�C�*�:�O�Hҕ�p�<K۝�(漚E0�k`M#��������F�����Θ/�{C����w͐o	���h�0���0'0k���*�d�;�4�U~F�<�Ci�Ʀ'�pv1�`}�G�W��s= .S���o�g�S��� ��yM��WwW����sv�-�h-3ZDy�=�ֲYG��C��O�#v�kg�7x߾�P�ET!E�À�fP..SD���d$��u���o��b42=�~�x�c�@'?܋	��2���A�C@Ff�]2���r����;Y�.��mr�M>M8HO�E]#����FX�̓O�C��8�.C�W`���=-[�
QY��΃+�9/sv��N2�"d��mm9�� td��0O2M��[*����;��x�ը���2�q��<�M��)��t�'�&�^ǻ�o5��v��a���-$��v+� y����5�
B�X=�+}`�_�]=x�y�/B���$�VB�m8%�g��؈l��  	d�j^cUyś)	������ _�s`�)%�{�u�n���f�krx�����{��q�i]� BzڟG��JR��v��2E&-�- ���Y�L���K`����/�IƝH��D�/��}�7?	:�4ݣ>�Iŗg-GWt@�=�