-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1PJBWS60mPOej7yp3hzneRoRHM5XFJUzTAhPtoaaIEeKrKB0YJh5p58XhAOCPHdilQYE7BzTjmBb
Lb4BXdrlvtYUaqnf5QChZymnwbF2DhFbcd76daVYmXidyOybO9sv7BAxoKI7JCmk0BTNINwY5Nhr
4tgZCIAYGOp+9dH/DYaeCEDOIkHnvARlUaC/kV9tdhNkrFaEsM7Qf0Mg1YjtLcIcPI/v+o3zFKVW
2dhk46sJFpTXiO+jA/W4OzSmuFwceSlrRSjbp2jyfgOveRHAfc/dqeVv/lznXkXOXhGyuN3knZz4
Ay89iI/HvbPxPkPAkskWhnebXbmYdz7vi4Rhjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
TF/ukevaYt7PadgP5/mUZioJb5q2a6d8jbVeVL7ncaNWpJyNXqkB12gLMU9nNnRGU/1NyCv0CGWX
CPsqfKmOT6lHrpJGLCDZIcU0uiGve1CKROkbpNanqtD5gS5u3KmAdevHLqV6g+B8HTkBJ/MeGNpO
1/36wm9Mr+71h0x4/sGrP7YcoCvaz7N6ro1k9XaYzCUtP/SbyCRnZ5BPMxJhxoWaskqB3n/7JnQB
T0SpU9pqplaIXlrlT8MaH5YrWMODyPnTn9mS1EiH9MTMHl47fpgEV/tpHmtF/5jBmiuY06ayo0fg
2uQRGntXaBDw3Y7zPHWFy+aN4FPqBWb6d1OZ817vhxaz0pw7HrOBPxUGnGlwLavRExhUXrXO2x0L
0mDRVSpWiajH7zeCbYiSPcTpHxC0cw7JlRTGT2KZDX4JSTwsUE5swwF9Wgwcgqcze54jl4eyt2nh
qj/0LI4Q9teBnQwEHe+aYRQhhIeg+gosJq3l4+HNeZ6hsbSa/Xupdx+Og7x2Gzw50WLqhNPYDtr2
zwQ8N5F8P81GBHRpZvvfe93CuCsjLdQSUv+dPUvGgrWh8jjUZwlXBHGfq0mJGAJkaEm0030yGGnK
PM62ETdG11skTzSW8ayHQQ2m3f0reuovS9OCmVoQeIxBF1nwSfk2P4QVcj7o0fqN6FxHz18Ch7TP
+20wKSJMH7D7Cjq3Bh1hk+YCoY9rKK//ImNm+XhVRBPbWENkNuhvfARvwuNkTG/R4Z16WVU3OWlo
KAdrHM7kvgotXPBBBW9O8H55lE60ITaThbQCQ5ZI3+rxaMSoTYBod626pQyYA67d8O5QnHXlHrIK
65AeAfzQMg3YyM+Iju4g4md0sWR+CH8f4J52A/19la56oVJtzHO4zD6m9H3QA0lD2fJigRskQSHL
VtSU0tnnw+i++TS4MoLCjt3S5lp9H7DdQ9vj20PlqkoDoLYQ+oZ+TxVNkCf21DYppDS6RAsvpKQ3
wgg+FkvXRwiB+PXcadkZExgqlOQCUba2GbVGUzIAlQGvQYdxGiFRf+D286LjMFxr2o4S7GvZTcl9
lx/R2/Tv8JiZlepSjX/797MWTka9T2B0h1Tx6BdzypDyn2NsqnYyyT34bJmj9y6xTqyNpHFQAPuv
XbWC8UQy6IgUzfnLIkYGS4UAfNJM7LYZe4AaQCuZHv7TvuFr3IALh1I+ZQOixA1hNVEXo/vVzK9d
vSICGi0rIY8r9XHVilO66K3PCGUwzLy7bic47LVZSE2Ovw/5JV8LOllpwvblzoC9OIglNenplMlV
dLhmGW9w8NYy3EmPdrgcYiKvOJFG0ZTzcheeKLLnqHLCWrfuMCYTYoa3T5vySr51bNq8I+dQaH2o
S5WwyaArfuT0jdyESx9wlmprPNsQmDxFV8L8CT3OkTugYrPSY3tDYYzJAR4niir2OaXIrmLNxXrj
fgVSX/nf6soUE8sRtAzCTg3RHcb6cW2N8ZGbs3gmmm+U/vjJ5hVLK8TdDiaB7v6EEPcUzqxeVfoF
fY8HjGaPukSjT3DQjDwbYHWPbkegoW7cTFHseI4HaIg9TvblmdY3lG4LFGgs3jdC2xoETXB3Swuz
y+KuzqsFoJ8mdqnUmcCohzcvABd9QIT6oIAtGaFToKVH2kY8BR9ohDtGofC893oqhP3ZKTgHkdhh
5zuGW6EOeK1x5YU5LqGtjDD0xlUHW+qrzDxcsKN9gMYb/sZgvJ9DaCKPz3Zv+4T51x+9uB3AEpVr
yFBRlYBeVpfDiv0mZIch/owmsATAOeaXQBetjmB+1DrrZaHo4eskmbCt2OtL4HjY3OOppzJQafl6
34cOY/EB2Pa/W3z8f/waXwcBuDhEs4jEa9YaGNQdwrqKiBIJHAyXewaAfTHYaNhDor9SmOyB7IOP
DbDUw/FTqFOjZmsvrTvXjNQXQ03m4mxjJXAY0BihvI/tSlRbYZmbSDltfRD+cU+oZYJgqTxBQG1A
P9+X0NQ+JMXEFlGBWtoMa+QecIMxX0ASGKIG0oXvyUxvihXo/jh0ogroXT4xN03cWV+wAIzmxmdt
QaZn0Eo0ichTzm/RwDjgwlTATYV2GbYvn+pyp8911axsrdSgelqPzieXPPlKuTYpD5m4pXDLnj0i
obagCuTuTB4DYksSy89NWwPaBOZBKL/mKCeFrwPZ4ocL9EnSy+XeKSV6NCOxkm6PUEksppR81jU5
425NIMVhWakdtj1K3+TVOOet/ny1iFvzwwmrMcmIhMrDQXbLT9YCeXeGdy85wY3l5hlbpAUpWonM
z3ik3+5fpHLqMcOB+S7QLGW6gjnktfLonEM+iL4WM5e/5RxkveU8YcwIR8JMyTknDMYs8FdhGBbW
qCpssfkWE43LO7cZMZe88GE4JFadz2eXq2W+iiEAUgGO/HEJKrbzGzOy2FQeaXyKaBRf5bi39uoa
3dRMwHU1/Uzv4sCgNvFDL/Xr2Y951rf6G+HlddWjFnIfDn1XtdE0FvEEDJ/jAXGoujzJ0Cv4n+pc
+5QvAcInJd/5M/CCeyAWUUrmWOpqOgSCBfxzcYOxHg2jJziNA7kQekC7XH571sFbXuZtui8c9dwX
IhSXHDPlbUOFhXfh0df0tNpLMb1RNyC0XewLjXOJTzfKOxe5bqUW2BT9eKC5bwObA0GncTKyzrvH
qy5WzRmCWJlSkt/QVFgRKF42eEEAHhC8hamxJJSYR5+pCeNbw+61zcMvOO+bG/GtPOHZXP7bTa3i
bBxdJzOHNcvTd161+KiXzdkUklUtWNslVGGSrrdQAw3zC3s+VoK/i0udD87W8GdFasRIAbn2rJae
nKm79FHypvpj1DE5A8au6oVQNlJp6uo/5pizkL0vlBFsN9fVvK+Y7Ev8XGmAz/B16qMCwxotjVim
3k/SLlwRtlO7vpZufVZ49zbjl6qIR3ZTkTA1xlEKcgFMW6sdElCyr4SpTrVoqMcavh/Be1xRYcy+
UyB3Utb2pG63jKFnN4AGxAgrT2J/bXANGJqkYzF35jhPtdCOtDGFvSsUDOoOvGanJ6zuDQdlT/fw
GAaa9r4CAcWu5xNbqfxjjyg9uKYDWVqZcGZL10rSrblboueqbfLcqa0AXSOSVNr+2ouJOrNWXOvJ
1gyiC/2PB68LvPbU9MKQ2z/mOKTDECmeaFCaY15DlTFMZxG7sTjcRyHkxu+AHV6f9Ill4NaLLsJH
TUMLbPxyweLGINjBT8JXvhb3JEu9t5Sbfm8wzfGJX1EMwh5JhKUBf3mZPHqyKJPAGdhPWu+JJ5qn
55B2Lj3WgTI4xoWCopio4FGPGniNxIIJyUkWGvgEr/94o4xwHhtDSWdIoKwVLxueF2aIYvS1kwWJ
Xpf1aYSVxpuGG4VDVRwADe8ft+u1Dk0WPUiJbyMP87fzOKTBikEB6abeaZ8AMrka2j1vJxd3B3Ny
6QyUa44HaIOLeDxGFfKiHIn3+Ozr7jR75s0FlDJEwjYiIbpYx8Sj4C2pkpoUXJrDJk2+qTNQk6R9
jl8paEtEOA7yzsVSX3/NYdqYXUajyEFQDRe7d5VGbJF5y7FVeShrH15EXqyyL+cz1jx6zLAEndwo
Zs1+I7p5DCjMhMcbWal6yBc0UPfstm2rgCJIJC1Dnj16R3MDmg7Yzw8oQ+/RUilGuNYCH8VarOb7
H0OLEFdmq8R8scHpiucfxgAfFWmATzYIUVyRoSqTkYV5VRQ9/A8irkuvXa2xY4Xj/RP6YnA8jAQf
unLz2Wi0PAcrzGjJYevPhcb0bgprZDAI5UaGQesbIJNV7osCAKvHB20yRENya730oPHEMy2xh6jC
s7kqg9UJGhHjpOcYHrqqOupHOrlUk2boOKdJoKyvBqe/TWBmOCnsJts27ldPAi0IiWXBDmjeHMx6
7/k9dRbWwrRLN7z37+NIgiCix2WZApfoI6aRqScd7jS7YVLKy34lYHZ4HZWQVzB/6YCdSn64MGVi
kITeFbXcAtunxB+BsH32ElB5otXUO8jwtVjtcK3116WDItD/mJilyUdq6Jc8FeTWtuir29zNnMpV
WBF6JfGcvlUy2fGRUnuyF6k/HXlvFFDxvKJJ81vNlRJztYs/ViKtziTWcH+DdvxMwH+a3eAPw+5J
/BOVTy4eIEfK7OHAYUzFSsyevhXxr4qh88fyULwgb9S8HBgWKZwvzLGh2EEyIF5fWIk38ur/fmr9
4I1sE3I7pq/HBzBB1ozojqwBef6ivxzVjSuyrCBXHPV19M7yd6n6TutaU+FZynIDjyf9wdDNoXWw
1FgGep9YWd12dTKCnVTTgTQ86nRTpVQn8quM3lCyN1KMdQ7RBVyat+gBgG/9xIxVjMFYUg0KhP/8
pDSujycxuo0YtFWr9r6zq+vEa7NGvj/PavW6lsQes6Jq8YcHmpJcYoGtP1czOCpM/kHQ4yacyVQP
8YQpYOan/SzshWJy5ovrZojcYawxMJcort84O0s2vqtCnsKZP5sy2ZIJ2EbrzX5UREin6nA4biSm
XuaMRqMqvGtMzQFqiIOvz/6dEYugzcWc42h7ZQZZ88mRg4mAm7JUfxT6gW/RqaqOyxGULFW5319C
HHRVYCOnwMQrEHOOc/sHqtCejzt+Sm7sW3e0jHkSUy+IBZy0H928usq8/vBjzManbXR08OnOb0GW
00o+6nikRuYB9UpVA37l7WSYlY/JdbxGdpFPG6wqn34mQ5+oI8bnRjZXUM/GrGUwS6/47cnv7hYR
UVFtdByHj3O/aCflAW3jdcZCymMtRoWW+zy/OUt5eL+1OJLyyyacFWIdeCGU4ZE8tZWAZupQHSqO
7IiqdbnPRJ676pUiPISvUvEeuBBO3MS/dFOahL5StndE07NjxlKn2mJsLrDmYtCZyMDZYGKNQtVu
FLZ5VhhgbwebckEnG0GotGYyOu8mCvrGijMkmFxesI1VnfTQliEzN5CcPzipTkSTpVEmOJv72JWm
Aj7pu4zD/Gj9ESsZwLhEpl/2CgIzgbblGxv+NPa7ROHRYqgpEuM8c7l7UWAztsIUIAYN26oq+C/L
mlpOZ0oIfCIu/eJa/+ZipJ6dUiCq54bm9bAdBYwOLbEh1Xmp3aDAfMgmsjbxLgQemkPAXFypxCY6
BBRQn6n55ZYfc5SCzEBxwLmDiD5dzOtZyY1y6/cSgsmkpTl7PzyvgS4bC1MewUojMkbLCXBp2rRz
LAwNiiv/5CpTzkMkfXfPLL8/+1+81NSy5DMIgc5zszA3VeLmS70DwxBn4+2/5pyLkIW6bMfAysYb
sUyv6eYk7ZHuTtzzH/bULzmmxzD9vCUNXwdtYwafz3LzyzDxAYD2B5blF8m2gDnBP9/hcr6/aekX
hZKD4nuzw87gpXpYYufsT8W/YHPV1hrQJOXRT3VrcarJ25Kt9d8I5SQELei/fI/wrhLPCVqYQKw6
aWSsPgwEUD0aCxxxnwd6bcGo9HqalgV9N8i5EsEP9KiHscAv2lN9YEfqjK/XOkLsiGOUoFLvLABf
tsFjsRcC4JKr+zpqo7GhScsHkYaHwi0JHmYRcfr+hmbJkOfmP84dkvzSKEjV665oEogY/JjoYDBT
82fagsXeHyOFYBIl1k34Uho/RzzYzjQrEjP8tkkLsVTqSD8slryyJ5F1izvaqXZyOI2K2CroEx4d
sGs4tEEZhsJsWJAvenalnReTFY1fP1p6PHa3BJuLJOUSlRT3G6eQkVN6x4FwIG0wzuAVXE5mLSol
47TQRgQs5gukTkxSz+5m95cSegjh0oh3wTuYOEVWI8xyLouvdOKL2kJByo/CSVNuYDZmzJeHJWqA
pmAOWZzW8wwEOA0QBdM38SeWzxVkjLGx+gH6rKl92EFRZONu4NpoZlazJkU9tWCJJsXbRcej79II
zLO64KQ3kckCa+TGtZxtnw3jt5qZXf1kWOQC530SHehYwIRQPEpAnTFm+llKPPiSyFli4Y4jU2Lc
4Qqpz2FdajfB/HaJnv4+8t4oTJOZKoAUfY5G7v64RDhaCPIuMpL1kfCyUvutG5UwAKE8U8q7A1Vb
FwOhcPOxEoLrX0KHA1Qcpw1V9bV5JFVwMzk6JrMGIc4eGDWbcFQv1M9maNBYZCMSx1Y1ij62ofHY
HZ4GVIHX7p1MV02WYy/QAAICiVcwQnkQToywZmkRL91sTCLxJ2hzH3h4JAMpg5VyvgNcfBZbqGqX
JsIUG1dhz3RN+6qV22J9UPXwFtKgTuyaZmYEbC6BXEhSRkOBvjqIo7qdrrBOM1soS9dVC7bAhgvR
JyKsNI0PQgvDVMMHe9kMKKl52H97A9k10jDR6nv30/CJZWQnt1+USxsX1uZNVVhrlSylVy3KFsZt
WEcoAPi1B2H9TnKePsIArPVKlGxjuPGsNiwgxq5P13Fj/3Aa6NEzDZvkDHzofh/T9puwHTjlWA0l
c1GCRnJjTOtB+dHQUQu71B+27OwnvbyS0KDaq2ZNIho6yhyavyBX68GU4zkltWhf0vNaWz2J9qN8
Bkgr9D/HYoc7eyuO9SjSIYSPJaFIojqU4SsNxhMr+Bsl81quhMAjmQqVaLCwQUb3Vpf9Dk7OnLAy
vDlwfVY/W2fbk58Efz1Sq0gOkT6VzqnND9SiUP3ul7ZKDQmbo1+KNJ1398CJ6acv7eOxDrwBIvMf
KZYn1/tzwm58C9jo/+mEiXPLEhHjLpxBessHHCXX8j2Gb3mElzoccAyCO4E+EGZ0F2Llh++fD8xx
2QEN8jybMAqE+LXim0KSOdIoKGxXwKA9PBPk12W3K8yoBWBVc22EANmokwxhFPZcCv4tNNNvzGZN
hxrNhNoT5WTqCvNK4JWz494wIebQA/tydwYc76oRpqFGvskQqMkSS9jZAEbmE9HzD5LNRXAPIgrS
aQes5JvL+8i8DLQ5tnPzHy85h7ZyrD3IhgSqAy2jxar3nC6IIlal4lecXQlcyv8fQ3D0NMkaDG7B
XW1bCezPAGeWTd8mUX/IpKMx3cnkJv+XI4NOotj7/OnOuOLTGuscUYfio1vmV2UObPJ1ONfLHYjI
9Pbr+I+jN8x6+hHORmxi2IfRwB6jFRSu5T/h0Ac0l6iVUgyHuoYLVsV2XTg/Imsz881YyJkZ7qk4
wC67KZH//ygFNJdAv22HiPo4/lPhh5YY4+WcXPkDe4f9zlyOzoTaTcM5Js0WFaZ4yaIua1OyOX94
mNq6Be1D5lBEskDWF2lhRX/R/yQmH7WELviD3LKzuqSioQ94VgyZEd5RpvnGASutSWzmGcn4+8sj
fJHJsNivHXgcrYh5Wj/MEY57EjJuHqzA7s6x5BSHcYMOchwIFciIHDOmY3dzinaIZ17hIYlIOmti
1alhccGu3U7hcW0A6CjC49xQUQ/3iTTAOmlvndLRA0hZm+pY/UjPtX2rh64VjWaQFqmdU4NKVLBn
v/d1eEbFMbyef1VxGHG2qyIbZ84aaLe6tWQMPIHdp3LJFEPXPAR2Al3DplXTqI7Y6ZiZj+egnNN8
RjLCWruVU+V8ECxdK7MG0tzfTQItGjsEf1XajnPFaEWYEnS6xxyJQaRNCUYtOfdnsvDEeCQbpaG9
f4/Lbw8ZOorUNJYF4Es5+FFiENTBvW38PU+l9RsgWAUXmpbvrb8HLXzYNuBotuXYdou1cqapBfqr
2SW8SEkWKNBHZRSuVoJ/pZf5RkBc6wnlgh3ctdrXKrXMGrpJd11ijNhJrRPwbu/VHnJpfFkiphEG
6TvDC2mnR1L8FziB/I0aQFnzPUq1K9aLwblZExMbnL31/h/i+sqzrdEnSZ5+tO2OwUysRgbVbhE9
jfftGCwfpelDe0QXw9wF1gQjeAEmcKw2qh9uXlOh21u3quj3WmOwhyVmKzxt7/jlH+c73WNxc0nA
a9QFClqPom/fH+Dm+grGq7dUYkbbqdqwWHAmJZjN23Hh+eAMFJXuXQKXtUkoLYHIYJRGU3fYQy1z
muAaZKMcZhEfVvPwJ+SBXAD4OFUpqx/nN3fz1JNUbx3cNauV+nvx6YR6kmw+KklnPQW8/M03x+oX
/pQ7E0k7S4slAlLkYxe3japD+0tXYpjRuCDSM1yiNHk/7mGzW4VtvNWm2BTt7m8wCXwAVU2SjyXf
nLoQ/gUaUpQxrpgmnOoPPYVfWlONg7VrAsvgHPHZQ/5zQFx2JuFOzc7Nx/pBfM9YnJSYAWYDHf6e
vA8gLZ8iXkqvLtgCaYN09Vzp/OvRfs5X3HtVbeoEjuhzmFwMTp0vHsyM3PMk81Meanog8mElo+U3
9y3rGBnoQdEF7DgnCx+ElPzN626rZPbF5mzmELQ07zbLpAblr6LM7TsJc96UuR5TwtbDU8cTCC7W
H7rR7j6VRRF2J9nA0C27h3vmmcmuysWSYXr8TmJQU+Yty4jkeE1qaiYJimhH7Uw+hR+7zFb9E9O9
FxuMqoaT4dBVgq0kddtOpJ+udWHMnWel3a9cNN6t2Pu50OrjoY+MQUrM3qJYkiQ7IW4fdjoA4Z3e
k0m0iehANNdeL+voi82ea5rXGq12IC/cTvIEA6JfmEzQCGlxVBTMQKXi9iQDI3J2hYkgvqJ7tzTA
/2pu9bQpsKxTWAi/+T2U6EdR+Cmtmi/ax4ct5leAgNJ5wQd2WMlt2hcNOv/hN0FxtB8489+y9lmr
P1ZydpVxduu6WsuZ1qBKituUK9VBbECzesOMq2W+1WL09KL/rUFSAaXD+RNeBISJ3DcjVPjFX5dp
cw5JKwFvSSTHSZd8P5RGvvzMtMItEIYIfPq7FkSTE77VtmGcYu9CNCR3P5cvvXXFsF3pIyLmP3Cm
1iDwd3pNvBvEYkZduvRi3aovsqNmyKwrzvdGxajLZIEQ10B7Z65PIegaoU5FXsZzRnxeD02ZWKv7
oYI2YcWby1T1qXkefkZzpoeXn130ZgUv1iv4LJmiZICZYDhyA1t70u3nscY=
`protect end_protected
