-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kvpvG8XtabnHAcKk5nUMpTF43WKMt9h+O63+1O3p+W77f9NcJR98RrE3+Ew+IK9Gcu6Xhm2yA4Kb
pJTAsm+PnshAPe0nnqUWuKa/z2oxOIAiK2+SdFRF07itVLcOI7qp4oT7MBmTRm/PAuo5whBIHx5A
eB7h8XuIzTnVCfMPzCogc6G8irJknCiBENK1+27RWQ5DxfobJ0XiTZFb4X/0RL33e7DFZ9DapgyG
HidUCdmEbQt44REjEJ9VuBeZRd/ZxdZ8Y0jFdLqZdIRUQWdoCWpd/KLA0BrYVU47FWQjZQDsemGs
4as/zUMkXtE2I7+dZTX7HqQIZH3Rjncbqcz3IA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
G5s0pK7EN6yRIjSVhLZdviF3AP3W+emWPlw+WkQVNZZgnyRmZ2p8OtidIEYE80Do1KioT3tcj1kD
JfWtgzdosTjRrwLI/yUK7mHfKKGRuwICMOooZd526NNmuGEUNYRFZ2Esa8qdhXtOTebv1xIb5Z7y
7AcnKGD44WIOtEPiPcKajOpzKRzdaFY6TBGWbLwvH7nN84fICsBRH0HJ2xOCxT177A8VNRleKAS0
XoYz6GkzKgnGBe54P4XM4EeOTv9YfwS6KMh8TYQ919SyDdc9cMG2mkUWodc+HlqG6++2JUa2XuAa
KwiNkSz666LgQqh2fMkI+DpyuIuVEOLLI50E+5fxz/cgGh6hzbliFVcDSzngFuP+8sks9ILiW1hJ
GyqPXIDpIkyWS3GXc5Ictx4zS8llK4AV5A+uQsqEdHJy2PNe/FQq5EFGnUkQm0GC1RiHiG8FJ7+s
VDNxFXdchEUfwvej8e5blRCe+fx5poplveExhzaZrG+uk1eZX6ABfcqZ4TdpZ1UQukm9DIBv37It
QHGzpNuD6N72RtUMggUks/ryYT4zk7b+trLwkV1qoDU6LsBoJzriY87gjVF9abp/QfMR4GD7jSCE
oMgS96zurzD6AUNaq/amtmXE75kwRdb3GUaWZ+DiepK2MGvd+E/DnsK5Kd5yFeeUitRucBwBrhd3
F9VdTqX1AJ9C9Kdl89Rw98BpwT2gGKg9D9FFwaVmnLgK10mnAxj3Snu7ijGiOApZAvDA8XCQCaT5
xcXNMbR4VHwKmgQ1NNGe/qof1uwxLKCn8pXoZ6zpvwaOAvOlzvLvQBdtbm7ddtzI0vy9CUCc5Oql
754xjUQ10Odm04loNd46DdRpfzkdPvuaI6vheEPCYU75Jlxaun3QZlkb6PARZOXmiBfbx0wZOTM4
hPHLhcoBT8macgcTE3royVNi15275czJHHazEMKnoAmpsWxkkdddGzQQYcLlXP0TpzoZgLumiojt
iuDcgKt2gBeLjAHufhuBFE8brcBH9OY7Q8ZXOHrgi7jnJe3vlZnUJTg1xAXpYwKkfPIuF22Zl5hX
cgw7FA4t3I4+m/WXP7z3Aem9122rJv+8+fDkNbtttKipgOdNBLHg78z6owOpLwk0jLAVJv8RUWXF
Bn68eszdmHvOXVvpRDc4HTLWRBbshZnvF/4/FR6MirJsTAOuYMtolwDkq49jznnDVdFZfozjlQmM
F2ZqkNrP1AzOZ9futk4AoMp0FrY+DqKXCfbAjLNvJShhnJDx6oYyHbpvMtiCPWy7dhuaNxVtvR5/
aCoYR9hHhqN70mth2N2oe1DbUkLooRd9uv/Axt5HS82EevT7tpdX5Ic2x8zbD0uzrPDV7uQE8vN5
3JmAeCYq6sVO/ITdBIKYhK/8IOctfL98gRoth8SE2aUOlI6FL7J5cLQqEHBpjwrZQFilvW0N/0g+
libe4vZslnp6lEOpbzdpOFGSpK+iMDJfdOC/mHP6cjSEPmefGkrAiivAQINutKBORpke1dQA618a
ZmJXKl2mx7/Xo3HaT+wdwteVRFGc7RqelXYek7CBn7df5sKcu/zNLsF7BF1p4po784jDqyhjMtdQ
n7tNbsmr716fiU62rVNWq5yhswNBY6c8sTH77TY2GKbpK1RpIwsI0zXmI3v5RMg8JgRlNIt+RA3p
pOfgbYeYZhDEngD6p3lt9xFFl0N8QaYdcXqmjzTcE6TXqH70oPwLwYNlBpyEdao8pqZHGi1uvNCn
Ujp3yMgw96y/vRxlF08p7YnYfyj/rM8IkkKT1OKdri+PTOIhAWY50I0msRXrajYKxQgaU5ZPF4z2
gle0h7GcnlCvtVinan/Z4EbNV1uMomaVsSkgVD8VZ2OMamAuHmyHMndh82cbihA446g1WPIy/Ddf
BeoU3zkRxwDFUsfscWEPNHqx+dwQw3Kh0trgRZlVMjDt2dUHuTWlphQH8830n0pdvznUCtnLBj+B
OXadLbi1W0C0wGIZuX/GAPDIP/QhGZHUEgYSCiBQ6YRgqFHS5obrh1ch+Nsr/Bm8As5Aq4su+4VE
qFy1pufFmZehrEsQMcPYL/A/lNpE49jo8y/MnD/w3EoY1Daz3uwUNYBHDwdPm2fl0Jw7XPUag57g
cMmTP02bRcPXWLrjdrKUE/B9WMoeXmywugHdNnrc/dO9AmIpokdiWu7oNtQnvEREYid8CRIxR7Ek
pYJpt/i6b2WVuAj2VxSqYyqMAx0FpseAfG1w4baKes0iyq+vsMMLkvQtPGX3p7PISvZcvFqpkoqD
b825ZuLhH1Uv4o+4/OOlIaRwDdKXtcvym5+iCTOGgOMSKsyh3S9fUyxfq6bcPZ4TkK41ilQD6Zt+
Enh6AY19YQdm+h8suqhji+6d+Hl2cRUWREd8YOci0H+hMs3oUXKgzZjkwPDOSZT/iz1YsRRKuHsU
4xHGnrQUeYFjj8Yb958fx5WR6+ZICFy28hsrG3fGqoALY8ZTFP/LG6NPRsAdcfcVhFlYKoQQirAi
/qTd8mGJ1PSUaPCf/z7iXdBI7y46+e9f/5y8Eh38trK158FTy5tvCq7jsSufU0BS2Po4HMPYwRPV
CNSOKZcLMFj8WtXYjoMnQKcraTQp6RHrHbmfPSeUSJnLhobfL3s6nTgLGpiqBtJsyg/vyzYbYc1u
epWXGBQf78c8yKI5SOJyTHGcALlOgEj2Sf/HK3AQntvT9tLt8QeF8GotqQeUY3uK0sMt4t1KinoR
y13xLl9YBYBV59IZxPd86vSBBqkNyAPYq+Ss/EGdKKNAZxosojVhgxTwrx8Jq4Ac0WDeGuKwBvge
7Xi6AxOFiR0203wqHfPVGAOLFXhbPSr8Hhx37ndd0MGLvr4N18B01ux+0MLO9Ab65PBYZT4fvuwx
KxPIulZbGIUPzNyo2EG1CZ77vpc+0yV6hIBBmK4BCIjhycI2d8BfLFstHlozV7S1FN8vQdJwFvwK
IPJT8f7Ribmc5DkD1lFWJRv3PkFMPL/tjJ0r/Up10WWokld8i+Xs5yHBH2+h1FpydeF9EqiOtall
9Qm7M12c6iskQqtVGuSSn8MUZC6oJyCM5aY02ts6RQuuuqhNHNf7Td1v7TPKSgSC8le8yqg/aV0l
KVA6gzrTpn/wSHb0c6UmWqTj/Xos0lgelNe0LDOA1+bJWMVTioS32GPv7AU60wH1NjXz2C07jeMk
mW/B3/xZ9dq06aw5IAQUybW95rwD9fhcLgGMfoULpamxGo7H8dT3APDuOT7ToZRvs8nBXs56iXwr
k1zzRzQ2Ba5qIdD8gMWzhovGNMyU0WHXpAisTv9VJqFpsH8q9u6dpTu1nUz7f3vYG0zZ+W2AZvPC
t6JekPmiaOxMI3fnuxgnW8rLC5sYJLO99IISAwYfvht1TH9cenOyNX5w/5dDSfLb6KE6kPJQLOGk
oXGH7b9szc3E223RVHkJ36aMYMcb4uzXN1HsmEPTdRXYG5w9yvaEXnGxvSeyC7SYgfb42YGVkFce
4Vzj9J4Fn0cgd4gDNpaLNYRRtMxT+svw20ltwkJcnY0zJYWicRcXenrebPl940YRy25GNkdUIVj+
fONU86XhJTLoVikULyksPUIMM5gklA7ziYYNXsWY+M0AWSpTl8NW3z5lnridlHWv8dGCKUv2DH6C
XTjJfiLYvPYVoVqBpkNAovNU3qpzxwBviaWnwZgKCIIeiEKPZzoTGaRDfzyF67yuIo5iUQ2s4afa
RHEun3hjjjLOGv+5FZnRdhMhX1EdPkVZX02t1n07S2hTJOzYmFBmcYUBsJwe1orxTWnETdbWUEOR
F70L7k87ZM21NZacPhYsgFoCnLHn4IAsi0Y8HT7jK0gmyQjABtcS10QBYLAtz+gtU3KxN6OmYTzV
Egp9Eto3v3EIG7hzHIp7TBb9jZk0p8YLazHEFS2P0zKLCRBm2cpuH1dUB0Sg3V7hCZeGxE3C54L6
lgwPU6vzM4IDSnV59P8WVHdG5HuNxjWnBKUan4r8WQrGrqd/oWzat/m9XLLphhA/PPokrEQ5UTlU
43akEHLmzoFI+pv8qCJn+LIyF2/2VE4dwEa+WdniD/z8XOZlZe1K0EXdi7VrVPMRtuSuTKxure+z
PL3V6n+XFR9C2uDYnCGQ5T0UDZLeVIzUY6v/pmOIWNV8Wyz1tc2CIuoVLm0pcU6YyXEx2zY8keef
DaYICpyuf8VvC3RyAj+V5872U3kLpzbAqxT89pM7lI8hVCbegjs2zguymjuUJatj+ywcCOn1rJU0
WIxd/XTQESeDZtgFJXqYtzokLGXShkbhdZVhtIbgykcUkYyBnW6lOZP5GnnY3E4Xchglt5N3+hHj
xAywouCQHoQbjiTTib3rIVo/Qw/13/dfVHx+716phmPrXfxJxphKgytIFrXeMEPAQSmhI0CrFiWz
ok0DsdK3QF2G6kfarzwYnHL8TQAvAREs6UBEecWfxVRHWPOfmzCC0y4pyHmqSHQcb5GueS5A/pUU
a66YENK79465L8oIwcToNs3C909rIX7qaAT3dKefuq6kDWq3V8ckUQuDugXloSl7cqOBe239HlkR
A2CuvEWuDnml6n2izRXG81RS9IgMg3wFE+VRFvh/hazaYXIgaPEHTSDTG2EJ7aEXVQTVKuCY+qUc
/ibYUC8EK1jZfizEjSNLqtckW22DAKnLwFpSN/xSf5uc0t73gBCCvYRPPdrwCn6udoEsoM9TXWHm
Bda7slHA++lQiRT4tWMcYHrbqLygaqwbw+k0GMPx8GFdMzIbrqkBb2Ptd3Q0n9LrXgGGXdJWf4D4
AeWTZzbVLZkiGXqnKxLs1XN+t33oUTGwPPkYA/pDMP2WuCMScsz22CJnw7LnzV94cJa4CgJzhiab
TZx0VTAFdtbv4QjYipByikucrMDqlXFaLufRfzlZ/+LWLb1GTIYahlt/UQWx2joGRIyNcRWNIc5v
cjmt8/pp7pp5pP+BcCk/qgjtVs8lUq957N6j6qtD5AUj6y8LuCP30AV1qSmXhZKZrtQEPo23ju30
PkfwrIHIA6O9YyQoUuG0qr/Mvy3s314spuPpnEKv01dJmNXf+gwd8rwRISi09RlWv+hWFnp0DDhH
HmMQSAR2vebEirVvArTCVBtI32ZstmjN+ljIRA1BlpfX6BveuzdaL1z6HymkNTjXF1FyCNfT1J0J
IZCHiXmJVPrRZjh6rQ5SXTRhOzOczHML5jK7WI0GuJ1iys/KBtVZ2t8ZvirQpyQ29ILNExs4NYAq
DQ/4b8ULLepAnvuEsLqxDTb9+WbifwSZzwYKy7m061tUAc8HGhvrnq1MZSpRVvmpfdhSrL3Hw3wb
Pd9L2XcpJiaHA0ClAu37xY5L8q+9hiDk7AcD5BtEzIIAlCR5BqOFz6jXwS/2kjJDWDhSJ9rUeTpP
+B22nTcVKeIczqHiRT5F1uQAgDxu5m8LA3oUtyQa2xtfPxS0hAEZWYiy7OrbfRaob2/ixlbe1WBr
DvMI+ScYoJpstPG3do0yyTYG0t9j1avrPGQoi9Dy4kQvx6QK7xB9mPx4T+EJ3/OkIyIvEiIwzj7c
RSG4kytd4f+cPmpyUCGtPvt3v04mD0QaD7BnWB6VhT4q91BRe4PBPQeR+Pz4292OgdColjd7F/82
O3V9SrT9t97Ay367HfO3mgehkHoddfXL31moxJ1+BTH64Tw0+fZKiYIGvdxPq1k32pAzphSEhs+9
tqKKKdKNfxH2lrizb/CTgrY89eOuO3Zcf/qbD53fmlLHIGRCUmvdM7+8o3Yt9pwvI9WGZSKAbb6l
TCD1yoe6b8xDj4E7wOy3m5F2UTmPpkqjEIV2qSpz822t10Cn/ieneqvdbcKdtZ2zx4KfCKBzVTnX
9OGjuuS6tH6p+cnyQUmM2GtTXTeyWop7S+vbmtrrNwgQGg0zOXGSzquWN+KbBwOQz+7H2SrHpXj9
3DR+fkay26hlaP+/+SKWsmj3eulO4kqYSfLSDbYIa0AZ8THeA4BwPViX6L7UXenQnRkpeLUKvjEM
EUUY12sx0drjpk3wSD4zJ1Q66qssp48XYRNE8wOYv45QjR39oTsCmsJVYby5PuON56MaFnXLVawS
DBw0X2YIFRHo3uMKmxyO+8C6seBXpuI+CVPd9Q1ckWbk43LnFNEIzXWAEgCqaSk5GR3CBT2mXr0N
c7kCE8gUkK3OkrwQ4Zu9PoRzrDoe3JStuYZnmthEjqE4JH8tu6YU9OsYAGpMpmfeesLKNmO9711f
w+tE0pEXO/MblpRoT7BlquaeRXHcLM1ReVgVXRCBaxVeq7+wpAbZIVuEpNp4Ez4BjfewLIICjFXE
j2gjp7jC6dUFTgWUXyXo43G6/YUIrBf9xq+pG2gR0iKIhxB5FxBWj1+XIOmIKp3Riv96BL2SJjcO
rz4gHspks04ZNxDPSMKp5IiN/ySKL5Uqp5ghrQXWWpVthEiKMXlmkGwAvBmvaAVwwT6cPc70epC+
NLO8Wpsxwi5xcswLGU5tkg9Bz6H+nDYO35a7eE3P0R6GwYAn7Hnf47q8IL2iSdzX6XGOQaBEmhJT
O4ZIjYus7BJkVdrRW4lCu22bpp2iq08RFMFpKFsqScOrR+5pLZ/XoPSSkFnE0htVDpPFTTCNbrr+
BzGJx66/mFEVxC2DbecEExhPu3h3CW/3dgBRS9TFyIsBVj86t8wzqtOmY0t84NvNR4nx+kJCtj8T
5dYW8pdpWoShOlgzNvmLauP7de3Svvvhw6bTgcaqi44YTRAb+0PA6ooIZoKZlJcbGbQ4xkdXeCSa
J/+r4XbFiDAe2/t2NhJHHzrga7JossjccErtPkdq4L5/VqFQxfnco3Zn6PKxAI6bNDL1/uMR0fDJ
eRQToF+0hTi/HaiI2R1dRNcs8VRtUKJ6XUhzOre2Q3eeDrCum4GoLuZc8TN1A9ettsWMEB7/LX4p
8IlGhB9VaC/ceFqDL9/9CGpS3nXLb3nEL8RUryQ6MvEYLhCVdXt5JSJSDeHaxQPJ7EybbSjE7PaI
lfVOCz3pMobRaR6ptmyN7NleE4YH+/WDclD0F87cwCRze4Emm+ZiPeVJrxwdavm0VUOJ0tWzJNfs
qH38s0PmsA7q1CdjzQPG6JAsbMUzJ7AdJxzX6d3yS0Oi5U8201o83TVHJos36bhxcCYI8q6/ZFl7
CRf1GUQwIGp8ue/dSaKjZ8KReXs5JLPm4XtJQAxXsyNPE9gofGPwx3H2JZXjRQMV1rjoHwmNJqOg
/aqnPL0UasTkV7YnjPVKiKXyaueZ+c8U63XVlEKZf9dMC4R+mzoMaRhuZRtPNOdlrVIslQoh6Lqh
qEcraGQcAQqQbc1OSlg19yBqZKoSrDk5eY3YIBqZczswbaq8dKODbEe2cCcMN391as0h/7L/nD60
/Zn5MziJdzE+/VUjwYlt3XL4jZAVTR0ZJeoVcQZ/Ty8uWq2C+f3Sy1wA4g6J6DgIMcRSAPVHNV0k
D1r3fwnDStbFKEGObCG8VV2sfqm9ZzPFMrmwdDMjJvVES6mS2RaPBqfIYpYbOBsHfcnVtn8nQXMh
vGR3iQSa7o9Atejwayr7q5HlpZFqfaSiXgQIs7x34BLLRx6+uDlmxfwpCge2QnPfi/zQi2KxKh/u
yfxL9QGh3azEN07qJLdZKL2qjdTMGXsh1D+HdqqQiIKd9i9/xtujsEu5pjXWL9rP2KTd9CRQJ+aC
iaOw+HwWr3ohU364hJCnIAHmSLVGC+w5ny48a/Nj/ZjfWLluDI+nPM7ppsfpzWmc6Sos/Jz0/77I
YZIBUpx89a92E+ZN3uORBK9scNkNDaKRpABZDkekJLMuCIpvyF5TaqJ1e6W7zSQaPQMTOCMI37u1
5pEQf1dxTzqk8QgPsAXIe0yOd2bGCI8ZMp0GqGSaUHlX8xIP+ELME97Ru7SjCxLmKBEYk5US6khE
grOo7v/iCekE1ZCoefrwISgIHzCi6qZIpK/HGPsmrTXRjrr95pPTtlCcl8JGIjX/d9c8/IBWmmE8
hYXPHfermaIV3JZ3gv9orLnusOJrkMffoGjLcosTJW6ogyvEGYnGk5/jnwvuJsbSIJ+oydFxYqqk
waNSHUG00U2iHvC4fHKPiREjf3zUqcR64wJ8Nkg+A3Rz6mnzwEBHVX9utSN/Dz+1Wt+1LM+HLiRo
rIxh/63667DlwKjNHFfYsA8GYTOcFVreArf7vslhpop+1pAMpOOeq6GXRjOdMJnaHQg4w9s3sgj1
if/5s/8NycGPUj/3KtCE7hihHhVlmjKmdF3N9xcmfT27iEj7IiwOaNzmkUqmjg3wPF9eqDYvz3tn
8aU5apcpmhLDSZ9r+239YN0WZa1UEudgko3qxAhcC7VZ1C1YVBtgnvjwogpwF3jwr0OdgxLtRita
nEveHuUpYWU45tXhJnAjim2dPyzXWEPZfNh7l6o5mrLkC6va/CGMu8UKGApyZm4UuCY/7r9x66Og
GKcd4mzFNhX0IFE1CI36lDWdUFNTsoPJUQjH81U/alyuj98O97j216aHzTyHpLe94JsouhAVKds5
lIVOAakCrtRii7g76cmlqOQUdi7nY49AXcFvcB3QZou5E2EEnRxYvE2/OzfQ3LGyh6a2D6Hpm6Yk
G98MoU0vNEpoFPJ/3TZ5/2yLtSp2AorHV9nZEKjsCxwieWd3ZZDQRAAfyTxU4Q2dA5xvmHdS2GJ6
SB0MDSZfTbmCSSA3dDHzbHIP3siTj36vevW3VLCfdxznUS9dYjaylbOwyenaUTdGiM1XDP36F1Tn
e3odQuGOhnUsrnnwg/5htjAXoKzkZUpZhWs2sTLbUqUA/hZEoClCHomaX+rVuRYiEgnYGKs7x/Qg
/xF/jJlLR9U6PObOrnTp6shT5H/t5UXB0ABtKo1kK0FNNoz3Pgxk8yhmp2tWZ896g+5mh2oCjLUE
rr1y9yobZYFkqOwQ3a62RZh2pGKvCjyeIRQWqCRetqIdglwTocxb8CNG1Wbr3lfnE881pXU5D3/h
AJHnU0mj55E1aCyZHGLrRSJyPTD71hK3Jcne2nihXe7JdfH0xQgVG7sU04BG/3NVYUs0KDN2tMLU
opRH2u+DFf8K2HhBFfTFq67mj1w5j24WCt5M4K/f0PTsNl813vdSwKl7OsP2MwQxS8cgnE5mtg6M
w+2eMY2y+BsxpVHb9COIb0ROm18B8TXNcr0vH1Xq1TgMAHSkRaII4UQ8xd+UVojwkdfwzCCIuPqr
nFmLiWfv4t2vig75Xr2NTY4gV6aCoYNhlZ4QUIKijLvjNyDDPkWQJ3/GgYFiFA02EZRvtUvGY7DJ
r1/K48Nz+ooeAnk4sUGUObgDJpkHKhq3plIvT0zs5hygC1HZ6BEuj5x1bXo0gzz8u3Jx7rP6kqWU
JN8TAkJmGtGDVBqQqvN0SOXQ9NUA/jv8ghZCXLCy0WwbjLw8nQ4+Ug0bROOvfINer9och3lXPNvq
hrYFzEFJRGYgAq2nEQ5cjTn9z7K3n3p+42v9V0BZsQWNEhzvHCLqkFkJ3tl4u4GUdDFANekFr0s0
HgnVsg1CyC9yuJqevOSuMsWuqOD8XfzlVSwWuYk+WzxYtLtDUZFLvtZ0pPVMAaWzHJW9oLDDke3d
rr8zwvHsKO9BYz6GweJhAG21yiHITU9XI8S89LhuAE8fO+sA8R42OHbSQ/EkMwpMmYJJWGT9GnH7
cgBHhPfdIx7lqCMPMbRZBRFKS0ATPmd+oAbLzBuVbSgyRgJp22zljZcZN4zPL+VuLqal257wdSSC
QlprnHylM60ceg0VFwoFAD+M7Ka8HPmFuGaxElS3u/7jib0NxDTtYwd49JjFHbn90+Kkb7VAjZHO
eWj7BNMyR2gGMcv6yfKnCfynr9/tMR621OqFMke+tSGGDpkmn6tPIxknPXOg9AbarT/cdACNg2ri
7guBD+MMlV18qjYDbDlZ5a+PSf3m3mK/P0X71hbM8aszrR8X3Pr5svE5lIG3MmfIQ8Bkp+muyfYn
m3XpUKwjtMaHDVJTf3luXXOMcUc1WNG0c3ySNvoQR0Dr/yC0Ip0nOPri/h+pYXA25N8K8pYB7CHX
fDa3bab85PjRU5qwqMnXClFMhMB0W8XVN3++bc2BQt42tdgMf/oZ75UT4VvaStCkHr3TnJ/TGw8X
Dt+3p4g3RoI7/SAdmNtrexDs8CefgJ1dgDqAJsvY6qR2JUz3d25l3p4D9hadT5kCCri42GXh50ny
uIN+gWREeDJ8cvPaeHVotAeQC3sWSDad9AZQrpyp2n2eMMpyg6D9wrc+U9wmEYD4nbveo7HPg76v
CI+ryF0PW4jxmD0++sN4mDIlKYmvjznnYiMoHc1HMcWgebHaX5jTjbJl5pw1jfpw/K+6UtSl7H8j
CNA6Q5DxDrGpTGUpJ7fZOztx7mmRzYiNjRy/rwAGHCtiqXuOb1yTqFxdSSb3/kmYexLHHuqrB25I
/tz+T0yumzuCf8/tsQ7Lz8vFX8TJ1ZnCyB6ljAp9JiAbjhX1TFsfeLHFPJBWZ9g3mYGV740P9g9c
Fk0MMqiohFMtf0Z4IFKC/g2KgGgfAzNgl+mU6SaGm5opNIpCC7gdw8JY/zmXJAD1r24kyaQosTni
WWeQLsHf3dpV3c9uo98Ceqj0nxe4NUf25egP4Rerg0sZ5GUFWeKxCUK6efG2OxLQtUXF8jpzLLAs
nWECkIAsqaoiMcFswf+CP57r6MRkLkSUFgWiRDFNeJRfa+yxs4OvfTzage5kIYLzeGlAO60BNWSn
lTnwtWsFUwZ4NwTgMOB6jEknwSJTjnh6b5XyFntQEpym5QHCnB7KHUbkyl9FnaN3N+IsDJiEWpho
Kkrxq8Oylu/fjBm+PW8t8bRRimgZuxvHWRWHYPFlhm9BX27dacW+HV8gxDRmwS67h5yDMMituX4i
P8Wn+NtIddrt9/FH9gkmnSPqZc/gQKfK1trvRNoQe1b2ZfIzcimUXNnv2aidDKznCSFP3Jdv2Mhm
FJF1o5g0O2hnx5v0VNxHmue/UQAF560T4fvRiOzcSMJum1nc1fHlqn/CJ3FmUShNnCMW8/NsX2v1
kSYOP22zjIBO8lQLENs+ohgjaFwGFOkCGiSK14IGNtRrSEs9S3ZvXj9Gdgawu9tvEK6SqPCYVCPn
m3yTdezEolun4AfhKPP1Ow2aFjbxeL7dn/N1AGBjRcd0q7xpornn+8KJQJh1TK6FM8FYDHD+i1Tk
QsYsouJ/kufUYH7CY+f0rl01jTRAR7aj5XObTq/lm0nLQL5ll63+A8Xiu2NUi53Qi5AcQTcWh6zj
U8y3Td0byyGDNuPGK12QIu6hIEUXiTLTIsYSj4CmMgDe8bQln7Jz7jX0L5jeNcfguG5xz2kgaoZN
hLpfI6Xi+E/zSQJtMLKx45F3kWsoqGHEa3rIc8NTxsa28ywTFd0RWAhVE6CFHw/cy0hU0KFVgAT6
tHS93Z7rfOSgd4Kc0IVnHQ0RLSkbbANkx4kvLYL5WsBM33N8dWqpXR64nVhGX4euV+uRi8uoz7SV
DtYp3l8qv1FSjAGE6NZLmExegFMjXIPdPGf08AENvsufgR1dvHfElmElas/3w49w0Qdt1Zxcylic
0U5vcrJKlliJ6gAxpSVujPuMmqdWej37AJZwvsg95TdLrn3uJOHkpDYU6bsNpUGEDYj1Xe/8gjxQ
YjllWumx+Bm3Mnr0qVvAOqcN/dcdxsppM4kWI/2GyPsoy0JoIIeI8YQmf4SzN4oESe/xzDVGg+jo
xMbn/y/EqIrgBtq8sa5Lf2WMW+leBVeS/tJehlH7GAfJkjkEO0DPziYLskVrNrMkk3pDa3gNz7eb
3vxAJbIvmYqre6ndDk6aGBh9VnVNtPRbVmGpn7UjDhMZkqsTOoq6eAhfyr+Cyg8TQqB95HTVnOWq
yX2APi0nX5R7d1J6UDZXCP/8/00QIB2Oei8DSP4y3FCRZ0BAcGkWCE7oREEAraWrZgIzfS2SG+gG
iXAYDLlsyahdJJBEnhihpe7pGEsMwJw7aQ9vl/GkBqNb7ivGzKoGxSSt9F8SXKAUbqeJNK9WSg8b
Ktiu1BKwSjZ1xxnbxqtY3zfyKZRmnccLbS5KFUX62ZiDiv4yvsPXYGEJWg563iyATHEAGrMG/KZX
Dkv5zu5a9hvhqCENahAQPvHkZ6gn9/SS4Kp+JoUlQ6T+aiKEqYVTDLI4Qm0O1GEiT/oEQBaRAogB
5X8r5SvoxlcuIhVqkt3125Gr4GRpbTQ1vV0ak9XoxGi3ygh7AJau8xb41hiOBr+yaSIme/XMYpVa
G1DbTr2re6Fi7U+j318GNGqPp8G17fK7Cs5i8hdMQ7l4FfWxpEoU7yoIKgf8STwEcJwdBn0rasQ7
UzUhkjxQeDO/8WIpPHy9gV+NJxG1s5SQtUvPehG655Ry9W2LpQj68XL2ertSij4ZUxG5v5JfhKf2
1+XGdxL60D0/xdGpbUhEhHoFxLwIB4flMdsWr9q4f+gIuAvLw8XE0tYy7KzCd7RdkE7/9F9WHCMD
BdEvK9aBKPWK/AgkFOQLoaWxUANZay8Y5ADsebx51oVFhdEdDgGpQMpwZcZsFfY/YO+Gmy/L3oBL
r84HCDXA1oGm1AYOEBMO1RFlNjE/CetqUddfClGEEPg/6s2H6P/ZQey2OQ8yAXNJE+Hkp6gbmKxt
gfob5xdIwjzwFZA6Dzv7jD/EnLyI6UARjNpe9fB25lDtc4sK+zOn0BEKPr6wQibd0CRCKFWja6o6
FIKwVIrIwMnqZ1QsC63oZWs9OsQLpjWwix140GgfAlDFIvsMllhVKjyd+mpJuGS1Re2/MH0i6tec
9EAcyfr2+NH7pBP5O1NnYKNWsg2jpTQAXG9JKtK+HQKbrbFRBJSir2B3+W9Zfu1Jc6zAqELk6Z/o
ewi2La8o5Jzig+5Db1ic/wnmxtFFRd6HLRUJ2yYuJjM0ujnU7QUyXGYEKcpUpujOlrMNy1ljRI6i
Ss5rsGWkln/eiGBX2uEFy5SHgP0AF6l1So7WQtAwba73UMBLpE9oJ/jUoG9ojEU21zYgwCZS9wpK
m80WKJYGmOBn0pmbJQvaeDXanKs1Vv0Qya0/lTwyb6/zxu/4jFNZSiAuHtrSOL85O3TIUvvXy/Ux
p6+UBWB4wu4vbunfiSwcxZuWpZhJPI/Elom0GrDCz+q/vQqPUeEkSYy517gjzJw/YomWAsFIBTMF
ynql5PCb4BmGZpZ19CUhksgSklzNHg8XMEwT58q4oGyDzaZLS6GLbUEwj3MphoFH8+4g7/bmoya/
rv97zWnQhMJGOnIA1Weo8Y6wPTB5lMSSwMJZOXQ8fyGbM55ddg1mXzGjUq/EWv++JykqlzIyXus1
WdZG5gjg2jMg3Kiww5J1sue3rqAn/q1RT8S7clocXii3aNEg6rKZPL0BoIiHJmB7KfgaKn5QASlR
d7PrutTUeNH1eNIMjc0vme940glTYRuUTBNP5yA/qi3570ZcUe8puWln7UyvzSSJqNUJDe8Ts2VB
QKvDIjZiJSUGa+1HeAw/+8b7qVE5zUZlEXyWd5NkkRp6YXZApDmHxOGdU6qKUnLPQfwyAg/7Ya6z
S9/fmPnWIFvApPd3KKikHOlZDp+taq/kPbIzG2akDG7uZNRz4M2C2ZmlHjoeMZAhuatDR/fw9uDT
7YQsMRLFWRktSs9kzJdzyf5MXgAnleRm7UuXTPjI0mdl8vpVFk2NOCX0e/+3WPQYOTGGU0VYBsH4
vhXGkuiYUSSTREnvqdL/ZQeHrZemtoP6aZJ9/IMDKyFKD/yFbFWVuUTQzOMEc5RKykeQx1FInBKD
BCYrGRr2LyoLDFwHtu/gyimWaDe9mO2FXFEZrpR1vgf0qWAndTXQZ+xSYrF0BJPAL0ybYLvQ/tKC
O5hOBY4LVmdk06/qK94W7CS0IlJNVMHorfB/JhiGz27cRaFv2MsO3jSNnQcsxGWmrGsBeocgYrJ9
dkd695lxlTb8Rd50fhWGjhaALBnHoA7UlAdYURRQmY9YRhGrtm5ROqQ1ANKpuLxFM6gzzfIf6vZb
J70QmI71WQ25DLtJryUVCzkt2XfNp40Wzx8JXWl9FTwbiGF5PNOSi9aeZrnyV0/zCWEvpoze3gRS
IXuUH0g4rl0YXaLSPC8ntlgnLTa8unGhTu7JB4mIEmYQqovyM/wF/W9WS4fJjrsbRaKv2pI0kMc5
dBLia7e7bkW4z9uZdi3fGEWGpoERTiriNLbs0Rq4Oh38jMJks5P3Jg6q4+V3PuDchYnFxtwvpXCp
isdshweiKhY0rcNbgtxymnLbLt3l+RRhBWgn8tTN1qiFn7C0mzJOA0DovDxoWcmhIu3iD3xYTNmh
cCGyZVHXOgT3pNYuuQH7nXP5BA0KcnpMxjDOyTHME+dlonWn/tIS7W+gMWp3RZTtR4So9GdvYm8n
foPfZkqaxujr2iEYPb155j4tj6CEb/iCEpIHA4CBLYB8GoLdgYR384J3aNvlxI/NLDMwnx8o8S0I
FAhAWu3bhYC43Xt013HXNOf95PA+nRBPFl3S6kRsWByRb67xyX0ygiFfjepisTqx8HNIP7QYbYPD
1Dqt4PaVHAwEpWwAQcOlBKobVHBQjnT1Ue66fwViU7dlo0fstdnnPtXjSsF8Aq8C22blRIteLACd
46CauJYtIVwZHITnQYKx1rNYGiQY3SLa08ILIZKSiIQta9pravdCxt+LU4xyb8MYKLWhWV9DWIIt
CElh7rHacF2M44xseeXRzs/ZwAtIreWWGahMTVBqUD0XeehAeo25fPnyXt3Dreh+Xl2VSTDhO20V
lQj1mRt3WW31X4fNr236flcPmdweXN5SDLP+RApbbhfWGChW1KjoqQpe45G492wVcPqDgAQ5WNjx
YWozhA2zgtUDV886J5dEVIX8L6GBuuu4Hb5rdiRrrYDgdRDaxH+6l4OP8f8yOnMAs//vqkFSr3Gi
EZ1TjU9YvnUBEFV09SIR+PGY2VxounjNvhapsZhwaTgiOV6sWkjASVEeUx0JzjsH5laYKQ1pI4kL
UDAFfdJPeeT1bmG8mhWHNbiwqA6nHJNp2qAmOP4xOQAE7GbxN1EFvRUQePVKMF4clhLqCreP2pFh
JwfxnKxZBH75COJR8SSIoaBbkgPNfUf5oTZPZ5virfzIM74rWZ7mP8Xhq1TbEvbAh4CDLPSgK4Fe
CK8nJ0PZ7UuSrGqpxDhgMRDQvGI6nySPTnowibRbM/xHhvhS4YvDpAsJKWwGFYtEFjNd4ggV6pqg
aerT7bh2K8huMOT19NpZbcvIoJqYNPdGFkle5I8csby/BHDBFg7EcNLvsMtQriQFPCHOMLO0AlCn
l67HH/23bWQJMHz5lm797e4EWP2zv9Cm5eEPLQSFzBAQcN2dj/To/44e6HMtfG9Ous5tXiEtP3Hm
GvG9eEJ6nxBh57i4/hzfTySJqiAC2Rz7Z909S9JxJNxcxska8eMizSBvB3sknifl/QVIkAu4oS0Z
XnG5gSHP6DImHWZmtdWaqXXAyS4M9j01QVZJOgc9UU1XVinkkxVvq9BwwTOdaBN9BpRmLERurTpq
+yNOY6kFoYji4/UDXuN/MJs/i9x/Jyg09Ac+byUGjksGHF6U+euEfi8Br/Xd3CCBae2PUeCBTmcU
PIync6fnqOTnl5LX5FF1f5fih5epCvhjtSIsdLAX2OCTwD4Hcbr4/VceZPotfOIJbVC9AmyMMoAb
d65iOkxUpcVDRd6jUUcU9UQqEXWdCUZo6BbpUyT8RndPawpwQt7X135d04ue37DAiA6MthdjJb0W
KyaQvn5QhfdjSsl/br7g8MnxE3WkSiCZhE6vruGTHgeNKhjbJ4dD9i79tHF4Sq2MrZ1AtduorJLI
vjRf0RrqgV59pfef8OH8b1qY3tZ5YKnuzSdCao2s9ttOw/aUznoxXHTqM4vRh2g7+gqJU9Dyk1LO
RzC1OtusIo/W4PFo+DXaNhXaP7AuEJF2BvQoBKeXzH7moLve2C4YKIfq+25Glec3wgX9aq+B0UCg
k+Q/k+RsgLVMtJMW6cDYKHhjR3Ij99LTCPxtzzoxP427/RPZVpqKzQ5M2v0T2Y95S2Rp3AAibatk
54AHPfnofNZBiVeklyOetw5KLepmSNdcouOQKWERDIdBc8yudlVwH7LXD1A3vJlGEzEZ7UAWWF26
TI90Y3Y9Cs16cbL4lcdnIHcb0Idj125EoHQqznox5JFBpnjmnGHPDjtdjlE0xhoKAgDxFKbfAEdt
FnRPTrk0HWy8rWEfJNVIxleCMjL0RySfS+E2NiIUr2TNj++HQx7jiBNS8o2vGRFIK+wDj9KIh8w7
j+dsVFVB2Dpzabx4TYiI2Gx+LXOkpHWzBlIbwr32deN0WW89SXQLv9W9dBAw2K+9qZbGRBej8+HA
JxDiKMAN3UR5eln37zqzdwR3X0QyWZ5rDSN6o1GvwWm8+OowZNMbnnTOuabm6YcL1LMoSd8uyEHZ
O+eg6SDFEaLGd5yGoyF7beShQoLuWUp8V2Ue+goGwEYKadEWT9XYE13ZY1wQgtWAOJI70wTqAcL+
Z1i/f0RlVvEyikW8Mg1qsEHnss+4fOxqHm666GG5d6nK39Ci3f64lg8oAFvBP+mldaAPEqBq0a1/
fxyuww5Br7A1J8ID/H2oUcHhC0JeuvemfHQ0klAX1iCqUq00USdtzy1BN3tjYoI5lWT+/R4LxJiH
wtB+p9XqUZwF3NWpoSQUwGrzQGkBSIOsKIVNYvYstCUkBpEBKFyZwsNUdXSIfdSa/IRHB85yd69E
CSK8yxRwwT68E318Pp2kQ809JYlE2BE5UGqLdvdJCWqtBxeH0yPMl8QPBQJOQejWlCO5vCSdWoOa
tPm0nXaOiY6j8Zpd/AXIsebaNGCka5upo3WzFAsChzjlVRtctWth4SzGZSwGdHA3S5tXuCRP++Co
nikPHdl8MkoDhVNKaqzj9JZZ0kU7rapxRu9n913GBAWo4ms438PjTmhaqhgjIxA2kpqcJSjsDq6X
dvNDtEqWkmzfFj8HYdr8BTFo4oJ1X/Hir3wM4mowA2Nmc17vrz4zfHnYKTw3rGLA5Z4DSHxke7Zi
gaDRvabTWGFKLuvEPDFl3ZFlxRlT4L1wJhMO/wrJF0uUmqmcQ+N3uvJunryqslP6YVCxRBT2gktp
Q6aPVp18ghjmnr86YC11OSri84nlbT6qQVj8k9I9WidldCuV59Yl0QnBE79WK0rwrJMbNUT9XEK0
CpulKUhlKz6rJZFWGbiGgjvfSA5pLYNkSQt2NiFn5cL8ZKukgwIt/qSdUrU6Qs+V1imCZjn6HWIc
8yg+TqqMx1EIJ3nIgdVtyBtALxN/YfWV8OID4VJquTfFezMY2UFaulonElVEVagPJTsUoM7lki5N
XBZVBuJ2MnCTMxSAgVrdpEilfp39YZBXpkPbR79T3BIXIYVAVnWzBVKGaiXzb7i5cGLsuOMIDFKP
qotf8BI2Tz24zj9bmQVLvnV73Ye3Dh4Ihfb1Pya8bLgwbrjsBC+2Dsl1Zsc1k6jQUCvwApztjaFZ
6g4QTGg/boLIjmaGHmdZ5f0GzTEN5xM1koVOixGSDJNonjZaKjgSpI9cMYDilGKOhLQrqHk2VCwB
GG59bwFEWCCakBh8vLzuP5Enm2s+8q7QtuqunjLqju2vqhz4TYiMjVcdatIfHqlGMJ3jAXfXqdiN
UmBCBzGZXf7hP8iw2/MUWtA9rc/t+FHoUF8kjQG0cHVXeOrtkvdR689+3tAZpgX3EnHssLVTe/9m
n/IimoVlIgEytKVF5J611Yet/XD3w+XOwsfcPAEWLm0c4GaMxOjarGzCipdhpwSeIbCSxUst5x0p
TJGfU3ImOJG2Fu2EG1GxLA/1FdYzOOo8zX0Y7GE3YIbew4eAXCR9dQ7M75uxwuNmxg8ktrD3c/xg
VUM2KNVvQFCaxtwxdLzAehrkRNfPWgU/LMU7TZzR5rxQzrIlEcIUj+o/sRMje+YgSpraV3YtbvPa
1wUtLaYTaAtW0Nk/FywBkP+369HM19Pn9ECGoFeS2B30MDlMBUUZZxA82Ana13KEyREMZOJkmotj
s26pvc/jH4w7VI8/RuSOSPMQN6cdPTkVWi1q2v2ZTRBR/NyeVeJt0MsjJYPkGco+feMfpRYnkzrb
BX73E7kH5LA40H37Z4VQd+/rAytUfJakYoGmKOfrSdFKhkLftC8x0NQBRt/qRUxQWxrHqnhQSFeQ
TidXB6Ud1Fsy2YF3JZ/Z8Jiyz5e5CxfWVURYSdGqSZnnYjMfSBr+vp23mjX0AOHElfLBMdq+kcIG
TGVaaRE2jJRzDmajaWcuE3D7MYylNyN2xIpvo08Ca98P8T1/WrMZT4KmDtEu3WS/KCtOiU5iq+29
Fd4JGWgC4lkdrc21oQ1TwR1o1BbpLZRMJiHePnDWoRTn+2z2eRothcmXA0NsR2M6FgWuZTlcsxMJ
zZpvFJtuNGlc6Bu7yWCayCTBXlNg9DN3cMrxjIv3rbwbS0LR1hObyg/i7SqAUhDOieXqGEBI/5Qu
V3pYqTuO/Y14w4GcK5NezZdFnNLp7TvVqGRtZ2vT1zcNwgSatUxB4+ZfcdRLQESFXG1WeRFeXv5h
eDsdCszgK6fZdgw6tFrWMu2+CH2B+SoKBzwc4xJfP+ndUuOdOT5NblEoKDhX6R9loqV/vf/G5xgg
8xZTy6YD1Q83MuhJTDxHIhHf2dO7HIt+euPAwiC8+0BIm6U/0BNFlHZdzo2G6nw3IXv56nYpUgHQ
qjjBOHoSkolMvb8MMEj5B9maNA6sn9Ylj6nSRIWDY0x18Yc598WTgg31MRipm2YRpZtPEn5sdsTP
1HZ7Oe6U074YCpqIpstT5MaS9v37CaPgw0qBwpvj6AJlANsION4a6xcVK9TerEs9IXR/UJRBqNZZ
Hag1S3k+Jvyeqoxy6Y0APWriw79dmJKcnYH6LlioG9XFGYIefsrsFOr2q8mD+foC7RuJySfRIo3c
uIgJ+IS3/S6A3q0loSBuI/xqxu+NTYQ0yYN7bIBQQdD7efjn46Eta/O8GwgzTGKDd2JQz2WUU7GM
vA4qedgRTx5KZUN9Kogo0Ridf/30/sLcqB8tz/L18nGh/z5jmS0HD+T2dTiUgVSpTClBsy8QUtpO
sK4aVvvAoUR+bErOSSba3OBisbG9pz9HGeeoH3sm1h4GqZ7oq1X/dMHonrf8iWMFn/G3e1yIplDw
DIGDjSu3CqssgjfCbBOHyTJT1fn1fYn0kPNL2zjc1b6AYNyCFz0PjL3Tz7UxLx3grWKpU/dICbsQ
d8ZscO8a8RfLuYfkyFnrmdddNhrES3DZo51ybQZUj/p0fVyLEtBMH3DRzvm52cpO8Tj9i/hSlbnX
R5vj+dGeyA1fSkFeTJ/fpKA7D7mb885DBQucAWU/GUF71dB1u7AiAy7iLOUUgkaIGO2D0fVh3Cbi
Kn71HhcX+U8GHff8egQ7m+PTHv+vwA8SWbRt+rYfvhty9qnZWf+ipe/kgo7R86njncemvFBz1K6j
jffuDrqhMGxnW3F12LiZ7lfy9kVlmhhX3RzLi2xEU3mirTRwr1pRB51FWg0Y6fj3Mkj3pbkQEUR/
Hgn6yYp0o2ydonMZVZM6uJUtmnO+MKPNcCoXOBChEI7p5d4V98oa+sRjJtmQz+R4aQWN8WQDl+jI
ySGEjxIhyLZ9vu3sCRHa9m8j3nO6SivizRbQqDqO1dRcK5YGjxaVfSnSirqBOxMatJPi1ijF+bPk
CHHOYTvo58MQyZF3hzxdYnKmEYcgE3TRHH2hh30mwkHkG0rZsUr2Z8zT2/d9I5KJZojhnJIs3nOd
8SbdeN3G47bR79YdC3LBEQHNZqyQsCmleTe0lov1XQz5DgWXYfNKl+2oAyYLHkFB8p1uKXh3FNaa
qJOAVLgW14aCk/wPDdfFM9ExO7FME+qln2XV1+ySaWeyn3MIcsE0W6yWoEF5cYZr8FTHioouGV4Q
/8HQE+RnSrVYHxJeH0kKDPhP5tE2gSnSjS8jFKHnGVoDLpYoVoewOPcwcumPICZBSQJqna2trX4Q
VChD0rx06lSrkwpFEJbyD+P62G1Mh5yfS95B0pPS3TiKWRSuhxkUX5lvAnuyZGT2Kh46uXHqiS2o
WOBc2nR8bQUStGeBOZnX4COvBhSYP3AT6pancnOZL/0ECTo+Re8FK+zmEeddKjdFXP4hSTilR7aH
3fWzTA+jKJhQStDwyxEziKk+hAFLMkoY9D6XtobwKULV3vAFZ5RuwrCdN2V7Yecf81E7RBi787/d
enOUvoiSSg26HTx49ErZ5awejBl802aE/EHBrLsKCvQzCmzRN2f0/jZgnpp/bLx4iCS87DVWxRMg
sqZ/SW/sOHCrdoS1hO5hINx1eg3rZzZEIWuMu8XnEEmFIK3v0qdhEHJGojSqDDBsudblvhCnlFbM
uWfKn0ZqWGUsOPPWKuShre5AyTO584ybDsSaTi6jjbIq1DAp2QRAmnQVgHDiFyP153PTALbJqni3
oMuiEZ2mJd21PhvM+lD67grU59gPSvXDvH6iZuR6vo/jM3bXT92FhjC/7yJkUIASZO6kK2ARYmF4
L2th7TSce6EAjgqiZkqNhNOnsZacbzNOvnhV+bxUWxE3JO+5Xf9RGAA/sGsXDoR3gdTSLtninx0d
3CIynceyMY6hMxt0roOXciywzbNH4GfTt8V09p30F4UtH8lr1ifI5ER5RQe+pW0Wvze39tk/qg75
enP6UL2S1uEYwVWuWJlNeH4okVBDd42NUlrzhRvOkGhvgkK2+ziDf3WR3o9e6hyvK9jZ/JEy+M6+
eQHACfQPTgTCzJYF4cBfCkJ7blM9GHw3m+/MtEmhUzx06tY1I6GXsUEzqKnzyoKpmzA1V4QrIvai
EufvrmVfodCNTRPou4IstfvOp3tMxJ4oiLGijOESOAe9zw+6s+gw/3KCvklrGhFWT09zvrXTu10w
bTXujfEj0PbVjVHpHUYyEFa+t68WKZUxlHdj2Sc2/HePWWuHtJXFv3fepbso7nhvadjx2z7s6fUR
iNJcInNQRtYjU0sagm4tCiTC8DvAonY2wGMno4qw+s9/3pOGY3+5ti3bSkqe+PtGPOSt37q6nM/J
xnhTxEudgupP6rKAuLVYgsAniASIbn1AHR0qd1pR3tTIcLYQ/6znEY5YuKPqyepQDMMYbX7f6Zqi
nUvEAWvNVAF9bMSoa6ZEtrHF/zvQ27dEWZuAeKEcjKCj5q2AiBYHTaeOuuo/1pTL4qymTxTR45wQ
qTc0zDrizqZxWxwz8zm8GpG+4rtTXc0zdICPgy4E+wRXdz9Fk1hSpcnvwVKEF/CwS358jBHCHeRt
unBVFd4JovC4HUNXV1fOoET4FdFpgt241agCfYT+R4D/5aBIU/Bqy+lvNwGRsMW9wRaTWNSph8zo
HEqsb51EwDTXRvMQk4MqV4XCEkM7kz/Q9+1c2ZPexGBLY2huSEdWPHYc0X1uSy4uFONzC9TtilqC
i5DEgs3x/MDiqjKmem266BD7lDWIeSrxf1MQVd3hmgMzZXaPPKwQVcAPSY0f6v+H/JBHFKaBusKw
Vrfhx5HTPd6dXAW1GKVL5Q8pQ0a8h9IM7iYDO/A20YP8cSY5ilvAL0qhSXh4/XJOPpNg5JE4xNiM
EQmaWKxt5lk7G/bgK5TL9jFC3mC3qXU4t4tA9VbtZ8M7GNXLnRqR3aJz5mQ8UTMMXEajXOArKhL6
3q5UUQx999au3RnyXdGWnWZaPZMG++ll/7yuPNf6QAzxMORsln8wRGw6Ln6TNIHxRZiY9mXYNos3
0src/nGnpKrZ+Lvi3RoAjAvTjuS1fQgZgwCrhowbeSoJtfH8ptUeCCKwW8e3sD2YfJRX0o5nrTV7
m9g5obFy6qKiIpwb5o9Gx4N3CDjX8ocj0ZyncjXDd7WqB0j6peUSGTg/VcF0uhZ3XvLBh4qR+DMJ
LDo4TagBrTN3DR2WHt7e4sKFeFtFYGXhCVx5ZGaQh70OIw0iJ98PnWWqRh4HZQiOxc3ZJhASWGp6
jzuq42QFuQTBpti70MjzuLGvRRa8fDvcMe4/fkeVxO9drYunRfH9RuGhugoKF6m1l6GHbo6mfBB1
dw/jKw4GgeXHOFesrl8uLS9gW/gAhnK52618tCAC5wah9mRTo69CW2dgJ1vJQebXDT1oqYuQZs4r
kNFrTESKYkEMjeFYawzCXuevX4biBGgexG/uO+xo4iBL6xdnwTF15tNtfr9hQy2VDTfbEn8rEX+o
OcT8EKZwwzlK88f1JqMJdSZzftdyg0HDcKk6V6t1HRo8sU7fexeB516UcAaMA7m5gFJterHhEVM5
F+tE5E+ZVBRp+C2SjotWK6kBV2gm1KgJVEXNCxsQ/2EpDAMI6Gv5wNv9HNhqNLlqgenjOSP1K7Rr
34MXd24hKb/fsh7ucrOkDu2pyAtlDBZu73jAM2dfqi3rQYqVajHP8kRMGCTB2gAqiMq0WExVzkiI
PEPx+ixrMm9J/3ABOTFx21t1okLZXXWLJEuSegdrGosgb6YNPAUyFvOdBIWxcCr7VvkLK+cpDbYS
pXeF7adsqRgx0zmd46ype3g4uTgNExS9AO4ChVl6ZEMqGK2/xb5wZvDjfBhInUwvhl0YK32/wAca
Sr/iTnaS+4zutasmVk/BWCuWF+pnItvYeDnUbuTTVo2uNy4bFapoYASYPvw2pHVAprvg/Z8WySOx
M1W0ucdCJRXTP0lor5ndaqf3xATa2YHE1X/drh9Gbb9PDG/K6YGo67U0EiqsdLb/2suij6auvOj5
yov6FaOnmq9B2SjrXVx8OeD9FAbw6I19WxxS1L7Cx19WIbBQC6Wn8ywWMrr6z5awqaR0GB7xZDNE
q06VCvCRlVI/yH93rTTSZ0UbJn+n16dRdp9G2Kb1hXMa84PDwAqkY3DRuFZnaht6wIarPMkhJWNt
zoIgtIgepguHRmCNjxNWdjC0j9im21SefiyJY6wXA7IgRZgJlNqU2PDyMFIfwR2SjcZE2W4oPMES
6SsiKxfE9xKTkVA1Yv22xR/FTlxZexO35JC25qlf2i97tomKtpPcCjmWIEYrWCt6x+GSi3IMm/y+
khtrfGI9kbLB+MAjkiBdE12R0k2XYE/RDkn8ASg+iEDDSBr9Ns9OSS9h4E4eqE7c0eD7GTX0gyMY
2gLb5GODfAN7AfSDmUqwR1KHPbHOjEppi2Uwpscmjw0rjQ6E6pUydgXUTuznCbcWE+B5MWW7CoEU
nv5pe7gGeZgTnKe5d7O31yqhy4ft+5o+5VoowPgFxZpzbQNoXk15rMxVwIIK/UcKs21I8Yoe6R3l
63FOTGUqubowR2JpCRzYhFcCvcafO2zf2VQqYt+9N3ygDmFGUDG9qcvtg/ZxdxKj96C1kZbQ58jk
2cf9P734QwJ7WUy+cNV4m7vV6wm7NrpNivgkk8em5XDBwkxdeiFDVPRgBMyrBggpyCooFUv+wcmb
axPw4ez51Krv13rzKru695MLRvdyNIaOlAq62WwPE1+fI7xqqmzQlnZ3pX84qZebOo85YFbk2jEw
bkPAT4v8eJX0yh7HRHANrkmc9JGPs8J8mxff1SYyuQyJrP4/sF/zD+O2yP8+wlfWf309x1HaUyzm
1jWSpxNWXyBdwjKxjiAiY8LlCaXs3RU6wSRvohIOlzDyN684Ev41oHUJQJCsbIm4Zw5kzQnnqP4X
8Ud1a9gqvCBSrJg+4Xo1a1Pe82mpc4SqbOQRb33W5J9Nnx4jqyGmyyUnPNRr3Z1ENaTJNKVp5NfI
GHsAwJQ2dSeYQ9KlIwAdLDo4wCaImn6+eenzuRra0DzwXnbfVPnta0TvIKDzGa0VQROVwr+pl2yM
SaYvL4b9AnPhMlNr1KKp7bqpX84LleqC3qKQd+4fmhd7a+L70916KwDITye3llDYS8FEKlORHmJj
mjrAeNLOcDu4m7IJbpJBdm27eRK5RVwbGchKJ1uje0zKm40n90oYSNJ8/wdXdNKj7sGPeXvuolzl
gDIJ0j+oXCHD6pT3NpRHciU2l8nu+1saHEI9l3ENmkgERVhhPKF8lpNEDlJPlf69ILYGGXxy/+W8
oGQLpxKJL2DYTHT1K845XYFGnlRm8zcv1PNGSj9YWbNlkhPoUz7dv/D+BLhdNBH+TLwxvv+2ylc3
sg82Okmaeqj/uk5Xab4IagRJ0UyIDAKbfldzOWdqnxjZk20rpfvljtH/nL4ny0B8IcAxPLEB4+q8
CsYD+EIGP1vAX9OjMGQorme19bM2GkHK6PVnRwTmH8exrw==
`protect end_protected
